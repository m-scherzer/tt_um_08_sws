MACRO digital_top
  CLASS BLOCK ;
  FOREIGN digital_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 131.150 BY 141.870 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.520 10.640 26.520 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.520 10.640 86.520 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.520 10.640 116.520 130.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.520 10.640 11.520 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.520 10.640 41.520 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 10.640 71.520 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.520 10.640 101.520 130.800 ;
    END
  END VPWR
  PIN i_dem_dis
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.000 123.040 ;
    END
  END i_dem_dis
  PIN i_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.000 52.320 ;
    END
  END i_reset
  PIN i_sys_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 2.000 87.680 ;
    END
  END i_sys_clk
  PIN o_cs_cell_hi[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 4.230 139.870 4.510 141.870 ;
    END
  END o_cs_cell_hi[0]
  PIN o_cs_cell_hi[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 10.670 139.870 10.950 141.870 ;
    END
  END o_cs_cell_hi[1]
  PIN o_cs_cell_hi[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 139.870 17.390 141.870 ;
    END
  END o_cs_cell_hi[2]
  PIN o_cs_cell_hi[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 23.550 139.870 23.830 141.870 ;
    END
  END o_cs_cell_hi[3]
  PIN o_cs_cell_hi[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 29.990 139.870 30.270 141.870 ;
    END
  END o_cs_cell_hi[4]
  PIN o_cs_cell_hi[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 139.870 36.710 141.870 ;
    END
  END o_cs_cell_hi[5]
  PIN o_cs_cell_hi[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 139.870 43.150 141.870 ;
    END
  END o_cs_cell_hi[6]
  PIN o_cs_cell_hi[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 49.310 139.870 49.590 141.870 ;
    END
  END o_cs_cell_hi[7]
  PIN o_cs_cell_hi[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 55.750 139.870 56.030 141.870 ;
    END
  END o_cs_cell_hi[8]
  PIN o_cs_cell_hi[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 139.870 62.470 141.870 ;
    END
  END o_cs_cell_hi[9]
  PIN o_cs_cell_lo[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 68.630 139.870 68.910 141.870 ;
    END
  END o_cs_cell_lo[0]
  PIN o_cs_cell_lo[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 75.070 139.870 75.350 141.870 ;
    END
  END o_cs_cell_lo[1]
  PIN o_cs_cell_lo[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 139.870 81.790 141.870 ;
    END
  END o_cs_cell_lo[2]
  PIN o_cs_cell_lo[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 87.950 139.870 88.230 141.870 ;
    END
  END o_cs_cell_lo[3]
  PIN o_cs_cell_lo[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 94.390 139.870 94.670 141.870 ;
    END
  END o_cs_cell_lo[4]
  PIN o_cs_cell_lo[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 100.830 139.870 101.110 141.870 ;
    END
  END o_cs_cell_lo[5]
  PIN o_cs_cell_lo[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 139.870 107.550 141.870 ;
    END
  END o_cs_cell_lo[6]
  PIN o_cs_cell_lo[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 113.710 139.870 113.990 141.870 ;
    END
  END o_cs_cell_lo[7]
  PIN o_cs_cell_lo[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 139.870 120.430 141.870 ;
    END
  END o_cs_cell_lo[8]
  PIN o_cs_cell_lo[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 139.870 126.870 141.870 ;
    END
  END o_cs_cell_lo[9]
  OBS
      LAYER pwell ;
        RECT 5.665 130.455 5.835 130.645 ;
        RECT 7.045 130.455 7.215 130.645 ;
        RECT 12.560 130.505 12.680 130.615 ;
        RECT 13.945 130.455 14.115 130.645 ;
        RECT 14.405 130.455 14.575 130.645 ;
        RECT 18.080 130.505 18.200 130.615 ;
        RECT 19.005 130.455 19.175 130.645 ;
        RECT 24.525 130.455 24.695 130.645 ;
        RECT 30.045 130.455 30.215 130.645 ;
        RECT 31.885 130.455 32.055 130.645 ;
        RECT 42.465 130.455 42.635 130.645 ;
        RECT 44.765 130.455 44.935 130.645 ;
        RECT 50.285 130.455 50.455 130.645 ;
        RECT 55.805 130.455 55.975 130.645 ;
        RECT 57.645 130.455 57.815 130.645 ;
        RECT 68.225 130.455 68.395 130.645 ;
        RECT 70.525 130.455 70.695 130.645 ;
        RECT 76.045 130.455 76.215 130.645 ;
        RECT 81.565 130.455 81.735 130.645 ;
        RECT 83.405 130.455 83.575 130.645 ;
        RECT 88.925 130.455 89.095 130.645 ;
        RECT 94.445 130.455 94.615 130.645 ;
        RECT 96.285 130.455 96.455 130.645 ;
        RECT 101.805 130.455 101.975 130.645 ;
        RECT 107.325 130.455 107.495 130.645 ;
        RECT 109.165 130.455 109.335 130.645 ;
        RECT 110.545 130.455 110.715 130.645 ;
        RECT 121.120 130.505 121.240 130.615 ;
        RECT 122.045 130.455 122.215 130.645 ;
        RECT 123.880 130.505 124.000 130.615 ;
        RECT 125.265 130.455 125.435 130.645 ;
        RECT 5.525 129.645 6.895 130.455 ;
        RECT 6.905 129.645 12.415 130.455 ;
        RECT 12.895 129.545 14.245 130.455 ;
        RECT 14.265 129.645 17.935 130.455 ;
        RECT 18.415 129.585 18.845 130.370 ;
        RECT 18.865 129.645 24.375 130.455 ;
        RECT 24.385 129.645 29.895 130.455 ;
        RECT 29.905 129.645 31.275 130.455 ;
        RECT 31.295 129.585 31.725 130.370 ;
        RECT 31.745 129.775 42.115 130.455 ;
        RECT 36.255 129.555 37.185 129.775 ;
        RECT 39.905 129.545 42.115 129.775 ;
        RECT 42.325 129.645 44.155 130.455 ;
        RECT 44.175 129.585 44.605 130.370 ;
        RECT 44.625 129.645 50.135 130.455 ;
        RECT 50.145 129.645 55.655 130.455 ;
        RECT 55.665 129.645 57.035 130.455 ;
        RECT 57.055 129.585 57.485 130.370 ;
        RECT 57.505 129.775 67.875 130.455 ;
        RECT 62.015 129.555 62.945 129.775 ;
        RECT 65.665 129.545 67.875 129.775 ;
        RECT 68.085 129.645 69.915 130.455 ;
        RECT 69.935 129.585 70.365 130.370 ;
        RECT 70.385 129.645 75.895 130.455 ;
        RECT 75.905 129.645 81.415 130.455 ;
        RECT 81.425 129.645 82.795 130.455 ;
        RECT 82.815 129.585 83.245 130.370 ;
        RECT 83.265 129.645 88.775 130.455 ;
        RECT 88.785 129.645 94.295 130.455 ;
        RECT 94.305 129.645 95.675 130.455 ;
        RECT 95.695 129.585 96.125 130.370 ;
        RECT 96.145 129.645 101.655 130.455 ;
        RECT 101.665 129.645 107.175 130.455 ;
        RECT 107.185 129.645 108.555 130.455 ;
        RECT 108.575 129.585 109.005 130.370 ;
        RECT 109.025 129.645 110.395 130.455 ;
        RECT 110.405 129.775 120.775 130.455 ;
        RECT 114.915 129.555 115.845 129.775 ;
        RECT 118.565 129.545 120.775 129.775 ;
        RECT 121.455 129.585 121.885 130.370 ;
        RECT 121.905 129.645 123.735 130.455 ;
        RECT 124.205 129.645 125.575 130.455 ;
      LAYER nwell ;
        RECT 5.330 126.425 125.770 129.255 ;
      LAYER pwell ;
        RECT 5.525 125.225 6.895 126.035 ;
        RECT 12.335 125.905 13.265 126.125 ;
        RECT 15.985 125.905 18.195 126.135 ;
        RECT 7.825 125.225 18.195 125.905 ;
        RECT 18.415 125.310 18.845 126.095 ;
        RECT 18.865 125.225 22.535 126.035 ;
        RECT 27.515 125.905 28.445 126.125 ;
        RECT 31.165 125.905 33.375 126.135 ;
        RECT 38.095 125.905 39.025 126.125 ;
        RECT 41.745 125.905 43.955 126.135 ;
        RECT 23.005 125.225 33.375 125.905 ;
        RECT 33.585 125.225 43.955 125.905 ;
        RECT 44.175 125.310 44.605 126.095 ;
        RECT 44.625 125.225 46.455 126.035 ;
        RECT 46.475 125.225 47.825 126.135 ;
        RECT 53.275 125.905 54.205 126.125 ;
        RECT 56.925 125.905 59.135 126.135 ;
        RECT 63.855 125.905 64.785 126.125 ;
        RECT 67.505 125.905 69.715 126.135 ;
        RECT 48.765 125.225 59.135 125.905 ;
        RECT 59.345 125.225 69.715 125.905 ;
        RECT 69.935 125.310 70.365 126.095 ;
        RECT 70.385 125.225 73.135 126.035 ;
        RECT 78.115 125.905 79.045 126.125 ;
        RECT 81.765 125.905 83.975 126.135 ;
        RECT 88.695 125.905 89.625 126.125 ;
        RECT 92.345 125.905 94.555 126.135 ;
        RECT 73.605 125.225 83.975 125.905 ;
        RECT 84.185 125.225 94.555 125.905 ;
        RECT 95.695 125.310 96.125 126.095 ;
        RECT 100.655 125.905 101.585 126.125 ;
        RECT 104.305 125.905 106.515 126.135 ;
        RECT 111.235 125.905 112.165 126.125 ;
        RECT 114.885 125.905 117.095 126.135 ;
        RECT 96.145 125.225 106.515 125.905 ;
        RECT 106.725 125.225 117.095 125.905 ;
        RECT 117.305 125.225 120.975 126.035 ;
        RECT 121.455 125.310 121.885 126.095 ;
        RECT 121.905 125.225 123.735 126.035 ;
        RECT 124.205 125.225 125.575 126.035 ;
        RECT 5.665 125.015 5.835 125.225 ;
        RECT 7.055 125.070 7.215 125.180 ;
        RECT 7.965 125.035 8.135 125.225 ;
        RECT 17.165 125.015 17.335 125.205 ;
        RECT 18.545 125.015 18.715 125.205 ;
        RECT 19.005 125.175 19.175 125.225 ;
        RECT 19.000 125.065 19.175 125.175 ;
        RECT 19.005 125.035 19.175 125.065 ;
        RECT 19.465 125.015 19.635 125.205 ;
        RECT 22.680 125.065 22.800 125.175 ;
        RECT 23.145 125.035 23.315 125.225 ;
        RECT 30.965 125.015 31.135 125.205 ;
        RECT 31.885 125.015 32.055 125.205 ;
        RECT 33.725 125.035 33.895 125.225 ;
        RECT 35.565 125.015 35.735 125.205 ;
        RECT 36.945 125.015 37.115 125.205 ;
        RECT 39.700 125.065 39.820 125.175 ;
        RECT 41.085 125.015 41.255 125.205 ;
        RECT 41.545 125.015 41.715 125.205 ;
        RECT 44.765 125.035 44.935 125.225 ;
        RECT 46.605 125.035 46.775 125.225 ;
        RECT 47.995 125.070 48.155 125.180 ;
        RECT 48.905 125.035 49.075 125.225 ;
        RECT 52.125 125.015 52.295 125.205 ;
        RECT 53.505 125.015 53.675 125.205 ;
        RECT 55.805 125.015 55.975 125.205 ;
        RECT 56.275 125.060 56.435 125.170 ;
        RECT 57.640 125.065 57.760 125.175 ;
        RECT 58.105 125.015 58.275 125.205 ;
        RECT 59.485 125.015 59.655 125.225 ;
        RECT 60.865 125.015 61.035 125.205 ;
        RECT 66.385 125.015 66.555 125.205 ;
        RECT 67.765 125.015 67.935 125.205 ;
        RECT 70.525 125.035 70.695 125.225 ;
        RECT 73.280 125.065 73.400 125.175 ;
        RECT 73.745 125.035 73.915 125.225 ;
        RECT 79.265 125.015 79.435 125.205 ;
        RECT 80.645 125.015 80.815 125.205 ;
        RECT 81.105 125.015 81.275 125.205 ;
        RECT 83.405 125.015 83.575 125.205 ;
        RECT 84.325 125.035 84.495 125.225 ;
        RECT 85.245 125.015 85.415 125.205 ;
        RECT 86.620 125.065 86.740 125.175 ;
        RECT 87.085 125.015 87.255 125.205 ;
        RECT 94.915 125.070 95.075 125.180 ;
        RECT 96.285 125.035 96.455 125.225 ;
        RECT 97.665 125.015 97.835 125.205 ;
        RECT 99.045 125.015 99.215 125.205 ;
        RECT 104.560 125.065 104.680 125.175 ;
        RECT 105.025 125.015 105.195 125.205 ;
        RECT 106.415 125.060 106.575 125.170 ;
        RECT 106.865 125.035 107.035 125.225 ;
        RECT 107.325 125.015 107.495 125.205 ;
        RECT 109.165 125.015 109.335 125.205 ;
        RECT 117.445 125.035 117.615 125.225 ;
        RECT 120.665 125.015 120.835 125.205 ;
        RECT 121.125 125.175 121.295 125.205 ;
        RECT 121.120 125.065 121.295 125.175 ;
        RECT 121.125 125.015 121.295 125.065 ;
        RECT 122.045 125.035 122.215 125.225 ;
        RECT 122.505 125.015 122.675 125.205 ;
        RECT 123.880 125.065 124.000 125.175 ;
        RECT 125.265 125.015 125.435 125.225 ;
        RECT 5.525 124.205 6.895 125.015 ;
        RECT 7.105 124.335 17.475 125.015 ;
        RECT 7.105 124.105 9.315 124.335 ;
        RECT 12.035 124.115 12.965 124.335 ;
        RECT 17.495 124.105 18.845 125.015 ;
        RECT 19.325 124.335 29.695 125.015 ;
        RECT 23.835 124.115 24.765 124.335 ;
        RECT 27.485 124.105 29.695 124.335 ;
        RECT 29.915 124.105 31.265 125.015 ;
        RECT 31.295 124.145 31.725 124.930 ;
        RECT 31.745 124.205 35.415 125.015 ;
        RECT 35.435 124.105 36.785 125.015 ;
        RECT 36.805 124.205 39.555 125.015 ;
        RECT 40.035 124.105 41.385 125.015 ;
        RECT 41.405 124.335 51.775 125.015 ;
        RECT 45.915 124.115 46.845 124.335 ;
        RECT 49.565 124.105 51.775 124.335 ;
        RECT 51.985 124.205 53.355 125.015 ;
        RECT 53.375 124.105 54.725 125.015 ;
        RECT 54.745 124.235 56.115 125.015 ;
        RECT 57.055 124.145 57.485 124.930 ;
        RECT 57.965 124.235 59.335 125.015 ;
        RECT 59.355 124.105 60.705 125.015 ;
        RECT 60.725 124.205 66.235 125.015 ;
        RECT 66.245 124.205 67.615 125.015 ;
        RECT 67.625 124.335 77.995 125.015 ;
        RECT 72.135 124.115 73.065 124.335 ;
        RECT 75.785 124.105 77.995 124.335 ;
        RECT 78.215 124.105 79.565 125.015 ;
        RECT 79.595 124.105 80.945 125.015 ;
        RECT 80.965 124.205 82.795 125.015 ;
        RECT 82.815 124.145 83.245 124.930 ;
        RECT 83.265 124.205 85.095 125.015 ;
        RECT 85.115 124.105 86.465 125.015 ;
        RECT 86.945 124.335 97.315 125.015 ;
        RECT 91.455 124.115 92.385 124.335 ;
        RECT 95.105 124.105 97.315 124.335 ;
        RECT 97.535 124.105 98.885 125.015 ;
        RECT 98.905 124.205 104.415 125.015 ;
        RECT 104.895 124.105 106.245 125.015 ;
        RECT 107.195 124.105 108.545 125.015 ;
        RECT 108.575 124.145 109.005 124.930 ;
        RECT 109.025 124.335 119.395 125.015 ;
        RECT 113.535 124.115 114.465 124.335 ;
        RECT 117.185 124.105 119.395 124.335 ;
        RECT 119.615 124.105 120.965 125.015 ;
        RECT 120.995 124.105 122.345 125.015 ;
        RECT 122.365 124.205 124.195 125.015 ;
        RECT 124.205 124.205 125.575 125.015 ;
      LAYER nwell ;
        RECT 5.330 120.985 125.770 123.815 ;
      LAYER pwell ;
        RECT 5.525 119.785 6.895 120.595 ;
        RECT 7.105 120.465 9.315 120.695 ;
        RECT 12.035 120.465 12.965 120.685 ;
        RECT 7.105 119.785 17.475 120.465 ;
        RECT 18.415 119.870 18.845 120.655 ;
        RECT 18.865 119.785 20.695 120.595 ;
        RECT 21.165 119.785 22.535 120.565 ;
        RECT 23.465 119.785 24.835 120.565 ;
        RECT 24.855 119.785 26.205 120.695 ;
        RECT 26.225 119.785 27.595 120.595 ;
        RECT 27.605 119.785 28.975 120.565 ;
        RECT 28.985 119.785 34.495 120.595 ;
        RECT 34.505 119.785 35.875 120.565 ;
        RECT 35.885 119.785 39.555 120.595 ;
        RECT 40.485 119.785 41.855 120.565 ;
        RECT 41.865 119.785 43.695 120.595 ;
        RECT 44.175 119.870 44.605 120.655 ;
        RECT 45.545 119.785 46.915 120.565 ;
        RECT 46.925 119.785 52.435 120.595 ;
        RECT 52.585 119.785 55.195 120.695 ;
        RECT 55.205 119.785 57.955 120.595 ;
        RECT 58.435 119.785 59.785 120.695 ;
        RECT 59.805 119.785 65.315 120.595 ;
        RECT 65.325 119.785 67.155 120.595 ;
        RECT 67.625 119.785 68.995 120.565 ;
        RECT 69.935 119.870 70.365 120.655 ;
        RECT 70.395 119.785 71.745 120.695 ;
        RECT 72.825 119.785 75.435 120.695 ;
        RECT 75.445 119.785 76.815 120.565 ;
        RECT 76.825 119.785 78.655 120.595 ;
        RECT 78.665 119.785 80.035 120.565 ;
        RECT 80.045 119.785 83.715 120.595 ;
        RECT 84.185 119.785 85.555 120.565 ;
        RECT 85.565 119.785 89.235 120.595 ;
        RECT 89.245 119.785 90.615 120.565 ;
        RECT 90.625 119.785 91.995 120.595 ;
        RECT 92.005 119.785 93.375 120.565 ;
        RECT 93.395 119.785 94.745 120.695 ;
        RECT 95.695 119.870 96.125 120.655 ;
        RECT 96.145 119.785 101.655 120.595 ;
        RECT 102.125 119.785 103.495 120.565 ;
        RECT 103.505 119.785 105.335 120.595 ;
        RECT 105.805 119.785 107.175 120.565 ;
        RECT 107.185 119.785 108.555 120.565 ;
        RECT 109.485 119.785 110.855 120.565 ;
        RECT 115.375 120.465 116.305 120.685 ;
        RECT 119.025 120.465 121.235 120.695 ;
        RECT 110.865 119.785 121.235 120.465 ;
        RECT 121.455 119.870 121.885 120.655 ;
        RECT 121.905 119.785 123.735 120.595 ;
        RECT 124.205 119.785 125.575 120.595 ;
        RECT 5.665 119.575 5.835 119.785 ;
        RECT 7.055 119.575 7.225 119.765 ;
        RECT 8.425 119.575 8.595 119.765 ;
        RECT 10.265 119.575 10.435 119.765 ;
        RECT 11.645 119.575 11.815 119.765 ;
        RECT 13.945 119.575 14.115 119.765 ;
        RECT 14.405 119.575 14.575 119.765 ;
        RECT 17.165 119.595 17.335 119.785 ;
        RECT 17.635 119.630 17.795 119.740 ;
        RECT 19.005 119.595 19.175 119.785 ;
        RECT 19.925 119.575 20.095 119.765 ;
        RECT 20.840 119.625 20.960 119.735 ;
        RECT 22.225 119.595 22.395 119.785 ;
        RECT 22.695 119.630 22.855 119.740 ;
        RECT 24.525 119.595 24.695 119.785 ;
        RECT 25.445 119.575 25.615 119.765 ;
        RECT 25.905 119.595 26.075 119.785 ;
        RECT 26.365 119.595 26.535 119.785 ;
        RECT 28.665 119.595 28.835 119.785 ;
        RECT 29.125 119.595 29.295 119.785 ;
        RECT 30.960 119.625 31.080 119.735 ;
        RECT 31.885 119.575 32.055 119.765 ;
        RECT 35.565 119.595 35.735 119.785 ;
        RECT 36.025 119.595 36.195 119.785 ;
        RECT 37.405 119.575 37.575 119.765 ;
        RECT 39.715 119.630 39.875 119.740 ;
        RECT 41.545 119.595 41.715 119.785 ;
        RECT 42.005 119.595 42.175 119.785 ;
        RECT 42.925 119.575 43.095 119.765 ;
        RECT 43.840 119.625 43.960 119.735 ;
        RECT 44.775 119.630 44.935 119.740 ;
        RECT 46.605 119.595 46.775 119.785 ;
        RECT 47.065 119.595 47.235 119.785 ;
        RECT 48.445 119.575 48.615 119.765 ;
        RECT 53.965 119.575 54.135 119.765 ;
        RECT 54.880 119.595 55.050 119.785 ;
        RECT 55.345 119.595 55.515 119.785 ;
        RECT 56.720 119.625 56.840 119.735 ;
        RECT 57.645 119.575 57.815 119.765 ;
        RECT 58.100 119.625 58.220 119.735 ;
        RECT 58.565 119.595 58.735 119.785 ;
        RECT 59.945 119.595 60.115 119.785 ;
        RECT 63.165 119.575 63.335 119.765 ;
        RECT 65.465 119.595 65.635 119.785 ;
        RECT 67.300 119.625 67.420 119.735 ;
        RECT 68.685 119.575 68.855 119.785 ;
        RECT 69.155 119.630 69.315 119.740 ;
        RECT 71.445 119.595 71.615 119.785 ;
        RECT 71.915 119.630 72.075 119.740 ;
        RECT 74.205 119.575 74.375 119.765 ;
        RECT 75.120 119.595 75.290 119.785 ;
        RECT 76.505 119.595 76.675 119.785 ;
        RECT 76.965 119.595 77.135 119.785 ;
        RECT 79.725 119.575 79.895 119.785 ;
        RECT 80.185 119.595 80.355 119.785 ;
        RECT 82.480 119.625 82.600 119.735 ;
        RECT 83.405 119.575 83.575 119.765 ;
        RECT 83.860 119.625 83.980 119.735 ;
        RECT 84.325 119.595 84.495 119.785 ;
        RECT 85.705 119.595 85.875 119.785 ;
        RECT 87.085 119.575 87.255 119.765 ;
        RECT 89.385 119.575 89.555 119.765 ;
        RECT 89.845 119.575 90.015 119.765 ;
        RECT 90.305 119.595 90.475 119.785 ;
        RECT 90.765 119.595 90.935 119.785 ;
        RECT 92.145 119.595 92.315 119.785 ;
        RECT 94.445 119.595 94.615 119.785 ;
        RECT 94.915 119.630 95.075 119.740 ;
        RECT 95.365 119.575 95.535 119.765 ;
        RECT 96.285 119.595 96.455 119.785 ;
        RECT 100.885 119.575 101.055 119.765 ;
        RECT 101.800 119.625 101.920 119.735 ;
        RECT 102.265 119.595 102.435 119.785 ;
        RECT 103.645 119.595 103.815 119.785 ;
        RECT 105.480 119.625 105.600 119.735 ;
        RECT 105.945 119.595 106.115 119.785 ;
        RECT 106.405 119.575 106.575 119.765 ;
        RECT 107.325 119.595 107.495 119.785 ;
        RECT 108.240 119.625 108.360 119.735 ;
        RECT 108.715 119.630 108.875 119.740 ;
        RECT 109.165 119.575 109.335 119.765 ;
        RECT 109.625 119.595 109.795 119.785 ;
        RECT 111.005 119.595 111.175 119.785 ;
        RECT 114.685 119.575 114.855 119.765 ;
        RECT 120.205 119.575 120.375 119.765 ;
        RECT 122.045 119.595 122.215 119.785 ;
        RECT 123.880 119.625 124.000 119.735 ;
        RECT 125.265 119.575 125.435 119.785 ;
        RECT 5.525 118.765 6.895 119.575 ;
        RECT 6.905 118.795 8.275 119.575 ;
        RECT 8.285 118.765 10.115 119.575 ;
        RECT 10.125 118.795 11.495 119.575 ;
        RECT 11.505 118.795 12.875 119.575 ;
        RECT 12.895 118.665 14.245 119.575 ;
        RECT 14.265 118.765 19.775 119.575 ;
        RECT 19.785 118.765 25.295 119.575 ;
        RECT 25.305 118.765 30.815 119.575 ;
        RECT 31.295 118.705 31.725 119.490 ;
        RECT 31.745 118.765 37.255 119.575 ;
        RECT 37.265 118.765 42.775 119.575 ;
        RECT 42.785 118.765 48.295 119.575 ;
        RECT 48.305 118.765 53.815 119.575 ;
        RECT 53.825 118.765 56.575 119.575 ;
        RECT 57.055 118.705 57.485 119.490 ;
        RECT 57.505 118.765 63.015 119.575 ;
        RECT 63.025 118.765 68.535 119.575 ;
        RECT 68.545 118.765 74.055 119.575 ;
        RECT 74.065 118.765 79.575 119.575 ;
        RECT 79.585 118.765 82.335 119.575 ;
        RECT 82.815 118.705 83.245 119.490 ;
        RECT 83.265 118.765 86.935 119.575 ;
        RECT 86.945 118.765 88.315 119.575 ;
        RECT 88.335 118.665 89.685 119.575 ;
        RECT 89.705 118.765 95.215 119.575 ;
        RECT 95.225 118.765 100.735 119.575 ;
        RECT 100.745 118.765 106.255 119.575 ;
        RECT 106.265 118.765 108.095 119.575 ;
        RECT 108.575 118.705 109.005 119.490 ;
        RECT 109.025 118.765 114.535 119.575 ;
        RECT 114.545 118.765 120.055 119.575 ;
        RECT 120.065 118.765 123.735 119.575 ;
        RECT 124.205 118.765 125.575 119.575 ;
      LAYER nwell ;
        RECT 5.330 115.545 125.770 118.375 ;
      LAYER pwell ;
        RECT 5.525 114.345 6.895 115.155 ;
        RECT 6.905 114.345 12.415 115.155 ;
        RECT 12.425 114.345 15.175 115.155 ;
        RECT 15.185 114.345 16.555 115.125 ;
        RECT 16.565 114.345 18.395 115.155 ;
        RECT 18.415 114.430 18.845 115.215 ;
        RECT 18.865 114.345 24.375 115.155 ;
        RECT 24.385 114.345 29.895 115.155 ;
        RECT 29.905 114.345 35.415 115.155 ;
        RECT 35.425 114.345 40.935 115.155 ;
        RECT 40.945 114.345 43.695 115.155 ;
        RECT 44.175 114.430 44.605 115.215 ;
        RECT 44.625 114.345 47.375 115.155 ;
        RECT 47.855 114.345 49.205 115.255 ;
        RECT 49.225 114.345 54.735 115.155 ;
        RECT 55.665 114.345 57.035 115.125 ;
        RECT 57.045 114.345 60.715 115.155 ;
        RECT 60.735 114.345 62.085 115.255 ;
        RECT 62.105 114.345 67.615 115.155 ;
        RECT 67.625 114.345 69.455 115.155 ;
        RECT 69.935 114.430 70.365 115.215 ;
        RECT 70.385 114.345 75.895 115.155 ;
        RECT 75.905 114.345 81.415 115.155 ;
        RECT 81.425 114.345 83.255 115.155 ;
        RECT 83.635 115.145 84.555 115.255 ;
        RECT 83.635 115.025 85.970 115.145 ;
        RECT 90.635 115.025 91.555 115.245 ;
        RECT 83.635 114.345 92.915 115.025 ;
        RECT 92.925 114.345 95.675 115.155 ;
        RECT 95.695 114.430 96.125 115.215 ;
        RECT 96.145 114.345 98.755 115.255 ;
        RECT 99.375 114.345 100.725 115.255 ;
        RECT 100.745 114.345 103.495 115.155 ;
        RECT 103.505 114.345 104.875 115.125 ;
        RECT 104.885 114.345 110.395 115.155 ;
        RECT 110.405 114.345 111.775 115.155 ;
        RECT 113.145 115.025 114.065 115.245 ;
        RECT 120.145 115.145 121.065 115.255 ;
        RECT 118.730 115.025 121.065 115.145 ;
        RECT 111.785 114.345 121.065 115.025 ;
        RECT 121.455 114.430 121.885 115.215 ;
        RECT 121.905 114.345 123.735 115.155 ;
        RECT 124.205 114.345 125.575 115.155 ;
        RECT 5.665 114.135 5.835 114.345 ;
        RECT 7.045 114.135 7.215 114.345 ;
        RECT 10.735 114.180 10.895 114.290 ;
        RECT 11.645 114.135 11.815 114.325 ;
        RECT 12.565 114.155 12.735 114.345 ;
        RECT 16.245 114.155 16.415 114.345 ;
        RECT 16.705 114.155 16.875 114.345 ;
        RECT 19.005 114.155 19.175 114.345 ;
        RECT 21.300 114.185 21.420 114.295 ;
        RECT 21.765 114.135 21.935 114.325 ;
        RECT 24.525 114.155 24.695 114.345 ;
        RECT 30.045 114.155 30.215 114.345 ;
        RECT 32.160 114.135 32.330 114.325 ;
        RECT 35.565 114.155 35.735 114.345 ;
        RECT 36.945 114.135 37.115 114.325 ;
        RECT 37.405 114.135 37.575 114.325 ;
        RECT 38.785 114.135 38.955 114.325 ;
        RECT 41.085 114.135 41.255 114.345 ;
        RECT 41.545 114.155 41.715 114.325 ;
        RECT 43.840 114.185 43.960 114.295 ;
        RECT 44.765 114.155 44.935 114.345 ;
        RECT 47.520 114.185 47.640 114.295 ;
        RECT 47.985 114.155 48.155 114.345 ;
        RECT 49.365 114.155 49.535 114.345 ;
        RECT 52.585 114.135 52.755 114.325 ;
        RECT 54.895 114.190 55.055 114.300 ;
        RECT 55.805 114.155 55.975 114.345 ;
        RECT 56.450 114.135 56.620 114.325 ;
        RECT 57.185 114.155 57.355 114.345 ;
        RECT 60.865 114.155 61.035 114.345 ;
        RECT 62.245 114.155 62.415 114.345 ;
        RECT 66.845 114.135 67.015 114.325 ;
        RECT 67.305 114.135 67.475 114.325 ;
        RECT 67.765 114.155 67.935 114.345 ;
        RECT 69.600 114.185 69.720 114.295 ;
        RECT 70.065 114.135 70.235 114.325 ;
        RECT 70.525 114.155 70.695 114.345 ;
        RECT 76.045 114.155 76.215 114.345 ;
        RECT 79.725 114.135 79.895 114.325 ;
        RECT 81.565 114.155 81.735 114.345 ;
        RECT 82.480 114.185 82.600 114.295 ;
        RECT 83.405 114.135 83.575 114.325 ;
        RECT 88.190 114.135 88.360 114.325 ;
        RECT 88.925 114.135 89.095 114.325 ;
        RECT 90.305 114.135 90.475 114.325 ;
        RECT 92.140 114.185 92.260 114.295 ;
        RECT 92.605 114.135 92.775 114.345 ;
        RECT 93.065 114.155 93.235 114.345 ;
        RECT 93.985 114.135 94.155 114.325 ;
        RECT 96.290 114.155 96.460 114.345 ;
        RECT 99.040 114.185 99.160 114.295 ;
        RECT 100.425 114.155 100.595 114.345 ;
        RECT 100.885 114.155 101.055 114.345 ;
        RECT 103.645 114.155 103.815 114.345 ;
        RECT 103.920 114.135 104.090 114.325 ;
        RECT 105.025 114.155 105.195 114.345 ;
        RECT 107.795 114.180 107.955 114.290 ;
        RECT 109.165 114.135 109.335 114.325 ;
        RECT 110.545 114.155 110.715 114.345 ;
        RECT 111.005 114.135 111.175 114.325 ;
        RECT 111.925 114.155 112.095 114.345 ;
        RECT 120.665 114.135 120.835 114.325 ;
        RECT 122.045 114.155 122.215 114.345 ;
        RECT 123.880 114.185 124.000 114.295 ;
        RECT 125.265 114.135 125.435 114.345 ;
        RECT 5.525 113.325 6.895 114.135 ;
        RECT 6.905 113.325 10.575 114.135 ;
        RECT 11.505 113.455 20.785 114.135 ;
        RECT 21.625 113.455 30.905 114.135 ;
        RECT 12.865 113.235 13.785 113.455 ;
        RECT 18.450 113.335 20.785 113.455 ;
        RECT 19.865 113.225 20.785 113.335 ;
        RECT 22.985 113.235 23.905 113.455 ;
        RECT 28.570 113.335 30.905 113.455 ;
        RECT 29.985 113.225 30.905 113.335 ;
        RECT 31.295 113.265 31.725 114.050 ;
        RECT 31.745 113.455 35.645 114.135 ;
        RECT 31.745 113.225 32.675 113.455 ;
        RECT 35.885 113.355 37.255 114.135 ;
        RECT 37.265 113.325 38.635 114.135 ;
        RECT 38.645 113.355 40.015 114.135 ;
        RECT 40.035 113.225 41.385 114.135 ;
        RECT 41.870 113.455 43.235 114.135 ;
        RECT 43.615 113.455 52.895 114.135 ;
        RECT 53.135 113.455 57.035 114.135 ;
        RECT 43.615 113.335 45.950 113.455 ;
        RECT 43.615 113.225 44.535 113.335 ;
        RECT 50.615 113.235 51.535 113.455 ;
        RECT 56.105 113.225 57.035 113.455 ;
        RECT 57.055 113.265 57.485 114.050 ;
        RECT 57.875 113.455 67.155 114.135 ;
        RECT 57.875 113.335 60.210 113.455 ;
        RECT 57.875 113.225 58.795 113.335 ;
        RECT 64.875 113.235 65.795 113.455 ;
        RECT 67.165 113.325 69.915 114.135 ;
        RECT 69.925 113.455 79.205 114.135 ;
        RECT 71.285 113.235 72.205 113.455 ;
        RECT 76.870 113.335 79.205 113.455 ;
        RECT 78.285 113.225 79.205 113.335 ;
        RECT 79.585 113.325 82.335 114.135 ;
        RECT 82.815 113.265 83.245 114.050 ;
        RECT 83.275 113.225 84.625 114.135 ;
        RECT 84.875 113.455 88.775 114.135 ;
        RECT 87.845 113.225 88.775 113.455 ;
        RECT 88.785 113.355 90.155 114.135 ;
        RECT 90.165 113.325 91.995 114.135 ;
        RECT 92.465 113.355 93.835 114.135 ;
        RECT 93.845 113.455 103.125 114.135 ;
        RECT 95.205 113.235 96.125 113.455 ;
        RECT 100.790 113.335 103.125 113.455 ;
        RECT 102.205 113.225 103.125 113.335 ;
        RECT 103.505 113.455 107.405 114.135 ;
        RECT 103.505 113.225 104.435 113.455 ;
        RECT 108.575 113.265 109.005 114.050 ;
        RECT 109.025 113.325 110.855 114.135 ;
        RECT 110.865 113.455 120.145 114.135 ;
        RECT 112.225 113.235 113.145 113.455 ;
        RECT 117.810 113.335 120.145 113.455 ;
        RECT 119.225 113.225 120.145 113.335 ;
        RECT 120.525 113.325 124.195 114.135 ;
        RECT 124.205 113.325 125.575 114.135 ;
      LAYER nwell ;
        RECT 5.330 110.105 125.770 112.935 ;
      LAYER pwell ;
        RECT 5.525 108.905 6.895 109.715 ;
        RECT 6.905 108.905 12.415 109.715 ;
        RECT 12.425 108.905 16.095 109.715 ;
        RECT 16.115 108.905 17.465 109.815 ;
        RECT 18.415 108.990 18.845 109.775 ;
        RECT 18.865 109.585 19.795 109.815 ;
        RECT 18.865 108.905 22.765 109.585 ;
        RECT 23.465 108.905 24.835 109.685 ;
        RECT 35.405 109.585 36.325 109.805 ;
        RECT 42.405 109.705 43.325 109.815 ;
        RECT 40.990 109.585 43.325 109.705 ;
        RECT 24.930 108.905 34.035 109.585 ;
        RECT 34.045 108.905 43.325 109.585 ;
        RECT 44.175 108.990 44.605 109.775 ;
        RECT 55.645 109.585 56.565 109.805 ;
        RECT 62.645 109.705 63.565 109.815 ;
        RECT 61.230 109.585 63.565 109.705 ;
        RECT 44.710 108.905 53.815 109.585 ;
        RECT 54.285 108.905 63.565 109.585 ;
        RECT 63.955 108.905 65.305 109.815 ;
        RECT 65.325 108.905 68.075 109.715 ;
        RECT 68.545 108.905 69.915 109.685 ;
        RECT 69.935 108.990 70.365 109.775 ;
        RECT 71.745 109.585 72.665 109.805 ;
        RECT 78.745 109.705 79.665 109.815 ;
        RECT 77.330 109.585 79.665 109.705 ;
        RECT 81.405 109.585 82.325 109.805 ;
        RECT 88.405 109.705 89.325 109.815 ;
        RECT 86.990 109.585 89.325 109.705 ;
        RECT 70.385 108.905 79.665 109.585 ;
        RECT 80.045 108.905 89.325 109.585 ;
        RECT 89.705 108.905 91.795 109.715 ;
        RECT 92.465 108.905 95.215 109.715 ;
        RECT 95.695 108.990 96.125 109.775 ;
        RECT 96.145 109.585 97.075 109.815 ;
        RECT 96.145 108.905 100.045 109.585 ;
        RECT 100.285 108.905 103.955 109.715 ;
        RECT 105.325 109.585 106.245 109.805 ;
        RECT 112.325 109.705 113.245 109.815 ;
        RECT 110.910 109.585 113.245 109.705 ;
        RECT 103.965 108.905 113.245 109.585 ;
        RECT 113.625 109.585 114.555 109.815 ;
        RECT 113.625 108.905 117.525 109.585 ;
        RECT 117.775 108.905 119.125 109.815 ;
        RECT 119.145 108.905 120.515 109.685 ;
        RECT 121.455 108.990 121.885 109.775 ;
        RECT 121.915 108.905 123.265 109.815 ;
        RECT 124.205 108.905 125.575 109.715 ;
        RECT 5.665 108.695 5.835 108.905 ;
        RECT 7.045 108.695 7.215 108.905 ;
        RECT 10.725 108.695 10.895 108.885 ;
        RECT 12.565 108.715 12.735 108.905 ;
        RECT 13.025 108.695 13.195 108.885 ;
        RECT 14.405 108.695 14.575 108.885 ;
        RECT 14.860 108.745 14.980 108.855 ;
        RECT 16.245 108.695 16.415 108.905 ;
        RECT 16.980 108.695 17.150 108.885 ;
        RECT 17.635 108.750 17.795 108.860 ;
        RECT 19.280 108.715 19.450 108.905 ;
        RECT 20.845 108.695 21.015 108.885 ;
        RECT 23.140 108.745 23.260 108.855 ;
        RECT 23.605 108.695 23.775 108.885 ;
        RECT 24.525 108.715 24.695 108.905 ;
        RECT 24.985 108.695 25.155 108.885 ;
        RECT 27.740 108.745 27.860 108.855 ;
        RECT 29.125 108.695 29.295 108.885 ;
        RECT 29.585 108.695 29.755 108.885 ;
        RECT 30.960 108.745 31.080 108.855 ;
        RECT 31.885 108.695 32.055 108.885 ;
        RECT 33.725 108.715 33.895 108.905 ;
        RECT 34.185 108.715 34.355 108.905 ;
        RECT 37.130 108.695 37.300 108.885 ;
        RECT 37.860 108.745 37.980 108.855 ;
        RECT 38.325 108.695 38.495 108.885 ;
        RECT 43.840 108.745 43.960 108.855 ;
        RECT 48.905 108.695 49.075 108.885 ;
        RECT 49.365 108.695 49.535 108.885 ;
        RECT 51.020 108.695 51.190 108.885 ;
        RECT 53.505 108.715 53.675 108.905 ;
        RECT 53.960 108.745 54.080 108.855 ;
        RECT 54.425 108.715 54.595 108.905 ;
        RECT 54.880 108.745 55.000 108.855 ;
        RECT 56.265 108.695 56.435 108.885 ;
        RECT 56.720 108.745 56.840 108.855 ;
        RECT 57.920 108.695 58.090 108.885 ;
        RECT 61.785 108.695 61.955 108.885 ;
        RECT 65.005 108.715 65.175 108.905 ;
        RECT 65.465 108.715 65.635 108.905 ;
        RECT 67.305 108.695 67.475 108.885 ;
        RECT 68.220 108.745 68.340 108.855 ;
        RECT 68.685 108.715 68.855 108.905 ;
        RECT 69.140 108.745 69.260 108.855 ;
        RECT 69.605 108.695 69.775 108.885 ;
        RECT 70.525 108.715 70.695 108.905 ;
        RECT 70.995 108.740 71.155 108.850 ;
        RECT 71.905 108.695 72.075 108.885 ;
        RECT 73.295 108.740 73.455 108.850 ;
        RECT 74.480 108.695 74.650 108.885 ;
        RECT 79.265 108.695 79.435 108.885 ;
        RECT 79.725 108.695 79.895 108.885 ;
        RECT 80.185 108.715 80.355 108.905 ;
        RECT 81.105 108.695 81.275 108.885 ;
        RECT 83.405 108.695 83.575 108.885 ;
        RECT 89.845 108.715 90.015 108.905 ;
        RECT 92.605 108.695 92.775 108.905 ;
        RECT 95.360 108.745 95.480 108.855 ;
        RECT 95.825 108.695 95.995 108.885 ;
        RECT 96.560 108.715 96.730 108.905 ;
        RECT 100.425 108.715 100.595 108.905 ;
        RECT 104.105 108.715 104.275 108.905 ;
        RECT 106.405 108.695 106.575 108.885 ;
        RECT 106.865 108.695 107.035 108.885 ;
        RECT 110.085 108.695 110.255 108.885 ;
        RECT 110.545 108.695 110.715 108.885 ;
        RECT 112.845 108.695 113.015 108.885 ;
        RECT 113.305 108.695 113.475 108.885 ;
        RECT 114.040 108.715 114.210 108.905 ;
        RECT 115.140 108.745 115.260 108.855 ;
        RECT 118.825 108.715 118.995 108.905 ;
        RECT 119.010 108.695 119.180 108.885 ;
        RECT 119.745 108.695 119.915 108.885 ;
        RECT 120.205 108.715 120.375 108.905 ;
        RECT 120.675 108.750 120.835 108.860 ;
        RECT 122.045 108.715 122.215 108.905 ;
        RECT 123.435 108.740 123.595 108.860 ;
        RECT 125.265 108.695 125.435 108.905 ;
        RECT 5.525 107.885 6.895 108.695 ;
        RECT 6.905 107.885 10.575 108.695 ;
        RECT 10.585 107.885 11.955 108.695 ;
        RECT 11.965 107.915 13.335 108.695 ;
        RECT 13.345 107.915 14.715 108.695 ;
        RECT 15.195 107.785 16.545 108.695 ;
        RECT 16.565 108.015 20.465 108.695 ;
        RECT 16.565 107.785 17.495 108.015 ;
        RECT 20.705 107.885 23.455 108.695 ;
        RECT 23.465 107.915 24.835 108.695 ;
        RECT 24.845 108.015 27.585 108.695 ;
        RECT 28.075 107.785 29.425 108.695 ;
        RECT 29.455 107.785 30.805 108.695 ;
        RECT 31.295 107.825 31.725 108.610 ;
        RECT 31.745 107.885 33.575 108.695 ;
        RECT 33.815 108.015 37.715 108.695 ;
        RECT 38.185 108.015 47.465 108.695 ;
        RECT 36.785 107.785 37.715 108.015 ;
        RECT 39.545 107.795 40.465 108.015 ;
        RECT 45.130 107.895 47.465 108.015 ;
        RECT 46.545 107.785 47.465 107.895 ;
        RECT 47.855 107.785 49.205 108.695 ;
        RECT 49.225 107.915 50.595 108.695 ;
        RECT 50.605 108.015 54.505 108.695 ;
        RECT 50.605 107.785 51.535 108.015 ;
        RECT 55.205 107.915 56.575 108.695 ;
        RECT 57.055 107.825 57.485 108.610 ;
        RECT 57.505 108.015 61.405 108.695 ;
        RECT 57.505 107.785 58.435 108.015 ;
        RECT 61.645 107.885 67.155 108.695 ;
        RECT 67.165 107.885 68.995 108.695 ;
        RECT 69.465 107.915 70.835 108.695 ;
        RECT 71.775 107.785 73.125 108.695 ;
        RECT 74.065 108.015 77.965 108.695 ;
        RECT 74.065 107.785 74.995 108.015 ;
        RECT 78.215 107.785 79.565 108.695 ;
        RECT 79.585 107.915 80.955 108.695 ;
        RECT 80.965 107.885 82.795 108.695 ;
        RECT 82.815 107.825 83.245 108.610 ;
        RECT 83.265 108.015 92.370 108.695 ;
        RECT 92.465 107.885 95.215 108.695 ;
        RECT 95.685 108.015 104.965 108.695 ;
        RECT 97.045 107.795 97.965 108.015 ;
        RECT 102.630 107.895 104.965 108.015 ;
        RECT 104.045 107.785 104.965 107.895 ;
        RECT 105.355 107.785 106.705 108.695 ;
        RECT 106.725 107.885 108.555 108.695 ;
        RECT 108.575 107.825 109.005 108.610 ;
        RECT 109.035 107.785 110.385 108.695 ;
        RECT 110.405 107.885 111.775 108.695 ;
        RECT 111.785 107.915 113.155 108.695 ;
        RECT 113.165 107.885 114.995 108.695 ;
        RECT 115.695 108.015 119.595 108.695 ;
        RECT 118.665 107.785 119.595 108.015 ;
        RECT 119.605 107.885 123.275 108.695 ;
        RECT 124.205 107.885 125.575 108.695 ;
      LAYER nwell ;
        RECT 5.330 104.665 125.770 107.495 ;
      LAYER pwell ;
        RECT 5.525 103.465 6.895 104.275 ;
        RECT 6.905 103.465 8.275 104.275 ;
        RECT 9.645 104.145 10.565 104.365 ;
        RECT 16.645 104.265 17.565 104.375 ;
        RECT 15.230 104.145 17.565 104.265 ;
        RECT 8.285 103.465 17.565 104.145 ;
        RECT 18.415 103.550 18.845 104.335 ;
        RECT 18.865 104.145 19.795 104.375 ;
        RECT 18.865 103.465 22.765 104.145 ;
        RECT 23.005 103.465 24.835 104.275 ;
        RECT 26.205 104.145 27.125 104.365 ;
        RECT 33.205 104.265 34.125 104.375 ;
        RECT 31.790 104.145 34.125 104.265 ;
        RECT 24.845 103.465 34.125 104.145 ;
        RECT 34.505 103.465 40.015 104.275 ;
        RECT 40.025 103.465 43.695 104.275 ;
        RECT 44.175 103.550 44.605 104.335 ;
        RECT 44.625 104.145 45.555 104.375 ;
        RECT 57.725 104.285 58.675 104.375 ;
        RECT 44.625 103.465 48.525 104.145 ;
        RECT 48.765 103.465 54.275 104.275 ;
        RECT 54.285 103.465 56.115 104.275 ;
        RECT 56.745 103.465 58.675 104.285 ;
        RECT 59.085 104.285 60.035 104.375 ;
        RECT 59.085 103.465 61.015 104.285 ;
        RECT 61.185 103.465 66.695 104.275 ;
        RECT 66.705 103.465 69.455 104.275 ;
        RECT 69.935 103.550 70.365 104.335 ;
        RECT 71.305 104.145 72.235 104.375 ;
        RECT 71.305 103.465 75.205 104.145 ;
        RECT 75.445 103.465 80.955 104.275 ;
        RECT 80.965 103.465 82.795 104.275 ;
        RECT 83.265 104.145 84.195 104.375 ;
        RECT 89.445 104.285 90.395 104.375 ;
        RECT 91.745 104.285 92.695 104.375 ;
        RECT 83.265 103.465 87.165 104.145 ;
        RECT 87.405 103.465 89.235 104.275 ;
        RECT 89.445 103.465 91.375 104.285 ;
        RECT 91.745 103.465 93.675 104.285 ;
        RECT 93.845 103.465 95.675 104.275 ;
        RECT 95.695 103.550 96.125 104.335 ;
        RECT 96.145 103.465 97.515 104.245 ;
        RECT 97.525 104.145 98.455 104.375 ;
        RECT 97.525 103.465 101.425 104.145 ;
        RECT 101.665 103.465 103.035 104.275 ;
        RECT 103.045 103.465 112.150 104.145 ;
        RECT 112.245 103.465 117.755 104.275 ;
        RECT 117.765 103.465 121.435 104.275 ;
        RECT 121.455 103.550 121.885 104.335 ;
        RECT 121.905 103.465 123.735 104.275 ;
        RECT 124.205 103.465 125.575 104.275 ;
        RECT 5.665 103.255 5.835 103.465 ;
        RECT 7.045 103.255 7.215 103.465 ;
        RECT 8.425 103.275 8.595 103.465 ;
        RECT 9.800 103.305 9.920 103.415 ;
        RECT 10.265 103.255 10.435 103.445 ;
        RECT 18.080 103.305 18.200 103.415 ;
        RECT 19.280 103.275 19.450 103.465 ;
        RECT 19.925 103.255 20.095 103.445 ;
        RECT 23.145 103.275 23.315 103.465 ;
        RECT 23.605 103.255 23.775 103.445 ;
        RECT 24.985 103.275 25.155 103.465 ;
        RECT 25.260 103.255 25.430 103.445 ;
        RECT 29.125 103.255 29.295 103.445 ;
        RECT 30.960 103.305 31.080 103.415 ;
        RECT 31.885 103.255 32.055 103.445 ;
        RECT 34.645 103.275 34.815 103.465 ;
        RECT 37.405 103.255 37.575 103.445 ;
        RECT 40.165 103.275 40.335 103.465 ;
        RECT 42.925 103.255 43.095 103.445 ;
        RECT 43.840 103.305 43.960 103.415 ;
        RECT 45.040 103.275 45.210 103.465 ;
        RECT 46.605 103.255 46.775 103.445 ;
        RECT 47.985 103.255 48.155 103.445 ;
        RECT 48.905 103.275 49.075 103.465 ;
        RECT 49.365 103.255 49.535 103.445 ;
        RECT 54.425 103.275 54.595 103.465 ;
        RECT 56.745 103.445 56.895 103.465 ;
        RECT 60.865 103.445 61.015 103.465 ;
        RECT 54.885 103.275 55.055 103.445 ;
        RECT 56.260 103.305 56.380 103.415 ;
        RECT 56.725 103.275 56.895 103.445 ;
        RECT 59.485 103.275 59.655 103.445 ;
        RECT 54.905 103.255 55.055 103.275 ;
        RECT 59.485 103.255 59.635 103.275 ;
        RECT 59.945 103.255 60.115 103.445 ;
        RECT 60.865 103.275 61.035 103.445 ;
        RECT 61.325 103.275 61.495 103.465 ;
        RECT 61.780 103.305 61.900 103.415 ;
        RECT 64.545 103.255 64.715 103.445 ;
        RECT 65.005 103.255 65.175 103.445 ;
        RECT 66.845 103.275 67.015 103.465 ;
        RECT 69.600 103.305 69.720 103.415 ;
        RECT 70.525 103.255 70.695 103.445 ;
        RECT 71.720 103.275 71.890 103.465 ;
        RECT 75.585 103.275 75.755 103.465 ;
        RECT 76.045 103.255 76.215 103.445 ;
        RECT 81.105 103.275 81.275 103.465 ;
        RECT 81.565 103.255 81.735 103.445 ;
        RECT 82.940 103.305 83.060 103.415 ;
        RECT 83.405 103.255 83.575 103.445 ;
        RECT 83.680 103.275 83.850 103.465 ;
        RECT 5.525 102.445 6.895 103.255 ;
        RECT 6.905 102.445 9.655 103.255 ;
        RECT 10.125 102.575 19.405 103.255 ;
        RECT 11.485 102.355 12.405 102.575 ;
        RECT 17.070 102.455 19.405 102.575 ;
        RECT 18.485 102.345 19.405 102.455 ;
        RECT 19.785 102.445 23.455 103.255 ;
        RECT 23.465 102.445 24.835 103.255 ;
        RECT 24.845 102.575 28.745 103.255 ;
        RECT 24.845 102.345 25.775 102.575 ;
        RECT 28.985 102.445 30.815 103.255 ;
        RECT 31.295 102.385 31.725 103.170 ;
        RECT 31.745 102.445 37.255 103.255 ;
        RECT 37.265 102.445 42.775 103.255 ;
        RECT 42.785 102.445 46.455 103.255 ;
        RECT 46.465 102.445 47.835 103.255 ;
        RECT 47.855 102.345 49.205 103.255 ;
        RECT 49.225 102.445 54.735 103.255 ;
        RECT 54.905 102.435 56.835 103.255 ;
        RECT 55.885 102.345 56.835 102.435 ;
        RECT 57.055 102.385 57.485 103.170 ;
        RECT 57.705 102.435 59.635 103.255 ;
        RECT 59.805 102.445 61.635 103.255 ;
        RECT 62.115 102.575 64.855 103.255 ;
        RECT 64.865 102.445 70.375 103.255 ;
        RECT 70.385 102.445 75.895 103.255 ;
        RECT 75.905 102.445 81.415 103.255 ;
        RECT 81.425 102.445 82.795 103.255 ;
        RECT 57.705 102.345 58.655 102.435 ;
        RECT 82.815 102.385 83.245 103.170 ;
        RECT 83.265 102.445 86.015 103.255 ;
        RECT 86.170 103.225 86.340 103.445 ;
        RECT 87.545 103.275 87.715 103.465 ;
        RECT 91.225 103.445 91.375 103.465 ;
        RECT 93.525 103.445 93.675 103.465 ;
        RECT 87.830 103.225 88.775 103.255 ;
        RECT 88.930 103.225 89.100 103.445 ;
        RECT 91.225 103.275 91.395 103.445 ;
        RECT 91.680 103.305 91.800 103.415 ;
        RECT 93.525 103.275 93.695 103.445 ;
        RECT 93.985 103.275 94.155 103.465 ;
        RECT 96.285 103.275 96.455 103.465 ;
        RECT 93.985 103.255 94.135 103.275 ;
        RECT 96.285 103.255 96.435 103.275 ;
        RECT 96.745 103.255 96.915 103.445 ;
        RECT 97.940 103.275 98.110 103.465 ;
        RECT 101.805 103.275 101.975 103.465 ;
        RECT 102.265 103.255 102.435 103.445 ;
        RECT 103.185 103.275 103.355 103.465 ;
        RECT 107.795 103.300 107.955 103.410 ;
        RECT 109.165 103.255 109.335 103.445 ;
        RECT 111.465 103.255 111.635 103.445 ;
        RECT 111.925 103.255 112.095 103.445 ;
        RECT 112.385 103.275 112.555 103.465 ;
        RECT 117.445 103.255 117.615 103.445 ;
        RECT 117.905 103.275 118.075 103.465 ;
        RECT 122.045 103.275 122.215 103.465 ;
        RECT 122.965 103.255 123.135 103.445 ;
        RECT 123.880 103.305 124.000 103.415 ;
        RECT 125.265 103.255 125.435 103.465 ;
        RECT 90.590 103.225 91.535 103.255 ;
        RECT 86.025 102.545 88.775 103.225 ;
        RECT 88.785 102.545 91.535 103.225 ;
        RECT 87.830 102.345 88.775 102.545 ;
        RECT 90.590 102.345 91.535 102.545 ;
        RECT 92.205 102.435 94.135 103.255 ;
        RECT 94.505 102.435 96.435 103.255 ;
        RECT 96.605 102.445 102.115 103.255 ;
        RECT 102.125 102.445 107.635 103.255 ;
        RECT 92.205 102.345 93.155 102.435 ;
        RECT 94.505 102.345 95.455 102.435 ;
        RECT 108.575 102.385 109.005 103.170 ;
        RECT 109.025 102.445 110.395 103.255 ;
        RECT 110.415 102.345 111.765 103.255 ;
        RECT 111.785 102.445 117.295 103.255 ;
        RECT 117.305 102.445 122.815 103.255 ;
        RECT 122.825 102.445 124.195 103.255 ;
        RECT 124.205 102.445 125.575 103.255 ;
      LAYER nwell ;
        RECT 5.330 99.225 125.770 102.055 ;
      LAYER pwell ;
        RECT 5.525 98.025 6.895 98.835 ;
        RECT 6.905 98.025 12.415 98.835 ;
        RECT 12.425 98.025 14.255 98.835 ;
        RECT 14.275 98.025 15.625 98.935 ;
        RECT 15.645 98.025 18.395 98.835 ;
        RECT 18.415 98.110 18.845 98.895 ;
        RECT 22.305 98.845 23.255 98.935 ;
        RECT 24.605 98.845 25.555 98.935 ;
        RECT 18.865 98.025 20.695 98.835 ;
        RECT 21.325 98.025 23.255 98.845 ;
        RECT 23.625 98.025 25.555 98.845 ;
        RECT 25.965 98.845 26.915 98.935 ;
        RECT 29.205 98.845 30.155 98.935 ;
        RECT 25.965 98.025 27.895 98.845 ;
        RECT 5.665 97.815 5.835 98.025 ;
        RECT 7.045 97.815 7.215 98.025 ;
        RECT 12.565 97.835 12.735 98.025 ;
        RECT 14.405 97.815 14.575 98.005 ;
        RECT 14.865 97.815 15.035 98.005 ;
        RECT 15.325 97.835 15.495 98.025 ;
        RECT 15.785 97.835 15.955 98.025 ;
        RECT 19.005 97.835 19.175 98.025 ;
        RECT 21.325 98.005 21.475 98.025 ;
        RECT 23.625 98.005 23.775 98.025 ;
        RECT 27.745 98.005 27.895 98.025 ;
        RECT 28.225 98.025 30.155 98.845 ;
        RECT 30.565 98.845 31.515 98.935 ;
        RECT 37.485 98.845 38.435 98.935 ;
        RECT 30.565 98.025 32.495 98.845 ;
        RECT 32.665 98.025 36.335 98.835 ;
        RECT 36.505 98.025 38.435 98.845 ;
        RECT 38.645 98.025 40.015 98.805 ;
        RECT 40.025 98.025 43.695 98.835 ;
        RECT 44.175 98.110 44.605 98.895 ;
        RECT 45.985 98.705 46.905 98.925 ;
        RECT 52.985 98.825 53.905 98.935 ;
        RECT 51.570 98.705 53.905 98.825 ;
        RECT 44.625 98.025 53.905 98.705 ;
        RECT 54.285 98.025 55.655 98.835 ;
        RECT 57.470 98.735 58.415 98.935 ;
        RECT 55.665 98.055 58.415 98.735 ;
        RECT 28.225 98.005 28.375 98.025 ;
        RECT 20.385 97.815 20.555 98.005 ;
        RECT 20.840 97.865 20.960 97.975 ;
        RECT 21.305 97.835 21.475 98.005 ;
        RECT 23.605 97.835 23.775 98.005 ;
        RECT 25.905 97.815 26.075 98.005 ;
        RECT 27.745 97.835 27.915 98.005 ;
        RECT 28.205 97.835 28.375 98.005 ;
        RECT 32.345 98.005 32.495 98.025 ;
        RECT 31.895 97.860 32.055 97.970 ;
        RECT 32.345 97.835 32.515 98.005 ;
        RECT 32.805 97.835 32.975 98.025 ;
        RECT 36.505 98.005 36.655 98.025 ;
        RECT 33.725 97.815 33.895 98.005 ;
        RECT 34.185 97.815 34.355 98.005 ;
        RECT 36.485 97.835 36.655 98.005 ;
        RECT 36.940 97.865 37.060 97.975 ;
        RECT 37.405 97.815 37.575 98.005 ;
        RECT 38.785 97.835 38.955 98.025 ;
        RECT 40.165 97.835 40.335 98.025 ;
        RECT 43.840 97.865 43.960 97.975 ;
        RECT 44.765 97.835 44.935 98.025 ;
        RECT 47.985 97.815 48.155 98.005 ;
        RECT 48.720 97.815 48.890 98.005 ;
        RECT 52.595 97.860 52.755 97.970 ;
        RECT 53.510 97.815 53.680 98.005 ;
        RECT 54.425 97.835 54.595 98.025 ;
        RECT 55.810 97.835 55.980 98.055 ;
        RECT 57.470 98.025 58.415 98.055 ;
        RECT 58.425 98.025 63.935 98.835 ;
        RECT 63.945 98.025 66.695 98.835 ;
        RECT 67.165 98.025 69.905 98.705 ;
        RECT 69.935 98.110 70.365 98.895 ;
        RECT 70.855 98.025 72.205 98.935 ;
        RECT 72.225 98.025 73.595 98.805 ;
        RECT 73.605 98.025 77.275 98.835 ;
        RECT 77.480 98.025 80.955 98.935 ;
        RECT 81.160 98.025 84.635 98.935 ;
        RECT 84.840 98.025 88.315 98.935 ;
        RECT 93.585 98.845 94.535 98.935 ;
        RECT 88.325 98.025 91.995 98.835 ;
        RECT 92.005 98.025 93.375 98.835 ;
        RECT 93.585 98.025 95.515 98.845 ;
        RECT 95.695 98.110 96.125 98.895 ;
        RECT 97.065 98.025 98.435 98.805 ;
        RECT 98.445 98.025 100.275 98.835 ;
        RECT 100.755 98.025 102.105 98.935 ;
        RECT 102.125 98.025 104.875 98.835 ;
        RECT 106.705 98.705 107.625 98.925 ;
        RECT 113.705 98.825 114.625 98.935 ;
        RECT 112.290 98.705 114.625 98.825 ;
        RECT 118.205 98.705 119.135 98.935 ;
        RECT 105.345 98.025 114.625 98.705 ;
        RECT 115.235 98.025 119.135 98.705 ;
        RECT 119.145 98.025 120.515 98.805 ;
        RECT 121.455 98.110 121.885 98.895 ;
        RECT 121.915 98.025 123.265 98.935 ;
        RECT 124.205 98.025 125.575 98.835 ;
        RECT 58.565 97.835 58.735 98.025 ;
        RECT 60.860 97.815 61.030 98.005 ;
        RECT 61.325 97.815 61.495 98.005 ;
        RECT 63.165 97.835 63.335 98.005 ;
        RECT 64.085 97.835 64.255 98.025 ;
        RECT 65.460 97.865 65.580 97.975 ;
        RECT 63.185 97.815 63.335 97.835 ;
        RECT 65.925 97.815 66.095 98.005 ;
        RECT 66.840 97.865 66.960 97.975 ;
        RECT 67.305 97.835 67.475 98.025 ;
        RECT 70.520 97.865 70.640 97.975 ;
        RECT 71.905 97.835 72.075 98.025 ;
        RECT 73.285 97.835 73.455 98.025 ;
        RECT 73.745 97.835 73.915 98.025 ;
        RECT 78.800 97.815 78.970 98.005 ;
        RECT 79.265 97.815 79.435 98.005 ;
        RECT 80.640 97.835 80.810 98.025 ;
        RECT 84.320 97.835 84.490 98.025 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.005 12.415 97.815 ;
        RECT 13.345 97.035 14.715 97.815 ;
        RECT 14.725 97.005 20.235 97.815 ;
        RECT 20.245 97.005 25.755 97.815 ;
        RECT 25.765 97.005 31.275 97.815 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 32.675 96.905 34.025 97.815 ;
        RECT 34.045 97.005 36.795 97.815 ;
        RECT 37.265 97.135 46.545 97.815 ;
        RECT 38.625 96.915 39.545 97.135 ;
        RECT 44.210 97.015 46.545 97.135 ;
        RECT 46.925 97.035 48.295 97.815 ;
        RECT 48.305 97.135 52.205 97.815 ;
        RECT 45.625 96.905 46.545 97.015 ;
        RECT 48.305 96.905 49.235 97.135 ;
        RECT 53.365 96.905 56.840 97.815 ;
        RECT 57.055 96.945 57.485 97.730 ;
        RECT 57.700 96.905 61.175 97.815 ;
        RECT 61.185 97.005 63.015 97.815 ;
        RECT 63.185 96.995 65.115 97.815 ;
        RECT 65.785 97.135 75.065 97.815 ;
        RECT 64.165 96.905 65.115 96.995 ;
        RECT 67.145 96.915 68.065 97.135 ;
        RECT 72.730 97.015 75.065 97.135 ;
        RECT 74.145 96.905 75.065 97.015 ;
        RECT 75.640 96.905 79.115 97.815 ;
        RECT 79.125 97.005 82.795 97.815 ;
        RECT 83.265 97.785 84.210 97.815 ;
        RECT 85.700 97.785 85.870 98.005 ;
        RECT 86.165 97.815 86.335 98.005 ;
        RECT 88.000 97.835 88.170 98.025 ;
        RECT 88.465 97.835 88.635 98.025 ;
        RECT 91.685 97.815 91.855 98.005 ;
        RECT 92.145 97.835 92.315 98.025 ;
        RECT 95.365 98.005 95.515 98.025 ;
        RECT 95.360 97.835 95.535 98.005 ;
        RECT 82.815 96.945 83.245 97.730 ;
        RECT 83.265 97.105 86.015 97.785 ;
        RECT 83.265 96.905 84.210 97.105 ;
        RECT 86.025 97.005 91.535 97.815 ;
        RECT 91.545 97.005 92.915 97.815 ;
        RECT 92.925 97.785 93.870 97.815 ;
        RECT 95.360 97.785 95.530 97.835 ;
        RECT 95.825 97.815 95.995 98.005 ;
        RECT 96.295 97.870 96.455 97.980 ;
        RECT 98.125 97.835 98.295 98.025 ;
        RECT 98.585 97.835 98.755 98.025 ;
        RECT 100.420 97.865 100.540 97.975 ;
        RECT 101.805 97.835 101.975 98.025 ;
        RECT 102.265 97.835 102.435 98.025 ;
        RECT 105.020 97.865 105.140 97.975 ;
        RECT 105.485 97.835 105.655 98.025 ;
        RECT 107.325 97.835 107.495 98.005 ;
        RECT 107.795 97.860 107.955 97.970 ;
        RECT 107.325 97.815 107.475 97.835 ;
        RECT 109.440 97.815 109.610 98.005 ;
        RECT 113.300 97.865 113.420 97.975 ;
        RECT 113.765 97.815 113.935 98.005 ;
        RECT 118.550 97.835 118.720 98.025 ;
        RECT 120.205 97.835 120.375 98.025 ;
        RECT 120.675 97.870 120.835 97.980 ;
        RECT 122.045 97.835 122.215 98.025 ;
        RECT 123.435 97.860 123.595 97.980 ;
        RECT 125.265 97.815 125.435 98.025 ;
        RECT 92.925 97.105 95.675 97.785 ;
        RECT 95.685 97.135 104.965 97.815 ;
        RECT 92.925 96.905 93.870 97.105 ;
        RECT 97.045 96.915 97.965 97.135 ;
        RECT 102.630 97.015 104.965 97.135 ;
        RECT 104.045 96.905 104.965 97.015 ;
        RECT 105.545 96.995 107.475 97.815 ;
        RECT 105.545 96.905 106.495 96.995 ;
        RECT 108.575 96.945 109.005 97.730 ;
        RECT 109.025 97.135 112.925 97.815 ;
        RECT 113.625 97.135 122.905 97.815 ;
        RECT 109.025 96.905 109.955 97.135 ;
        RECT 114.985 96.915 115.905 97.135 ;
        RECT 120.570 97.015 122.905 97.135 ;
        RECT 121.985 96.905 122.905 97.015 ;
        RECT 124.205 97.005 125.575 97.815 ;
      LAYER nwell ;
        RECT 5.330 93.785 125.770 96.615 ;
      LAYER pwell ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 8.735 93.395 ;
        RECT 10.105 93.265 11.025 93.485 ;
        RECT 17.105 93.385 18.025 93.495 ;
        RECT 15.690 93.265 18.025 93.385 ;
        RECT 8.745 92.585 18.025 93.265 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 18.865 92.585 24.375 93.395 ;
        RECT 24.385 92.585 26.215 93.395 ;
        RECT 26.225 92.585 27.595 93.365 ;
        RECT 28.965 93.265 29.885 93.485 ;
        RECT 35.965 93.385 36.885 93.495 ;
        RECT 34.550 93.265 36.885 93.385 ;
        RECT 27.605 92.585 36.885 93.265 ;
        RECT 38.185 93.265 39.115 93.495 ;
        RECT 38.185 92.585 42.085 93.265 ;
        RECT 42.335 92.585 43.685 93.495 ;
        RECT 44.175 92.670 44.605 93.455 ;
        RECT 44.625 92.585 50.135 93.395 ;
        RECT 50.145 92.585 55.655 93.395 ;
        RECT 56.585 93.295 57.530 93.495 ;
        RECT 56.585 92.615 59.335 93.295 ;
        RECT 56.585 92.585 57.530 92.615 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.535 7.215 92.585 ;
        RECT 7.040 92.425 7.215 92.535 ;
        RECT 7.045 92.395 7.215 92.425 ;
        RECT 7.505 92.375 7.675 92.565 ;
        RECT 8.885 92.395 9.055 92.585 ;
        RECT 17.440 92.375 17.610 92.565 ;
        RECT 19.005 92.395 19.175 92.585 ;
        RECT 24.525 92.565 24.695 92.585 ;
        RECT 22.225 92.375 22.395 92.565 ;
        RECT 22.685 92.375 22.855 92.565 ;
        RECT 24.525 92.395 24.700 92.565 ;
        RECT 26.365 92.395 26.535 92.585 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 7.365 91.695 16.645 92.375 ;
        RECT 8.725 91.475 9.645 91.695 ;
        RECT 14.310 91.575 16.645 91.695 ;
        RECT 15.725 91.465 16.645 91.575 ;
        RECT 17.025 91.695 20.925 92.375 ;
        RECT 17.025 91.465 17.955 91.695 ;
        RECT 21.175 91.465 22.525 92.375 ;
        RECT 22.545 91.565 24.375 92.375 ;
        RECT 24.530 92.345 24.700 92.395 ;
        RECT 27.285 92.375 27.455 92.565 ;
        RECT 27.745 92.395 27.915 92.585 ;
        RECT 26.190 92.345 27.135 92.375 ;
        RECT 24.385 91.665 27.135 92.345 ;
        RECT 26.190 91.465 27.135 91.665 ;
        RECT 27.145 91.565 28.515 92.375 ;
        RECT 28.525 92.345 29.470 92.375 ;
        RECT 30.960 92.345 31.130 92.565 ;
        RECT 32.160 92.375 32.330 92.565 ;
        RECT 36.025 92.375 36.195 92.565 ;
        RECT 37.415 92.430 37.575 92.540 ;
        RECT 38.600 92.395 38.770 92.585 ;
        RECT 41.545 92.375 41.715 92.565 ;
        RECT 43.385 92.395 43.555 92.585 ;
        RECT 43.840 92.425 43.960 92.535 ;
        RECT 44.765 92.395 44.935 92.585 ;
        RECT 47.065 92.375 47.235 92.565 ;
        RECT 50.285 92.395 50.455 92.585 ;
        RECT 52.585 92.375 52.755 92.565 ;
        RECT 55.815 92.430 55.975 92.540 ;
        RECT 56.275 92.420 56.435 92.530 ;
        RECT 28.525 91.665 31.275 92.345 ;
        RECT 28.525 91.465 29.470 91.665 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 31.745 91.695 35.645 92.375 ;
        RECT 31.745 91.465 32.675 91.695 ;
        RECT 35.885 91.565 41.395 92.375 ;
        RECT 41.405 91.565 46.915 92.375 ;
        RECT 46.925 91.565 52.435 92.375 ;
        RECT 52.445 91.565 56.115 92.375 ;
        RECT 57.650 92.345 57.820 92.565 ;
        RECT 59.020 92.395 59.190 92.615 ;
        RECT 59.345 92.585 63.015 93.395 ;
        RECT 63.945 92.585 65.775 93.265 ;
        RECT 65.785 92.585 69.455 93.395 ;
        RECT 69.935 92.670 70.365 93.455 ;
        RECT 73.585 93.265 74.515 93.495 ;
        RECT 70.615 92.585 74.515 93.265 ;
        RECT 74.525 92.585 78.195 93.395 ;
        RECT 78.205 93.295 79.150 93.495 ;
        RECT 78.205 92.615 80.955 93.295 ;
        RECT 78.205 92.585 79.150 92.615 ;
        RECT 59.485 92.395 59.655 92.585 ;
        RECT 60.405 92.375 60.575 92.565 ;
        RECT 63.175 92.535 63.335 92.540 ;
        RECT 63.160 92.430 63.335 92.535 ;
        RECT 63.160 92.425 63.280 92.430 ;
        RECT 64.085 92.395 64.255 92.585 ;
        RECT 65.005 92.375 65.175 92.565 ;
        RECT 65.465 92.375 65.635 92.565 ;
        RECT 65.925 92.395 66.095 92.585 ;
        RECT 69.600 92.425 69.720 92.535 ;
        RECT 73.930 92.395 74.100 92.585 ;
        RECT 74.665 92.395 74.835 92.585 ;
        RECT 77.885 92.375 78.055 92.565 ;
        RECT 80.640 92.395 80.810 92.615 ;
        RECT 80.965 92.585 83.715 93.395 ;
        RECT 84.380 92.585 87.855 93.495 ;
        RECT 93.585 93.405 94.535 93.495 ;
        RECT 87.865 92.585 93.375 93.395 ;
        RECT 93.585 92.585 95.515 93.405 ;
        RECT 95.695 92.670 96.125 93.455 ;
        RECT 96.145 92.585 97.515 93.395 ;
        RECT 97.525 93.265 98.455 93.495 ;
        RECT 97.525 92.585 101.425 93.265 ;
        RECT 101.665 92.585 105.335 93.395 ;
        RECT 105.345 92.585 106.715 93.395 ;
        RECT 106.725 92.585 108.095 93.365 ;
        RECT 108.105 92.585 113.615 93.395 ;
        RECT 113.625 92.585 117.295 93.395 ;
        RECT 117.775 92.585 119.125 93.495 ;
        RECT 119.145 92.585 120.975 93.395 ;
        RECT 121.455 92.670 121.885 93.455 ;
        RECT 121.905 92.585 123.735 93.395 ;
        RECT 124.205 92.585 125.575 93.395 ;
        RECT 81.105 92.395 81.275 92.585 ;
        RECT 81.560 92.375 81.730 92.565 ;
        RECT 82.035 92.420 82.195 92.530 ;
        RECT 83.860 92.425 83.980 92.535 ;
        RECT 59.310 92.345 60.255 92.375 ;
        RECT 57.055 91.505 57.485 92.290 ;
        RECT 57.505 91.665 60.255 92.345 ;
        RECT 59.310 91.465 60.255 91.665 ;
        RECT 60.265 91.565 63.015 92.375 ;
        RECT 63.485 91.695 65.315 92.375 ;
        RECT 65.325 91.695 74.515 92.375 ;
        RECT 69.835 91.475 70.765 91.695 ;
        RECT 73.595 91.465 74.515 91.695 ;
        RECT 74.620 91.695 78.085 92.375 ;
        RECT 74.620 91.465 75.540 91.695 ;
        RECT 78.400 91.465 81.875 92.375 ;
        RECT 83.265 92.345 84.210 92.375 ;
        RECT 85.700 92.345 85.870 92.565 ;
        RECT 86.165 92.375 86.335 92.565 ;
        RECT 87.540 92.395 87.710 92.585 ;
        RECT 88.005 92.395 88.175 92.585 ;
        RECT 95.365 92.565 95.515 92.585 ;
        RECT 90.950 92.375 91.120 92.565 ;
        RECT 92.605 92.375 92.775 92.565 ;
        RECT 93.985 92.375 94.155 92.565 ;
        RECT 94.445 92.375 94.615 92.565 ;
        RECT 95.365 92.395 95.535 92.565 ;
        RECT 96.285 92.395 96.455 92.585 ;
        RECT 97.940 92.395 98.110 92.585 ;
        RECT 99.965 92.375 100.135 92.565 ;
        RECT 101.805 92.395 101.975 92.585 ;
        RECT 105.485 92.375 105.655 92.585 ;
        RECT 107.785 92.395 107.955 92.585 ;
        RECT 108.245 92.535 108.415 92.585 ;
        RECT 108.240 92.425 108.415 92.535 ;
        RECT 108.245 92.395 108.415 92.425 ;
        RECT 109.165 92.375 109.335 92.565 ;
        RECT 112.845 92.375 113.015 92.565 ;
        RECT 113.765 92.395 113.935 92.585 ;
        RECT 114.500 92.375 114.670 92.565 ;
        RECT 117.440 92.425 117.560 92.535 ;
        RECT 118.825 92.395 118.995 92.585 ;
        RECT 119.285 92.395 119.455 92.585 ;
        RECT 121.120 92.425 121.240 92.535 ;
        RECT 121.770 92.375 121.940 92.565 ;
        RECT 122.045 92.395 122.215 92.585 ;
        RECT 122.505 92.375 122.675 92.565 ;
        RECT 123.880 92.425 124.000 92.535 ;
        RECT 125.265 92.375 125.435 92.585 ;
        RECT 82.815 91.505 83.245 92.290 ;
        RECT 83.265 91.665 86.015 92.345 ;
        RECT 83.265 91.465 84.210 91.665 ;
        RECT 86.025 91.565 87.395 92.375 ;
        RECT 87.635 91.695 91.535 92.375 ;
        RECT 90.605 91.465 91.535 91.695 ;
        RECT 91.545 91.595 92.915 92.375 ;
        RECT 92.935 91.465 94.285 92.375 ;
        RECT 94.305 91.565 99.815 92.375 ;
        RECT 99.825 91.565 105.335 92.375 ;
        RECT 105.345 91.565 108.095 92.375 ;
        RECT 108.575 91.505 109.005 92.290 ;
        RECT 109.025 91.565 112.695 92.375 ;
        RECT 112.705 91.565 114.075 92.375 ;
        RECT 114.085 91.695 117.985 92.375 ;
        RECT 118.455 91.695 122.355 92.375 ;
        RECT 114.085 91.465 115.015 91.695 ;
        RECT 121.425 91.465 122.355 91.695 ;
        RECT 122.365 91.565 124.195 92.375 ;
        RECT 124.205 91.565 125.575 92.375 ;
      LAYER nwell ;
        RECT 5.330 88.345 125.770 91.175 ;
      LAYER pwell ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 6.905 87.145 10.575 87.955 ;
        RECT 10.585 87.145 11.955 87.925 ;
        RECT 12.435 87.145 13.785 88.055 ;
        RECT 13.805 87.825 14.735 88.055 ;
        RECT 13.805 87.145 17.705 87.825 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 18.865 87.145 20.695 87.955 ;
        RECT 21.360 87.145 24.835 88.055 ;
        RECT 25.960 87.145 29.435 88.055 ;
        RECT 29.445 87.145 33.115 87.955 ;
        RECT 33.780 87.145 37.255 88.055 ;
        RECT 39.070 87.855 40.015 88.055 ;
        RECT 37.265 87.175 40.015 87.855 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.045 86.935 7.215 87.145 ;
        RECT 11.645 86.955 11.815 87.145 ;
        RECT 12.100 86.985 12.220 87.095 ;
        RECT 12.565 86.935 12.735 87.125 ;
        RECT 13.485 86.955 13.655 87.145 ;
        RECT 14.220 86.955 14.390 87.145 ;
        RECT 18.085 87.095 18.255 87.125 ;
        RECT 18.080 86.985 18.255 87.095 ;
        RECT 18.085 86.935 18.255 86.985 ;
        RECT 19.005 86.955 19.175 87.145 ;
        RECT 20.840 86.985 20.960 87.095 ;
        RECT 21.765 86.935 21.935 87.125 ;
        RECT 24.520 86.955 24.690 87.145 ;
        RECT 24.995 86.990 25.155 87.100 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 6.905 86.125 12.415 86.935 ;
        RECT 12.425 86.125 17.935 86.935 ;
        RECT 17.945 86.125 21.615 86.935 ;
        RECT 21.625 86.125 22.995 86.935 ;
        RECT 23.005 86.905 23.950 86.935 ;
        RECT 25.440 86.905 25.610 87.125 ;
        RECT 25.905 86.935 26.075 87.125 ;
        RECT 29.120 86.955 29.290 87.145 ;
        RECT 29.585 86.955 29.755 87.145 ;
        RECT 31.885 86.935 32.055 87.125 ;
        RECT 33.260 86.985 33.380 87.095 ;
        RECT 36.940 86.955 37.110 87.145 ;
        RECT 37.410 87.125 37.580 87.175 ;
        RECT 39.070 87.145 40.015 87.175 ;
        RECT 40.025 87.145 43.695 87.955 ;
        RECT 44.175 87.230 44.605 88.015 ;
        RECT 44.625 87.145 45.995 87.955 ;
        RECT 46.005 87.145 47.375 87.925 ;
        RECT 47.385 87.145 48.755 87.925 ;
        RECT 49.225 87.825 50.155 88.055 ;
        RECT 53.365 87.825 54.295 88.055 ;
        RECT 49.225 87.145 53.125 87.825 ;
        RECT 53.365 87.145 57.265 87.825 ;
        RECT 57.505 87.145 60.980 88.055 ;
        RECT 61.185 87.145 66.695 87.955 ;
        RECT 67.625 87.145 68.995 87.925 ;
        RECT 69.935 87.230 70.365 88.015 ;
        RECT 70.385 87.825 71.315 88.055 ;
        RECT 70.385 87.145 74.285 87.825 ;
        RECT 74.535 87.145 75.885 88.055 ;
        RECT 75.905 87.145 81.415 87.955 ;
        RECT 81.425 87.145 85.095 87.955 ;
        RECT 87.385 87.825 88.305 88.045 ;
        RECT 94.385 87.945 95.305 88.055 ;
        RECT 92.970 87.825 95.305 87.945 ;
        RECT 86.025 87.145 95.305 87.825 ;
        RECT 95.695 87.230 96.125 88.015 ;
        RECT 105.085 87.965 106.035 88.055 ;
        RECT 107.385 87.965 108.335 88.055 ;
        RECT 96.145 87.145 101.655 87.955 ;
        RECT 101.665 87.145 104.415 87.955 ;
        RECT 105.085 87.145 107.015 87.965 ;
        RECT 107.385 87.145 109.315 87.965 ;
        RECT 110.405 87.145 111.775 87.925 ;
        RECT 113.145 87.825 114.065 88.045 ;
        RECT 120.145 87.945 121.065 88.055 ;
        RECT 118.730 87.825 121.065 87.945 ;
        RECT 111.785 87.145 121.065 87.825 ;
        RECT 121.455 87.230 121.885 88.015 ;
        RECT 121.905 87.145 123.275 87.925 ;
        RECT 124.205 87.145 125.575 87.955 ;
        RECT 37.405 86.955 37.580 87.125 ;
        RECT 40.165 86.955 40.335 87.145 ;
        RECT 37.405 86.935 37.575 86.955 ;
        RECT 42.925 86.935 43.095 87.125 ;
        RECT 43.840 86.985 43.960 87.095 ;
        RECT 44.305 86.935 44.475 87.125 ;
        RECT 44.765 86.955 44.935 87.145 ;
        RECT 45.685 86.935 45.855 87.125 ;
        RECT 46.145 86.955 46.315 87.145 ;
        RECT 48.445 86.955 48.615 87.145 ;
        RECT 48.900 86.985 49.020 87.095 ;
        RECT 49.640 86.955 49.810 87.145 ;
        RECT 53.780 86.955 53.950 87.145 ;
        RECT 55.345 86.935 55.515 87.125 ;
        RECT 57.650 86.935 57.820 87.145 ;
        RECT 61.325 86.935 61.495 87.145 ;
        RECT 63.160 86.985 63.280 87.095 ;
        RECT 65.005 86.935 65.175 87.125 ;
        RECT 65.465 86.935 65.635 87.125 ;
        RECT 66.855 86.990 67.015 87.100 ;
        RECT 68.685 86.955 68.855 87.145 ;
        RECT 69.155 86.990 69.315 87.100 ;
        RECT 70.800 86.955 70.970 87.145 ;
        RECT 70.985 86.935 71.155 87.125 ;
        RECT 75.585 86.955 75.755 87.145 ;
        RECT 76.045 86.955 76.215 87.145 ;
        RECT 77.425 86.935 77.595 87.125 ;
        RECT 78.805 86.935 78.975 87.125 ;
        RECT 79.265 86.935 79.435 87.125 ;
        RECT 81.565 86.955 81.735 87.145 ;
        RECT 83.405 86.935 83.575 87.125 ;
        RECT 85.255 86.990 85.415 87.100 ;
        RECT 86.165 86.955 86.335 87.145 ;
        RECT 87.095 86.980 87.255 87.090 ;
        RECT 88.925 86.935 89.095 87.125 ;
        RECT 89.385 86.935 89.555 87.125 ;
        RECT 95.360 86.935 95.530 87.125 ;
        RECT 95.825 86.935 95.995 87.125 ;
        RECT 96.285 86.955 96.455 87.145 ;
        RECT 101.355 86.980 101.515 87.090 ;
        RECT 101.805 86.955 101.975 87.145 ;
        RECT 106.865 87.125 107.015 87.145 ;
        RECT 109.165 87.125 109.315 87.145 ;
        RECT 23.005 86.225 25.755 86.905 ;
        RECT 23.005 86.025 23.950 86.225 ;
        RECT 25.765 86.125 31.275 86.935 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 31.745 86.125 37.255 86.935 ;
        RECT 37.265 86.125 42.775 86.935 ;
        RECT 42.785 86.125 44.155 86.935 ;
        RECT 44.175 86.025 45.525 86.935 ;
        RECT 45.545 86.255 54.825 86.935 ;
        RECT 46.905 86.035 47.825 86.255 ;
        RECT 52.490 86.135 54.825 86.255 ;
        RECT 53.905 86.025 54.825 86.135 ;
        RECT 55.205 86.125 57.035 86.935 ;
        RECT 57.055 86.065 57.485 86.850 ;
        RECT 57.505 86.025 60.980 86.935 ;
        RECT 61.185 86.125 63.015 86.935 ;
        RECT 63.485 86.255 65.315 86.935 ;
        RECT 63.485 86.025 64.830 86.255 ;
        RECT 65.325 86.125 70.835 86.935 ;
        RECT 70.845 86.125 76.355 86.935 ;
        RECT 76.365 86.155 77.735 86.935 ;
        RECT 77.755 86.025 79.105 86.935 ;
        RECT 79.125 86.125 82.795 86.935 ;
        RECT 82.815 86.065 83.245 86.850 ;
        RECT 83.265 86.125 86.935 86.935 ;
        RECT 87.865 86.155 89.235 86.935 ;
        RECT 89.245 86.125 91.995 86.935 ;
        RECT 92.200 86.025 95.675 86.935 ;
        RECT 95.685 86.125 101.195 86.935 ;
        RECT 102.270 86.905 102.440 87.125 ;
        RECT 104.560 86.985 104.680 87.095 ;
        RECT 106.865 86.955 107.035 87.125 ;
        RECT 106.865 86.935 107.015 86.955 ;
        RECT 107.325 86.935 107.495 87.125 ;
        RECT 109.165 86.935 109.335 87.125 ;
        RECT 109.635 86.990 109.795 87.100 ;
        RECT 110.545 86.955 110.715 87.145 ;
        RECT 111.925 86.955 112.095 87.145 ;
        RECT 112.845 86.935 113.015 87.125 ;
        RECT 122.505 86.935 122.675 87.125 ;
        RECT 122.965 86.955 123.135 87.145 ;
        RECT 123.435 86.990 123.595 87.100 ;
        RECT 125.265 86.935 125.435 87.145 ;
        RECT 103.930 86.905 104.875 86.935 ;
        RECT 102.125 86.225 104.875 86.905 ;
        RECT 103.930 86.025 104.875 86.225 ;
        RECT 105.085 86.115 107.015 86.935 ;
        RECT 107.185 86.125 108.555 86.935 ;
        RECT 105.085 86.025 106.035 86.115 ;
        RECT 108.575 86.065 109.005 86.850 ;
        RECT 109.025 86.125 112.695 86.935 ;
        RECT 112.705 86.255 121.985 86.935 ;
        RECT 114.065 86.035 114.985 86.255 ;
        RECT 119.650 86.135 121.985 86.255 ;
        RECT 121.065 86.025 121.985 86.135 ;
        RECT 122.365 86.125 124.195 86.935 ;
        RECT 124.205 86.125 125.575 86.935 ;
      LAYER nwell ;
        RECT 5.330 82.905 125.770 85.735 ;
      LAYER pwell ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 6.905 81.705 12.415 82.515 ;
        RECT 12.425 81.705 17.935 82.515 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 18.865 81.705 20.695 82.515 ;
        RECT 20.900 81.705 24.375 82.615 ;
        RECT 25.500 81.705 28.975 82.615 ;
        RECT 29.080 82.385 30.000 82.615 ;
        RECT 37.175 82.385 38.105 82.605 ;
        RECT 40.935 82.385 41.855 82.615 ;
        RECT 29.080 81.705 32.545 82.385 ;
        RECT 32.665 81.705 41.855 82.385 ;
        RECT 41.875 81.705 43.225 82.615 ;
        RECT 44.175 81.790 44.605 82.575 ;
        RECT 45.985 82.385 46.905 82.605 ;
        RECT 52.985 82.505 53.905 82.615 ;
        RECT 51.570 82.385 53.905 82.505 ;
        RECT 44.625 81.705 53.905 82.385 ;
        RECT 54.285 82.415 55.230 82.615 ;
        RECT 54.285 81.735 57.035 82.415 ;
        RECT 54.285 81.705 55.230 81.735 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 9.805 81.495 9.975 81.685 ;
        RECT 11.185 81.495 11.355 81.685 ;
        RECT 11.920 81.495 12.090 81.685 ;
        RECT 12.565 81.515 12.735 81.705 ;
        RECT 16.060 81.495 16.230 81.685 ;
        RECT 18.080 81.545 18.200 81.655 ;
        RECT 19.005 81.515 19.175 81.705 ;
        RECT 19.925 81.495 20.095 81.685 ;
        RECT 24.060 81.515 24.230 81.705 ;
        RECT 24.520 81.660 24.690 81.685 ;
        RECT 24.520 81.550 24.695 81.660 ;
        RECT 24.520 81.495 24.690 81.550 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.685 8.735 81.495 ;
        RECT 8.745 80.715 10.115 81.495 ;
        RECT 10.125 80.715 11.495 81.495 ;
        RECT 11.505 80.815 15.405 81.495 ;
        RECT 15.645 80.815 19.545 81.495 ;
        RECT 11.505 80.585 12.435 80.815 ;
        RECT 15.645 80.585 16.575 80.815 ;
        RECT 19.785 80.685 21.155 81.495 ;
        RECT 21.360 80.585 24.835 81.495 ;
        RECT 24.990 81.465 25.160 81.685 ;
        RECT 28.660 81.515 28.830 81.705 ;
        RECT 26.650 81.465 27.595 81.495 ;
        RECT 24.845 80.785 27.595 81.465 ;
        RECT 26.650 80.585 27.595 80.785 ;
        RECT 27.605 81.465 28.550 81.495 ;
        RECT 30.040 81.465 30.210 81.685 ;
        RECT 30.515 81.540 30.675 81.650 ;
        RECT 31.885 81.495 32.055 81.685 ;
        RECT 32.345 81.515 32.515 81.705 ;
        RECT 32.805 81.515 32.975 81.705 ;
        RECT 36.485 81.495 36.655 81.685 ;
        RECT 36.940 81.545 37.060 81.655 ;
        RECT 37.680 81.495 37.850 81.685 ;
        RECT 41.545 81.495 41.715 81.685 ;
        RECT 42.925 81.515 43.095 81.705 ;
        RECT 43.395 81.550 43.555 81.660 ;
        RECT 44.765 81.515 44.935 81.705 ;
        RECT 47.075 81.540 47.235 81.650 ;
        RECT 47.985 81.495 48.155 81.685 ;
        RECT 49.365 81.495 49.535 81.685 ;
        RECT 54.885 81.495 55.055 81.685 ;
        RECT 56.720 81.515 56.890 81.735 ;
        RECT 57.045 81.705 58.875 82.515 ;
        RECT 63.025 82.385 64.370 82.615 ;
        RECT 68.570 82.385 69.915 82.615 ;
        RECT 59.355 81.705 62.095 82.385 ;
        RECT 63.025 81.705 64.855 82.385 ;
        RECT 65.325 81.705 68.065 82.385 ;
        RECT 68.085 81.705 69.915 82.385 ;
        RECT 69.935 81.790 70.365 82.575 ;
        RECT 70.385 81.705 73.595 82.615 ;
        RECT 73.615 81.705 74.965 82.615 ;
        RECT 75.540 82.385 76.460 82.615 ;
        RECT 75.540 81.705 79.005 82.385 ;
        RECT 80.240 81.705 83.715 82.615 ;
        RECT 83.725 81.705 85.555 82.515 ;
        RECT 87.385 82.385 88.305 82.605 ;
        RECT 94.385 82.505 95.305 82.615 ;
        RECT 92.970 82.385 95.305 82.505 ;
        RECT 86.025 81.705 95.305 82.385 ;
        RECT 95.695 81.790 96.125 82.575 ;
        RECT 96.340 81.705 99.815 82.615 ;
        RECT 99.825 81.705 101.655 82.515 ;
        RECT 103.930 82.415 104.875 82.615 ;
        RECT 106.690 82.415 107.635 82.615 ;
        RECT 102.125 81.735 104.875 82.415 ;
        RECT 104.885 81.735 107.635 82.415 ;
        RECT 57.185 81.515 57.355 81.705 ;
        RECT 57.645 81.495 57.815 81.685 ;
        RECT 59.020 81.545 59.140 81.655 ;
        RECT 61.785 81.515 61.955 81.705 ;
        RECT 62.255 81.550 62.415 81.660 ;
        RECT 63.625 81.495 63.795 81.685 ;
        RECT 64.545 81.515 64.715 81.705 ;
        RECT 65.000 81.545 65.120 81.655 ;
        RECT 65.465 81.495 65.635 81.705 ;
        RECT 65.925 81.495 66.095 81.685 ;
        RECT 67.775 81.540 67.935 81.650 ;
        RECT 68.225 81.515 68.395 81.705 ;
        RECT 68.685 81.495 68.855 81.685 ;
        RECT 73.285 81.515 73.455 81.705 ;
        RECT 74.665 81.515 74.835 81.705 ;
        RECT 75.120 81.545 75.240 81.655 ;
        RECT 78.355 81.540 78.515 81.650 ;
        RECT 78.805 81.515 78.975 81.705 ;
        RECT 79.270 81.495 79.440 81.685 ;
        RECT 83.400 81.515 83.570 81.705 ;
        RECT 83.680 81.495 83.850 81.685 ;
        RECT 83.865 81.515 84.035 81.705 ;
        RECT 85.700 81.545 85.820 81.655 ;
        RECT 86.165 81.515 86.335 81.705 ;
        RECT 99.500 81.685 99.670 81.705 ;
        RECT 87.540 81.545 87.660 81.655 ;
        RECT 88.280 81.495 88.450 81.685 ;
        RECT 93.065 81.495 93.235 81.685 ;
        RECT 93.525 81.495 93.695 81.685 ;
        RECT 96.280 81.545 96.400 81.655 ;
        RECT 27.605 80.785 30.355 81.465 ;
        RECT 27.605 80.585 28.550 80.785 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 31.745 80.685 35.415 81.495 ;
        RECT 35.425 80.715 36.795 81.495 ;
        RECT 37.265 80.815 41.165 81.495 ;
        RECT 37.265 80.585 38.195 80.815 ;
        RECT 41.405 80.685 46.915 81.495 ;
        RECT 47.855 80.585 49.205 81.495 ;
        RECT 49.225 80.685 54.735 81.495 ;
        RECT 54.745 80.685 56.575 81.495 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 57.505 80.685 61.175 81.495 ;
        RECT 61.215 80.585 63.935 81.495 ;
        RECT 63.945 80.815 65.775 81.495 ;
        RECT 65.785 80.815 67.615 81.495 ;
        RECT 68.545 80.815 77.825 81.495 ;
        RECT 63.945 80.585 65.290 80.815 ;
        RECT 66.270 80.585 67.615 80.815 ;
        RECT 69.905 80.595 70.825 80.815 ;
        RECT 75.490 80.695 77.825 80.815 ;
        RECT 76.905 80.585 77.825 80.695 ;
        RECT 79.125 80.585 82.600 81.495 ;
        RECT 82.815 80.625 83.245 81.410 ;
        RECT 83.265 80.815 87.165 81.495 ;
        RECT 87.865 80.815 91.765 81.495 ;
        RECT 83.265 80.585 84.195 80.815 ;
        RECT 87.865 80.585 88.795 80.815 ;
        RECT 92.015 80.585 93.365 81.495 ;
        RECT 93.385 80.685 96.135 81.495 ;
        RECT 96.750 81.465 96.920 81.685 ;
        RECT 99.500 81.515 99.675 81.685 ;
        RECT 99.965 81.515 100.135 81.705 ;
        RECT 101.800 81.545 101.920 81.655 ;
        RECT 102.270 81.515 102.440 81.735 ;
        RECT 103.930 81.705 104.875 81.735 ;
        RECT 105.030 81.685 105.200 81.735 ;
        RECT 106.690 81.705 107.635 81.735 ;
        RECT 107.645 81.705 113.155 82.515 ;
        RECT 113.165 81.705 116.835 82.515 ;
        RECT 117.315 81.705 118.665 82.615 ;
        RECT 118.685 81.705 121.435 82.515 ;
        RECT 121.455 81.790 121.885 82.575 ;
        RECT 121.905 81.705 123.735 82.515 ;
        RECT 124.205 81.705 125.575 82.515 ;
        RECT 105.025 81.515 105.200 81.685 ;
        RECT 107.785 81.515 107.955 81.705 ;
        RECT 99.505 81.495 99.675 81.515 ;
        RECT 105.025 81.495 105.195 81.515 ;
        RECT 109.165 81.495 109.335 81.685 ;
        RECT 113.305 81.515 113.475 81.705 ;
        RECT 114.685 81.495 114.855 81.685 ;
        RECT 116.980 81.545 117.100 81.655 ;
        RECT 118.365 81.515 118.535 81.705 ;
        RECT 118.825 81.515 118.995 81.705 ;
        RECT 120.205 81.495 120.375 81.685 ;
        RECT 122.045 81.515 122.215 81.705 ;
        RECT 123.880 81.545 124.000 81.655 ;
        RECT 125.265 81.495 125.435 81.705 ;
        RECT 98.410 81.465 99.355 81.495 ;
        RECT 96.605 80.785 99.355 81.465 ;
        RECT 98.410 80.585 99.355 80.785 ;
        RECT 99.365 80.685 104.875 81.495 ;
        RECT 104.885 80.685 108.555 81.495 ;
        RECT 108.575 80.625 109.005 81.410 ;
        RECT 109.025 80.685 114.535 81.495 ;
        RECT 114.545 80.685 120.055 81.495 ;
        RECT 120.065 80.685 123.735 81.495 ;
        RECT 124.205 80.685 125.575 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 125.770 80.295 ;
      LAYER pwell ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 8.725 76.945 9.645 77.165 ;
        RECT 15.725 77.065 16.645 77.175 ;
        RECT 14.310 76.945 16.645 77.065 ;
        RECT 7.365 76.265 16.645 76.945 ;
        RECT 17.035 76.265 18.385 77.175 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 18.960 76.945 19.880 77.175 ;
        RECT 18.960 76.265 22.425 76.945 ;
        RECT 22.555 76.265 23.905 77.175 ;
        RECT 23.925 76.265 29.435 77.075 ;
        RECT 29.445 76.265 34.955 77.075 ;
        RECT 34.965 76.265 40.475 77.075 ;
        RECT 40.485 76.265 44.155 77.075 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 44.625 76.265 50.135 77.075 ;
        RECT 50.145 76.265 55.655 77.075 ;
        RECT 55.665 76.265 61.175 77.075 ;
        RECT 61.185 76.265 63.015 77.075 ;
        RECT 63.510 76.945 64.855 77.175 ;
        RECT 63.025 76.265 64.855 76.945 ;
        RECT 64.865 76.265 68.535 77.075 ;
        RECT 68.545 76.265 69.915 77.075 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 70.385 76.265 72.215 77.075 ;
        RECT 74.045 76.945 74.965 77.165 ;
        RECT 81.045 77.065 81.965 77.175 ;
        RECT 79.630 76.945 81.965 77.065 ;
        RECT 72.685 76.265 81.965 76.945 ;
        RECT 82.345 76.265 87.855 77.075 ;
        RECT 87.865 76.265 93.375 77.075 ;
        RECT 93.385 76.265 95.215 77.075 ;
        RECT 95.695 76.350 96.125 77.135 ;
        RECT 96.145 76.265 99.815 77.075 ;
        RECT 99.825 76.265 101.195 77.075 ;
        RECT 101.400 76.265 104.875 77.175 ;
        RECT 104.885 76.265 108.360 77.175 ;
        RECT 108.565 76.265 110.395 77.075 ;
        RECT 110.405 76.265 111.775 77.045 ;
        RECT 113.145 76.945 114.065 77.165 ;
        RECT 120.145 77.065 121.065 77.175 ;
        RECT 118.730 76.945 121.065 77.065 ;
        RECT 111.785 76.265 121.065 76.945 ;
        RECT 121.455 76.350 121.885 77.135 ;
        RECT 121.905 76.265 123.735 77.075 ;
        RECT 124.205 76.265 125.575 77.075 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.215 7.215 76.245 ;
        RECT 7.040 76.105 7.215 76.215 ;
        RECT 7.045 76.055 7.215 76.105 ;
        RECT 7.505 76.075 7.675 76.265 ;
        RECT 8.425 76.055 8.595 76.245 ;
        RECT 18.085 76.075 18.255 76.265 ;
        RECT 19.920 76.055 20.090 76.245 ;
        RECT 22.225 76.075 22.395 76.265 ;
        RECT 23.605 76.245 23.775 76.265 ;
        RECT 23.600 76.075 23.775 76.245 ;
        RECT 24.065 76.075 24.235 76.265 ;
        RECT 23.600 76.055 23.770 76.075 ;
        RECT 27.280 76.055 27.450 76.245 ;
        RECT 29.585 76.075 29.755 76.265 ;
        RECT 30.960 76.055 31.130 76.245 ;
        RECT 31.885 76.055 32.055 76.245 ;
        RECT 35.105 76.075 35.275 76.265 ;
        RECT 37.860 76.055 38.030 76.245 ;
        RECT 38.600 76.055 38.770 76.245 ;
        RECT 40.625 76.075 40.795 76.265 ;
        RECT 42.465 76.055 42.635 76.245 ;
        RECT 44.765 76.075 44.935 76.265 ;
        RECT 47.985 76.055 48.155 76.245 ;
        RECT 49.365 76.055 49.535 76.245 ;
        RECT 50.285 76.075 50.455 76.265 ;
        RECT 50.745 76.055 50.915 76.245 ;
        RECT 55.805 76.075 55.975 76.265 ;
        RECT 56.720 76.055 56.890 76.245 ;
        RECT 57.650 76.055 57.820 76.245 ;
        RECT 61.325 76.055 61.495 76.265 ;
        RECT 63.165 76.075 63.335 76.265 ;
        RECT 65.005 76.055 65.175 76.265 ;
        RECT 68.685 76.075 68.855 76.265 ;
        RECT 70.525 76.075 70.695 76.265 ;
        RECT 72.360 76.105 72.480 76.215 ;
        RECT 72.825 76.075 72.995 76.265 ;
        RECT 74.205 76.055 74.375 76.245 ;
        RECT 79.725 76.055 79.895 76.245 ;
        RECT 82.485 76.215 82.655 76.265 ;
        RECT 82.480 76.105 82.655 76.215 ;
        RECT 82.485 76.075 82.655 76.105 ;
        RECT 83.405 76.055 83.575 76.245 ;
        RECT 88.005 76.075 88.175 76.265 ;
        RECT 88.925 76.055 89.095 76.245 ;
        RECT 90.760 76.105 90.880 76.215 ;
        RECT 93.525 76.075 93.695 76.265 ;
        RECT 94.440 76.055 94.610 76.245 ;
        RECT 94.905 76.055 95.075 76.245 ;
        RECT 95.360 76.105 95.480 76.215 ;
        RECT 96.285 76.075 96.455 76.265 ;
        RECT 99.965 76.055 100.135 76.265 ;
        RECT 100.425 76.055 100.595 76.245 ;
        RECT 102.260 76.105 102.380 76.215 ;
        RECT 104.560 76.075 104.730 76.265 ;
        RECT 105.030 76.075 105.200 76.265 ;
        RECT 105.940 76.055 106.110 76.245 ;
        RECT 106.405 76.055 106.575 76.245 ;
        RECT 108.240 76.105 108.360 76.215 ;
        RECT 108.705 76.075 108.875 76.265 ;
        RECT 109.160 76.105 109.280 76.215 ;
        RECT 110.545 76.075 110.715 76.265 ;
        RECT 111.925 76.075 112.095 76.265 ;
        RECT 113.030 76.055 113.200 76.245 ;
        RECT 113.765 76.055 113.935 76.245 ;
        RECT 116.525 76.055 116.695 76.245 ;
        RECT 118.825 76.055 118.995 76.245 ;
        RECT 119.285 76.055 119.455 76.245 ;
        RECT 122.045 76.075 122.215 76.265 ;
        RECT 122.965 76.055 123.135 76.245 ;
        RECT 123.880 76.105 124.000 76.215 ;
        RECT 125.265 76.055 125.435 76.265 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 6.905 75.245 8.275 76.055 ;
        RECT 8.285 75.375 17.475 76.055 ;
        RECT 12.795 75.155 13.725 75.375 ;
        RECT 16.555 75.145 17.475 75.375 ;
        RECT 17.625 75.145 20.235 76.055 ;
        RECT 20.440 75.145 23.915 76.055 ;
        RECT 24.120 75.145 27.595 76.055 ;
        RECT 27.800 75.145 31.275 76.055 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 31.745 75.245 34.495 76.055 ;
        RECT 34.700 75.145 38.175 76.055 ;
        RECT 38.185 75.375 42.085 76.055 ;
        RECT 38.185 75.145 39.115 75.375 ;
        RECT 42.325 75.245 47.835 76.055 ;
        RECT 47.845 75.245 49.215 76.055 ;
        RECT 49.235 75.145 50.585 76.055 ;
        RECT 50.605 75.245 53.355 76.055 ;
        RECT 53.560 75.145 57.035 76.055 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.505 75.145 60.980 76.055 ;
        RECT 61.185 75.245 64.855 76.055 ;
        RECT 64.865 75.375 73.970 76.055 ;
        RECT 74.065 75.245 79.575 76.055 ;
        RECT 79.585 75.245 82.335 76.055 ;
        RECT 82.815 75.185 83.245 75.970 ;
        RECT 83.265 75.245 88.775 76.055 ;
        RECT 88.785 75.245 90.615 76.055 ;
        RECT 91.280 75.145 94.755 76.055 ;
        RECT 94.765 75.245 96.595 76.055 ;
        RECT 96.700 75.375 100.165 76.055 ;
        RECT 96.700 75.145 97.620 75.375 ;
        RECT 100.285 75.245 102.115 76.055 ;
        RECT 102.780 75.145 106.255 76.055 ;
        RECT 106.265 75.245 108.095 76.055 ;
        RECT 108.575 75.185 109.005 75.970 ;
        RECT 109.715 75.375 113.615 76.055 ;
        RECT 112.685 75.145 113.615 75.375 ;
        RECT 113.625 75.245 116.375 76.055 ;
        RECT 116.395 75.145 117.745 76.055 ;
        RECT 117.765 75.275 119.135 76.055 ;
        RECT 119.145 75.245 122.815 76.055 ;
        RECT 122.825 75.245 124.195 76.055 ;
        RECT 124.205 75.245 125.575 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 125.770 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 6.905 70.825 12.415 71.635 ;
        RECT 12.425 70.825 17.935 71.635 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 18.865 70.825 20.235 71.635 ;
        RECT 20.440 70.825 23.915 71.735 ;
        RECT 24.120 70.825 27.595 71.735 ;
        RECT 27.605 70.825 33.115 71.635 ;
        RECT 33.125 70.825 34.495 71.605 ;
        RECT 35.865 71.505 36.785 71.725 ;
        RECT 42.865 71.625 43.785 71.735 ;
        RECT 41.450 71.505 43.785 71.625 ;
        RECT 34.505 70.825 43.785 71.505 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.635 70.825 45.985 71.735 ;
        RECT 47.365 71.505 48.285 71.725 ;
        RECT 54.365 71.625 55.285 71.735 ;
        RECT 52.950 71.505 55.285 71.625 ;
        RECT 46.005 70.825 55.285 71.505 ;
        RECT 55.860 70.825 59.335 71.735 ;
        RECT 59.345 70.825 62.820 71.735 ;
        RECT 63.510 71.505 64.855 71.735 ;
        RECT 63.025 70.825 64.855 71.505 ;
        RECT 64.865 70.825 68.535 71.635 ;
        RECT 68.545 70.825 69.915 71.635 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 70.385 70.825 72.995 71.735 ;
        RECT 73.145 70.825 75.895 71.635 ;
        RECT 76.560 70.825 80.035 71.735 ;
        RECT 80.240 70.825 83.715 71.735 ;
        RECT 83.725 70.825 87.200 71.735 ;
        RECT 87.405 70.825 90.880 71.735 ;
        RECT 91.085 70.825 94.560 71.735 ;
        RECT 95.695 70.910 96.125 71.695 ;
        RECT 96.145 70.825 99.620 71.735 ;
        RECT 99.825 70.825 101.195 71.605 ;
        RECT 102.565 71.505 103.485 71.725 ;
        RECT 109.565 71.625 110.485 71.735 ;
        RECT 108.150 71.505 110.485 71.625 ;
        RECT 113.145 71.505 114.065 71.725 ;
        RECT 120.145 71.625 121.065 71.735 ;
        RECT 118.730 71.505 121.065 71.625 ;
        RECT 101.205 70.825 110.485 71.505 ;
        RECT 111.785 70.825 121.065 71.505 ;
        RECT 121.455 70.910 121.885 71.695 ;
        RECT 121.915 70.825 123.265 71.735 ;
        RECT 124.205 70.825 125.575 71.635 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.615 7.215 70.825 ;
        RECT 12.565 70.615 12.735 70.825 ;
        RECT 13.950 70.615 14.120 70.805 ;
        RECT 16.705 70.615 16.875 70.805 ;
        RECT 18.080 70.665 18.200 70.775 ;
        RECT 19.005 70.635 19.175 70.825 ;
        RECT 22.225 70.615 22.395 70.805 ;
        RECT 23.600 70.635 23.770 70.825 ;
        RECT 27.280 70.635 27.450 70.825 ;
        RECT 27.745 70.615 27.915 70.825 ;
        RECT 29.580 70.665 29.700 70.775 ;
        RECT 30.045 70.615 30.215 70.805 ;
        RECT 31.885 70.615 32.055 70.805 ;
        RECT 33.265 70.635 33.435 70.825 ;
        RECT 34.645 70.635 34.815 70.825 ;
        RECT 41.545 70.615 41.715 70.805 ;
        RECT 45.685 70.635 45.855 70.825 ;
        RECT 46.145 70.635 46.315 70.825 ;
        RECT 47.065 70.615 47.235 70.805 ;
        RECT 49.825 70.615 49.995 70.805 ;
        RECT 50.560 70.615 50.730 70.805 ;
        RECT 54.425 70.615 54.595 70.805 ;
        RECT 57.645 70.615 57.815 70.805 ;
        RECT 59.020 70.635 59.190 70.825 ;
        RECT 59.490 70.635 59.660 70.825 ;
        RECT 61.335 70.660 61.495 70.770 ;
        RECT 63.165 70.635 63.335 70.825 ;
        RECT 63.625 70.615 63.795 70.805 ;
        RECT 65.005 70.635 65.175 70.825 ;
        RECT 65.465 70.615 65.635 70.805 ;
        RECT 65.925 70.615 66.095 70.805 ;
        RECT 67.765 70.615 67.935 70.805 ;
        RECT 68.685 70.635 68.855 70.825 ;
        RECT 69.605 70.615 69.775 70.805 ;
        RECT 70.530 70.635 70.700 70.825 ;
        RECT 73.285 70.775 73.455 70.825 ;
        RECT 73.280 70.665 73.455 70.775 ;
        RECT 73.285 70.635 73.455 70.665 ;
        RECT 74.020 70.615 74.190 70.805 ;
        RECT 76.040 70.665 76.160 70.775 ;
        RECT 77.885 70.615 78.055 70.805 ;
        RECT 79.720 70.635 79.890 70.825 ;
        RECT 81.565 70.615 81.735 70.805 ;
        RECT 83.400 70.635 83.570 70.825 ;
        RECT 83.870 70.635 84.040 70.825 ;
        RECT 86.625 70.615 86.795 70.805 ;
        RECT 87.550 70.635 87.720 70.825 ;
        RECT 90.305 70.615 90.475 70.805 ;
        RECT 90.765 70.615 90.935 70.805 ;
        RECT 91.230 70.635 91.400 70.825 ;
        RECT 94.915 70.670 95.075 70.780 ;
        RECT 96.290 70.635 96.460 70.825 ;
        RECT 97.850 70.615 98.020 70.805 ;
        RECT 99.505 70.615 99.675 70.805 ;
        RECT 99.965 70.615 100.135 70.825 ;
        RECT 101.345 70.635 101.515 70.825 ;
        RECT 101.620 70.615 101.790 70.805 ;
        RECT 105.495 70.660 105.655 70.770 ;
        RECT 107.325 70.615 107.495 70.805 ;
        RECT 107.795 70.660 107.955 70.770 ;
        RECT 109.165 70.615 109.335 70.805 ;
        RECT 111.015 70.670 111.175 70.780 ;
        RECT 111.925 70.635 112.095 70.825 ;
        RECT 114.680 70.665 114.800 70.775 ;
        RECT 118.550 70.615 118.720 70.805 ;
        RECT 119.285 70.615 119.455 70.805 ;
        RECT 122.045 70.635 122.215 70.825 ;
        RECT 122.965 70.615 123.135 70.805 ;
        RECT 123.435 70.670 123.595 70.780 ;
        RECT 125.265 70.615 125.435 70.825 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 6.905 69.805 12.415 70.615 ;
        RECT 12.425 69.805 13.795 70.615 ;
        RECT 13.805 69.705 16.415 70.615 ;
        RECT 16.565 69.805 22.075 70.615 ;
        RECT 22.085 69.805 27.595 70.615 ;
        RECT 27.605 69.805 29.435 70.615 ;
        RECT 29.905 69.835 31.275 70.615 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 31.745 69.935 41.025 70.615 ;
        RECT 33.105 69.715 34.025 69.935 ;
        RECT 38.690 69.815 41.025 69.935 ;
        RECT 40.105 69.705 41.025 69.815 ;
        RECT 41.405 69.805 46.915 70.615 ;
        RECT 46.925 69.805 48.755 70.615 ;
        RECT 48.765 69.835 50.135 70.615 ;
        RECT 50.145 69.935 54.045 70.615 ;
        RECT 50.145 69.705 51.075 69.935 ;
        RECT 54.285 69.805 57.035 70.615 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.505 69.805 61.175 70.615 ;
        RECT 62.105 69.935 63.935 70.615 ;
        RECT 63.945 69.935 65.775 70.615 ;
        RECT 65.785 69.935 67.615 70.615 ;
        RECT 67.625 69.935 69.455 70.615 ;
        RECT 62.105 69.705 63.450 69.935 ;
        RECT 63.945 69.705 65.290 69.935 ;
        RECT 66.270 69.705 67.615 69.935 ;
        RECT 68.110 69.705 69.455 69.935 ;
        RECT 69.465 69.805 73.135 70.615 ;
        RECT 73.605 69.935 77.505 70.615 ;
        RECT 73.605 69.705 74.535 69.935 ;
        RECT 77.745 69.805 81.415 70.615 ;
        RECT 81.425 69.805 82.795 70.615 ;
        RECT 82.815 69.745 83.245 70.530 ;
        RECT 83.360 69.935 86.825 70.615 ;
        RECT 87.040 69.935 90.505 70.615 ;
        RECT 83.360 69.705 84.280 69.935 ;
        RECT 87.040 69.705 87.960 69.935 ;
        RECT 90.625 69.805 94.295 70.615 ;
        RECT 94.535 69.935 98.435 70.615 ;
        RECT 97.505 69.705 98.435 69.935 ;
        RECT 98.445 69.835 99.815 70.615 ;
        RECT 99.825 69.805 101.195 70.615 ;
        RECT 101.205 69.935 105.105 70.615 ;
        RECT 101.205 69.705 102.135 69.935 ;
        RECT 106.275 69.705 107.625 70.615 ;
        RECT 108.575 69.745 109.005 70.530 ;
        RECT 109.025 69.805 114.535 70.615 ;
        RECT 115.235 69.935 119.135 70.615 ;
        RECT 118.205 69.705 119.135 69.935 ;
        RECT 119.145 69.805 122.815 70.615 ;
        RECT 122.825 69.805 124.195 70.615 ;
        RECT 124.205 69.805 125.575 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 125.770 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 6.905 65.385 10.575 66.195 ;
        RECT 10.680 66.065 11.600 66.295 ;
        RECT 14.265 66.065 15.195 66.295 ;
        RECT 10.680 65.385 14.145 66.065 ;
        RECT 14.265 65.385 18.165 66.065 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 18.865 66.065 19.795 66.295 ;
        RECT 26.580 66.065 27.500 66.295 ;
        RECT 30.260 66.065 31.180 66.295 ;
        RECT 18.865 65.385 22.765 66.065 ;
        RECT 24.035 65.385 27.500 66.065 ;
        RECT 27.715 65.385 31.180 66.065 ;
        RECT 31.285 66.065 32.215 66.295 ;
        RECT 31.285 65.385 35.185 66.065 ;
        RECT 35.435 65.385 36.785 66.295 ;
        RECT 36.805 65.385 42.315 66.195 ;
        RECT 42.325 65.385 44.155 66.195 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.635 65.385 45.985 66.295 ;
        RECT 46.005 65.385 47.375 66.195 ;
        RECT 47.395 65.385 48.745 66.295 ;
        RECT 48.765 65.385 50.135 66.165 ;
        RECT 51.065 66.065 51.995 66.295 ;
        RECT 51.065 65.385 54.965 66.065 ;
        RECT 55.205 65.385 60.715 66.195 ;
        RECT 61.670 66.065 63.015 66.295 ;
        RECT 61.185 65.385 63.015 66.065 ;
        RECT 63.025 65.385 65.635 66.295 ;
        RECT 65.785 65.385 68.525 66.065 ;
        RECT 68.545 65.385 69.915 66.165 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 74.895 66.065 75.825 66.285 ;
        RECT 78.655 66.065 79.575 66.295 ;
        RECT 70.385 65.385 79.575 66.065 ;
        RECT 79.585 66.065 80.515 66.295 ;
        RECT 83.820 66.065 84.740 66.295 ;
        RECT 90.605 66.065 91.535 66.295 ;
        RECT 94.200 66.065 95.120 66.295 ;
        RECT 79.585 65.385 83.485 66.065 ;
        RECT 83.820 65.385 87.285 66.065 ;
        RECT 87.635 65.385 91.535 66.065 ;
        RECT 91.655 65.385 95.120 66.065 ;
        RECT 95.695 65.470 96.125 66.255 ;
        RECT 97.505 66.065 98.425 66.285 ;
        RECT 104.505 66.185 105.425 66.295 ;
        RECT 103.090 66.065 105.425 66.185 ;
        RECT 96.145 65.385 105.425 66.065 ;
        RECT 105.805 65.385 111.315 66.195 ;
        RECT 111.325 65.385 114.075 66.195 ;
        RECT 117.745 66.065 118.675 66.295 ;
        RECT 114.775 65.385 118.675 66.065 ;
        RECT 118.685 65.385 120.055 66.165 ;
        RECT 120.075 65.385 121.425 66.295 ;
        RECT 121.455 65.470 121.885 66.255 ;
        RECT 121.905 65.385 123.735 66.195 ;
        RECT 124.205 65.385 125.575 66.195 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.175 7.215 65.385 ;
        RECT 10.725 65.175 10.895 65.365 ;
        RECT 11.185 65.175 11.355 65.365 ;
        RECT 12.565 65.175 12.735 65.365 ;
        RECT 13.945 65.195 14.115 65.385 ;
        RECT 14.680 65.195 14.850 65.385 ;
        RECT 19.280 65.195 19.450 65.385 ;
        RECT 21.765 65.195 21.935 65.365 ;
        RECT 23.155 65.230 23.315 65.340 ;
        RECT 23.615 65.220 23.775 65.330 ;
        RECT 24.065 65.195 24.235 65.385 ;
        RECT 27.745 65.195 27.915 65.385 ;
        RECT 27.930 65.175 28.100 65.365 ;
        RECT 29.585 65.175 29.755 65.365 ;
        RECT 30.045 65.175 30.215 65.365 ;
        RECT 31.700 65.195 31.870 65.385 ;
        RECT 31.885 65.175 32.055 65.365 ;
        RECT 35.565 65.195 35.735 65.385 ;
        RECT 36.485 65.175 36.655 65.365 ;
        RECT 36.945 65.175 37.115 65.385 ;
        RECT 40.635 65.220 40.795 65.330 ;
        RECT 42.465 65.195 42.635 65.385 ;
        RECT 44.765 65.175 44.935 65.385 ;
        RECT 45.235 65.220 45.395 65.330 ;
        RECT 46.145 65.175 46.315 65.385 ;
        RECT 47.525 65.195 47.695 65.385 ;
        RECT 49.825 65.195 49.995 65.385 ;
        RECT 50.295 65.230 50.455 65.340 ;
        RECT 51.480 65.195 51.650 65.385 ;
        RECT 55.345 65.195 55.515 65.385 ;
        RECT 55.805 65.175 55.975 65.365 ;
        RECT 57.920 65.175 58.090 65.365 ;
        RECT 60.860 65.225 60.980 65.335 ;
        RECT 61.325 65.195 61.495 65.385 ;
        RECT 63.170 65.195 63.340 65.385 ;
        RECT 64.085 65.175 64.255 65.365 ;
        RECT 64.545 65.175 64.715 65.365 ;
        RECT 65.925 65.195 66.095 65.385 ;
        RECT 68.685 65.195 68.855 65.385 ;
        RECT 70.075 65.220 70.235 65.330 ;
        RECT 70.525 65.195 70.695 65.385 ;
        RECT 71.905 65.175 72.075 65.365 ;
        RECT 72.365 65.175 72.535 65.365 ;
        RECT 80.000 65.195 80.170 65.385 ;
        RECT 82.485 65.175 82.655 65.365 ;
        RECT 83.680 65.175 83.850 65.365 ;
        RECT 87.085 65.195 87.255 65.385 ;
        RECT 87.540 65.225 87.660 65.335 ;
        RECT 88.005 65.175 88.175 65.365 ;
        RECT 90.950 65.195 91.120 65.385 ;
        RECT 91.685 65.195 91.855 65.385 ;
        RECT 95.360 65.225 95.480 65.335 ;
        RECT 96.285 65.195 96.455 65.385 ;
        RECT 97.205 65.175 97.375 65.365 ;
        RECT 100.885 65.175 101.055 65.365 ;
        RECT 102.265 65.175 102.435 65.365 ;
        RECT 105.945 65.175 106.115 65.385 ;
        RECT 107.325 65.175 107.495 65.365 ;
        RECT 109.440 65.175 109.610 65.365 ;
        RECT 111.465 65.195 111.635 65.385 ;
        RECT 113.305 65.175 113.475 65.365 ;
        RECT 114.220 65.225 114.340 65.335 ;
        RECT 118.090 65.195 118.260 65.385 ;
        RECT 119.745 65.195 119.915 65.385 ;
        RECT 121.125 65.195 121.295 65.385 ;
        RECT 122.045 65.195 122.215 65.385 ;
        RECT 122.965 65.175 123.135 65.365 ;
        RECT 123.880 65.225 124.000 65.335 ;
        RECT 125.265 65.175 125.435 65.385 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.365 9.655 65.175 ;
        RECT 9.665 64.395 11.035 65.175 ;
        RECT 11.045 64.395 12.415 65.175 ;
        RECT 12.425 64.495 21.615 65.175 ;
        RECT 22.090 64.495 23.455 65.175 ;
        RECT 24.615 64.495 28.515 65.175 ;
        RECT 16.935 64.275 17.865 64.495 ;
        RECT 20.695 64.265 21.615 64.495 ;
        RECT 27.585 64.265 28.515 64.495 ;
        RECT 28.525 64.395 29.895 65.175 ;
        RECT 29.905 64.365 31.275 65.175 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 31.745 64.365 33.115 65.175 ;
        RECT 33.220 64.495 36.685 65.175 ;
        RECT 33.220 64.265 34.140 64.495 ;
        RECT 36.805 64.365 40.475 65.175 ;
        RECT 41.500 64.495 44.965 65.175 ;
        RECT 46.005 64.495 55.285 65.175 ;
        RECT 41.500 64.265 42.420 64.495 ;
        RECT 47.365 64.275 48.285 64.495 ;
        RECT 52.950 64.375 55.285 64.495 ;
        RECT 54.365 64.265 55.285 64.375 ;
        RECT 55.665 64.365 57.035 65.175 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.505 64.495 61.405 65.175 ;
        RECT 57.505 64.265 58.435 64.495 ;
        RECT 61.675 64.265 64.395 65.175 ;
        RECT 64.405 64.365 69.915 65.175 ;
        RECT 70.855 64.265 72.205 65.175 ;
        RECT 72.225 64.495 81.415 65.175 ;
        RECT 76.735 64.275 77.665 64.495 ;
        RECT 80.495 64.265 81.415 64.495 ;
        RECT 81.425 64.395 82.795 65.175 ;
        RECT 82.815 64.305 83.245 65.090 ;
        RECT 83.265 64.495 87.165 65.175 ;
        RECT 87.865 64.495 97.055 65.175 ;
        RECT 97.175 64.495 100.640 65.175 ;
        RECT 83.265 64.265 84.195 64.495 ;
        RECT 92.375 64.275 93.305 64.495 ;
        RECT 96.135 64.265 97.055 64.495 ;
        RECT 99.720 64.265 100.640 64.495 ;
        RECT 100.755 64.265 102.105 65.175 ;
        RECT 102.125 64.365 105.795 65.175 ;
        RECT 105.805 64.365 107.175 65.175 ;
        RECT 107.185 64.395 108.555 65.175 ;
        RECT 108.575 64.305 109.005 65.090 ;
        RECT 109.025 64.495 112.925 65.175 ;
        RECT 113.165 64.495 122.445 65.175 ;
        RECT 109.025 64.265 109.955 64.495 ;
        RECT 114.525 64.275 115.445 64.495 ;
        RECT 120.110 64.375 122.445 64.495 ;
        RECT 121.525 64.265 122.445 64.375 ;
        RECT 122.825 64.365 124.195 65.175 ;
        RECT 124.205 64.365 125.575 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 125.770 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 6.905 59.945 8.275 60.755 ;
        RECT 12.795 60.625 13.725 60.845 ;
        RECT 16.555 60.625 17.475 60.855 ;
        RECT 8.285 59.945 17.475 60.625 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 18.865 60.625 19.795 60.855 ;
        RECT 28.435 60.625 29.365 60.845 ;
        RECT 32.195 60.625 33.115 60.855 ;
        RECT 18.865 59.945 22.765 60.625 ;
        RECT 23.925 59.945 33.115 60.625 ;
        RECT 33.135 59.945 34.485 60.855 ;
        RECT 34.505 59.945 38.175 60.755 ;
        RECT 38.185 60.625 39.115 60.855 ;
        RECT 38.185 59.945 42.085 60.625 ;
        RECT 42.325 59.945 44.155 60.755 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 45.985 60.625 46.905 60.845 ;
        RECT 52.985 60.745 53.905 60.855 ;
        RECT 51.570 60.625 53.905 60.745 ;
        RECT 44.625 59.945 53.905 60.625 ;
        RECT 54.285 59.945 57.955 60.755 ;
        RECT 57.965 59.945 59.335 60.755 ;
        RECT 59.355 59.945 62.095 60.625 ;
        RECT 62.105 59.945 65.775 60.755 ;
        RECT 65.785 59.945 68.395 60.855 ;
        RECT 68.545 59.945 69.915 60.755 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 74.055 60.755 ;
        RECT 74.065 59.945 75.435 60.725 ;
        RECT 75.445 59.945 77.275 60.755 ;
        RECT 77.295 59.945 78.645 60.855 ;
        RECT 83.635 60.625 84.565 60.845 ;
        RECT 87.395 60.625 88.315 60.855 ;
        RECT 79.125 59.945 88.315 60.625 ;
        RECT 88.880 60.625 89.800 60.855 ;
        RECT 88.880 59.945 92.345 60.625 ;
        RECT 92.475 59.945 93.825 60.855 ;
        RECT 93.845 59.945 95.215 60.725 ;
        RECT 95.695 60.030 96.125 60.815 ;
        RECT 96.155 59.945 97.505 60.855 ;
        RECT 97.525 59.945 103.035 60.755 ;
        RECT 103.045 59.945 105.795 60.755 ;
        RECT 106.265 60.625 107.185 60.855 ;
        RECT 110.015 60.625 110.945 60.845 ;
        RECT 106.265 59.945 115.455 60.625 ;
        RECT 115.465 59.945 120.975 60.755 ;
        RECT 121.455 60.030 121.885 60.815 ;
        RECT 121.905 59.945 123.735 60.755 ;
        RECT 124.205 59.945 125.575 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.045 59.735 7.215 59.945 ;
        RECT 8.425 59.755 8.595 59.945 ;
        RECT 11.645 59.735 11.815 59.925 ;
        RECT 13.025 59.735 13.195 59.925 ;
        RECT 16.705 59.735 16.875 59.925 ;
        RECT 17.635 59.790 17.795 59.900 ;
        RECT 19.280 59.755 19.450 59.945 ;
        RECT 20.385 59.735 20.555 59.925 ;
        RECT 21.765 59.735 21.935 59.925 ;
        RECT 23.155 59.790 23.315 59.900 ;
        RECT 24.065 59.755 24.235 59.945 ;
        RECT 30.965 59.735 31.135 59.925 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 33.265 59.735 33.435 59.925 ;
        RECT 34.185 59.755 34.355 59.945 ;
        RECT 34.645 59.755 34.815 59.945 ;
        RECT 38.600 59.755 38.770 59.945 ;
        RECT 42.465 59.735 42.635 59.945 ;
        RECT 44.765 59.755 44.935 59.945 ;
        RECT 46.155 59.780 46.315 59.890 ;
        RECT 47.985 59.735 48.155 59.925 ;
        RECT 48.445 59.735 48.615 59.925 ;
        RECT 53.965 59.735 54.135 59.925 ;
        RECT 54.425 59.755 54.595 59.945 ;
        RECT 56.720 59.785 56.840 59.895 ;
        RECT 57.645 59.735 57.815 59.925 ;
        RECT 58.105 59.755 58.275 59.945 ;
        RECT 61.325 59.735 61.495 59.925 ;
        RECT 61.785 59.755 61.955 59.945 ;
        RECT 62.245 59.755 62.415 59.945 ;
        RECT 62.705 59.735 62.875 59.925 ;
        RECT 65.465 59.735 65.635 59.925 ;
        RECT 65.930 59.755 66.100 59.945 ;
        RECT 68.685 59.755 68.855 59.945 ;
        RECT 70.525 59.755 70.695 59.945 ;
        RECT 70.990 59.735 71.160 59.925 ;
        RECT 73.745 59.735 73.915 59.925 ;
        RECT 75.125 59.755 75.295 59.945 ;
        RECT 75.585 59.755 75.755 59.945 ;
        RECT 77.425 59.755 77.595 59.945 ;
        RECT 78.800 59.785 78.920 59.895 ;
        RECT 79.265 59.735 79.435 59.945 ;
        RECT 81.105 59.755 81.275 59.925 ;
        RECT 88.460 59.785 88.580 59.895 ;
        RECT 92.145 59.735 92.315 59.945 ;
        RECT 92.605 59.735 92.775 59.925 ;
        RECT 93.525 59.755 93.695 59.945 ;
        RECT 94.905 59.755 95.075 59.945 ;
        RECT 95.360 59.785 95.480 59.895 ;
        RECT 97.205 59.755 97.375 59.945 ;
        RECT 97.665 59.755 97.835 59.945 ;
        RECT 98.125 59.735 98.295 59.925 ;
        RECT 100.880 59.785 101.000 59.895 ;
        RECT 101.345 59.735 101.515 59.925 ;
        RECT 103.185 59.755 103.355 59.945 ;
        RECT 105.940 59.785 106.060 59.895 ;
        RECT 107.320 59.735 107.490 59.925 ;
        RECT 107.795 59.780 107.955 59.890 ;
        RECT 109.165 59.735 109.335 59.925 ;
        RECT 111.465 59.735 111.635 59.925 ;
        RECT 111.925 59.735 112.095 59.925 ;
        RECT 115.145 59.755 115.315 59.945 ;
        RECT 115.605 59.755 115.775 59.945 ;
        RECT 117.445 59.735 117.615 59.925 ;
        RECT 121.120 59.785 121.240 59.895 ;
        RECT 122.045 59.755 122.215 59.945 ;
        RECT 122.965 59.735 123.135 59.925 ;
        RECT 123.880 59.785 124.000 59.895 ;
        RECT 125.265 59.735 125.435 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 58.925 10.575 59.735 ;
        RECT 10.585 58.955 11.955 59.735 ;
        RECT 11.975 58.825 13.325 59.735 ;
        RECT 13.440 59.055 16.905 59.735 ;
        RECT 17.120 59.055 20.585 59.735 ;
        RECT 13.440 58.825 14.360 59.055 ;
        RECT 17.120 58.825 18.040 59.055 ;
        RECT 20.715 58.825 22.065 59.735 ;
        RECT 22.170 59.055 31.275 59.735 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 58.925 33.115 59.735 ;
        RECT 33.125 59.055 42.315 59.735 ;
        RECT 37.635 58.835 38.565 59.055 ;
        RECT 41.395 58.825 42.315 59.055 ;
        RECT 42.325 58.925 45.995 59.735 ;
        RECT 46.925 58.955 48.295 59.735 ;
        RECT 48.305 58.925 53.815 59.735 ;
        RECT 53.825 58.925 56.575 59.735 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 57.505 58.925 61.175 59.735 ;
        RECT 61.185 58.925 62.555 59.735 ;
        RECT 62.565 59.055 65.305 59.735 ;
        RECT 65.325 58.925 70.835 59.735 ;
        RECT 70.845 58.825 73.455 59.735 ;
        RECT 73.605 58.925 79.115 59.735 ;
        RECT 79.125 58.925 80.955 59.735 ;
        RECT 81.430 59.055 82.795 59.735 ;
        RECT 82.815 58.865 83.245 59.650 ;
        RECT 83.350 59.055 92.455 59.735 ;
        RECT 92.465 58.925 97.975 59.735 ;
        RECT 97.985 58.925 100.735 59.735 ;
        RECT 101.205 58.925 103.295 59.735 ;
        RECT 104.160 58.825 107.635 59.735 ;
        RECT 108.575 58.865 109.005 59.650 ;
        RECT 109.025 58.925 110.395 59.735 ;
        RECT 110.415 58.825 111.765 59.735 ;
        RECT 111.785 58.925 117.295 59.735 ;
        RECT 117.305 58.925 122.815 59.735 ;
        RECT 122.825 58.925 124.195 59.735 ;
        RECT 124.205 58.925 125.575 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 125.770 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 54.505 8.275 55.315 ;
        RECT 12.795 55.185 13.725 55.405 ;
        RECT 16.555 55.185 17.475 55.415 ;
        RECT 8.285 54.505 17.475 55.185 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 21.980 55.185 22.900 55.415 ;
        RECT 19.435 54.505 22.900 55.185 ;
        RECT 23.200 54.505 26.675 55.415 ;
        RECT 26.685 54.505 32.195 55.315 ;
        RECT 32.205 54.505 35.875 55.315 ;
        RECT 35.885 54.505 37.255 55.285 ;
        RECT 38.195 54.505 39.545 55.415 ;
        RECT 40.490 54.505 41.855 55.185 ;
        RECT 41.865 54.505 43.695 55.315 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 44.625 54.505 46.455 55.315 ;
        RECT 47.065 54.505 49.675 55.415 ;
        RECT 49.695 54.505 52.435 55.185 ;
        RECT 52.445 54.505 57.955 55.315 ;
        RECT 57.965 54.505 61.635 55.315 ;
        RECT 62.135 54.505 64.855 55.415 ;
        RECT 65.325 55.185 66.670 55.415 ;
        RECT 67.650 55.185 68.995 55.415 ;
        RECT 65.325 54.505 67.155 55.185 ;
        RECT 67.165 54.505 68.995 55.185 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 70.385 54.505 75.895 55.315 ;
        RECT 75.905 54.505 81.415 55.315 ;
        RECT 81.425 54.505 86.935 55.315 ;
        RECT 86.945 54.505 89.695 55.315 ;
        RECT 89.900 54.505 93.375 55.415 ;
        RECT 93.385 54.505 95.215 55.315 ;
        RECT 95.695 54.590 96.125 55.375 ;
        RECT 96.145 54.505 97.975 55.315 ;
        RECT 98.640 54.505 102.115 55.415 ;
        RECT 102.125 54.505 111.230 55.185 ;
        RECT 111.335 54.505 112.685 55.415 ;
        RECT 112.705 54.505 118.215 55.315 ;
        RECT 118.225 54.505 120.975 55.315 ;
        RECT 121.455 54.590 121.885 55.375 ;
        RECT 121.905 54.505 123.735 55.315 ;
        RECT 124.205 54.505 125.575 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.045 54.295 7.215 54.505 ;
        RECT 8.425 54.315 8.595 54.505 ;
        RECT 9.800 54.345 9.920 54.455 ;
        RECT 10.265 54.295 10.435 54.485 ;
        RECT 12.105 54.295 12.275 54.485 ;
        RECT 13.940 54.345 14.060 54.455 ;
        RECT 15.325 54.295 15.495 54.485 ;
        RECT 15.785 54.295 15.955 54.485 ;
        RECT 17.635 54.350 17.795 54.460 ;
        RECT 19.000 54.345 19.120 54.455 ;
        RECT 19.465 54.315 19.635 54.505 ;
        RECT 22.680 54.295 22.850 54.485 ;
        RECT 26.360 54.295 26.530 54.505 ;
        RECT 26.825 54.315 26.995 54.505 ;
        RECT 30.040 54.295 30.210 54.485 ;
        RECT 30.515 54.340 30.675 54.450 ;
        RECT 31.885 54.295 32.055 54.485 ;
        RECT 32.345 54.315 32.515 54.505 ;
        RECT 36.480 54.295 36.650 54.485 ;
        RECT 36.945 54.295 37.115 54.505 ;
        RECT 37.415 54.350 37.575 54.460 ;
        RECT 38.325 54.315 38.495 54.505 ;
        RECT 39.700 54.345 39.820 54.455 ;
        RECT 40.165 54.315 40.335 54.485 ;
        RECT 42.005 54.315 42.175 54.505 ;
        RECT 43.840 54.345 43.960 54.455 ;
        RECT 44.765 54.315 44.935 54.505 ;
        RECT 49.360 54.485 49.530 54.505 ;
        RECT 46.600 54.345 46.720 54.455 ;
        RECT 48.905 54.295 49.075 54.485 ;
        RECT 49.360 54.315 49.535 54.485 ;
        RECT 51.200 54.345 51.320 54.455 ;
        RECT 52.125 54.315 52.295 54.505 ;
        RECT 52.585 54.315 52.755 54.505 ;
        RECT 49.365 54.295 49.535 54.315 ;
        RECT 54.880 54.295 55.050 54.485 ;
        RECT 55.345 54.295 55.515 54.485 ;
        RECT 57.655 54.340 57.815 54.450 ;
        RECT 58.105 54.315 58.275 54.505 ;
        RECT 59.945 54.295 60.115 54.485 ;
        RECT 61.785 54.455 61.955 54.485 ;
        RECT 61.780 54.345 61.955 54.455 ;
        RECT 61.785 54.295 61.955 54.345 ;
        RECT 62.245 54.295 62.415 54.485 ;
        RECT 64.545 54.315 64.715 54.505 ;
        RECT 65.000 54.345 65.120 54.455 ;
        RECT 66.845 54.315 67.015 54.505 ;
        RECT 67.305 54.315 67.475 54.505 ;
        RECT 69.155 54.350 69.315 54.460 ;
        RECT 69.605 54.315 69.775 54.485 ;
        RECT 69.605 54.295 69.675 54.315 ;
        RECT 70.065 54.295 70.235 54.485 ;
        RECT 70.525 54.315 70.695 54.505 ;
        RECT 71.905 54.295 72.075 54.485 ;
        RECT 76.045 54.315 76.215 54.505 ;
        RECT 77.425 54.295 77.595 54.485 ;
        RECT 81.565 54.315 81.735 54.505 ;
        RECT 83.405 54.295 83.575 54.485 ;
        RECT 87.085 54.315 87.255 54.505 ;
        RECT 88.000 54.295 88.170 54.485 ;
        RECT 88.470 54.295 88.640 54.485 ;
        RECT 93.060 54.315 93.230 54.505 ;
        RECT 93.525 54.315 93.695 54.505 ;
        RECT 95.360 54.295 95.530 54.485 ;
        RECT 95.825 54.295 95.995 54.485 ;
        RECT 96.285 54.315 96.455 54.505 ;
        RECT 98.120 54.345 98.240 54.455 ;
        RECT 99.505 54.295 99.675 54.485 ;
        RECT 101.800 54.315 101.970 54.505 ;
        RECT 102.265 54.315 102.435 54.505 ;
        RECT 112.385 54.295 112.555 54.505 ;
        RECT 112.845 54.485 113.015 54.505 ;
        RECT 112.845 54.315 113.020 54.485 ;
        RECT 112.850 54.295 113.020 54.315 ;
        RECT 116.525 54.295 116.695 54.485 ;
        RECT 118.365 54.315 118.535 54.505 ;
        RECT 121.120 54.345 121.240 54.455 ;
        RECT 122.045 54.295 122.215 54.505 ;
        RECT 123.880 54.345 124.000 54.455 ;
        RECT 125.265 54.295 125.435 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.485 9.655 54.295 ;
        RECT 10.125 53.615 11.955 54.295 ;
        RECT 11.965 53.485 13.795 54.295 ;
        RECT 14.275 53.385 15.625 54.295 ;
        RECT 15.645 53.485 19.315 54.295 ;
        RECT 19.520 53.385 22.995 54.295 ;
        RECT 23.200 53.385 26.675 54.295 ;
        RECT 26.880 53.385 30.355 54.295 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.745 53.485 33.115 54.295 ;
        RECT 33.320 53.385 36.795 54.295 ;
        RECT 36.805 53.485 39.555 54.295 ;
        RECT 40.110 53.615 49.215 54.295 ;
        RECT 49.225 53.485 51.055 54.295 ;
        RECT 51.720 53.385 55.195 54.295 ;
        RECT 55.205 53.485 57.035 54.295 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 58.425 53.615 60.255 54.295 ;
        RECT 60.265 53.615 62.095 54.295 ;
        RECT 62.105 54.065 63.675 54.295 ;
        RECT 65.765 54.255 66.685 54.295 ;
        RECT 65.765 54.065 66.695 54.255 ;
        RECT 67.405 54.065 69.675 54.295 ;
        RECT 62.105 53.705 66.695 54.065 ;
        RECT 62.105 53.615 66.685 53.705 ;
        RECT 58.425 53.385 59.770 53.615 ;
        RECT 60.265 53.385 61.610 53.615 ;
        RECT 63.685 53.385 66.685 53.615 ;
        RECT 66.920 53.385 69.675 54.065 ;
        RECT 69.925 53.615 71.755 54.295 ;
        RECT 70.410 53.385 71.755 53.615 ;
        RECT 71.765 53.485 77.275 54.295 ;
        RECT 77.285 53.485 82.795 54.295 ;
        RECT 82.815 53.425 83.245 54.210 ;
        RECT 83.265 53.485 84.635 54.295 ;
        RECT 84.840 53.385 88.315 54.295 ;
        RECT 88.325 53.385 91.800 54.295 ;
        RECT 92.200 53.385 95.675 54.295 ;
        RECT 95.795 53.615 99.260 54.295 ;
        RECT 99.365 53.615 108.555 54.295 ;
        RECT 98.340 53.385 99.260 53.615 ;
        RECT 103.875 53.395 104.805 53.615 ;
        RECT 107.635 53.385 108.555 53.615 ;
        RECT 108.575 53.425 109.005 54.210 ;
        RECT 109.120 53.615 112.585 54.295 ;
        RECT 109.120 53.385 110.040 53.615 ;
        RECT 112.705 53.385 116.180 54.295 ;
        RECT 116.385 53.485 121.895 54.295 ;
        RECT 121.905 53.485 123.735 54.295 ;
        RECT 124.205 53.485 125.575 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 125.770 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 6.905 49.065 12.415 49.875 ;
        RECT 12.885 49.065 14.255 49.845 ;
        RECT 14.265 49.065 15.635 49.845 ;
        RECT 15.645 49.065 18.395 49.875 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 18.865 49.065 21.615 49.875 ;
        RECT 24.740 49.745 25.660 49.975 ;
        RECT 22.195 49.065 25.660 49.745 ;
        RECT 25.960 49.065 29.435 49.975 ;
        RECT 29.540 49.745 30.460 49.975 ;
        RECT 29.540 49.065 33.005 49.745 ;
        RECT 33.125 49.065 34.495 49.875 ;
        RECT 37.705 49.745 38.635 49.975 ;
        RECT 34.735 49.065 38.635 49.745 ;
        RECT 38.740 49.745 39.660 49.975 ;
        RECT 38.740 49.065 42.205 49.745 ;
        RECT 42.785 49.065 44.155 49.845 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 45.640 49.745 46.560 49.975 ;
        RECT 45.640 49.065 49.105 49.745 ;
        RECT 49.365 49.065 51.975 49.975 ;
        RECT 52.640 49.065 56.115 49.975 ;
        RECT 56.125 49.065 59.600 49.975 ;
        RECT 59.805 49.065 61.635 49.875 ;
        RECT 61.860 49.295 64.615 49.975 ;
        RECT 65.080 49.295 67.835 49.975 ;
        RECT 62.345 49.065 64.615 49.295 ;
        RECT 65.565 49.065 67.835 49.295 ;
        RECT 68.095 49.065 69.445 49.975 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 70.385 49.065 74.055 49.875 ;
        RECT 74.065 49.065 76.805 49.745 ;
        RECT 77.020 49.065 80.495 49.975 ;
        RECT 80.600 49.745 81.520 49.975 ;
        RECT 80.600 49.065 84.065 49.745 ;
        RECT 85.105 49.065 86.475 49.845 ;
        RECT 90.995 49.745 91.925 49.965 ;
        RECT 94.755 49.745 95.675 49.975 ;
        RECT 86.485 49.065 95.675 49.745 ;
        RECT 95.695 49.150 96.125 49.935 ;
        RECT 96.155 49.065 97.505 49.975 ;
        RECT 97.985 49.745 98.915 49.975 ;
        RECT 97.985 49.065 101.885 49.745 ;
        RECT 102.125 49.065 103.495 49.845 ;
        RECT 106.705 49.745 107.635 49.975 ;
        RECT 112.155 49.745 113.085 49.965 ;
        RECT 115.915 49.745 116.835 49.975 ;
        RECT 103.735 49.065 107.635 49.745 ;
        RECT 107.645 49.065 116.835 49.745 ;
        RECT 116.845 49.065 120.515 49.875 ;
        RECT 121.455 49.150 121.885 49.935 ;
        RECT 121.905 49.065 123.735 49.875 ;
        RECT 124.205 49.065 125.575 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.045 48.855 7.215 49.065 ;
        RECT 10.735 48.900 10.895 49.010 ;
        RECT 11.645 48.855 11.815 49.045 ;
        RECT 12.560 48.905 12.680 49.015 ;
        RECT 13.945 48.875 14.115 49.065 ;
        RECT 15.325 48.875 15.495 49.065 ;
        RECT 15.785 48.875 15.955 49.065 ;
        RECT 19.005 48.875 19.175 49.065 ;
        RECT 21.120 48.855 21.290 49.045 ;
        RECT 21.760 48.905 21.880 49.015 ;
        RECT 22.225 48.875 22.395 49.065 ;
        RECT 24.985 48.855 25.155 49.045 ;
        RECT 29.120 48.875 29.290 49.065 ;
        RECT 30.230 48.855 30.400 49.045 ;
        RECT 30.960 48.905 31.080 49.015 ;
        RECT 31.895 48.900 32.055 49.010 ;
        RECT 32.805 48.855 32.975 49.065 ;
        RECT 33.265 48.875 33.435 49.065 ;
        RECT 38.050 48.875 38.220 49.065 ;
        RECT 42.005 48.875 42.175 49.065 ;
        RECT 42.460 48.905 42.580 49.015 ;
        RECT 42.925 48.855 43.095 49.065 ;
        RECT 44.775 48.910 44.935 49.020 ;
        RECT 48.905 48.875 49.075 49.065 ;
        RECT 51.660 48.875 51.830 49.065 ;
        RECT 55.800 49.045 55.970 49.065 ;
        RECT 52.120 48.905 52.240 49.015 ;
        RECT 55.340 48.855 55.510 49.045 ;
        RECT 55.800 48.875 55.975 49.045 ;
        RECT 56.270 48.875 56.440 49.065 ;
        RECT 55.805 48.855 55.975 48.875 ;
        RECT 57.645 48.855 57.815 49.045 ;
        RECT 59.945 48.875 60.115 49.065 ;
        RECT 64.545 49.045 64.615 49.065 ;
        RECT 67.765 49.045 67.835 49.065 ;
        RECT 61.335 48.900 61.495 49.010 ;
        RECT 64.545 48.875 64.715 49.045 ;
        RECT 65.005 48.875 65.175 49.045 ;
        RECT 65.005 48.855 65.075 48.875 ;
        RECT 65.465 48.855 65.635 49.045 ;
        RECT 67.765 48.875 67.935 49.045 ;
        RECT 69.145 48.875 69.315 49.065 ;
        RECT 69.600 48.905 69.720 49.015 ;
        RECT 70.525 48.875 70.695 49.065 ;
        RECT 70.985 48.855 71.155 49.045 ;
        RECT 74.205 48.875 74.375 49.065 ;
        RECT 74.675 48.900 74.835 49.010 ;
        RECT 76.505 48.855 76.675 49.045 ;
        RECT 80.180 48.875 80.350 49.065 ;
        RECT 80.370 48.855 80.540 49.045 ;
        RECT 81.105 48.855 81.275 49.045 ;
        RECT 83.410 48.855 83.580 49.045 ;
        RECT 83.865 48.875 84.035 49.065 ;
        RECT 84.335 48.910 84.495 49.020 ;
        RECT 85.245 48.875 85.415 49.065 ;
        RECT 86.625 48.875 86.795 49.065 ;
        RECT 87.085 48.855 87.255 49.045 ;
        RECT 90.120 48.855 90.290 49.045 ;
        RECT 93.985 48.855 94.155 49.045 ;
        RECT 97.205 48.875 97.375 49.065 ;
        RECT 97.660 48.905 97.780 49.015 ;
        RECT 98.125 48.855 98.295 49.045 ;
        RECT 98.400 48.875 98.570 49.065 ;
        RECT 101.805 48.855 101.975 49.045 ;
        RECT 103.185 48.875 103.355 49.065 ;
        RECT 107.050 48.875 107.220 49.065 ;
        RECT 107.325 48.855 107.495 49.045 ;
        RECT 107.785 48.875 107.955 49.065 ;
        RECT 112.385 48.855 112.555 49.045 ;
        RECT 116.065 48.855 116.235 49.045 ;
        RECT 116.525 48.855 116.695 49.045 ;
        RECT 116.985 48.875 117.155 49.065 ;
        RECT 120.675 48.910 120.835 49.020 ;
        RECT 122.045 48.855 122.215 49.065 ;
        RECT 123.880 48.905 124.000 49.015 ;
        RECT 125.265 48.855 125.435 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.045 10.575 48.855 ;
        RECT 11.505 48.175 20.695 48.855 ;
        RECT 16.015 47.955 16.945 48.175 ;
        RECT 19.775 47.945 20.695 48.175 ;
        RECT 20.705 48.175 24.605 48.855 ;
        RECT 20.705 47.945 21.635 48.175 ;
        RECT 24.845 48.045 26.675 48.855 ;
        RECT 26.915 48.175 30.815 48.855 ;
        RECT 29.885 47.945 30.815 48.175 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 32.665 48.175 41.855 48.855 ;
        RECT 42.785 48.175 51.975 48.855 ;
        RECT 37.175 47.955 38.105 48.175 ;
        RECT 40.935 47.945 41.855 48.175 ;
        RECT 47.295 47.955 48.225 48.175 ;
        RECT 51.055 47.945 51.975 48.175 ;
        RECT 52.180 47.945 55.655 48.855 ;
        RECT 55.675 47.945 57.025 48.855 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.505 48.045 61.175 48.855 ;
        RECT 62.805 48.625 65.075 48.855 ;
        RECT 62.320 47.945 65.075 48.625 ;
        RECT 65.325 48.045 70.835 48.855 ;
        RECT 70.845 48.045 74.515 48.855 ;
        RECT 75.445 48.075 76.815 48.855 ;
        RECT 77.055 48.175 80.955 48.855 ;
        RECT 80.025 47.945 80.955 48.175 ;
        RECT 80.965 48.045 82.795 48.855 ;
        RECT 82.815 47.985 83.245 48.770 ;
        RECT 83.265 47.945 86.740 48.855 ;
        RECT 86.945 48.045 89.695 48.855 ;
        RECT 89.705 48.175 93.605 48.855 ;
        RECT 89.705 47.945 90.635 48.175 ;
        RECT 93.845 48.045 97.515 48.855 ;
        RECT 98.095 48.175 101.560 48.855 ;
        RECT 100.640 47.945 101.560 48.175 ;
        RECT 101.665 48.045 107.175 48.855 ;
        RECT 107.185 48.075 108.555 48.855 ;
        RECT 108.575 47.985 109.005 48.770 ;
        RECT 109.120 48.175 112.585 48.855 ;
        RECT 112.800 48.175 116.265 48.855 ;
        RECT 109.120 47.945 110.040 48.175 ;
        RECT 112.800 47.945 113.720 48.175 ;
        RECT 116.385 48.045 121.895 48.855 ;
        RECT 121.905 48.045 123.735 48.855 ;
        RECT 124.205 48.045 125.575 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 125.770 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 8.735 44.435 ;
        RECT 13.715 44.305 14.645 44.525 ;
        RECT 17.475 44.305 18.395 44.535 ;
        RECT 9.205 43.625 18.395 44.305 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 18.865 44.305 19.795 44.535 ;
        RECT 18.865 43.625 22.765 44.305 ;
        RECT 23.005 43.625 24.375 44.435 ;
        RECT 24.385 43.625 25.755 44.405 ;
        RECT 30.275 44.305 31.205 44.525 ;
        RECT 34.035 44.305 34.955 44.535 ;
        RECT 38.540 44.305 39.460 44.535 ;
        RECT 25.765 43.625 34.955 44.305 ;
        RECT 35.995 43.625 39.460 44.305 ;
        RECT 39.575 43.625 40.925 44.535 ;
        RECT 40.945 43.625 43.695 44.435 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 45.545 44.305 46.475 44.535 ;
        RECT 49.685 44.305 50.615 44.535 ;
        RECT 53.920 44.305 54.840 44.535 ;
        RECT 45.545 43.625 49.445 44.305 ;
        RECT 49.685 43.625 53.585 44.305 ;
        RECT 53.920 43.625 57.385 44.305 ;
        RECT 57.505 43.625 63.015 44.435 ;
        RECT 63.025 43.625 68.535 44.435 ;
        RECT 68.545 43.625 69.915 44.435 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 70.385 43.625 73.135 44.435 ;
        RECT 78.115 44.305 79.045 44.525 ;
        RECT 81.875 44.305 82.795 44.535 ;
        RECT 73.605 43.625 82.795 44.305 ;
        RECT 82.900 44.305 83.820 44.535 ;
        RECT 82.900 43.625 86.365 44.305 ;
        RECT 86.485 43.625 89.960 44.535 ;
        RECT 90.260 44.305 91.180 44.535 ;
        RECT 90.260 43.625 93.725 44.305 ;
        RECT 93.845 43.625 95.675 44.435 ;
        RECT 95.695 43.710 96.125 44.495 ;
        RECT 96.145 43.625 101.655 44.435 ;
        RECT 101.665 43.625 103.495 44.435 ;
        RECT 106.705 44.305 107.635 44.535 ;
        RECT 103.735 43.625 107.635 44.305 ;
        RECT 107.740 44.305 108.660 44.535 ;
        RECT 107.740 43.625 111.205 44.305 ;
        RECT 111.335 43.625 112.685 44.535 ;
        RECT 112.705 43.625 118.215 44.435 ;
        RECT 118.225 43.625 120.975 44.435 ;
        RECT 121.455 43.710 121.885 44.495 ;
        RECT 121.905 43.625 123.735 44.435 ;
        RECT 124.205 43.625 125.575 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.625 ;
        RECT 8.880 43.465 9.000 43.575 ;
        RECT 9.345 43.435 9.515 43.625 ;
        RECT 12.565 43.415 12.735 43.605 ;
        RECT 16.255 43.460 16.415 43.570 ;
        RECT 18.085 43.415 18.255 43.605 ;
        RECT 19.280 43.435 19.450 43.625 ;
        RECT 19.465 43.415 19.635 43.605 ;
        RECT 19.935 43.460 20.095 43.570 ;
        RECT 20.845 43.415 21.015 43.605 ;
        RECT 23.145 43.435 23.315 43.625 ;
        RECT 24.525 43.435 24.695 43.625 ;
        RECT 25.905 43.435 26.075 43.625 ;
        RECT 27.745 43.415 27.915 43.605 ;
        RECT 28.205 43.415 28.375 43.605 ;
        RECT 30.960 43.465 31.080 43.575 ;
        RECT 32.805 43.415 32.975 43.605 ;
        RECT 33.265 43.415 33.435 43.605 ;
        RECT 35.115 43.470 35.275 43.580 ;
        RECT 36.025 43.415 36.195 43.625 ;
        RECT 36.485 43.415 36.655 43.605 ;
        RECT 40.625 43.435 40.795 43.625 ;
        RECT 41.085 43.435 41.255 43.625 ;
        RECT 42.005 43.415 42.175 43.605 ;
        RECT 43.845 43.575 44.015 43.605 ;
        RECT 43.840 43.465 44.015 43.575 ;
        RECT 44.775 43.470 44.935 43.580 ;
        RECT 43.845 43.415 44.015 43.465 ;
        RECT 45.235 43.460 45.395 43.570 ;
        RECT 45.960 43.435 46.130 43.625 ;
        RECT 46.145 43.415 46.315 43.605 ;
        RECT 47.525 43.415 47.695 43.605 ;
        RECT 50.100 43.435 50.270 43.625 ;
        RECT 53.045 43.415 53.215 43.605 ;
        RECT 56.720 43.465 56.840 43.575 ;
        RECT 57.185 43.435 57.355 43.625 ;
        RECT 57.645 43.415 57.815 43.625 ;
        RECT 61.320 43.465 61.440 43.575 ;
        RECT 61.785 43.415 61.955 43.605 ;
        RECT 63.165 43.435 63.335 43.625 ;
        RECT 67.305 43.415 67.475 43.605 ;
        RECT 67.765 43.415 67.935 43.605 ;
        RECT 68.685 43.435 68.855 43.625 ;
        RECT 70.525 43.435 70.695 43.625 ;
        RECT 73.285 43.575 73.455 43.605 ;
        RECT 73.280 43.465 73.455 43.575 ;
        RECT 73.285 43.415 73.455 43.465 ;
        RECT 73.745 43.435 73.915 43.625 ;
        RECT 76.965 43.415 77.135 43.605 ;
        RECT 78.345 43.415 78.515 43.605 ;
        RECT 79.725 43.415 79.895 43.605 ;
        RECT 82.480 43.465 82.600 43.575 ;
        RECT 83.680 43.415 83.850 43.605 ;
        RECT 86.165 43.435 86.335 43.625 ;
        RECT 86.630 43.435 86.800 43.625 ;
        RECT 90.765 43.415 90.935 43.605 ;
        RECT 91.225 43.415 91.395 43.605 ;
        RECT 93.525 43.435 93.695 43.625 ;
        RECT 93.985 43.435 94.155 43.625 ;
        RECT 95.825 43.415 95.995 43.605 ;
        RECT 96.285 43.435 96.455 43.625 ;
        RECT 96.560 43.415 96.730 43.605 ;
        RECT 100.420 43.465 100.540 43.575 ;
        RECT 101.160 43.415 101.330 43.605 ;
        RECT 101.805 43.435 101.975 43.625 ;
        RECT 105.025 43.415 105.195 43.605 ;
        RECT 106.405 43.415 106.575 43.605 ;
        RECT 107.050 43.435 107.220 43.625 ;
        RECT 108.240 43.465 108.360 43.575 ;
        RECT 111.005 43.435 111.175 43.625 ;
        RECT 111.465 43.435 111.635 43.625 ;
        RECT 112.385 43.415 112.555 43.605 ;
        RECT 112.845 43.415 113.015 43.625 ;
        RECT 114.225 43.415 114.395 43.605 ;
        RECT 118.365 43.435 118.535 43.625 ;
        RECT 119.745 43.415 119.915 43.605 ;
        RECT 121.120 43.465 121.240 43.575 ;
        RECT 122.045 43.435 122.215 43.625 ;
        RECT 123.435 43.460 123.595 43.570 ;
        RECT 123.880 43.465 124.000 43.575 ;
        RECT 125.265 43.415 125.435 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 12.415 43.415 ;
        RECT 12.425 42.605 16.095 43.415 ;
        RECT 17.035 42.505 18.385 43.415 ;
        RECT 18.415 42.505 19.765 43.415 ;
        RECT 20.815 42.735 24.280 43.415 ;
        RECT 23.360 42.505 24.280 42.735 ;
        RECT 24.480 42.735 27.945 43.415 ;
        RECT 24.480 42.505 25.400 42.735 ;
        RECT 28.065 42.605 30.815 43.415 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.755 42.505 33.105 43.415 ;
        RECT 33.125 42.605 34.955 43.415 ;
        RECT 34.965 42.635 36.335 43.415 ;
        RECT 36.345 42.605 41.855 43.415 ;
        RECT 41.865 42.605 43.695 43.415 ;
        RECT 43.705 42.635 45.075 43.415 ;
        RECT 46.015 42.505 47.365 43.415 ;
        RECT 47.385 42.605 52.895 43.415 ;
        RECT 52.905 42.605 56.575 43.415 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 57.505 42.605 61.175 43.415 ;
        RECT 61.645 43.185 63.215 43.415 ;
        RECT 65.305 43.375 66.225 43.415 ;
        RECT 65.305 43.185 66.235 43.375 ;
        RECT 61.645 42.825 66.235 43.185 ;
        RECT 61.645 42.735 66.225 42.825 ;
        RECT 63.225 42.505 66.225 42.735 ;
        RECT 66.255 42.505 67.605 43.415 ;
        RECT 67.625 42.605 73.135 43.415 ;
        RECT 73.145 42.605 76.815 43.415 ;
        RECT 76.825 42.605 78.195 43.415 ;
        RECT 78.215 42.505 79.565 43.415 ;
        RECT 79.585 42.605 82.335 43.415 ;
        RECT 82.815 42.545 83.245 43.330 ;
        RECT 83.265 42.735 87.165 43.415 ;
        RECT 87.500 42.735 90.965 43.415 ;
        RECT 83.265 42.505 84.195 42.735 ;
        RECT 87.500 42.505 88.420 42.735 ;
        RECT 91.095 42.505 92.445 43.415 ;
        RECT 92.560 42.735 96.025 43.415 ;
        RECT 96.145 42.735 100.045 43.415 ;
        RECT 100.745 42.735 104.645 43.415 ;
        RECT 92.560 42.505 93.480 42.735 ;
        RECT 96.145 42.505 97.075 42.735 ;
        RECT 100.745 42.505 101.675 42.735 ;
        RECT 104.885 42.635 106.255 43.415 ;
        RECT 106.265 42.605 108.095 43.415 ;
        RECT 108.575 42.545 109.005 43.330 ;
        RECT 109.120 42.735 112.585 43.415 ;
        RECT 109.120 42.505 110.040 42.735 ;
        RECT 112.715 42.505 114.065 43.415 ;
        RECT 114.085 42.605 119.595 43.415 ;
        RECT 119.605 42.605 123.275 43.415 ;
        RECT 124.205 42.605 125.575 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 125.770 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 6.905 38.185 12.415 38.995 ;
        RECT 12.425 38.185 17.935 38.995 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.185 24.375 38.995 ;
        RECT 24.385 38.185 29.895 38.995 ;
        RECT 33.480 38.865 34.400 39.095 ;
        RECT 30.935 38.185 34.400 38.865 ;
        RECT 34.505 38.185 38.175 38.995 ;
        RECT 38.185 38.185 39.555 38.995 ;
        RECT 39.565 38.185 40.935 38.965 ;
        RECT 40.945 38.185 43.695 38.995 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 45.985 38.865 46.905 39.085 ;
        RECT 52.985 38.985 53.905 39.095 ;
        RECT 51.570 38.865 53.905 38.985 ;
        RECT 44.625 38.185 53.905 38.865 ;
        RECT 54.285 38.185 57.955 38.995 ;
        RECT 62.475 38.865 63.405 39.085 ;
        RECT 66.235 38.865 67.155 39.095 ;
        RECT 57.965 38.185 67.155 38.865 ;
        RECT 67.165 38.865 68.510 39.095 ;
        RECT 67.165 38.185 68.995 38.865 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 75.355 38.865 76.285 39.085 ;
        RECT 79.115 38.865 80.035 39.095 ;
        RECT 70.845 38.185 80.035 38.865 ;
        RECT 80.965 38.185 82.335 38.965 ;
        RECT 82.440 38.865 83.360 39.095 ;
        RECT 89.225 38.865 90.155 39.095 ;
        RECT 92.820 38.865 93.740 39.095 ;
        RECT 82.440 38.185 85.905 38.865 ;
        RECT 86.255 38.185 90.155 38.865 ;
        RECT 90.275 38.185 93.740 38.865 ;
        RECT 93.845 38.185 95.215 38.965 ;
        RECT 95.695 38.270 96.125 39.055 ;
        RECT 96.155 38.185 97.505 39.095 ;
        RECT 99.805 38.865 100.725 39.085 ;
        RECT 106.805 38.985 107.725 39.095 ;
        RECT 105.390 38.865 107.725 38.985 ;
        RECT 112.615 38.865 113.545 39.085 ;
        RECT 116.375 38.865 117.295 39.095 ;
        RECT 98.445 38.185 107.725 38.865 ;
        RECT 108.105 38.185 117.295 38.865 ;
        RECT 117.305 38.185 120.975 38.995 ;
        RECT 121.455 38.270 121.885 39.055 ;
        RECT 121.905 38.185 123.735 38.995 ;
        RECT 124.205 38.185 125.575 38.995 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.975 7.215 38.185 ;
        RECT 12.565 37.975 12.735 38.185 ;
        RECT 14.405 37.975 14.575 38.165 ;
        RECT 18.080 38.025 18.200 38.135 ;
        RECT 19.005 37.995 19.175 38.185 ;
        RECT 23.880 37.975 24.050 38.165 ;
        RECT 24.525 37.995 24.695 38.185 ;
        RECT 27.745 37.975 27.915 38.165 ;
        RECT 30.055 38.030 30.215 38.140 ;
        RECT 30.965 37.995 31.135 38.185 ;
        RECT 34.645 37.995 34.815 38.185 ;
        RECT 35.290 37.975 35.460 38.165 ;
        RECT 36.020 38.025 36.140 38.135 ;
        RECT 36.485 37.975 36.655 38.165 ;
        RECT 38.325 37.995 38.495 38.185 ;
        RECT 40.625 37.995 40.795 38.185 ;
        RECT 41.085 37.995 41.255 38.185 ;
        RECT 43.840 38.025 43.960 38.135 ;
        RECT 44.765 37.995 44.935 38.185 ;
        RECT 46.420 37.975 46.590 38.165 ;
        RECT 50.285 37.975 50.455 38.165 ;
        RECT 54.425 37.995 54.595 38.185 ;
        RECT 55.805 37.975 55.975 38.165 ;
        RECT 58.105 37.995 58.275 38.185 ;
        RECT 58.565 37.975 58.735 38.165 ;
        RECT 59.020 38.025 59.140 38.135 ;
        RECT 60.405 37.975 60.575 38.165 ;
        RECT 60.860 38.025 60.980 38.135 ;
        RECT 61.325 37.975 61.495 38.165 ;
        RECT 65.005 37.975 65.175 38.165 ;
        RECT 66.840 38.025 66.960 38.135 ;
        RECT 67.305 37.975 67.475 38.165 ;
        RECT 68.685 37.995 68.855 38.185 ;
        RECT 69.155 38.030 69.315 38.140 ;
        RECT 70.520 38.025 70.640 38.135 ;
        RECT 70.985 37.975 71.155 38.185 ;
        RECT 74.665 37.975 74.835 38.165 ;
        RECT 75.120 38.025 75.240 38.135 ;
        RECT 75.860 37.975 76.030 38.165 ;
        RECT 80.195 38.030 80.355 38.140 ;
        RECT 80.645 37.975 80.815 38.165 ;
        RECT 81.105 38.135 81.275 38.185 ;
        RECT 81.100 38.025 81.275 38.135 ;
        RECT 81.105 37.995 81.275 38.025 ;
        RECT 81.565 37.975 81.735 38.165 ;
        RECT 83.405 37.975 83.575 38.165 ;
        RECT 85.705 37.995 85.875 38.185 ;
        RECT 89.570 37.995 89.740 38.185 ;
        RECT 90.305 37.995 90.475 38.185 ;
        RECT 94.905 37.995 95.075 38.185 ;
        RECT 95.360 38.025 95.480 38.135 ;
        RECT 96.285 37.995 96.455 38.185 ;
        RECT 97.675 38.030 97.835 38.140 ;
        RECT 98.585 37.995 98.755 38.185 ;
        RECT 101.345 37.975 101.515 38.165 ;
        RECT 101.805 37.975 101.975 38.165 ;
        RECT 103.640 38.025 103.760 38.135 ;
        RECT 105.025 37.975 105.195 38.165 ;
        RECT 105.485 37.975 105.655 38.165 ;
        RECT 108.245 38.135 108.415 38.185 ;
        RECT 108.240 38.025 108.415 38.135 ;
        RECT 108.245 37.995 108.415 38.025 ;
        RECT 109.165 37.975 109.335 38.165 ;
        RECT 114.685 37.975 114.855 38.165 ;
        RECT 117.445 37.995 117.615 38.185 ;
        RECT 120.205 37.975 120.375 38.165 ;
        RECT 121.120 38.025 121.240 38.135 ;
        RECT 122.045 37.995 122.215 38.185 ;
        RECT 123.880 38.025 124.000 38.135 ;
        RECT 125.265 37.975 125.435 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.165 12.415 37.975 ;
        RECT 12.425 37.165 14.255 37.975 ;
        RECT 14.265 37.295 23.455 37.975 ;
        RECT 18.775 37.075 19.705 37.295 ;
        RECT 22.535 37.065 23.455 37.295 ;
        RECT 23.465 37.295 27.365 37.975 ;
        RECT 23.465 37.065 24.395 37.295 ;
        RECT 27.605 37.165 31.275 37.975 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.975 37.295 35.875 37.975 ;
        RECT 36.345 37.295 45.625 37.975 ;
        RECT 34.945 37.065 35.875 37.295 ;
        RECT 37.705 37.075 38.625 37.295 ;
        RECT 43.290 37.175 45.625 37.295 ;
        RECT 44.705 37.065 45.625 37.175 ;
        RECT 46.005 37.295 49.905 37.975 ;
        RECT 46.005 37.065 46.935 37.295 ;
        RECT 50.145 37.165 55.655 37.975 ;
        RECT 55.665 37.165 57.035 37.975 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 57.515 37.065 58.865 37.975 ;
        RECT 59.355 37.065 60.705 37.975 ;
        RECT 61.185 37.295 64.855 37.975 ;
        RECT 64.865 37.295 66.695 37.975 ;
        RECT 67.275 37.295 70.740 37.975 ;
        RECT 63.925 37.065 64.855 37.295 ;
        RECT 69.820 37.065 70.740 37.295 ;
        RECT 70.845 37.165 73.595 37.975 ;
        RECT 73.605 37.195 74.975 37.975 ;
        RECT 75.445 37.295 79.345 37.975 ;
        RECT 75.445 37.065 76.375 37.295 ;
        RECT 79.595 37.065 80.945 37.975 ;
        RECT 81.435 37.065 82.785 37.975 ;
        RECT 82.815 37.105 83.245 37.890 ;
        RECT 83.265 37.295 92.455 37.975 ;
        RECT 87.775 37.075 88.705 37.295 ;
        RECT 91.535 37.065 92.455 37.295 ;
        RECT 92.465 37.295 101.655 37.975 ;
        RECT 92.465 37.065 93.385 37.295 ;
        RECT 96.215 37.075 97.145 37.295 ;
        RECT 101.665 37.165 103.495 37.975 ;
        RECT 103.975 37.065 105.325 37.975 ;
        RECT 105.345 37.165 108.095 37.975 ;
        RECT 108.575 37.105 109.005 37.890 ;
        RECT 109.025 37.165 114.535 37.975 ;
        RECT 114.545 37.165 120.055 37.975 ;
        RECT 120.065 37.165 123.735 37.975 ;
        RECT 124.205 37.165 125.575 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 125.770 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 12.415 33.555 ;
        RECT 13.345 32.745 14.715 33.525 ;
        RECT 14.820 33.425 15.740 33.655 ;
        RECT 14.820 32.745 18.285 33.425 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 19.785 33.425 20.715 33.655 ;
        RECT 19.785 32.745 23.685 33.425 ;
        RECT 23.925 32.745 25.295 33.525 ;
        RECT 25.305 32.745 27.135 33.555 ;
        RECT 27.145 33.425 28.065 33.655 ;
        RECT 30.895 33.425 31.825 33.645 ;
        RECT 27.145 32.745 36.335 33.425 ;
        RECT 36.345 32.745 40.015 33.555 ;
        RECT 40.495 32.745 41.845 33.655 ;
        RECT 41.865 32.745 43.695 33.555 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 44.625 32.745 50.135 33.555 ;
        RECT 50.145 32.745 51.975 33.555 ;
        RECT 56.495 33.425 57.425 33.645 ;
        RECT 60.255 33.425 61.175 33.655 ;
        RECT 61.670 33.425 63.015 33.655 ;
        RECT 51.985 32.745 61.175 33.425 ;
        RECT 61.185 32.745 63.015 33.425 ;
        RECT 63.025 32.745 68.535 33.555 ;
        RECT 68.545 32.745 69.915 33.555 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 70.385 32.745 75.895 33.555 ;
        RECT 75.905 32.745 81.415 33.555 ;
        RECT 81.425 32.745 84.175 33.555 ;
        RECT 88.695 33.425 89.625 33.645 ;
        RECT 92.455 33.425 93.375 33.655 ;
        RECT 84.185 32.745 93.375 33.425 ;
        RECT 93.845 32.745 95.215 33.525 ;
        RECT 95.695 32.830 96.125 33.615 ;
        RECT 97.065 32.745 98.435 33.525 ;
        RECT 98.445 32.745 103.955 33.555 ;
        RECT 103.965 32.745 109.475 33.555 ;
        RECT 109.485 32.745 114.995 33.555 ;
        RECT 115.005 32.745 120.515 33.555 ;
        RECT 121.455 32.830 121.885 33.615 ;
        RECT 121.905 32.745 123.735 33.555 ;
        RECT 124.205 32.745 125.575 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.535 7.215 32.745 ;
        RECT 12.565 32.535 12.735 32.725 ;
        RECT 13.485 32.555 13.655 32.745 ;
        RECT 16.255 32.580 16.415 32.690 ;
        RECT 18.085 32.535 18.255 32.745 ;
        RECT 18.545 32.535 18.715 32.725 ;
        RECT 19.015 32.590 19.175 32.700 ;
        RECT 20.200 32.555 20.370 32.745 ;
        RECT 24.985 32.555 25.155 32.745 ;
        RECT 25.445 32.555 25.615 32.745 ;
        RECT 30.965 32.535 31.135 32.725 ;
        RECT 32.805 32.535 32.975 32.725 ;
        RECT 33.265 32.535 33.435 32.725 ;
        RECT 34.645 32.535 34.815 32.725 ;
        RECT 36.025 32.555 36.195 32.745 ;
        RECT 36.485 32.555 36.655 32.745 ;
        RECT 40.165 32.695 40.335 32.725 ;
        RECT 40.160 32.585 40.335 32.695 ;
        RECT 40.165 32.535 40.335 32.585 ;
        RECT 40.625 32.555 40.795 32.745 ;
        RECT 42.005 32.555 42.175 32.745 ;
        RECT 43.840 32.585 43.960 32.695 ;
        RECT 44.765 32.555 44.935 32.745 ;
        RECT 45.685 32.535 45.855 32.725 ;
        RECT 50.285 32.555 50.455 32.745 ;
        RECT 51.205 32.535 51.375 32.725 ;
        RECT 52.125 32.555 52.295 32.745 ;
        RECT 53.040 32.585 53.160 32.695 ;
        RECT 53.505 32.535 53.675 32.725 ;
        RECT 54.880 32.585 55.000 32.695 ;
        RECT 56.265 32.535 56.435 32.725 ;
        RECT 56.720 32.585 56.840 32.695 ;
        RECT 59.485 32.535 59.655 32.725 ;
        RECT 59.955 32.580 60.115 32.690 ;
        RECT 60.865 32.535 61.035 32.725 ;
        RECT 61.325 32.555 61.495 32.745 ;
        RECT 63.165 32.725 63.335 32.745 ;
        RECT 63.165 32.555 63.340 32.725 ;
        RECT 63.170 32.535 63.340 32.555 ;
        RECT 66.385 32.535 66.555 32.725 ;
        RECT 68.685 32.555 68.855 32.745 ;
        RECT 70.525 32.555 70.695 32.745 ;
        RECT 72.365 32.535 72.535 32.725 ;
        RECT 72.825 32.535 72.995 32.725 ;
        RECT 74.205 32.535 74.375 32.725 ;
        RECT 76.045 32.555 76.215 32.745 ;
        RECT 79.725 32.535 79.895 32.725 ;
        RECT 81.565 32.555 81.735 32.745 ;
        RECT 82.480 32.585 82.600 32.695 ;
        RECT 83.405 32.535 83.575 32.725 ;
        RECT 84.325 32.555 84.495 32.745 ;
        RECT 88.925 32.535 89.095 32.725 ;
        RECT 93.520 32.585 93.640 32.695 ;
        RECT 93.985 32.555 94.155 32.745 ;
        RECT 94.445 32.535 94.615 32.725 ;
        RECT 95.360 32.585 95.480 32.695 ;
        RECT 96.295 32.590 96.455 32.700 ;
        RECT 97.205 32.555 97.375 32.745 ;
        RECT 98.585 32.555 98.755 32.745 ;
        RECT 99.965 32.535 100.135 32.725 ;
        RECT 104.105 32.555 104.275 32.745 ;
        RECT 105.485 32.535 105.655 32.725 ;
        RECT 108.240 32.585 108.360 32.695 ;
        RECT 109.165 32.535 109.335 32.725 ;
        RECT 109.625 32.555 109.795 32.745 ;
        RECT 114.685 32.535 114.855 32.725 ;
        RECT 115.145 32.555 115.315 32.745 ;
        RECT 120.205 32.535 120.375 32.725 ;
        RECT 120.675 32.590 120.835 32.700 ;
        RECT 122.045 32.555 122.215 32.745 ;
        RECT 123.880 32.585 124.000 32.695 ;
        RECT 125.265 32.535 125.435 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.725 12.415 32.535 ;
        RECT 12.425 31.725 16.095 32.535 ;
        RECT 17.035 31.625 18.385 32.535 ;
        RECT 18.405 31.855 27.595 32.535 ;
        RECT 22.915 31.635 23.845 31.855 ;
        RECT 26.675 31.625 27.595 31.855 ;
        RECT 27.700 31.855 31.165 32.535 ;
        RECT 27.700 31.625 28.620 31.855 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.755 31.625 33.105 32.535 ;
        RECT 33.125 31.755 34.495 32.535 ;
        RECT 34.505 31.725 40.015 32.535 ;
        RECT 40.025 31.725 45.535 32.535 ;
        RECT 45.545 31.725 51.055 32.535 ;
        RECT 51.065 31.725 52.895 32.535 ;
        RECT 53.375 31.625 54.725 32.535 ;
        RECT 55.205 31.755 56.575 32.535 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 57.505 31.855 59.795 32.535 ;
        RECT 60.725 31.855 63.015 32.535 ;
        RECT 57.505 31.625 58.425 31.855 ;
        RECT 62.095 31.625 63.015 31.855 ;
        RECT 63.025 31.625 65.945 32.535 ;
        RECT 66.245 31.725 68.995 32.535 ;
        RECT 69.100 31.855 72.565 32.535 ;
        RECT 69.100 31.625 70.020 31.855 ;
        RECT 72.695 31.625 74.045 32.535 ;
        RECT 74.065 31.725 79.575 32.535 ;
        RECT 79.585 31.725 82.335 32.535 ;
        RECT 82.815 31.665 83.245 32.450 ;
        RECT 83.265 31.725 88.775 32.535 ;
        RECT 88.785 31.725 94.295 32.535 ;
        RECT 94.305 31.725 99.815 32.535 ;
        RECT 99.825 31.725 105.335 32.535 ;
        RECT 105.345 31.725 108.095 32.535 ;
        RECT 108.575 31.665 109.005 32.450 ;
        RECT 109.025 31.725 114.535 32.535 ;
        RECT 114.545 31.725 120.055 32.535 ;
        RECT 120.065 31.725 123.735 32.535 ;
        RECT 124.205 31.725 125.575 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 125.770 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 12.415 28.115 ;
        RECT 12.425 27.305 17.935 28.115 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.865 27.305 24.375 28.115 ;
        RECT 24.385 27.305 27.135 28.115 ;
        RECT 27.615 27.305 28.965 28.215 ;
        RECT 28.985 27.305 34.495 28.115 ;
        RECT 34.505 27.305 40.015 28.115 ;
        RECT 40.025 27.305 43.695 28.115 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.625 27.305 48.295 28.115 ;
        RECT 53.735 27.985 54.665 28.205 ;
        RECT 57.495 27.985 58.415 28.215 ;
        RECT 49.225 27.305 58.415 27.985 ;
        RECT 58.425 27.305 59.775 28.215 ;
        RECT 60.265 27.305 62.555 28.215 ;
        RECT 62.565 28.015 63.510 28.215 ;
        RECT 64.845 28.015 65.775 28.215 ;
        RECT 62.565 27.535 65.775 28.015 ;
        RECT 62.565 27.335 65.635 27.535 ;
        RECT 62.565 27.305 63.510 27.335 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.095 7.215 27.305 ;
        RECT 12.565 27.095 12.735 27.305 ;
        RECT 18.085 27.255 18.255 27.285 ;
        RECT 18.080 27.145 18.255 27.255 ;
        RECT 18.085 27.095 18.255 27.145 ;
        RECT 19.005 27.115 19.175 27.305 ;
        RECT 23.605 27.095 23.775 27.285 ;
        RECT 24.525 27.115 24.695 27.305 ;
        RECT 27.280 27.145 27.400 27.255 ;
        RECT 28.665 27.115 28.835 27.305 ;
        RECT 29.125 27.095 29.295 27.305 ;
        RECT 30.960 27.145 31.080 27.255 ;
        RECT 31.885 27.095 32.055 27.285 ;
        RECT 34.645 27.115 34.815 27.305 ;
        RECT 37.405 27.095 37.575 27.285 ;
        RECT 40.165 27.115 40.335 27.305 ;
        RECT 42.925 27.095 43.095 27.285 ;
        RECT 43.840 27.145 43.960 27.255 ;
        RECT 44.765 27.115 44.935 27.305 ;
        RECT 48.445 27.095 48.615 27.285 ;
        RECT 49.365 27.115 49.535 27.305 ;
        RECT 52.120 27.145 52.240 27.255 ;
        RECT 55.345 27.095 55.515 27.285 ;
        RECT 55.805 27.095 55.975 27.285 ;
        RECT 57.655 27.140 57.815 27.250 ;
        RECT 59.490 27.115 59.660 27.305 ;
        RECT 59.940 27.145 60.060 27.255 ;
        RECT 60.405 27.115 60.575 27.285 ;
        RECT 60.860 27.145 60.980 27.255 ;
        RECT 62.240 27.115 62.410 27.305 ;
        RECT 60.405 27.095 60.570 27.115 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 6.905 26.285 12.415 27.095 ;
        RECT 12.425 26.285 17.935 27.095 ;
        RECT 17.945 26.285 23.455 27.095 ;
        RECT 23.465 26.285 28.975 27.095 ;
        RECT 28.985 26.285 30.815 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.745 26.285 37.255 27.095 ;
        RECT 37.265 26.285 42.775 27.095 ;
        RECT 42.785 26.285 48.295 27.095 ;
        RECT 48.305 26.285 51.975 27.095 ;
        RECT 52.445 26.185 55.555 27.095 ;
        RECT 55.665 26.285 57.035 27.095 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 58.735 26.415 60.570 27.095 ;
        RECT 61.185 27.065 62.130 27.095 ;
        RECT 64.085 27.065 64.255 27.285 ;
        RECT 64.545 27.095 64.715 27.285 ;
        RECT 65.465 27.115 65.635 27.335 ;
        RECT 65.885 27.305 68.995 28.215 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 70.425 27.985 71.765 28.215 ;
        RECT 74.595 27.985 75.525 28.205 ;
        RECT 70.425 27.305 80.035 27.985 ;
        RECT 80.045 27.305 85.555 28.115 ;
        RECT 85.565 27.305 91.075 28.115 ;
        RECT 91.085 27.305 94.755 28.115 ;
        RECT 95.695 27.390 96.125 28.175 ;
        RECT 96.145 27.305 101.655 28.115 ;
        RECT 101.665 27.305 107.175 28.115 ;
        RECT 107.185 27.305 112.695 28.115 ;
        RECT 112.705 27.305 118.215 28.115 ;
        RECT 118.225 27.305 120.975 28.115 ;
        RECT 121.455 27.390 121.885 28.175 ;
        RECT 121.905 27.305 123.735 28.115 ;
        RECT 124.205 27.305 125.575 28.115 ;
        RECT 65.925 27.115 66.095 27.305 ;
        RECT 69.155 27.150 69.315 27.260 ;
        RECT 75.125 27.095 75.295 27.285 ;
        RECT 79.725 27.115 79.895 27.305 ;
        RECT 80.185 27.115 80.355 27.305 ;
        RECT 80.645 27.095 80.815 27.285 ;
        RECT 82.480 27.145 82.600 27.255 ;
        RECT 83.405 27.095 83.575 27.285 ;
        RECT 85.705 27.115 85.875 27.305 ;
        RECT 88.925 27.095 89.095 27.285 ;
        RECT 91.225 27.115 91.395 27.305 ;
        RECT 94.445 27.095 94.615 27.285 ;
        RECT 94.915 27.150 95.075 27.260 ;
        RECT 96.285 27.115 96.455 27.305 ;
        RECT 99.965 27.095 100.135 27.285 ;
        RECT 101.805 27.115 101.975 27.305 ;
        RECT 105.485 27.095 105.655 27.285 ;
        RECT 107.325 27.115 107.495 27.305 ;
        RECT 108.240 27.145 108.360 27.255 ;
        RECT 109.165 27.095 109.335 27.285 ;
        RECT 112.845 27.115 113.015 27.305 ;
        RECT 114.685 27.095 114.855 27.285 ;
        RECT 118.365 27.115 118.535 27.305 ;
        RECT 120.205 27.095 120.375 27.285 ;
        RECT 121.120 27.145 121.240 27.255 ;
        RECT 122.045 27.115 122.215 27.305 ;
        RECT 123.880 27.145 124.000 27.255 ;
        RECT 125.265 27.095 125.435 27.305 ;
        RECT 61.185 26.865 64.255 27.065 ;
        RECT 58.735 26.185 59.665 26.415 ;
        RECT 61.185 26.385 64.395 26.865 ;
        RECT 64.405 26.415 74.775 27.095 ;
        RECT 61.185 26.185 62.130 26.385 ;
        RECT 63.465 26.185 64.395 26.385 ;
        RECT 68.915 26.195 69.845 26.415 ;
        RECT 72.565 26.185 74.775 26.415 ;
        RECT 74.985 26.285 80.495 27.095 ;
        RECT 80.505 26.285 82.335 27.095 ;
        RECT 82.815 26.225 83.245 27.010 ;
        RECT 83.265 26.285 88.775 27.095 ;
        RECT 88.785 26.285 94.295 27.095 ;
        RECT 94.305 26.285 99.815 27.095 ;
        RECT 99.825 26.285 105.335 27.095 ;
        RECT 105.345 26.285 108.095 27.095 ;
        RECT 108.575 26.225 109.005 27.010 ;
        RECT 109.025 26.285 114.535 27.095 ;
        RECT 114.545 26.285 120.055 27.095 ;
        RECT 120.065 26.285 123.735 27.095 ;
        RECT 124.205 26.285 125.575 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 125.770 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 21.865 12.415 22.675 ;
        RECT 12.425 21.865 17.935 22.675 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 18.865 21.865 24.375 22.675 ;
        RECT 24.385 21.865 29.895 22.675 ;
        RECT 29.905 21.865 35.415 22.675 ;
        RECT 35.425 21.865 40.935 22.675 ;
        RECT 40.945 21.865 43.695 22.675 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 50.135 22.675 ;
        RECT 50.145 21.865 55.655 22.675 ;
        RECT 55.665 21.865 61.175 22.675 ;
        RECT 61.185 21.865 66.695 22.675 ;
        RECT 67.165 21.865 68.535 22.645 ;
        RECT 68.545 21.865 69.915 22.675 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.395 21.865 71.745 22.775 ;
        RECT 71.765 21.865 77.275 22.675 ;
        RECT 77.285 21.865 82.795 22.675 ;
        RECT 82.805 21.865 88.315 22.675 ;
        RECT 88.325 21.865 93.835 22.675 ;
        RECT 93.845 21.865 95.675 22.675 ;
        RECT 95.695 21.950 96.125 22.735 ;
        RECT 96.145 21.865 101.655 22.675 ;
        RECT 101.665 21.865 107.175 22.675 ;
        RECT 107.185 21.865 112.695 22.675 ;
        RECT 112.705 21.865 118.215 22.675 ;
        RECT 118.225 21.865 120.975 22.675 ;
        RECT 121.455 21.950 121.885 22.735 ;
        RECT 121.905 21.865 123.735 22.675 ;
        RECT 124.205 21.865 125.575 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.655 7.215 21.865 ;
        RECT 12.565 21.655 12.735 21.865 ;
        RECT 18.085 21.815 18.255 21.845 ;
        RECT 18.080 21.705 18.255 21.815 ;
        RECT 18.085 21.655 18.255 21.705 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 23.605 21.655 23.775 21.845 ;
        RECT 24.525 21.675 24.695 21.865 ;
        RECT 29.125 21.655 29.295 21.845 ;
        RECT 30.045 21.675 30.215 21.865 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 35.565 21.675 35.735 21.865 ;
        RECT 37.405 21.655 37.575 21.845 ;
        RECT 41.085 21.675 41.255 21.865 ;
        RECT 42.925 21.655 43.095 21.845 ;
        RECT 43.840 21.705 43.960 21.815 ;
        RECT 44.765 21.675 44.935 21.865 ;
        RECT 48.445 21.655 48.615 21.845 ;
        RECT 50.285 21.675 50.455 21.865 ;
        RECT 53.965 21.655 54.135 21.845 ;
        RECT 55.805 21.675 55.975 21.865 ;
        RECT 56.720 21.705 56.840 21.815 ;
        RECT 57.645 21.655 57.815 21.845 ;
        RECT 61.325 21.675 61.495 21.865 ;
        RECT 63.165 21.655 63.335 21.845 ;
        RECT 66.840 21.705 66.960 21.815 ;
        RECT 68.225 21.675 68.395 21.865 ;
        RECT 68.685 21.655 68.855 21.865 ;
        RECT 71.445 21.675 71.615 21.865 ;
        RECT 71.905 21.675 72.075 21.865 ;
        RECT 74.205 21.655 74.375 21.845 ;
        RECT 77.425 21.675 77.595 21.865 ;
        RECT 79.725 21.655 79.895 21.845 ;
        RECT 82.480 21.705 82.600 21.815 ;
        RECT 82.945 21.675 83.115 21.865 ;
        RECT 83.405 21.655 83.575 21.845 ;
        RECT 88.465 21.675 88.635 21.865 ;
        RECT 88.925 21.655 89.095 21.845 ;
        RECT 93.985 21.675 94.155 21.865 ;
        RECT 94.445 21.655 94.615 21.845 ;
        RECT 96.285 21.675 96.455 21.865 ;
        RECT 99.965 21.655 100.135 21.845 ;
        RECT 101.805 21.675 101.975 21.865 ;
        RECT 105.485 21.655 105.655 21.845 ;
        RECT 107.325 21.675 107.495 21.865 ;
        RECT 108.240 21.705 108.360 21.815 ;
        RECT 109.165 21.655 109.335 21.845 ;
        RECT 112.845 21.675 113.015 21.865 ;
        RECT 114.685 21.655 114.855 21.845 ;
        RECT 118.365 21.675 118.535 21.865 ;
        RECT 120.205 21.655 120.375 21.845 ;
        RECT 121.120 21.705 121.240 21.815 ;
        RECT 122.045 21.675 122.215 21.865 ;
        RECT 123.880 21.705 124.000 21.815 ;
        RECT 125.265 21.655 125.435 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.845 12.415 21.655 ;
        RECT 12.425 20.845 17.935 21.655 ;
        RECT 17.945 20.845 23.455 21.655 ;
        RECT 23.465 20.845 28.975 21.655 ;
        RECT 28.985 20.845 30.815 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.265 20.845 42.775 21.655 ;
        RECT 42.785 20.845 48.295 21.655 ;
        RECT 48.305 20.845 53.815 21.655 ;
        RECT 53.825 20.845 56.575 21.655 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.505 20.845 63.015 21.655 ;
        RECT 63.025 20.845 68.535 21.655 ;
        RECT 68.545 20.845 74.055 21.655 ;
        RECT 74.065 20.845 79.575 21.655 ;
        RECT 79.585 20.845 82.335 21.655 ;
        RECT 82.815 20.785 83.245 21.570 ;
        RECT 83.265 20.845 88.775 21.655 ;
        RECT 88.785 20.845 94.295 21.655 ;
        RECT 94.305 20.845 99.815 21.655 ;
        RECT 99.825 20.845 105.335 21.655 ;
        RECT 105.345 20.845 108.095 21.655 ;
        RECT 108.575 20.785 109.005 21.570 ;
        RECT 109.025 20.845 114.535 21.655 ;
        RECT 114.545 20.845 120.055 21.655 ;
        RECT 120.065 20.845 123.735 21.655 ;
        RECT 124.205 20.845 125.575 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 125.770 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 12.415 17.235 ;
        RECT 12.425 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 24.375 17.235 ;
        RECT 24.385 16.425 29.895 17.235 ;
        RECT 29.905 16.425 35.415 17.235 ;
        RECT 35.425 16.425 40.935 17.235 ;
        RECT 40.945 16.425 43.695 17.235 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 44.625 16.425 50.135 17.235 ;
        RECT 50.145 16.425 55.655 17.235 ;
        RECT 55.665 16.425 61.175 17.235 ;
        RECT 61.185 16.425 66.695 17.235 ;
        RECT 66.705 16.425 69.455 17.235 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 70.385 16.425 75.895 17.235 ;
        RECT 75.905 16.425 81.415 17.235 ;
        RECT 81.425 16.425 86.935 17.235 ;
        RECT 86.945 16.425 92.455 17.235 ;
        RECT 92.465 16.425 95.215 17.235 ;
        RECT 95.695 16.510 96.125 17.295 ;
        RECT 96.145 16.425 101.655 17.235 ;
        RECT 101.665 16.425 107.175 17.235 ;
        RECT 107.185 16.425 112.695 17.235 ;
        RECT 112.705 16.425 118.215 17.235 ;
        RECT 118.225 16.425 120.975 17.235 ;
        RECT 121.455 16.510 121.885 17.295 ;
        RECT 121.905 16.425 123.735 17.235 ;
        RECT 124.205 16.425 125.575 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 12.565 16.215 12.735 16.425 ;
        RECT 18.085 16.375 18.255 16.405 ;
        RECT 18.080 16.265 18.255 16.375 ;
        RECT 18.085 16.215 18.255 16.265 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.605 16.215 23.775 16.405 ;
        RECT 24.525 16.235 24.695 16.425 ;
        RECT 29.125 16.215 29.295 16.405 ;
        RECT 30.045 16.235 30.215 16.425 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 35.565 16.235 35.735 16.425 ;
        RECT 37.405 16.215 37.575 16.405 ;
        RECT 41.085 16.235 41.255 16.425 ;
        RECT 42.925 16.215 43.095 16.405 ;
        RECT 43.840 16.265 43.960 16.375 ;
        RECT 44.765 16.235 44.935 16.425 ;
        RECT 48.445 16.215 48.615 16.405 ;
        RECT 50.285 16.235 50.455 16.425 ;
        RECT 53.965 16.215 54.135 16.405 ;
        RECT 55.805 16.235 55.975 16.425 ;
        RECT 56.720 16.265 56.840 16.375 ;
        RECT 57.645 16.215 57.815 16.405 ;
        RECT 61.325 16.235 61.495 16.425 ;
        RECT 63.165 16.215 63.335 16.405 ;
        RECT 66.845 16.235 67.015 16.425 ;
        RECT 68.685 16.215 68.855 16.405 ;
        RECT 69.600 16.265 69.720 16.375 ;
        RECT 70.525 16.235 70.695 16.425 ;
        RECT 74.205 16.215 74.375 16.405 ;
        RECT 76.045 16.235 76.215 16.425 ;
        RECT 79.725 16.215 79.895 16.405 ;
        RECT 81.565 16.235 81.735 16.425 ;
        RECT 82.480 16.265 82.600 16.375 ;
        RECT 83.405 16.215 83.575 16.405 ;
        RECT 87.085 16.235 87.255 16.425 ;
        RECT 88.925 16.215 89.095 16.405 ;
        RECT 92.605 16.235 92.775 16.425 ;
        RECT 94.445 16.215 94.615 16.405 ;
        RECT 95.360 16.265 95.480 16.375 ;
        RECT 96.285 16.235 96.455 16.425 ;
        RECT 99.965 16.215 100.135 16.405 ;
        RECT 101.805 16.235 101.975 16.425 ;
        RECT 105.485 16.215 105.655 16.405 ;
        RECT 107.325 16.235 107.495 16.425 ;
        RECT 108.240 16.265 108.360 16.375 ;
        RECT 109.165 16.215 109.335 16.405 ;
        RECT 112.845 16.235 113.015 16.425 ;
        RECT 114.685 16.215 114.855 16.405 ;
        RECT 118.365 16.235 118.535 16.425 ;
        RECT 120.205 16.215 120.375 16.405 ;
        RECT 121.120 16.265 121.240 16.375 ;
        RECT 122.045 16.235 122.215 16.425 ;
        RECT 123.880 16.265 124.000 16.375 ;
        RECT 125.265 16.215 125.435 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 23.455 16.215 ;
        RECT 23.465 15.405 28.975 16.215 ;
        RECT 28.985 15.405 30.815 16.215 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.745 15.405 37.255 16.215 ;
        RECT 37.265 15.405 42.775 16.215 ;
        RECT 42.785 15.405 48.295 16.215 ;
        RECT 48.305 15.405 53.815 16.215 ;
        RECT 53.825 15.405 56.575 16.215 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.405 63.015 16.215 ;
        RECT 63.025 15.405 68.535 16.215 ;
        RECT 68.545 15.405 74.055 16.215 ;
        RECT 74.065 15.405 79.575 16.215 ;
        RECT 79.585 15.405 82.335 16.215 ;
        RECT 82.815 15.345 83.245 16.130 ;
        RECT 83.265 15.405 88.775 16.215 ;
        RECT 88.785 15.405 94.295 16.215 ;
        RECT 94.305 15.405 99.815 16.215 ;
        RECT 99.825 15.405 105.335 16.215 ;
        RECT 105.345 15.405 108.095 16.215 ;
        RECT 108.575 15.345 109.005 16.130 ;
        RECT 109.025 15.405 114.535 16.215 ;
        RECT 114.545 15.405 120.055 16.215 ;
        RECT 120.065 15.405 123.735 16.215 ;
        RECT 124.205 15.405 125.575 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 125.770 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 12.425 10.985 17.935 11.795 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 18.865 10.985 24.375 11.795 ;
        RECT 24.385 10.985 29.895 11.795 ;
        RECT 29.905 10.985 31.275 11.795 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 31.745 10.985 37.255 11.795 ;
        RECT 37.265 10.985 42.775 11.795 ;
        RECT 42.785 10.985 44.155 11.795 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 44.625 10.985 50.135 11.795 ;
        RECT 50.145 10.985 55.655 11.795 ;
        RECT 55.665 10.985 57.035 11.795 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 57.505 10.985 63.015 11.795 ;
        RECT 63.025 10.985 68.535 11.795 ;
        RECT 68.545 10.985 69.915 11.795 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 70.385 10.985 75.895 11.795 ;
        RECT 75.905 10.985 81.415 11.795 ;
        RECT 81.425 10.985 82.795 11.795 ;
        RECT 82.815 11.070 83.245 11.855 ;
        RECT 83.265 10.985 88.775 11.795 ;
        RECT 88.785 10.985 94.295 11.795 ;
        RECT 94.305 10.985 95.675 11.795 ;
        RECT 95.695 11.070 96.125 11.855 ;
        RECT 96.145 10.985 101.655 11.795 ;
        RECT 101.665 10.985 107.175 11.795 ;
        RECT 107.185 10.985 108.555 11.795 ;
        RECT 108.575 11.070 109.005 11.855 ;
        RECT 109.025 10.985 114.535 11.795 ;
        RECT 114.545 10.985 120.055 11.795 ;
        RECT 120.065 10.985 121.435 11.795 ;
        RECT 121.455 11.070 121.885 11.855 ;
        RECT 121.905 10.985 123.735 11.795 ;
        RECT 124.205 10.985 125.575 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.565 10.795 12.735 10.985 ;
        RECT 18.080 10.825 18.200 10.935 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 31.885 10.795 32.055 10.985 ;
        RECT 37.405 10.795 37.575 10.985 ;
        RECT 42.925 10.795 43.095 10.985 ;
        RECT 44.765 10.795 44.935 10.985 ;
        RECT 50.285 10.795 50.455 10.985 ;
        RECT 55.805 10.795 55.975 10.985 ;
        RECT 57.645 10.795 57.815 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 68.685 10.795 68.855 10.985 ;
        RECT 70.525 10.795 70.695 10.985 ;
        RECT 76.045 10.795 76.215 10.985 ;
        RECT 81.565 10.795 81.735 10.985 ;
        RECT 83.405 10.795 83.575 10.985 ;
        RECT 88.925 10.795 89.095 10.985 ;
        RECT 94.445 10.795 94.615 10.985 ;
        RECT 96.285 10.795 96.455 10.985 ;
        RECT 101.805 10.795 101.975 10.985 ;
        RECT 107.325 10.795 107.495 10.985 ;
        RECT 109.165 10.795 109.335 10.985 ;
        RECT 114.685 10.795 114.855 10.985 ;
        RECT 120.205 10.795 120.375 10.985 ;
        RECT 122.045 10.795 122.215 10.985 ;
        RECT 123.880 10.825 124.000 10.935 ;
        RECT 125.265 10.795 125.435 10.985 ;
      LAYER li1 ;
        RECT 5.520 130.475 125.580 130.645 ;
        RECT 5.605 129.725 6.815 130.475 ;
        RECT 6.985 129.930 12.330 130.475 ;
        RECT 5.605 129.185 6.125 129.725 ;
        RECT 6.295 129.015 6.815 129.555 ;
        RECT 8.570 129.100 8.910 129.930 ;
        RECT 13.025 129.655 13.235 130.475 ;
        RECT 13.405 129.675 13.735 130.305 ;
        RECT 5.605 127.925 6.815 129.015 ;
        RECT 10.390 128.360 10.740 129.610 ;
        RECT 13.405 129.075 13.655 129.675 ;
        RECT 13.905 129.655 14.135 130.475 ;
        RECT 14.345 129.705 17.855 130.475 ;
        RECT 18.485 129.750 18.775 130.475 ;
        RECT 18.945 129.930 24.290 130.475 ;
        RECT 24.465 129.930 29.810 130.475 ;
        RECT 13.825 129.235 14.155 129.485 ;
        RECT 14.345 129.185 15.995 129.705 ;
        RECT 6.985 127.925 12.330 128.360 ;
        RECT 13.025 127.925 13.235 129.065 ;
        RECT 13.405 128.095 13.735 129.075 ;
        RECT 13.905 127.925 14.135 129.065 ;
        RECT 16.165 129.015 17.855 129.535 ;
        RECT 20.530 129.100 20.870 129.930 ;
        RECT 14.345 127.925 17.855 129.015 ;
        RECT 18.485 127.925 18.775 129.090 ;
        RECT 22.350 128.360 22.700 129.610 ;
        RECT 26.050 129.100 26.390 129.930 ;
        RECT 29.985 129.725 31.195 130.475 ;
        RECT 31.365 129.750 31.655 130.475 ;
        RECT 31.830 129.925 32.085 130.215 ;
        RECT 32.255 130.095 32.585 130.475 ;
        RECT 31.830 129.755 32.580 129.925 ;
        RECT 27.870 128.360 28.220 129.610 ;
        RECT 29.985 129.185 30.505 129.725 ;
        RECT 30.675 129.015 31.195 129.555 ;
        RECT 18.945 127.925 24.290 128.360 ;
        RECT 24.465 127.925 29.810 128.360 ;
        RECT 29.985 127.925 31.195 129.015 ;
        RECT 31.365 127.925 31.655 129.090 ;
        RECT 31.830 128.935 32.180 129.585 ;
        RECT 32.350 128.765 32.580 129.755 ;
        RECT 31.830 128.595 32.580 128.765 ;
        RECT 31.830 128.095 32.085 128.595 ;
        RECT 32.255 127.925 32.585 128.425 ;
        RECT 32.755 128.095 32.925 130.215 ;
        RECT 33.285 130.115 33.615 130.475 ;
        RECT 33.785 130.085 34.280 130.255 ;
        RECT 34.485 130.085 35.340 130.255 ;
        RECT 33.155 128.895 33.615 129.945 ;
        RECT 33.095 128.110 33.420 128.895 ;
        RECT 33.785 128.725 33.955 130.085 ;
        RECT 34.125 129.175 34.475 129.795 ;
        RECT 34.645 129.575 35.000 129.795 ;
        RECT 34.645 128.985 34.815 129.575 ;
        RECT 35.170 129.375 35.340 130.085 ;
        RECT 36.215 130.015 36.545 130.475 ;
        RECT 36.755 130.115 37.105 130.285 ;
        RECT 35.545 129.545 36.335 129.795 ;
        RECT 36.755 129.725 37.015 130.115 ;
        RECT 37.325 130.025 38.275 130.305 ;
        RECT 38.445 130.035 38.635 130.475 ;
        RECT 38.805 130.095 39.875 130.265 ;
        RECT 36.505 129.375 36.675 129.555 ;
        RECT 33.785 128.555 34.180 128.725 ;
        RECT 34.350 128.595 34.815 128.985 ;
        RECT 34.985 129.205 36.675 129.375 ;
        RECT 34.010 128.425 34.180 128.555 ;
        RECT 34.985 128.425 35.155 129.205 ;
        RECT 36.845 129.035 37.015 129.725 ;
        RECT 35.515 128.865 37.015 129.035 ;
        RECT 37.205 129.065 37.415 129.855 ;
        RECT 37.585 129.235 37.935 129.855 ;
        RECT 38.105 129.245 38.275 130.025 ;
        RECT 38.805 129.865 38.975 130.095 ;
        RECT 38.445 129.695 38.975 129.865 ;
        RECT 38.445 129.415 38.665 129.695 ;
        RECT 39.145 129.525 39.385 129.925 ;
        RECT 38.105 129.075 38.510 129.245 ;
        RECT 38.845 129.155 39.385 129.525 ;
        RECT 39.555 129.740 39.875 130.095 ;
        RECT 39.555 129.485 39.880 129.740 ;
        RECT 40.075 129.665 40.245 130.475 ;
        RECT 40.415 129.825 40.745 130.305 ;
        RECT 40.915 130.005 41.085 130.475 ;
        RECT 41.255 129.825 41.585 130.305 ;
        RECT 41.755 130.005 41.925 130.475 ;
        RECT 40.415 129.655 42.180 129.825 ;
        RECT 39.555 129.275 41.585 129.485 ;
        RECT 39.555 129.265 39.900 129.275 ;
        RECT 37.205 128.905 37.880 129.065 ;
        RECT 38.340 128.985 38.510 129.075 ;
        RECT 37.205 128.895 38.170 128.905 ;
        RECT 36.845 128.725 37.015 128.865 ;
        RECT 33.590 127.925 33.840 128.385 ;
        RECT 34.010 128.095 34.260 128.425 ;
        RECT 34.475 128.095 35.155 128.425 ;
        RECT 35.325 128.525 36.400 128.695 ;
        RECT 36.845 128.555 37.405 128.725 ;
        RECT 37.710 128.605 38.170 128.895 ;
        RECT 38.340 128.815 39.560 128.985 ;
        RECT 35.325 128.185 35.495 128.525 ;
        RECT 35.730 127.925 36.060 128.355 ;
        RECT 36.230 128.185 36.400 128.525 ;
        RECT 36.695 127.925 37.065 128.385 ;
        RECT 37.235 128.095 37.405 128.555 ;
        RECT 38.340 128.435 38.510 128.815 ;
        RECT 39.730 128.645 39.900 129.265 ;
        RECT 41.770 129.105 42.180 129.655 ;
        RECT 42.405 129.705 44.075 130.475 ;
        RECT 44.245 129.750 44.535 130.475 ;
        RECT 44.705 129.930 50.050 130.475 ;
        RECT 50.225 129.930 55.570 130.475 ;
        RECT 42.405 129.185 43.155 129.705 ;
        RECT 37.640 128.095 38.510 128.435 ;
        RECT 39.100 128.475 39.900 128.645 ;
        RECT 38.680 127.925 38.930 128.385 ;
        RECT 39.100 128.185 39.270 128.475 ;
        RECT 39.450 127.925 39.780 128.305 ;
        RECT 40.075 127.925 40.245 128.985 ;
        RECT 40.455 128.935 42.180 129.105 ;
        RECT 43.325 129.015 44.075 129.535 ;
        RECT 46.290 129.100 46.630 129.930 ;
        RECT 40.455 128.095 40.745 128.935 ;
        RECT 40.915 127.925 41.085 128.765 ;
        RECT 41.295 128.095 41.545 128.935 ;
        RECT 41.755 127.925 41.925 128.765 ;
        RECT 42.405 127.925 44.075 129.015 ;
        RECT 44.245 127.925 44.535 129.090 ;
        RECT 48.110 128.360 48.460 129.610 ;
        RECT 51.810 129.100 52.150 129.930 ;
        RECT 55.745 129.725 56.955 130.475 ;
        RECT 57.125 129.750 57.415 130.475 ;
        RECT 57.590 129.925 57.845 130.215 ;
        RECT 58.015 130.095 58.345 130.475 ;
        RECT 57.590 129.755 58.340 129.925 ;
        RECT 53.630 128.360 53.980 129.610 ;
        RECT 55.745 129.185 56.265 129.725 ;
        RECT 56.435 129.015 56.955 129.555 ;
        RECT 44.705 127.925 50.050 128.360 ;
        RECT 50.225 127.925 55.570 128.360 ;
        RECT 55.745 127.925 56.955 129.015 ;
        RECT 57.125 127.925 57.415 129.090 ;
        RECT 57.590 128.935 57.940 129.585 ;
        RECT 58.110 128.765 58.340 129.755 ;
        RECT 57.590 128.595 58.340 128.765 ;
        RECT 57.590 128.095 57.845 128.595 ;
        RECT 58.015 127.925 58.345 128.425 ;
        RECT 58.515 128.095 58.685 130.215 ;
        RECT 59.045 130.115 59.375 130.475 ;
        RECT 59.545 130.085 60.040 130.255 ;
        RECT 60.245 130.085 61.100 130.255 ;
        RECT 58.915 128.895 59.375 129.945 ;
        RECT 58.855 128.110 59.180 128.895 ;
        RECT 59.545 128.725 59.715 130.085 ;
        RECT 59.885 129.175 60.235 129.795 ;
        RECT 60.405 129.575 60.760 129.795 ;
        RECT 60.405 128.985 60.575 129.575 ;
        RECT 60.930 129.375 61.100 130.085 ;
        RECT 61.975 130.015 62.305 130.475 ;
        RECT 62.515 130.115 62.865 130.285 ;
        RECT 61.305 129.545 62.095 129.795 ;
        RECT 62.515 129.725 62.775 130.115 ;
        RECT 63.085 130.025 64.035 130.305 ;
        RECT 64.205 130.035 64.395 130.475 ;
        RECT 64.565 130.095 65.635 130.265 ;
        RECT 62.265 129.375 62.435 129.555 ;
        RECT 59.545 128.555 59.940 128.725 ;
        RECT 60.110 128.595 60.575 128.985 ;
        RECT 60.745 129.205 62.435 129.375 ;
        RECT 59.770 128.425 59.940 128.555 ;
        RECT 60.745 128.425 60.915 129.205 ;
        RECT 62.605 129.035 62.775 129.725 ;
        RECT 61.275 128.865 62.775 129.035 ;
        RECT 62.965 129.065 63.175 129.855 ;
        RECT 63.345 129.235 63.695 129.855 ;
        RECT 63.865 129.245 64.035 130.025 ;
        RECT 64.565 129.865 64.735 130.095 ;
        RECT 64.205 129.695 64.735 129.865 ;
        RECT 64.205 129.415 64.425 129.695 ;
        RECT 64.905 129.525 65.145 129.925 ;
        RECT 63.865 129.075 64.270 129.245 ;
        RECT 64.605 129.155 65.145 129.525 ;
        RECT 65.315 129.740 65.635 130.095 ;
        RECT 65.315 129.485 65.640 129.740 ;
        RECT 65.835 129.665 66.005 130.475 ;
        RECT 66.175 129.825 66.505 130.305 ;
        RECT 66.675 130.005 66.845 130.475 ;
        RECT 67.015 129.825 67.345 130.305 ;
        RECT 67.515 130.005 67.685 130.475 ;
        RECT 66.175 129.655 67.940 129.825 ;
        RECT 65.315 129.275 67.345 129.485 ;
        RECT 65.315 129.265 65.660 129.275 ;
        RECT 62.965 128.905 63.640 129.065 ;
        RECT 64.100 128.985 64.270 129.075 ;
        RECT 62.965 128.895 63.930 128.905 ;
        RECT 62.605 128.725 62.775 128.865 ;
        RECT 59.350 127.925 59.600 128.385 ;
        RECT 59.770 128.095 60.020 128.425 ;
        RECT 60.235 128.095 60.915 128.425 ;
        RECT 61.085 128.525 62.160 128.695 ;
        RECT 62.605 128.555 63.165 128.725 ;
        RECT 63.470 128.605 63.930 128.895 ;
        RECT 64.100 128.815 65.320 128.985 ;
        RECT 61.085 128.185 61.255 128.525 ;
        RECT 61.490 127.925 61.820 128.355 ;
        RECT 61.990 128.185 62.160 128.525 ;
        RECT 62.455 127.925 62.825 128.385 ;
        RECT 62.995 128.095 63.165 128.555 ;
        RECT 64.100 128.435 64.270 128.815 ;
        RECT 65.490 128.645 65.660 129.265 ;
        RECT 67.530 129.105 67.940 129.655 ;
        RECT 68.165 129.705 69.835 130.475 ;
        RECT 70.005 129.750 70.295 130.475 ;
        RECT 70.465 129.930 75.810 130.475 ;
        RECT 75.985 129.930 81.330 130.475 ;
        RECT 68.165 129.185 68.915 129.705 ;
        RECT 63.400 128.095 64.270 128.435 ;
        RECT 64.860 128.475 65.660 128.645 ;
        RECT 64.440 127.925 64.690 128.385 ;
        RECT 64.860 128.185 65.030 128.475 ;
        RECT 65.210 127.925 65.540 128.305 ;
        RECT 65.835 127.925 66.005 128.985 ;
        RECT 66.215 128.935 67.940 129.105 ;
        RECT 69.085 129.015 69.835 129.535 ;
        RECT 72.050 129.100 72.390 129.930 ;
        RECT 66.215 128.095 66.505 128.935 ;
        RECT 66.675 127.925 66.845 128.765 ;
        RECT 67.055 128.095 67.305 128.935 ;
        RECT 67.515 127.925 67.685 128.765 ;
        RECT 68.165 127.925 69.835 129.015 ;
        RECT 70.005 127.925 70.295 129.090 ;
        RECT 73.870 128.360 74.220 129.610 ;
        RECT 77.570 129.100 77.910 129.930 ;
        RECT 81.505 129.725 82.715 130.475 ;
        RECT 82.885 129.750 83.175 130.475 ;
        RECT 83.345 129.930 88.690 130.475 ;
        RECT 88.865 129.930 94.210 130.475 ;
        RECT 79.390 128.360 79.740 129.610 ;
        RECT 81.505 129.185 82.025 129.725 ;
        RECT 82.195 129.015 82.715 129.555 ;
        RECT 84.930 129.100 85.270 129.930 ;
        RECT 70.465 127.925 75.810 128.360 ;
        RECT 75.985 127.925 81.330 128.360 ;
        RECT 81.505 127.925 82.715 129.015 ;
        RECT 82.885 127.925 83.175 129.090 ;
        RECT 86.750 128.360 87.100 129.610 ;
        RECT 90.450 129.100 90.790 129.930 ;
        RECT 94.385 129.725 95.595 130.475 ;
        RECT 95.765 129.750 96.055 130.475 ;
        RECT 96.225 129.930 101.570 130.475 ;
        RECT 101.745 129.930 107.090 130.475 ;
        RECT 92.270 128.360 92.620 129.610 ;
        RECT 94.385 129.185 94.905 129.725 ;
        RECT 95.075 129.015 95.595 129.555 ;
        RECT 97.810 129.100 98.150 129.930 ;
        RECT 83.345 127.925 88.690 128.360 ;
        RECT 88.865 127.925 94.210 128.360 ;
        RECT 94.385 127.925 95.595 129.015 ;
        RECT 95.765 127.925 96.055 129.090 ;
        RECT 99.630 128.360 99.980 129.610 ;
        RECT 103.330 129.100 103.670 129.930 ;
        RECT 107.265 129.725 108.475 130.475 ;
        RECT 108.645 129.750 108.935 130.475 ;
        RECT 109.105 129.725 110.315 130.475 ;
        RECT 110.490 129.925 110.745 130.215 ;
        RECT 110.915 130.095 111.245 130.475 ;
        RECT 110.490 129.755 111.240 129.925 ;
        RECT 105.150 128.360 105.500 129.610 ;
        RECT 107.265 129.185 107.785 129.725 ;
        RECT 107.955 129.015 108.475 129.555 ;
        RECT 109.105 129.185 109.625 129.725 ;
        RECT 96.225 127.925 101.570 128.360 ;
        RECT 101.745 127.925 107.090 128.360 ;
        RECT 107.265 127.925 108.475 129.015 ;
        RECT 108.645 127.925 108.935 129.090 ;
        RECT 109.795 129.015 110.315 129.555 ;
        RECT 109.105 127.925 110.315 129.015 ;
        RECT 110.490 128.935 110.840 129.585 ;
        RECT 111.010 128.765 111.240 129.755 ;
        RECT 110.490 128.595 111.240 128.765 ;
        RECT 110.490 128.095 110.745 128.595 ;
        RECT 110.915 127.925 111.245 128.425 ;
        RECT 111.415 128.095 111.585 130.215 ;
        RECT 111.945 130.115 112.275 130.475 ;
        RECT 112.445 130.085 112.940 130.255 ;
        RECT 113.145 130.085 114.000 130.255 ;
        RECT 111.815 128.895 112.275 129.945 ;
        RECT 111.755 128.110 112.080 128.895 ;
        RECT 112.445 128.725 112.615 130.085 ;
        RECT 112.785 129.175 113.135 129.795 ;
        RECT 113.305 129.575 113.660 129.795 ;
        RECT 113.305 128.985 113.475 129.575 ;
        RECT 113.830 129.375 114.000 130.085 ;
        RECT 114.875 130.015 115.205 130.475 ;
        RECT 115.415 130.115 115.765 130.285 ;
        RECT 114.205 129.545 114.995 129.795 ;
        RECT 115.415 129.725 115.675 130.115 ;
        RECT 115.985 130.025 116.935 130.305 ;
        RECT 117.105 130.035 117.295 130.475 ;
        RECT 117.465 130.095 118.535 130.265 ;
        RECT 115.165 129.375 115.335 129.555 ;
        RECT 112.445 128.555 112.840 128.725 ;
        RECT 113.010 128.595 113.475 128.985 ;
        RECT 113.645 129.205 115.335 129.375 ;
        RECT 112.670 128.425 112.840 128.555 ;
        RECT 113.645 128.425 113.815 129.205 ;
        RECT 115.505 129.035 115.675 129.725 ;
        RECT 114.175 128.865 115.675 129.035 ;
        RECT 115.865 129.065 116.075 129.855 ;
        RECT 116.245 129.235 116.595 129.855 ;
        RECT 116.765 129.245 116.935 130.025 ;
        RECT 117.465 129.865 117.635 130.095 ;
        RECT 117.105 129.695 117.635 129.865 ;
        RECT 117.105 129.415 117.325 129.695 ;
        RECT 117.805 129.525 118.045 129.925 ;
        RECT 116.765 129.075 117.170 129.245 ;
        RECT 117.505 129.155 118.045 129.525 ;
        RECT 118.215 129.740 118.535 130.095 ;
        RECT 118.215 129.485 118.540 129.740 ;
        RECT 118.735 129.665 118.905 130.475 ;
        RECT 119.075 129.825 119.405 130.305 ;
        RECT 119.575 130.005 119.745 130.475 ;
        RECT 119.915 129.825 120.245 130.305 ;
        RECT 120.415 130.005 120.585 130.475 ;
        RECT 119.075 129.655 120.840 129.825 ;
        RECT 121.525 129.750 121.815 130.475 ;
        RECT 118.215 129.275 120.245 129.485 ;
        RECT 118.215 129.265 118.560 129.275 ;
        RECT 115.865 128.905 116.540 129.065 ;
        RECT 117.000 128.985 117.170 129.075 ;
        RECT 115.865 128.895 116.830 128.905 ;
        RECT 115.505 128.725 115.675 128.865 ;
        RECT 112.250 127.925 112.500 128.385 ;
        RECT 112.670 128.095 112.920 128.425 ;
        RECT 113.135 128.095 113.815 128.425 ;
        RECT 113.985 128.525 115.060 128.695 ;
        RECT 115.505 128.555 116.065 128.725 ;
        RECT 116.370 128.605 116.830 128.895 ;
        RECT 117.000 128.815 118.220 128.985 ;
        RECT 113.985 128.185 114.155 128.525 ;
        RECT 114.390 127.925 114.720 128.355 ;
        RECT 114.890 128.185 115.060 128.525 ;
        RECT 115.355 127.925 115.725 128.385 ;
        RECT 115.895 128.095 116.065 128.555 ;
        RECT 117.000 128.435 117.170 128.815 ;
        RECT 118.390 128.645 118.560 129.265 ;
        RECT 120.430 129.105 120.840 129.655 ;
        RECT 121.985 129.705 123.655 130.475 ;
        RECT 124.285 129.725 125.495 130.475 ;
        RECT 121.985 129.185 122.735 129.705 ;
        RECT 116.300 128.095 117.170 128.435 ;
        RECT 117.760 128.475 118.560 128.645 ;
        RECT 117.340 127.925 117.590 128.385 ;
        RECT 117.760 128.185 117.930 128.475 ;
        RECT 118.110 127.925 118.440 128.305 ;
        RECT 118.735 127.925 118.905 128.985 ;
        RECT 119.115 128.935 120.840 129.105 ;
        RECT 119.115 128.095 119.405 128.935 ;
        RECT 119.575 127.925 119.745 128.765 ;
        RECT 119.955 128.095 120.205 128.935 ;
        RECT 120.415 127.925 120.585 128.765 ;
        RECT 121.525 127.925 121.815 129.090 ;
        RECT 122.905 129.015 123.655 129.535 ;
        RECT 121.985 127.925 123.655 129.015 ;
        RECT 124.285 129.015 124.805 129.555 ;
        RECT 124.975 129.185 125.495 129.725 ;
        RECT 124.285 127.925 125.495 129.015 ;
        RECT 5.520 127.755 125.580 127.925 ;
        RECT 5.605 126.665 6.815 127.755 ;
        RECT 7.910 127.085 8.165 127.585 ;
        RECT 8.335 127.255 8.665 127.755 ;
        RECT 7.910 126.915 8.660 127.085 ;
        RECT 5.605 125.955 6.125 126.495 ;
        RECT 6.295 126.125 6.815 126.665 ;
        RECT 7.910 126.095 8.260 126.745 ;
        RECT 5.605 125.205 6.815 125.955 ;
        RECT 8.430 125.925 8.660 126.915 ;
        RECT 7.910 125.755 8.660 125.925 ;
        RECT 7.910 125.465 8.165 125.755 ;
        RECT 8.335 125.205 8.665 125.585 ;
        RECT 8.835 125.465 9.005 127.585 ;
        RECT 9.175 126.785 9.500 127.570 ;
        RECT 9.670 127.295 9.920 127.755 ;
        RECT 10.090 127.255 10.340 127.585 ;
        RECT 10.555 127.255 11.235 127.585 ;
        RECT 10.090 127.125 10.260 127.255 ;
        RECT 9.865 126.955 10.260 127.125 ;
        RECT 9.235 125.735 9.695 126.785 ;
        RECT 9.865 125.595 10.035 126.955 ;
        RECT 10.430 126.695 10.895 127.085 ;
        RECT 10.205 125.885 10.555 126.505 ;
        RECT 10.725 126.105 10.895 126.695 ;
        RECT 11.065 126.475 11.235 127.255 ;
        RECT 11.405 127.155 11.575 127.495 ;
        RECT 11.810 127.325 12.140 127.755 ;
        RECT 12.310 127.155 12.480 127.495 ;
        RECT 12.775 127.295 13.145 127.755 ;
        RECT 11.405 126.985 12.480 127.155 ;
        RECT 13.315 127.125 13.485 127.585 ;
        RECT 13.720 127.245 14.590 127.585 ;
        RECT 14.760 127.295 15.010 127.755 ;
        RECT 12.925 126.955 13.485 127.125 ;
        RECT 12.925 126.815 13.095 126.955 ;
        RECT 11.595 126.645 13.095 126.815 ;
        RECT 13.790 126.785 14.250 127.075 ;
        RECT 11.065 126.305 12.755 126.475 ;
        RECT 10.725 125.885 11.080 126.105 ;
        RECT 11.250 125.595 11.420 126.305 ;
        RECT 11.625 125.885 12.415 126.135 ;
        RECT 12.585 126.125 12.755 126.305 ;
        RECT 12.925 125.955 13.095 126.645 ;
        RECT 9.365 125.205 9.695 125.565 ;
        RECT 9.865 125.425 10.360 125.595 ;
        RECT 10.565 125.425 11.420 125.595 ;
        RECT 12.295 125.205 12.625 125.665 ;
        RECT 12.835 125.565 13.095 125.955 ;
        RECT 13.285 126.775 14.250 126.785 ;
        RECT 14.420 126.865 14.590 127.245 ;
        RECT 15.180 127.205 15.350 127.495 ;
        RECT 15.530 127.375 15.860 127.755 ;
        RECT 15.180 127.035 15.980 127.205 ;
        RECT 13.285 126.615 13.960 126.775 ;
        RECT 14.420 126.695 15.640 126.865 ;
        RECT 13.285 125.825 13.495 126.615 ;
        RECT 14.420 126.605 14.590 126.695 ;
        RECT 13.665 125.825 14.015 126.445 ;
        RECT 14.185 126.435 14.590 126.605 ;
        RECT 14.185 125.655 14.355 126.435 ;
        RECT 14.525 125.985 14.745 126.265 ;
        RECT 14.925 126.155 15.465 126.525 ;
        RECT 15.810 126.415 15.980 127.035 ;
        RECT 16.155 126.695 16.325 127.755 ;
        RECT 16.535 126.745 16.825 127.585 ;
        RECT 16.995 126.915 17.165 127.755 ;
        RECT 17.375 126.745 17.625 127.585 ;
        RECT 17.835 126.915 18.005 127.755 ;
        RECT 16.535 126.575 18.260 126.745 ;
        RECT 18.485 126.590 18.775 127.755 ;
        RECT 18.945 126.665 22.455 127.755 ;
        RECT 23.090 127.085 23.345 127.585 ;
        RECT 23.515 127.255 23.845 127.755 ;
        RECT 23.090 126.915 23.840 127.085 ;
        RECT 14.525 125.815 15.055 125.985 ;
        RECT 12.835 125.395 13.185 125.565 ;
        RECT 13.405 125.375 14.355 125.655 ;
        RECT 14.525 125.205 14.715 125.645 ;
        RECT 14.885 125.585 15.055 125.815 ;
        RECT 15.225 125.755 15.465 126.155 ;
        RECT 15.635 126.405 15.980 126.415 ;
        RECT 15.635 126.195 17.665 126.405 ;
        RECT 15.635 125.940 15.960 126.195 ;
        RECT 17.850 126.025 18.260 126.575 ;
        RECT 15.635 125.585 15.955 125.940 ;
        RECT 14.885 125.415 15.955 125.585 ;
        RECT 16.155 125.205 16.325 126.015 ;
        RECT 16.495 125.855 18.260 126.025 ;
        RECT 18.945 125.975 20.595 126.495 ;
        RECT 20.765 126.145 22.455 126.665 ;
        RECT 23.090 126.095 23.440 126.745 ;
        RECT 16.495 125.375 16.825 125.855 ;
        RECT 16.995 125.205 17.165 125.675 ;
        RECT 17.335 125.375 17.665 125.855 ;
        RECT 17.835 125.205 18.005 125.675 ;
        RECT 18.485 125.205 18.775 125.930 ;
        RECT 18.945 125.205 22.455 125.975 ;
        RECT 23.610 125.925 23.840 126.915 ;
        RECT 23.090 125.755 23.840 125.925 ;
        RECT 23.090 125.465 23.345 125.755 ;
        RECT 23.515 125.205 23.845 125.585 ;
        RECT 24.015 125.465 24.185 127.585 ;
        RECT 24.355 126.785 24.680 127.570 ;
        RECT 24.850 127.295 25.100 127.755 ;
        RECT 25.270 127.255 25.520 127.585 ;
        RECT 25.735 127.255 26.415 127.585 ;
        RECT 25.270 127.125 25.440 127.255 ;
        RECT 25.045 126.955 25.440 127.125 ;
        RECT 24.415 125.735 24.875 126.785 ;
        RECT 25.045 125.595 25.215 126.955 ;
        RECT 25.610 126.695 26.075 127.085 ;
        RECT 25.385 125.885 25.735 126.505 ;
        RECT 25.905 126.105 26.075 126.695 ;
        RECT 26.245 126.475 26.415 127.255 ;
        RECT 26.585 127.155 26.755 127.495 ;
        RECT 26.990 127.325 27.320 127.755 ;
        RECT 27.490 127.155 27.660 127.495 ;
        RECT 27.955 127.295 28.325 127.755 ;
        RECT 26.585 126.985 27.660 127.155 ;
        RECT 28.495 127.125 28.665 127.585 ;
        RECT 28.900 127.245 29.770 127.585 ;
        RECT 29.940 127.295 30.190 127.755 ;
        RECT 28.105 126.955 28.665 127.125 ;
        RECT 28.105 126.815 28.275 126.955 ;
        RECT 26.775 126.645 28.275 126.815 ;
        RECT 28.970 126.785 29.430 127.075 ;
        RECT 26.245 126.305 27.935 126.475 ;
        RECT 25.905 125.885 26.260 126.105 ;
        RECT 26.430 125.595 26.600 126.305 ;
        RECT 26.805 125.885 27.595 126.135 ;
        RECT 27.765 126.125 27.935 126.305 ;
        RECT 28.105 125.955 28.275 126.645 ;
        RECT 24.545 125.205 24.875 125.565 ;
        RECT 25.045 125.425 25.540 125.595 ;
        RECT 25.745 125.425 26.600 125.595 ;
        RECT 27.475 125.205 27.805 125.665 ;
        RECT 28.015 125.565 28.275 125.955 ;
        RECT 28.465 126.775 29.430 126.785 ;
        RECT 29.600 126.865 29.770 127.245 ;
        RECT 30.360 127.205 30.530 127.495 ;
        RECT 30.710 127.375 31.040 127.755 ;
        RECT 30.360 127.035 31.160 127.205 ;
        RECT 28.465 126.615 29.140 126.775 ;
        RECT 29.600 126.695 30.820 126.865 ;
        RECT 28.465 125.825 28.675 126.615 ;
        RECT 29.600 126.605 29.770 126.695 ;
        RECT 28.845 125.825 29.195 126.445 ;
        RECT 29.365 126.435 29.770 126.605 ;
        RECT 29.365 125.655 29.535 126.435 ;
        RECT 29.705 125.985 29.925 126.265 ;
        RECT 30.105 126.155 30.645 126.525 ;
        RECT 30.990 126.415 31.160 127.035 ;
        RECT 31.335 126.695 31.505 127.755 ;
        RECT 31.715 126.745 32.005 127.585 ;
        RECT 32.175 126.915 32.345 127.755 ;
        RECT 32.555 126.745 32.805 127.585 ;
        RECT 33.015 126.915 33.185 127.755 ;
        RECT 33.670 127.085 33.925 127.585 ;
        RECT 34.095 127.255 34.425 127.755 ;
        RECT 33.670 126.915 34.420 127.085 ;
        RECT 31.715 126.575 33.440 126.745 ;
        RECT 29.705 125.815 30.235 125.985 ;
        RECT 28.015 125.395 28.365 125.565 ;
        RECT 28.585 125.375 29.535 125.655 ;
        RECT 29.705 125.205 29.895 125.645 ;
        RECT 30.065 125.585 30.235 125.815 ;
        RECT 30.405 125.755 30.645 126.155 ;
        RECT 30.815 126.405 31.160 126.415 ;
        RECT 30.815 126.195 32.845 126.405 ;
        RECT 30.815 125.940 31.140 126.195 ;
        RECT 33.030 126.025 33.440 126.575 ;
        RECT 33.670 126.095 34.020 126.745 ;
        RECT 30.815 125.585 31.135 125.940 ;
        RECT 30.065 125.415 31.135 125.585 ;
        RECT 31.335 125.205 31.505 126.015 ;
        RECT 31.675 125.855 33.440 126.025 ;
        RECT 34.190 125.925 34.420 126.915 ;
        RECT 31.675 125.375 32.005 125.855 ;
        RECT 32.175 125.205 32.345 125.675 ;
        RECT 32.515 125.375 32.845 125.855 ;
        RECT 33.670 125.755 34.420 125.925 ;
        RECT 33.015 125.205 33.185 125.675 ;
        RECT 33.670 125.465 33.925 125.755 ;
        RECT 34.095 125.205 34.425 125.585 ;
        RECT 34.595 125.465 34.765 127.585 ;
        RECT 34.935 126.785 35.260 127.570 ;
        RECT 35.430 127.295 35.680 127.755 ;
        RECT 35.850 127.255 36.100 127.585 ;
        RECT 36.315 127.255 36.995 127.585 ;
        RECT 35.850 127.125 36.020 127.255 ;
        RECT 35.625 126.955 36.020 127.125 ;
        RECT 34.995 125.735 35.455 126.785 ;
        RECT 35.625 125.595 35.795 126.955 ;
        RECT 36.190 126.695 36.655 127.085 ;
        RECT 35.965 125.885 36.315 126.505 ;
        RECT 36.485 126.105 36.655 126.695 ;
        RECT 36.825 126.475 36.995 127.255 ;
        RECT 37.165 127.155 37.335 127.495 ;
        RECT 37.570 127.325 37.900 127.755 ;
        RECT 38.070 127.155 38.240 127.495 ;
        RECT 38.535 127.295 38.905 127.755 ;
        RECT 37.165 126.985 38.240 127.155 ;
        RECT 39.075 127.125 39.245 127.585 ;
        RECT 39.480 127.245 40.350 127.585 ;
        RECT 40.520 127.295 40.770 127.755 ;
        RECT 38.685 126.955 39.245 127.125 ;
        RECT 38.685 126.815 38.855 126.955 ;
        RECT 37.355 126.645 38.855 126.815 ;
        RECT 39.550 126.785 40.010 127.075 ;
        RECT 36.825 126.305 38.515 126.475 ;
        RECT 36.485 125.885 36.840 126.105 ;
        RECT 37.010 125.595 37.180 126.305 ;
        RECT 37.385 125.885 38.175 126.135 ;
        RECT 38.345 126.125 38.515 126.305 ;
        RECT 38.685 125.955 38.855 126.645 ;
        RECT 35.125 125.205 35.455 125.565 ;
        RECT 35.625 125.425 36.120 125.595 ;
        RECT 36.325 125.425 37.180 125.595 ;
        RECT 38.055 125.205 38.385 125.665 ;
        RECT 38.595 125.565 38.855 125.955 ;
        RECT 39.045 126.775 40.010 126.785 ;
        RECT 40.180 126.865 40.350 127.245 ;
        RECT 40.940 127.205 41.110 127.495 ;
        RECT 41.290 127.375 41.620 127.755 ;
        RECT 40.940 127.035 41.740 127.205 ;
        RECT 39.045 126.615 39.720 126.775 ;
        RECT 40.180 126.695 41.400 126.865 ;
        RECT 39.045 125.825 39.255 126.615 ;
        RECT 40.180 126.605 40.350 126.695 ;
        RECT 39.425 125.825 39.775 126.445 ;
        RECT 39.945 126.435 40.350 126.605 ;
        RECT 39.945 125.655 40.115 126.435 ;
        RECT 40.285 125.985 40.505 126.265 ;
        RECT 40.685 126.155 41.225 126.525 ;
        RECT 41.570 126.415 41.740 127.035 ;
        RECT 41.915 126.695 42.085 127.755 ;
        RECT 42.295 126.745 42.585 127.585 ;
        RECT 42.755 126.915 42.925 127.755 ;
        RECT 43.135 126.745 43.385 127.585 ;
        RECT 43.595 126.915 43.765 127.755 ;
        RECT 42.295 126.575 44.020 126.745 ;
        RECT 44.245 126.590 44.535 127.755 ;
        RECT 44.705 126.665 46.375 127.755 ;
        RECT 40.285 125.815 40.815 125.985 ;
        RECT 38.595 125.395 38.945 125.565 ;
        RECT 39.165 125.375 40.115 125.655 ;
        RECT 40.285 125.205 40.475 125.645 ;
        RECT 40.645 125.585 40.815 125.815 ;
        RECT 40.985 125.755 41.225 126.155 ;
        RECT 41.395 126.405 41.740 126.415 ;
        RECT 41.395 126.195 43.425 126.405 ;
        RECT 41.395 125.940 41.720 126.195 ;
        RECT 43.610 126.025 44.020 126.575 ;
        RECT 41.395 125.585 41.715 125.940 ;
        RECT 40.645 125.415 41.715 125.585 ;
        RECT 41.915 125.205 42.085 126.015 ;
        RECT 42.255 125.855 44.020 126.025 ;
        RECT 44.705 125.975 45.455 126.495 ;
        RECT 45.625 126.145 46.375 126.665 ;
        RECT 46.585 126.615 46.815 127.755 ;
        RECT 46.985 126.605 47.315 127.585 ;
        RECT 47.485 126.615 47.695 127.755 ;
        RECT 48.850 127.085 49.105 127.585 ;
        RECT 49.275 127.255 49.605 127.755 ;
        RECT 48.850 126.915 49.600 127.085 ;
        RECT 46.565 126.195 46.895 126.445 ;
        RECT 42.255 125.375 42.585 125.855 ;
        RECT 42.755 125.205 42.925 125.675 ;
        RECT 43.095 125.375 43.425 125.855 ;
        RECT 43.595 125.205 43.765 125.675 ;
        RECT 44.245 125.205 44.535 125.930 ;
        RECT 44.705 125.205 46.375 125.975 ;
        RECT 46.585 125.205 46.815 126.025 ;
        RECT 47.065 126.005 47.315 126.605 ;
        RECT 48.850 126.095 49.200 126.745 ;
        RECT 46.985 125.375 47.315 126.005 ;
        RECT 47.485 125.205 47.695 126.025 ;
        RECT 49.370 125.925 49.600 126.915 ;
        RECT 48.850 125.755 49.600 125.925 ;
        RECT 48.850 125.465 49.105 125.755 ;
        RECT 49.275 125.205 49.605 125.585 ;
        RECT 49.775 125.465 49.945 127.585 ;
        RECT 50.115 126.785 50.440 127.570 ;
        RECT 50.610 127.295 50.860 127.755 ;
        RECT 51.030 127.255 51.280 127.585 ;
        RECT 51.495 127.255 52.175 127.585 ;
        RECT 51.030 127.125 51.200 127.255 ;
        RECT 50.805 126.955 51.200 127.125 ;
        RECT 50.175 125.735 50.635 126.785 ;
        RECT 50.805 125.595 50.975 126.955 ;
        RECT 51.370 126.695 51.835 127.085 ;
        RECT 51.145 125.885 51.495 126.505 ;
        RECT 51.665 126.105 51.835 126.695 ;
        RECT 52.005 126.475 52.175 127.255 ;
        RECT 52.345 127.155 52.515 127.495 ;
        RECT 52.750 127.325 53.080 127.755 ;
        RECT 53.250 127.155 53.420 127.495 ;
        RECT 53.715 127.295 54.085 127.755 ;
        RECT 52.345 126.985 53.420 127.155 ;
        RECT 54.255 127.125 54.425 127.585 ;
        RECT 54.660 127.245 55.530 127.585 ;
        RECT 55.700 127.295 55.950 127.755 ;
        RECT 53.865 126.955 54.425 127.125 ;
        RECT 53.865 126.815 54.035 126.955 ;
        RECT 52.535 126.645 54.035 126.815 ;
        RECT 54.730 126.785 55.190 127.075 ;
        RECT 52.005 126.305 53.695 126.475 ;
        RECT 51.665 125.885 52.020 126.105 ;
        RECT 52.190 125.595 52.360 126.305 ;
        RECT 52.565 125.885 53.355 126.135 ;
        RECT 53.525 126.125 53.695 126.305 ;
        RECT 53.865 125.955 54.035 126.645 ;
        RECT 50.305 125.205 50.635 125.565 ;
        RECT 50.805 125.425 51.300 125.595 ;
        RECT 51.505 125.425 52.360 125.595 ;
        RECT 53.235 125.205 53.565 125.665 ;
        RECT 53.775 125.565 54.035 125.955 ;
        RECT 54.225 126.775 55.190 126.785 ;
        RECT 55.360 126.865 55.530 127.245 ;
        RECT 56.120 127.205 56.290 127.495 ;
        RECT 56.470 127.375 56.800 127.755 ;
        RECT 56.120 127.035 56.920 127.205 ;
        RECT 54.225 126.615 54.900 126.775 ;
        RECT 55.360 126.695 56.580 126.865 ;
        RECT 54.225 125.825 54.435 126.615 ;
        RECT 55.360 126.605 55.530 126.695 ;
        RECT 54.605 125.825 54.955 126.445 ;
        RECT 55.125 126.435 55.530 126.605 ;
        RECT 55.125 125.655 55.295 126.435 ;
        RECT 55.465 125.985 55.685 126.265 ;
        RECT 55.865 126.155 56.405 126.525 ;
        RECT 56.750 126.415 56.920 127.035 ;
        RECT 57.095 126.695 57.265 127.755 ;
        RECT 57.475 126.745 57.765 127.585 ;
        RECT 57.935 126.915 58.105 127.755 ;
        RECT 58.315 126.745 58.565 127.585 ;
        RECT 58.775 126.915 58.945 127.755 ;
        RECT 59.430 127.085 59.685 127.585 ;
        RECT 59.855 127.255 60.185 127.755 ;
        RECT 59.430 126.915 60.180 127.085 ;
        RECT 57.475 126.575 59.200 126.745 ;
        RECT 55.465 125.815 55.995 125.985 ;
        RECT 53.775 125.395 54.125 125.565 ;
        RECT 54.345 125.375 55.295 125.655 ;
        RECT 55.465 125.205 55.655 125.645 ;
        RECT 55.825 125.585 55.995 125.815 ;
        RECT 56.165 125.755 56.405 126.155 ;
        RECT 56.575 126.405 56.920 126.415 ;
        RECT 56.575 126.195 58.605 126.405 ;
        RECT 56.575 125.940 56.900 126.195 ;
        RECT 58.790 126.025 59.200 126.575 ;
        RECT 59.430 126.095 59.780 126.745 ;
        RECT 56.575 125.585 56.895 125.940 ;
        RECT 55.825 125.415 56.895 125.585 ;
        RECT 57.095 125.205 57.265 126.015 ;
        RECT 57.435 125.855 59.200 126.025 ;
        RECT 59.950 125.925 60.180 126.915 ;
        RECT 57.435 125.375 57.765 125.855 ;
        RECT 57.935 125.205 58.105 125.675 ;
        RECT 58.275 125.375 58.605 125.855 ;
        RECT 59.430 125.755 60.180 125.925 ;
        RECT 58.775 125.205 58.945 125.675 ;
        RECT 59.430 125.465 59.685 125.755 ;
        RECT 59.855 125.205 60.185 125.585 ;
        RECT 60.355 125.465 60.525 127.585 ;
        RECT 60.695 126.785 61.020 127.570 ;
        RECT 61.190 127.295 61.440 127.755 ;
        RECT 61.610 127.255 61.860 127.585 ;
        RECT 62.075 127.255 62.755 127.585 ;
        RECT 61.610 127.125 61.780 127.255 ;
        RECT 61.385 126.955 61.780 127.125 ;
        RECT 60.755 125.735 61.215 126.785 ;
        RECT 61.385 125.595 61.555 126.955 ;
        RECT 61.950 126.695 62.415 127.085 ;
        RECT 61.725 125.885 62.075 126.505 ;
        RECT 62.245 126.105 62.415 126.695 ;
        RECT 62.585 126.475 62.755 127.255 ;
        RECT 62.925 127.155 63.095 127.495 ;
        RECT 63.330 127.325 63.660 127.755 ;
        RECT 63.830 127.155 64.000 127.495 ;
        RECT 64.295 127.295 64.665 127.755 ;
        RECT 62.925 126.985 64.000 127.155 ;
        RECT 64.835 127.125 65.005 127.585 ;
        RECT 65.240 127.245 66.110 127.585 ;
        RECT 66.280 127.295 66.530 127.755 ;
        RECT 64.445 126.955 65.005 127.125 ;
        RECT 64.445 126.815 64.615 126.955 ;
        RECT 63.115 126.645 64.615 126.815 ;
        RECT 65.310 126.785 65.770 127.075 ;
        RECT 62.585 126.305 64.275 126.475 ;
        RECT 62.245 125.885 62.600 126.105 ;
        RECT 62.770 125.595 62.940 126.305 ;
        RECT 63.145 125.885 63.935 126.135 ;
        RECT 64.105 126.125 64.275 126.305 ;
        RECT 64.445 125.955 64.615 126.645 ;
        RECT 60.885 125.205 61.215 125.565 ;
        RECT 61.385 125.425 61.880 125.595 ;
        RECT 62.085 125.425 62.940 125.595 ;
        RECT 63.815 125.205 64.145 125.665 ;
        RECT 64.355 125.565 64.615 125.955 ;
        RECT 64.805 126.775 65.770 126.785 ;
        RECT 65.940 126.865 66.110 127.245 ;
        RECT 66.700 127.205 66.870 127.495 ;
        RECT 67.050 127.375 67.380 127.755 ;
        RECT 66.700 127.035 67.500 127.205 ;
        RECT 64.805 126.615 65.480 126.775 ;
        RECT 65.940 126.695 67.160 126.865 ;
        RECT 64.805 125.825 65.015 126.615 ;
        RECT 65.940 126.605 66.110 126.695 ;
        RECT 65.185 125.825 65.535 126.445 ;
        RECT 65.705 126.435 66.110 126.605 ;
        RECT 65.705 125.655 65.875 126.435 ;
        RECT 66.045 125.985 66.265 126.265 ;
        RECT 66.445 126.155 66.985 126.525 ;
        RECT 67.330 126.415 67.500 127.035 ;
        RECT 67.675 126.695 67.845 127.755 ;
        RECT 68.055 126.745 68.345 127.585 ;
        RECT 68.515 126.915 68.685 127.755 ;
        RECT 68.895 126.745 69.145 127.585 ;
        RECT 69.355 126.915 69.525 127.755 ;
        RECT 68.055 126.575 69.780 126.745 ;
        RECT 70.005 126.590 70.295 127.755 ;
        RECT 70.465 126.665 73.055 127.755 ;
        RECT 73.690 127.085 73.945 127.585 ;
        RECT 74.115 127.255 74.445 127.755 ;
        RECT 73.690 126.915 74.440 127.085 ;
        RECT 66.045 125.815 66.575 125.985 ;
        RECT 64.355 125.395 64.705 125.565 ;
        RECT 64.925 125.375 65.875 125.655 ;
        RECT 66.045 125.205 66.235 125.645 ;
        RECT 66.405 125.585 66.575 125.815 ;
        RECT 66.745 125.755 66.985 126.155 ;
        RECT 67.155 126.405 67.500 126.415 ;
        RECT 67.155 126.195 69.185 126.405 ;
        RECT 67.155 125.940 67.480 126.195 ;
        RECT 69.370 126.025 69.780 126.575 ;
        RECT 67.155 125.585 67.475 125.940 ;
        RECT 66.405 125.415 67.475 125.585 ;
        RECT 67.675 125.205 67.845 126.015 ;
        RECT 68.015 125.855 69.780 126.025 ;
        RECT 70.465 125.975 71.675 126.495 ;
        RECT 71.845 126.145 73.055 126.665 ;
        RECT 73.690 126.095 74.040 126.745 ;
        RECT 68.015 125.375 68.345 125.855 ;
        RECT 68.515 125.205 68.685 125.675 ;
        RECT 68.855 125.375 69.185 125.855 ;
        RECT 69.355 125.205 69.525 125.675 ;
        RECT 70.005 125.205 70.295 125.930 ;
        RECT 70.465 125.205 73.055 125.975 ;
        RECT 74.210 125.925 74.440 126.915 ;
        RECT 73.690 125.755 74.440 125.925 ;
        RECT 73.690 125.465 73.945 125.755 ;
        RECT 74.115 125.205 74.445 125.585 ;
        RECT 74.615 125.465 74.785 127.585 ;
        RECT 74.955 126.785 75.280 127.570 ;
        RECT 75.450 127.295 75.700 127.755 ;
        RECT 75.870 127.255 76.120 127.585 ;
        RECT 76.335 127.255 77.015 127.585 ;
        RECT 75.870 127.125 76.040 127.255 ;
        RECT 75.645 126.955 76.040 127.125 ;
        RECT 75.015 125.735 75.475 126.785 ;
        RECT 75.645 125.595 75.815 126.955 ;
        RECT 76.210 126.695 76.675 127.085 ;
        RECT 75.985 125.885 76.335 126.505 ;
        RECT 76.505 126.105 76.675 126.695 ;
        RECT 76.845 126.475 77.015 127.255 ;
        RECT 77.185 127.155 77.355 127.495 ;
        RECT 77.590 127.325 77.920 127.755 ;
        RECT 78.090 127.155 78.260 127.495 ;
        RECT 78.555 127.295 78.925 127.755 ;
        RECT 77.185 126.985 78.260 127.155 ;
        RECT 79.095 127.125 79.265 127.585 ;
        RECT 79.500 127.245 80.370 127.585 ;
        RECT 80.540 127.295 80.790 127.755 ;
        RECT 78.705 126.955 79.265 127.125 ;
        RECT 78.705 126.815 78.875 126.955 ;
        RECT 77.375 126.645 78.875 126.815 ;
        RECT 79.570 126.785 80.030 127.075 ;
        RECT 76.845 126.305 78.535 126.475 ;
        RECT 76.505 125.885 76.860 126.105 ;
        RECT 77.030 125.595 77.200 126.305 ;
        RECT 77.405 125.885 78.195 126.135 ;
        RECT 78.365 126.125 78.535 126.305 ;
        RECT 78.705 125.955 78.875 126.645 ;
        RECT 75.145 125.205 75.475 125.565 ;
        RECT 75.645 125.425 76.140 125.595 ;
        RECT 76.345 125.425 77.200 125.595 ;
        RECT 78.075 125.205 78.405 125.665 ;
        RECT 78.615 125.565 78.875 125.955 ;
        RECT 79.065 126.775 80.030 126.785 ;
        RECT 80.200 126.865 80.370 127.245 ;
        RECT 80.960 127.205 81.130 127.495 ;
        RECT 81.310 127.375 81.640 127.755 ;
        RECT 80.960 127.035 81.760 127.205 ;
        RECT 79.065 126.615 79.740 126.775 ;
        RECT 80.200 126.695 81.420 126.865 ;
        RECT 79.065 125.825 79.275 126.615 ;
        RECT 80.200 126.605 80.370 126.695 ;
        RECT 79.445 125.825 79.795 126.445 ;
        RECT 79.965 126.435 80.370 126.605 ;
        RECT 79.965 125.655 80.135 126.435 ;
        RECT 80.305 125.985 80.525 126.265 ;
        RECT 80.705 126.155 81.245 126.525 ;
        RECT 81.590 126.415 81.760 127.035 ;
        RECT 81.935 126.695 82.105 127.755 ;
        RECT 82.315 126.745 82.605 127.585 ;
        RECT 82.775 126.915 82.945 127.755 ;
        RECT 83.155 126.745 83.405 127.585 ;
        RECT 83.615 126.915 83.785 127.755 ;
        RECT 84.270 127.085 84.525 127.585 ;
        RECT 84.695 127.255 85.025 127.755 ;
        RECT 84.270 126.915 85.020 127.085 ;
        RECT 82.315 126.575 84.040 126.745 ;
        RECT 80.305 125.815 80.835 125.985 ;
        RECT 78.615 125.395 78.965 125.565 ;
        RECT 79.185 125.375 80.135 125.655 ;
        RECT 80.305 125.205 80.495 125.645 ;
        RECT 80.665 125.585 80.835 125.815 ;
        RECT 81.005 125.755 81.245 126.155 ;
        RECT 81.415 126.405 81.760 126.415 ;
        RECT 81.415 126.195 83.445 126.405 ;
        RECT 81.415 125.940 81.740 126.195 ;
        RECT 83.630 126.025 84.040 126.575 ;
        RECT 84.270 126.095 84.620 126.745 ;
        RECT 81.415 125.585 81.735 125.940 ;
        RECT 80.665 125.415 81.735 125.585 ;
        RECT 81.935 125.205 82.105 126.015 ;
        RECT 82.275 125.855 84.040 126.025 ;
        RECT 84.790 125.925 85.020 126.915 ;
        RECT 82.275 125.375 82.605 125.855 ;
        RECT 82.775 125.205 82.945 125.675 ;
        RECT 83.115 125.375 83.445 125.855 ;
        RECT 84.270 125.755 85.020 125.925 ;
        RECT 83.615 125.205 83.785 125.675 ;
        RECT 84.270 125.465 84.525 125.755 ;
        RECT 84.695 125.205 85.025 125.585 ;
        RECT 85.195 125.465 85.365 127.585 ;
        RECT 85.535 126.785 85.860 127.570 ;
        RECT 86.030 127.295 86.280 127.755 ;
        RECT 86.450 127.255 86.700 127.585 ;
        RECT 86.915 127.255 87.595 127.585 ;
        RECT 86.450 127.125 86.620 127.255 ;
        RECT 86.225 126.955 86.620 127.125 ;
        RECT 85.595 125.735 86.055 126.785 ;
        RECT 86.225 125.595 86.395 126.955 ;
        RECT 86.790 126.695 87.255 127.085 ;
        RECT 86.565 125.885 86.915 126.505 ;
        RECT 87.085 126.105 87.255 126.695 ;
        RECT 87.425 126.475 87.595 127.255 ;
        RECT 87.765 127.155 87.935 127.495 ;
        RECT 88.170 127.325 88.500 127.755 ;
        RECT 88.670 127.155 88.840 127.495 ;
        RECT 89.135 127.295 89.505 127.755 ;
        RECT 87.765 126.985 88.840 127.155 ;
        RECT 89.675 127.125 89.845 127.585 ;
        RECT 90.080 127.245 90.950 127.585 ;
        RECT 91.120 127.295 91.370 127.755 ;
        RECT 89.285 126.955 89.845 127.125 ;
        RECT 89.285 126.815 89.455 126.955 ;
        RECT 87.955 126.645 89.455 126.815 ;
        RECT 90.150 126.785 90.610 127.075 ;
        RECT 87.425 126.305 89.115 126.475 ;
        RECT 87.085 125.885 87.440 126.105 ;
        RECT 87.610 125.595 87.780 126.305 ;
        RECT 87.985 125.885 88.775 126.135 ;
        RECT 88.945 126.125 89.115 126.305 ;
        RECT 89.285 125.955 89.455 126.645 ;
        RECT 85.725 125.205 86.055 125.565 ;
        RECT 86.225 125.425 86.720 125.595 ;
        RECT 86.925 125.425 87.780 125.595 ;
        RECT 88.655 125.205 88.985 125.665 ;
        RECT 89.195 125.565 89.455 125.955 ;
        RECT 89.645 126.775 90.610 126.785 ;
        RECT 90.780 126.865 90.950 127.245 ;
        RECT 91.540 127.205 91.710 127.495 ;
        RECT 91.890 127.375 92.220 127.755 ;
        RECT 91.540 127.035 92.340 127.205 ;
        RECT 89.645 126.615 90.320 126.775 ;
        RECT 90.780 126.695 92.000 126.865 ;
        RECT 89.645 125.825 89.855 126.615 ;
        RECT 90.780 126.605 90.950 126.695 ;
        RECT 90.025 125.825 90.375 126.445 ;
        RECT 90.545 126.435 90.950 126.605 ;
        RECT 90.545 125.655 90.715 126.435 ;
        RECT 90.885 125.985 91.105 126.265 ;
        RECT 91.285 126.155 91.825 126.525 ;
        RECT 92.170 126.415 92.340 127.035 ;
        RECT 92.515 126.695 92.685 127.755 ;
        RECT 92.895 126.745 93.185 127.585 ;
        RECT 93.355 126.915 93.525 127.755 ;
        RECT 93.735 126.745 93.985 127.585 ;
        RECT 94.195 126.915 94.365 127.755 ;
        RECT 92.895 126.575 94.620 126.745 ;
        RECT 95.765 126.590 96.055 127.755 ;
        RECT 96.230 127.085 96.485 127.585 ;
        RECT 96.655 127.255 96.985 127.755 ;
        RECT 96.230 126.915 96.980 127.085 ;
        RECT 90.885 125.815 91.415 125.985 ;
        RECT 89.195 125.395 89.545 125.565 ;
        RECT 89.765 125.375 90.715 125.655 ;
        RECT 90.885 125.205 91.075 125.645 ;
        RECT 91.245 125.585 91.415 125.815 ;
        RECT 91.585 125.755 91.825 126.155 ;
        RECT 91.995 126.405 92.340 126.415 ;
        RECT 91.995 126.195 94.025 126.405 ;
        RECT 91.995 125.940 92.320 126.195 ;
        RECT 94.210 126.025 94.620 126.575 ;
        RECT 96.230 126.095 96.580 126.745 ;
        RECT 91.995 125.585 92.315 125.940 ;
        RECT 91.245 125.415 92.315 125.585 ;
        RECT 92.515 125.205 92.685 126.015 ;
        RECT 92.855 125.855 94.620 126.025 ;
        RECT 92.855 125.375 93.185 125.855 ;
        RECT 93.355 125.205 93.525 125.675 ;
        RECT 93.695 125.375 94.025 125.855 ;
        RECT 94.195 125.205 94.365 125.675 ;
        RECT 95.765 125.205 96.055 125.930 ;
        RECT 96.750 125.925 96.980 126.915 ;
        RECT 96.230 125.755 96.980 125.925 ;
        RECT 96.230 125.465 96.485 125.755 ;
        RECT 96.655 125.205 96.985 125.585 ;
        RECT 97.155 125.465 97.325 127.585 ;
        RECT 97.495 126.785 97.820 127.570 ;
        RECT 97.990 127.295 98.240 127.755 ;
        RECT 98.410 127.255 98.660 127.585 ;
        RECT 98.875 127.255 99.555 127.585 ;
        RECT 98.410 127.125 98.580 127.255 ;
        RECT 98.185 126.955 98.580 127.125 ;
        RECT 97.555 125.735 98.015 126.785 ;
        RECT 98.185 125.595 98.355 126.955 ;
        RECT 98.750 126.695 99.215 127.085 ;
        RECT 98.525 125.885 98.875 126.505 ;
        RECT 99.045 126.105 99.215 126.695 ;
        RECT 99.385 126.475 99.555 127.255 ;
        RECT 99.725 127.155 99.895 127.495 ;
        RECT 100.130 127.325 100.460 127.755 ;
        RECT 100.630 127.155 100.800 127.495 ;
        RECT 101.095 127.295 101.465 127.755 ;
        RECT 99.725 126.985 100.800 127.155 ;
        RECT 101.635 127.125 101.805 127.585 ;
        RECT 102.040 127.245 102.910 127.585 ;
        RECT 103.080 127.295 103.330 127.755 ;
        RECT 101.245 126.955 101.805 127.125 ;
        RECT 101.245 126.815 101.415 126.955 ;
        RECT 99.915 126.645 101.415 126.815 ;
        RECT 102.110 126.785 102.570 127.075 ;
        RECT 99.385 126.305 101.075 126.475 ;
        RECT 99.045 125.885 99.400 126.105 ;
        RECT 99.570 125.595 99.740 126.305 ;
        RECT 99.945 125.885 100.735 126.135 ;
        RECT 100.905 126.125 101.075 126.305 ;
        RECT 101.245 125.955 101.415 126.645 ;
        RECT 97.685 125.205 98.015 125.565 ;
        RECT 98.185 125.425 98.680 125.595 ;
        RECT 98.885 125.425 99.740 125.595 ;
        RECT 100.615 125.205 100.945 125.665 ;
        RECT 101.155 125.565 101.415 125.955 ;
        RECT 101.605 126.775 102.570 126.785 ;
        RECT 102.740 126.865 102.910 127.245 ;
        RECT 103.500 127.205 103.670 127.495 ;
        RECT 103.850 127.375 104.180 127.755 ;
        RECT 103.500 127.035 104.300 127.205 ;
        RECT 101.605 126.615 102.280 126.775 ;
        RECT 102.740 126.695 103.960 126.865 ;
        RECT 101.605 125.825 101.815 126.615 ;
        RECT 102.740 126.605 102.910 126.695 ;
        RECT 101.985 125.825 102.335 126.445 ;
        RECT 102.505 126.435 102.910 126.605 ;
        RECT 102.505 125.655 102.675 126.435 ;
        RECT 102.845 125.985 103.065 126.265 ;
        RECT 103.245 126.155 103.785 126.525 ;
        RECT 104.130 126.415 104.300 127.035 ;
        RECT 104.475 126.695 104.645 127.755 ;
        RECT 104.855 126.745 105.145 127.585 ;
        RECT 105.315 126.915 105.485 127.755 ;
        RECT 105.695 126.745 105.945 127.585 ;
        RECT 106.155 126.915 106.325 127.755 ;
        RECT 106.810 127.085 107.065 127.585 ;
        RECT 107.235 127.255 107.565 127.755 ;
        RECT 106.810 126.915 107.560 127.085 ;
        RECT 104.855 126.575 106.580 126.745 ;
        RECT 102.845 125.815 103.375 125.985 ;
        RECT 101.155 125.395 101.505 125.565 ;
        RECT 101.725 125.375 102.675 125.655 ;
        RECT 102.845 125.205 103.035 125.645 ;
        RECT 103.205 125.585 103.375 125.815 ;
        RECT 103.545 125.755 103.785 126.155 ;
        RECT 103.955 126.405 104.300 126.415 ;
        RECT 103.955 126.195 105.985 126.405 ;
        RECT 103.955 125.940 104.280 126.195 ;
        RECT 106.170 126.025 106.580 126.575 ;
        RECT 106.810 126.095 107.160 126.745 ;
        RECT 103.955 125.585 104.275 125.940 ;
        RECT 103.205 125.415 104.275 125.585 ;
        RECT 104.475 125.205 104.645 126.015 ;
        RECT 104.815 125.855 106.580 126.025 ;
        RECT 107.330 125.925 107.560 126.915 ;
        RECT 104.815 125.375 105.145 125.855 ;
        RECT 105.315 125.205 105.485 125.675 ;
        RECT 105.655 125.375 105.985 125.855 ;
        RECT 106.810 125.755 107.560 125.925 ;
        RECT 106.155 125.205 106.325 125.675 ;
        RECT 106.810 125.465 107.065 125.755 ;
        RECT 107.235 125.205 107.565 125.585 ;
        RECT 107.735 125.465 107.905 127.585 ;
        RECT 108.075 126.785 108.400 127.570 ;
        RECT 108.570 127.295 108.820 127.755 ;
        RECT 108.990 127.255 109.240 127.585 ;
        RECT 109.455 127.255 110.135 127.585 ;
        RECT 108.990 127.125 109.160 127.255 ;
        RECT 108.765 126.955 109.160 127.125 ;
        RECT 108.135 125.735 108.595 126.785 ;
        RECT 108.765 125.595 108.935 126.955 ;
        RECT 109.330 126.695 109.795 127.085 ;
        RECT 109.105 125.885 109.455 126.505 ;
        RECT 109.625 126.105 109.795 126.695 ;
        RECT 109.965 126.475 110.135 127.255 ;
        RECT 110.305 127.155 110.475 127.495 ;
        RECT 110.710 127.325 111.040 127.755 ;
        RECT 111.210 127.155 111.380 127.495 ;
        RECT 111.675 127.295 112.045 127.755 ;
        RECT 110.305 126.985 111.380 127.155 ;
        RECT 112.215 127.125 112.385 127.585 ;
        RECT 112.620 127.245 113.490 127.585 ;
        RECT 113.660 127.295 113.910 127.755 ;
        RECT 111.825 126.955 112.385 127.125 ;
        RECT 111.825 126.815 111.995 126.955 ;
        RECT 110.495 126.645 111.995 126.815 ;
        RECT 112.690 126.785 113.150 127.075 ;
        RECT 109.965 126.305 111.655 126.475 ;
        RECT 109.625 125.885 109.980 126.105 ;
        RECT 110.150 125.595 110.320 126.305 ;
        RECT 110.525 125.885 111.315 126.135 ;
        RECT 111.485 126.125 111.655 126.305 ;
        RECT 111.825 125.955 111.995 126.645 ;
        RECT 108.265 125.205 108.595 125.565 ;
        RECT 108.765 125.425 109.260 125.595 ;
        RECT 109.465 125.425 110.320 125.595 ;
        RECT 111.195 125.205 111.525 125.665 ;
        RECT 111.735 125.565 111.995 125.955 ;
        RECT 112.185 126.775 113.150 126.785 ;
        RECT 113.320 126.865 113.490 127.245 ;
        RECT 114.080 127.205 114.250 127.495 ;
        RECT 114.430 127.375 114.760 127.755 ;
        RECT 114.080 127.035 114.880 127.205 ;
        RECT 112.185 126.615 112.860 126.775 ;
        RECT 113.320 126.695 114.540 126.865 ;
        RECT 112.185 125.825 112.395 126.615 ;
        RECT 113.320 126.605 113.490 126.695 ;
        RECT 112.565 125.825 112.915 126.445 ;
        RECT 113.085 126.435 113.490 126.605 ;
        RECT 113.085 125.655 113.255 126.435 ;
        RECT 113.425 125.985 113.645 126.265 ;
        RECT 113.825 126.155 114.365 126.525 ;
        RECT 114.710 126.415 114.880 127.035 ;
        RECT 115.055 126.695 115.225 127.755 ;
        RECT 115.435 126.745 115.725 127.585 ;
        RECT 115.895 126.915 116.065 127.755 ;
        RECT 116.275 126.745 116.525 127.585 ;
        RECT 116.735 126.915 116.905 127.755 ;
        RECT 115.435 126.575 117.160 126.745 ;
        RECT 117.385 126.665 120.895 127.755 ;
        RECT 113.425 125.815 113.955 125.985 ;
        RECT 111.735 125.395 112.085 125.565 ;
        RECT 112.305 125.375 113.255 125.655 ;
        RECT 113.425 125.205 113.615 125.645 ;
        RECT 113.785 125.585 113.955 125.815 ;
        RECT 114.125 125.755 114.365 126.155 ;
        RECT 114.535 126.405 114.880 126.415 ;
        RECT 114.535 126.195 116.565 126.405 ;
        RECT 114.535 125.940 114.860 126.195 ;
        RECT 116.750 126.025 117.160 126.575 ;
        RECT 114.535 125.585 114.855 125.940 ;
        RECT 113.785 125.415 114.855 125.585 ;
        RECT 115.055 125.205 115.225 126.015 ;
        RECT 115.395 125.855 117.160 126.025 ;
        RECT 117.385 125.975 119.035 126.495 ;
        RECT 119.205 126.145 120.895 126.665 ;
        RECT 121.525 126.590 121.815 127.755 ;
        RECT 121.985 126.665 123.655 127.755 ;
        RECT 121.985 125.975 122.735 126.495 ;
        RECT 122.905 126.145 123.655 126.665 ;
        RECT 124.285 126.665 125.495 127.755 ;
        RECT 124.285 126.125 124.805 126.665 ;
        RECT 115.395 125.375 115.725 125.855 ;
        RECT 115.895 125.205 116.065 125.675 ;
        RECT 116.235 125.375 116.565 125.855 ;
        RECT 116.735 125.205 116.905 125.675 ;
        RECT 117.385 125.205 120.895 125.975 ;
        RECT 121.525 125.205 121.815 125.930 ;
        RECT 121.985 125.205 123.655 125.975 ;
        RECT 124.975 125.955 125.495 126.495 ;
        RECT 124.285 125.205 125.495 125.955 ;
        RECT 5.520 125.035 125.580 125.205 ;
        RECT 5.605 124.285 6.815 125.035 ;
        RECT 7.295 124.565 7.465 125.035 ;
        RECT 7.635 124.385 7.965 124.865 ;
        RECT 8.135 124.565 8.305 125.035 ;
        RECT 8.475 124.385 8.805 124.865 ;
        RECT 5.605 123.745 6.125 124.285 ;
        RECT 7.040 124.215 8.805 124.385 ;
        RECT 8.975 124.225 9.145 125.035 ;
        RECT 9.345 124.655 10.415 124.825 ;
        RECT 9.345 124.300 9.665 124.655 ;
        RECT 6.295 123.575 6.815 124.115 ;
        RECT 5.605 122.485 6.815 123.575 ;
        RECT 7.040 123.665 7.450 124.215 ;
        RECT 9.340 124.045 9.665 124.300 ;
        RECT 7.635 123.835 9.665 124.045 ;
        RECT 9.320 123.825 9.665 123.835 ;
        RECT 9.835 124.085 10.075 124.485 ;
        RECT 10.245 124.425 10.415 124.655 ;
        RECT 10.585 124.595 10.775 125.035 ;
        RECT 10.945 124.585 11.895 124.865 ;
        RECT 12.115 124.675 12.465 124.845 ;
        RECT 10.245 124.255 10.775 124.425 ;
        RECT 7.040 123.495 8.765 123.665 ;
        RECT 7.295 122.485 7.465 123.325 ;
        RECT 7.675 122.655 7.925 123.495 ;
        RECT 8.135 122.485 8.305 123.325 ;
        RECT 8.475 122.655 8.765 123.495 ;
        RECT 8.975 122.485 9.145 123.545 ;
        RECT 9.320 123.205 9.490 123.825 ;
        RECT 9.835 123.715 10.375 124.085 ;
        RECT 10.555 123.975 10.775 124.255 ;
        RECT 10.945 123.805 11.115 124.585 ;
        RECT 10.710 123.635 11.115 123.805 ;
        RECT 11.285 123.795 11.635 124.415 ;
        RECT 10.710 123.545 10.880 123.635 ;
        RECT 11.805 123.625 12.015 124.415 ;
        RECT 9.660 123.375 10.880 123.545 ;
        RECT 11.340 123.465 12.015 123.625 ;
        RECT 9.320 123.035 10.120 123.205 ;
        RECT 9.440 122.485 9.770 122.865 ;
        RECT 9.950 122.745 10.120 123.035 ;
        RECT 10.710 122.995 10.880 123.375 ;
        RECT 11.050 123.455 12.015 123.465 ;
        RECT 12.205 124.285 12.465 124.675 ;
        RECT 12.675 124.575 13.005 125.035 ;
        RECT 13.880 124.645 14.735 124.815 ;
        RECT 14.940 124.645 15.435 124.815 ;
        RECT 15.605 124.675 15.935 125.035 ;
        RECT 12.205 123.595 12.375 124.285 ;
        RECT 12.545 123.935 12.715 124.115 ;
        RECT 12.885 124.105 13.675 124.355 ;
        RECT 13.880 123.935 14.050 124.645 ;
        RECT 14.220 124.135 14.575 124.355 ;
        RECT 12.545 123.765 14.235 123.935 ;
        RECT 11.050 123.165 11.510 123.455 ;
        RECT 12.205 123.425 13.705 123.595 ;
        RECT 12.205 123.285 12.375 123.425 ;
        RECT 11.815 123.115 12.375 123.285 ;
        RECT 10.290 122.485 10.540 122.945 ;
        RECT 10.710 122.655 11.580 122.995 ;
        RECT 11.815 122.655 11.985 123.115 ;
        RECT 12.820 123.085 13.895 123.255 ;
        RECT 12.155 122.485 12.525 122.945 ;
        RECT 12.820 122.745 12.990 123.085 ;
        RECT 13.160 122.485 13.490 122.915 ;
        RECT 13.725 122.745 13.895 123.085 ;
        RECT 14.065 122.985 14.235 123.765 ;
        RECT 14.405 123.545 14.575 124.135 ;
        RECT 14.745 123.735 15.095 124.355 ;
        RECT 14.405 123.155 14.870 123.545 ;
        RECT 15.265 123.285 15.435 124.645 ;
        RECT 15.605 123.455 16.065 124.505 ;
        RECT 15.040 123.115 15.435 123.285 ;
        RECT 15.040 122.985 15.210 123.115 ;
        RECT 14.065 122.655 14.745 122.985 ;
        RECT 14.960 122.655 15.210 122.985 ;
        RECT 15.380 122.485 15.630 122.945 ;
        RECT 15.800 122.670 16.125 123.455 ;
        RECT 16.295 122.655 16.465 124.775 ;
        RECT 16.635 124.655 16.965 125.035 ;
        RECT 17.135 124.485 17.390 124.775 ;
        RECT 16.640 124.315 17.390 124.485 ;
        RECT 16.640 123.325 16.870 124.315 ;
        RECT 17.625 124.215 17.835 125.035 ;
        RECT 18.005 124.235 18.335 124.865 ;
        RECT 17.040 123.495 17.390 124.145 ;
        RECT 18.005 123.635 18.255 124.235 ;
        RECT 18.505 124.215 18.735 125.035 ;
        RECT 19.410 124.485 19.665 124.775 ;
        RECT 19.835 124.655 20.165 125.035 ;
        RECT 19.410 124.315 20.160 124.485 ;
        RECT 18.425 123.795 18.755 124.045 ;
        RECT 16.640 123.155 17.390 123.325 ;
        RECT 16.635 122.485 16.965 122.985 ;
        RECT 17.135 122.655 17.390 123.155 ;
        RECT 17.625 122.485 17.835 123.625 ;
        RECT 18.005 122.655 18.335 123.635 ;
        RECT 18.505 122.485 18.735 123.625 ;
        RECT 19.410 123.495 19.760 124.145 ;
        RECT 19.930 123.325 20.160 124.315 ;
        RECT 19.410 123.155 20.160 123.325 ;
        RECT 19.410 122.655 19.665 123.155 ;
        RECT 19.835 122.485 20.165 122.985 ;
        RECT 20.335 122.655 20.505 124.775 ;
        RECT 20.865 124.675 21.195 125.035 ;
        RECT 21.365 124.645 21.860 124.815 ;
        RECT 22.065 124.645 22.920 124.815 ;
        RECT 20.735 123.455 21.195 124.505 ;
        RECT 20.675 122.670 21.000 123.455 ;
        RECT 21.365 123.285 21.535 124.645 ;
        RECT 21.705 123.735 22.055 124.355 ;
        RECT 22.225 124.135 22.580 124.355 ;
        RECT 22.225 123.545 22.395 124.135 ;
        RECT 22.750 123.935 22.920 124.645 ;
        RECT 23.795 124.575 24.125 125.035 ;
        RECT 24.335 124.675 24.685 124.845 ;
        RECT 23.125 124.105 23.915 124.355 ;
        RECT 24.335 124.285 24.595 124.675 ;
        RECT 24.905 124.585 25.855 124.865 ;
        RECT 26.025 124.595 26.215 125.035 ;
        RECT 26.385 124.655 27.455 124.825 ;
        RECT 24.085 123.935 24.255 124.115 ;
        RECT 21.365 123.115 21.760 123.285 ;
        RECT 21.930 123.155 22.395 123.545 ;
        RECT 22.565 123.765 24.255 123.935 ;
        RECT 21.590 122.985 21.760 123.115 ;
        RECT 22.565 122.985 22.735 123.765 ;
        RECT 24.425 123.595 24.595 124.285 ;
        RECT 23.095 123.425 24.595 123.595 ;
        RECT 24.785 123.625 24.995 124.415 ;
        RECT 25.165 123.795 25.515 124.415 ;
        RECT 25.685 123.805 25.855 124.585 ;
        RECT 26.385 124.425 26.555 124.655 ;
        RECT 26.025 124.255 26.555 124.425 ;
        RECT 26.025 123.975 26.245 124.255 ;
        RECT 26.725 124.085 26.965 124.485 ;
        RECT 25.685 123.635 26.090 123.805 ;
        RECT 26.425 123.715 26.965 124.085 ;
        RECT 27.135 124.300 27.455 124.655 ;
        RECT 27.135 124.045 27.460 124.300 ;
        RECT 27.655 124.225 27.825 125.035 ;
        RECT 27.995 124.385 28.325 124.865 ;
        RECT 28.495 124.565 28.665 125.035 ;
        RECT 28.835 124.385 29.165 124.865 ;
        RECT 29.335 124.565 29.505 125.035 ;
        RECT 27.995 124.215 29.760 124.385 ;
        RECT 30.045 124.215 30.255 125.035 ;
        RECT 30.425 124.235 30.755 124.865 ;
        RECT 27.135 123.835 29.165 124.045 ;
        RECT 27.135 123.825 27.480 123.835 ;
        RECT 24.785 123.465 25.460 123.625 ;
        RECT 25.920 123.545 26.090 123.635 ;
        RECT 24.785 123.455 25.750 123.465 ;
        RECT 24.425 123.285 24.595 123.425 ;
        RECT 21.170 122.485 21.420 122.945 ;
        RECT 21.590 122.655 21.840 122.985 ;
        RECT 22.055 122.655 22.735 122.985 ;
        RECT 22.905 123.085 23.980 123.255 ;
        RECT 24.425 123.115 24.985 123.285 ;
        RECT 25.290 123.165 25.750 123.455 ;
        RECT 25.920 123.375 27.140 123.545 ;
        RECT 22.905 122.745 23.075 123.085 ;
        RECT 23.310 122.485 23.640 122.915 ;
        RECT 23.810 122.745 23.980 123.085 ;
        RECT 24.275 122.485 24.645 122.945 ;
        RECT 24.815 122.655 24.985 123.115 ;
        RECT 25.920 122.995 26.090 123.375 ;
        RECT 27.310 123.205 27.480 123.825 ;
        RECT 29.350 123.665 29.760 124.215 ;
        RECT 25.220 122.655 26.090 122.995 ;
        RECT 26.680 123.035 27.480 123.205 ;
        RECT 26.260 122.485 26.510 122.945 ;
        RECT 26.680 122.745 26.850 123.035 ;
        RECT 27.030 122.485 27.360 122.865 ;
        RECT 27.655 122.485 27.825 123.545 ;
        RECT 28.035 123.495 29.760 123.665 ;
        RECT 30.425 123.635 30.675 124.235 ;
        RECT 30.925 124.215 31.155 125.035 ;
        RECT 31.365 124.310 31.655 125.035 ;
        RECT 31.825 124.265 35.335 125.035 ;
        RECT 30.845 123.795 31.175 124.045 ;
        RECT 31.825 123.745 33.475 124.265 ;
        RECT 35.545 124.215 35.775 125.035 ;
        RECT 35.945 124.235 36.275 124.865 ;
        RECT 28.035 122.655 28.325 123.495 ;
        RECT 28.495 122.485 28.665 123.325 ;
        RECT 28.875 122.655 29.125 123.495 ;
        RECT 29.335 122.485 29.505 123.325 ;
        RECT 30.045 122.485 30.255 123.625 ;
        RECT 30.425 122.655 30.755 123.635 ;
        RECT 30.925 122.485 31.155 123.625 ;
        RECT 31.365 122.485 31.655 123.650 ;
        RECT 33.645 123.575 35.335 124.095 ;
        RECT 35.525 123.795 35.855 124.045 ;
        RECT 36.025 123.635 36.275 124.235 ;
        RECT 36.445 124.215 36.655 125.035 ;
        RECT 36.885 124.265 39.475 125.035 ;
        RECT 36.885 123.745 38.095 124.265 ;
        RECT 40.165 124.215 40.375 125.035 ;
        RECT 40.545 124.235 40.875 124.865 ;
        RECT 31.825 122.485 35.335 123.575 ;
        RECT 35.545 122.485 35.775 123.625 ;
        RECT 35.945 122.655 36.275 123.635 ;
        RECT 36.445 122.485 36.655 123.625 ;
        RECT 38.265 123.575 39.475 124.095 ;
        RECT 40.545 123.635 40.795 124.235 ;
        RECT 41.045 124.215 41.275 125.035 ;
        RECT 41.490 124.485 41.745 124.775 ;
        RECT 41.915 124.655 42.245 125.035 ;
        RECT 41.490 124.315 42.240 124.485 ;
        RECT 40.965 123.795 41.295 124.045 ;
        RECT 36.885 122.485 39.475 123.575 ;
        RECT 40.165 122.485 40.375 123.625 ;
        RECT 40.545 122.655 40.875 123.635 ;
        RECT 41.045 122.485 41.275 123.625 ;
        RECT 41.490 123.495 41.840 124.145 ;
        RECT 42.010 123.325 42.240 124.315 ;
        RECT 41.490 123.155 42.240 123.325 ;
        RECT 41.490 122.655 41.745 123.155 ;
        RECT 41.915 122.485 42.245 122.985 ;
        RECT 42.415 122.655 42.585 124.775 ;
        RECT 42.945 124.675 43.275 125.035 ;
        RECT 43.445 124.645 43.940 124.815 ;
        RECT 44.145 124.645 45.000 124.815 ;
        RECT 42.815 123.455 43.275 124.505 ;
        RECT 42.755 122.670 43.080 123.455 ;
        RECT 43.445 123.285 43.615 124.645 ;
        RECT 43.785 123.735 44.135 124.355 ;
        RECT 44.305 124.135 44.660 124.355 ;
        RECT 44.305 123.545 44.475 124.135 ;
        RECT 44.830 123.935 45.000 124.645 ;
        RECT 45.875 124.575 46.205 125.035 ;
        RECT 46.415 124.675 46.765 124.845 ;
        RECT 45.205 124.105 45.995 124.355 ;
        RECT 46.415 124.285 46.675 124.675 ;
        RECT 46.985 124.585 47.935 124.865 ;
        RECT 48.105 124.595 48.295 125.035 ;
        RECT 48.465 124.655 49.535 124.825 ;
        RECT 46.165 123.935 46.335 124.115 ;
        RECT 43.445 123.115 43.840 123.285 ;
        RECT 44.010 123.155 44.475 123.545 ;
        RECT 44.645 123.765 46.335 123.935 ;
        RECT 43.670 122.985 43.840 123.115 ;
        RECT 44.645 122.985 44.815 123.765 ;
        RECT 46.505 123.595 46.675 124.285 ;
        RECT 45.175 123.425 46.675 123.595 ;
        RECT 46.865 123.625 47.075 124.415 ;
        RECT 47.245 123.795 47.595 124.415 ;
        RECT 47.765 123.805 47.935 124.585 ;
        RECT 48.465 124.425 48.635 124.655 ;
        RECT 48.105 124.255 48.635 124.425 ;
        RECT 48.105 123.975 48.325 124.255 ;
        RECT 48.805 124.085 49.045 124.485 ;
        RECT 47.765 123.635 48.170 123.805 ;
        RECT 48.505 123.715 49.045 124.085 ;
        RECT 49.215 124.300 49.535 124.655 ;
        RECT 49.215 124.045 49.540 124.300 ;
        RECT 49.735 124.225 49.905 125.035 ;
        RECT 50.075 124.385 50.405 124.865 ;
        RECT 50.575 124.565 50.745 125.035 ;
        RECT 50.915 124.385 51.245 124.865 ;
        RECT 51.415 124.565 51.585 125.035 ;
        RECT 50.075 124.215 51.840 124.385 ;
        RECT 49.215 123.835 51.245 124.045 ;
        RECT 49.215 123.825 49.560 123.835 ;
        RECT 46.865 123.465 47.540 123.625 ;
        RECT 48.000 123.545 48.170 123.635 ;
        RECT 46.865 123.455 47.830 123.465 ;
        RECT 46.505 123.285 46.675 123.425 ;
        RECT 43.250 122.485 43.500 122.945 ;
        RECT 43.670 122.655 43.920 122.985 ;
        RECT 44.135 122.655 44.815 122.985 ;
        RECT 44.985 123.085 46.060 123.255 ;
        RECT 46.505 123.115 47.065 123.285 ;
        RECT 47.370 123.165 47.830 123.455 ;
        RECT 48.000 123.375 49.220 123.545 ;
        RECT 44.985 122.745 45.155 123.085 ;
        RECT 45.390 122.485 45.720 122.915 ;
        RECT 45.890 122.745 46.060 123.085 ;
        RECT 46.355 122.485 46.725 122.945 ;
        RECT 46.895 122.655 47.065 123.115 ;
        RECT 48.000 122.995 48.170 123.375 ;
        RECT 49.390 123.205 49.560 123.825 ;
        RECT 51.430 123.665 51.840 124.215 ;
        RECT 52.065 124.285 53.275 125.035 ;
        RECT 52.065 123.745 52.585 124.285 ;
        RECT 53.485 124.215 53.715 125.035 ;
        RECT 53.885 124.235 54.215 124.865 ;
        RECT 47.300 122.655 48.170 122.995 ;
        RECT 48.760 123.035 49.560 123.205 ;
        RECT 48.340 122.485 48.590 122.945 ;
        RECT 48.760 122.745 48.930 123.035 ;
        RECT 49.110 122.485 49.440 122.865 ;
        RECT 49.735 122.485 49.905 123.545 ;
        RECT 50.115 123.495 51.840 123.665 ;
        RECT 52.755 123.575 53.275 124.115 ;
        RECT 53.465 123.795 53.795 124.045 ;
        RECT 53.965 123.635 54.215 124.235 ;
        RECT 54.385 124.215 54.595 125.035 ;
        RECT 54.825 124.360 55.085 124.865 ;
        RECT 55.265 124.655 55.595 125.035 ;
        RECT 55.775 124.485 55.945 124.865 ;
        RECT 50.115 122.655 50.405 123.495 ;
        RECT 50.575 122.485 50.745 123.325 ;
        RECT 50.955 122.655 51.205 123.495 ;
        RECT 51.415 122.485 51.585 123.325 ;
        RECT 52.065 122.485 53.275 123.575 ;
        RECT 53.485 122.485 53.715 123.625 ;
        RECT 53.885 122.655 54.215 123.635 ;
        RECT 54.385 122.485 54.595 123.625 ;
        RECT 54.825 123.560 54.995 124.360 ;
        RECT 55.280 124.315 55.945 124.485 ;
        RECT 55.280 124.060 55.450 124.315 ;
        RECT 57.125 124.310 57.415 125.035 ;
        RECT 58.135 124.485 58.305 124.865 ;
        RECT 58.485 124.655 58.815 125.035 ;
        RECT 58.135 124.315 58.800 124.485 ;
        RECT 58.995 124.360 59.255 124.865 ;
        RECT 55.165 123.730 55.450 124.060 ;
        RECT 55.685 123.765 56.015 124.135 ;
        RECT 58.065 123.765 58.395 124.135 ;
        RECT 58.630 124.060 58.800 124.315 ;
        RECT 55.280 123.585 55.450 123.730 ;
        RECT 58.630 123.730 58.915 124.060 ;
        RECT 54.825 122.655 55.095 123.560 ;
        RECT 55.280 123.415 55.945 123.585 ;
        RECT 55.265 122.485 55.595 123.245 ;
        RECT 55.775 122.655 55.945 123.415 ;
        RECT 57.125 122.485 57.415 123.650 ;
        RECT 58.630 123.585 58.800 123.730 ;
        RECT 58.135 123.415 58.800 123.585 ;
        RECT 59.085 123.560 59.255 124.360 ;
        RECT 59.465 124.215 59.695 125.035 ;
        RECT 59.865 124.235 60.195 124.865 ;
        RECT 59.445 123.795 59.775 124.045 ;
        RECT 59.945 123.635 60.195 124.235 ;
        RECT 60.365 124.215 60.575 125.035 ;
        RECT 60.805 124.490 66.150 125.035 ;
        RECT 62.390 123.660 62.730 124.490 ;
        RECT 66.325 124.285 67.535 125.035 ;
        RECT 67.710 124.485 67.965 124.775 ;
        RECT 68.135 124.655 68.465 125.035 ;
        RECT 67.710 124.315 68.460 124.485 ;
        RECT 58.135 122.655 58.305 123.415 ;
        RECT 58.485 122.485 58.815 123.245 ;
        RECT 58.985 122.655 59.255 123.560 ;
        RECT 59.465 122.485 59.695 123.625 ;
        RECT 59.865 122.655 60.195 123.635 ;
        RECT 60.365 122.485 60.575 123.625 ;
        RECT 64.210 122.920 64.560 124.170 ;
        RECT 66.325 123.745 66.845 124.285 ;
        RECT 67.015 123.575 67.535 124.115 ;
        RECT 60.805 122.485 66.150 122.920 ;
        RECT 66.325 122.485 67.535 123.575 ;
        RECT 67.710 123.495 68.060 124.145 ;
        RECT 68.230 123.325 68.460 124.315 ;
        RECT 67.710 123.155 68.460 123.325 ;
        RECT 67.710 122.655 67.965 123.155 ;
        RECT 68.135 122.485 68.465 122.985 ;
        RECT 68.635 122.655 68.805 124.775 ;
        RECT 69.165 124.675 69.495 125.035 ;
        RECT 69.665 124.645 70.160 124.815 ;
        RECT 70.365 124.645 71.220 124.815 ;
        RECT 69.035 123.455 69.495 124.505 ;
        RECT 68.975 122.670 69.300 123.455 ;
        RECT 69.665 123.285 69.835 124.645 ;
        RECT 70.005 123.735 70.355 124.355 ;
        RECT 70.525 124.135 70.880 124.355 ;
        RECT 70.525 123.545 70.695 124.135 ;
        RECT 71.050 123.935 71.220 124.645 ;
        RECT 72.095 124.575 72.425 125.035 ;
        RECT 72.635 124.675 72.985 124.845 ;
        RECT 71.425 124.105 72.215 124.355 ;
        RECT 72.635 124.285 72.895 124.675 ;
        RECT 73.205 124.585 74.155 124.865 ;
        RECT 74.325 124.595 74.515 125.035 ;
        RECT 74.685 124.655 75.755 124.825 ;
        RECT 72.385 123.935 72.555 124.115 ;
        RECT 69.665 123.115 70.060 123.285 ;
        RECT 70.230 123.155 70.695 123.545 ;
        RECT 70.865 123.765 72.555 123.935 ;
        RECT 69.890 122.985 70.060 123.115 ;
        RECT 70.865 122.985 71.035 123.765 ;
        RECT 72.725 123.595 72.895 124.285 ;
        RECT 71.395 123.425 72.895 123.595 ;
        RECT 73.085 123.625 73.295 124.415 ;
        RECT 73.465 123.795 73.815 124.415 ;
        RECT 73.985 123.805 74.155 124.585 ;
        RECT 74.685 124.425 74.855 124.655 ;
        RECT 74.325 124.255 74.855 124.425 ;
        RECT 74.325 123.975 74.545 124.255 ;
        RECT 75.025 124.085 75.265 124.485 ;
        RECT 73.985 123.635 74.390 123.805 ;
        RECT 74.725 123.715 75.265 124.085 ;
        RECT 75.435 124.300 75.755 124.655 ;
        RECT 75.435 124.045 75.760 124.300 ;
        RECT 75.955 124.225 76.125 125.035 ;
        RECT 76.295 124.385 76.625 124.865 ;
        RECT 76.795 124.565 76.965 125.035 ;
        RECT 77.135 124.385 77.465 124.865 ;
        RECT 77.635 124.565 77.805 125.035 ;
        RECT 76.295 124.215 78.060 124.385 ;
        RECT 78.345 124.215 78.555 125.035 ;
        RECT 78.725 124.235 79.055 124.865 ;
        RECT 75.435 123.835 77.465 124.045 ;
        RECT 75.435 123.825 75.780 123.835 ;
        RECT 73.085 123.465 73.760 123.625 ;
        RECT 74.220 123.545 74.390 123.635 ;
        RECT 73.085 123.455 74.050 123.465 ;
        RECT 72.725 123.285 72.895 123.425 ;
        RECT 69.470 122.485 69.720 122.945 ;
        RECT 69.890 122.655 70.140 122.985 ;
        RECT 70.355 122.655 71.035 122.985 ;
        RECT 71.205 123.085 72.280 123.255 ;
        RECT 72.725 123.115 73.285 123.285 ;
        RECT 73.590 123.165 74.050 123.455 ;
        RECT 74.220 123.375 75.440 123.545 ;
        RECT 71.205 122.745 71.375 123.085 ;
        RECT 71.610 122.485 71.940 122.915 ;
        RECT 72.110 122.745 72.280 123.085 ;
        RECT 72.575 122.485 72.945 122.945 ;
        RECT 73.115 122.655 73.285 123.115 ;
        RECT 74.220 122.995 74.390 123.375 ;
        RECT 75.610 123.205 75.780 123.825 ;
        RECT 77.650 123.665 78.060 124.215 ;
        RECT 73.520 122.655 74.390 122.995 ;
        RECT 74.980 123.035 75.780 123.205 ;
        RECT 74.560 122.485 74.810 122.945 ;
        RECT 74.980 122.745 75.150 123.035 ;
        RECT 75.330 122.485 75.660 122.865 ;
        RECT 75.955 122.485 76.125 123.545 ;
        RECT 76.335 123.495 78.060 123.665 ;
        RECT 78.725 123.635 78.975 124.235 ;
        RECT 79.225 124.215 79.455 125.035 ;
        RECT 79.725 124.215 79.935 125.035 ;
        RECT 80.105 124.235 80.435 124.865 ;
        RECT 79.145 123.795 79.475 124.045 ;
        RECT 80.105 123.635 80.355 124.235 ;
        RECT 80.605 124.215 80.835 125.035 ;
        RECT 81.045 124.265 82.715 125.035 ;
        RECT 82.885 124.310 83.175 125.035 ;
        RECT 83.345 124.265 85.015 125.035 ;
        RECT 80.525 123.795 80.855 124.045 ;
        RECT 81.045 123.745 81.795 124.265 ;
        RECT 76.335 122.655 76.625 123.495 ;
        RECT 76.795 122.485 76.965 123.325 ;
        RECT 77.175 122.655 77.425 123.495 ;
        RECT 77.635 122.485 77.805 123.325 ;
        RECT 78.345 122.485 78.555 123.625 ;
        RECT 78.725 122.655 79.055 123.635 ;
        RECT 79.225 122.485 79.455 123.625 ;
        RECT 79.725 122.485 79.935 123.625 ;
        RECT 80.105 122.655 80.435 123.635 ;
        RECT 80.605 122.485 80.835 123.625 ;
        RECT 81.965 123.575 82.715 124.095 ;
        RECT 83.345 123.745 84.095 124.265 ;
        RECT 85.225 124.215 85.455 125.035 ;
        RECT 85.625 124.235 85.955 124.865 ;
        RECT 81.045 122.485 82.715 123.575 ;
        RECT 82.885 122.485 83.175 123.650 ;
        RECT 84.265 123.575 85.015 124.095 ;
        RECT 85.205 123.795 85.535 124.045 ;
        RECT 85.705 123.635 85.955 124.235 ;
        RECT 86.125 124.215 86.335 125.035 ;
        RECT 87.030 124.485 87.285 124.775 ;
        RECT 87.455 124.655 87.785 125.035 ;
        RECT 87.030 124.315 87.780 124.485 ;
        RECT 83.345 122.485 85.015 123.575 ;
        RECT 85.225 122.485 85.455 123.625 ;
        RECT 85.625 122.655 85.955 123.635 ;
        RECT 86.125 122.485 86.335 123.625 ;
        RECT 87.030 123.495 87.380 124.145 ;
        RECT 87.550 123.325 87.780 124.315 ;
        RECT 87.030 123.155 87.780 123.325 ;
        RECT 87.030 122.655 87.285 123.155 ;
        RECT 87.455 122.485 87.785 122.985 ;
        RECT 87.955 122.655 88.125 124.775 ;
        RECT 88.485 124.675 88.815 125.035 ;
        RECT 88.985 124.645 89.480 124.815 ;
        RECT 89.685 124.645 90.540 124.815 ;
        RECT 88.355 123.455 88.815 124.505 ;
        RECT 88.295 122.670 88.620 123.455 ;
        RECT 88.985 123.285 89.155 124.645 ;
        RECT 89.325 123.735 89.675 124.355 ;
        RECT 89.845 124.135 90.200 124.355 ;
        RECT 89.845 123.545 90.015 124.135 ;
        RECT 90.370 123.935 90.540 124.645 ;
        RECT 91.415 124.575 91.745 125.035 ;
        RECT 91.955 124.675 92.305 124.845 ;
        RECT 90.745 124.105 91.535 124.355 ;
        RECT 91.955 124.285 92.215 124.675 ;
        RECT 92.525 124.585 93.475 124.865 ;
        RECT 93.645 124.595 93.835 125.035 ;
        RECT 94.005 124.655 95.075 124.825 ;
        RECT 91.705 123.935 91.875 124.115 ;
        RECT 88.985 123.115 89.380 123.285 ;
        RECT 89.550 123.155 90.015 123.545 ;
        RECT 90.185 123.765 91.875 123.935 ;
        RECT 89.210 122.985 89.380 123.115 ;
        RECT 90.185 122.985 90.355 123.765 ;
        RECT 92.045 123.595 92.215 124.285 ;
        RECT 90.715 123.425 92.215 123.595 ;
        RECT 92.405 123.625 92.615 124.415 ;
        RECT 92.785 123.795 93.135 124.415 ;
        RECT 93.305 123.805 93.475 124.585 ;
        RECT 94.005 124.425 94.175 124.655 ;
        RECT 93.645 124.255 94.175 124.425 ;
        RECT 93.645 123.975 93.865 124.255 ;
        RECT 94.345 124.085 94.585 124.485 ;
        RECT 93.305 123.635 93.710 123.805 ;
        RECT 94.045 123.715 94.585 124.085 ;
        RECT 94.755 124.300 95.075 124.655 ;
        RECT 94.755 124.045 95.080 124.300 ;
        RECT 95.275 124.225 95.445 125.035 ;
        RECT 95.615 124.385 95.945 124.865 ;
        RECT 96.115 124.565 96.285 125.035 ;
        RECT 96.455 124.385 96.785 124.865 ;
        RECT 96.955 124.565 97.125 125.035 ;
        RECT 95.615 124.215 97.380 124.385 ;
        RECT 97.645 124.215 97.875 125.035 ;
        RECT 98.045 124.235 98.375 124.865 ;
        RECT 94.755 123.835 96.785 124.045 ;
        RECT 94.755 123.825 95.100 123.835 ;
        RECT 92.405 123.465 93.080 123.625 ;
        RECT 93.540 123.545 93.710 123.635 ;
        RECT 92.405 123.455 93.370 123.465 ;
        RECT 92.045 123.285 92.215 123.425 ;
        RECT 88.790 122.485 89.040 122.945 ;
        RECT 89.210 122.655 89.460 122.985 ;
        RECT 89.675 122.655 90.355 122.985 ;
        RECT 90.525 123.085 91.600 123.255 ;
        RECT 92.045 123.115 92.605 123.285 ;
        RECT 92.910 123.165 93.370 123.455 ;
        RECT 93.540 123.375 94.760 123.545 ;
        RECT 90.525 122.745 90.695 123.085 ;
        RECT 90.930 122.485 91.260 122.915 ;
        RECT 91.430 122.745 91.600 123.085 ;
        RECT 91.895 122.485 92.265 122.945 ;
        RECT 92.435 122.655 92.605 123.115 ;
        RECT 93.540 122.995 93.710 123.375 ;
        RECT 94.930 123.205 95.100 123.825 ;
        RECT 96.970 123.665 97.380 124.215 ;
        RECT 97.625 123.795 97.955 124.045 ;
        RECT 92.840 122.655 93.710 122.995 ;
        RECT 94.300 123.035 95.100 123.205 ;
        RECT 93.880 122.485 94.130 122.945 ;
        RECT 94.300 122.745 94.470 123.035 ;
        RECT 94.650 122.485 94.980 122.865 ;
        RECT 95.275 122.485 95.445 123.545 ;
        RECT 95.655 123.495 97.380 123.665 ;
        RECT 98.125 123.635 98.375 124.235 ;
        RECT 98.545 124.215 98.755 125.035 ;
        RECT 98.985 124.490 104.330 125.035 ;
        RECT 100.570 123.660 100.910 124.490 ;
        RECT 105.005 124.215 105.235 125.035 ;
        RECT 105.405 124.235 105.735 124.865 ;
        RECT 95.655 122.655 95.945 123.495 ;
        RECT 96.115 122.485 96.285 123.325 ;
        RECT 96.495 122.655 96.745 123.495 ;
        RECT 96.955 122.485 97.125 123.325 ;
        RECT 97.645 122.485 97.875 123.625 ;
        RECT 98.045 122.655 98.375 123.635 ;
        RECT 98.545 122.485 98.755 123.625 ;
        RECT 102.390 122.920 102.740 124.170 ;
        RECT 104.985 123.795 105.315 124.045 ;
        RECT 105.485 123.635 105.735 124.235 ;
        RECT 105.905 124.215 106.115 125.035 ;
        RECT 107.305 124.215 107.535 125.035 ;
        RECT 107.705 124.235 108.035 124.865 ;
        RECT 107.285 123.795 107.615 124.045 ;
        RECT 107.785 123.635 108.035 124.235 ;
        RECT 108.205 124.215 108.415 125.035 ;
        RECT 108.645 124.310 108.935 125.035 ;
        RECT 109.110 124.485 109.365 124.775 ;
        RECT 109.535 124.655 109.865 125.035 ;
        RECT 109.110 124.315 109.860 124.485 ;
        RECT 98.985 122.485 104.330 122.920 ;
        RECT 105.005 122.485 105.235 123.625 ;
        RECT 105.405 122.655 105.735 123.635 ;
        RECT 105.905 122.485 106.115 123.625 ;
        RECT 107.305 122.485 107.535 123.625 ;
        RECT 107.705 122.655 108.035 123.635 ;
        RECT 108.205 122.485 108.415 123.625 ;
        RECT 108.645 122.485 108.935 123.650 ;
        RECT 109.110 123.495 109.460 124.145 ;
        RECT 109.630 123.325 109.860 124.315 ;
        RECT 109.110 123.155 109.860 123.325 ;
        RECT 109.110 122.655 109.365 123.155 ;
        RECT 109.535 122.485 109.865 122.985 ;
        RECT 110.035 122.655 110.205 124.775 ;
        RECT 110.565 124.675 110.895 125.035 ;
        RECT 111.065 124.645 111.560 124.815 ;
        RECT 111.765 124.645 112.620 124.815 ;
        RECT 110.435 123.455 110.895 124.505 ;
        RECT 110.375 122.670 110.700 123.455 ;
        RECT 111.065 123.285 111.235 124.645 ;
        RECT 111.405 123.735 111.755 124.355 ;
        RECT 111.925 124.135 112.280 124.355 ;
        RECT 111.925 123.545 112.095 124.135 ;
        RECT 112.450 123.935 112.620 124.645 ;
        RECT 113.495 124.575 113.825 125.035 ;
        RECT 114.035 124.675 114.385 124.845 ;
        RECT 112.825 124.105 113.615 124.355 ;
        RECT 114.035 124.285 114.295 124.675 ;
        RECT 114.605 124.585 115.555 124.865 ;
        RECT 115.725 124.595 115.915 125.035 ;
        RECT 116.085 124.655 117.155 124.825 ;
        RECT 113.785 123.935 113.955 124.115 ;
        RECT 111.065 123.115 111.460 123.285 ;
        RECT 111.630 123.155 112.095 123.545 ;
        RECT 112.265 123.765 113.955 123.935 ;
        RECT 111.290 122.985 111.460 123.115 ;
        RECT 112.265 122.985 112.435 123.765 ;
        RECT 114.125 123.595 114.295 124.285 ;
        RECT 112.795 123.425 114.295 123.595 ;
        RECT 114.485 123.625 114.695 124.415 ;
        RECT 114.865 123.795 115.215 124.415 ;
        RECT 115.385 123.805 115.555 124.585 ;
        RECT 116.085 124.425 116.255 124.655 ;
        RECT 115.725 124.255 116.255 124.425 ;
        RECT 115.725 123.975 115.945 124.255 ;
        RECT 116.425 124.085 116.665 124.485 ;
        RECT 115.385 123.635 115.790 123.805 ;
        RECT 116.125 123.715 116.665 124.085 ;
        RECT 116.835 124.300 117.155 124.655 ;
        RECT 116.835 124.045 117.160 124.300 ;
        RECT 117.355 124.225 117.525 125.035 ;
        RECT 117.695 124.385 118.025 124.865 ;
        RECT 118.195 124.565 118.365 125.035 ;
        RECT 118.535 124.385 118.865 124.865 ;
        RECT 119.035 124.565 119.205 125.035 ;
        RECT 117.695 124.215 119.460 124.385 ;
        RECT 119.745 124.215 119.955 125.035 ;
        RECT 120.125 124.235 120.455 124.865 ;
        RECT 116.835 123.835 118.865 124.045 ;
        RECT 116.835 123.825 117.180 123.835 ;
        RECT 114.485 123.465 115.160 123.625 ;
        RECT 115.620 123.545 115.790 123.635 ;
        RECT 114.485 123.455 115.450 123.465 ;
        RECT 114.125 123.285 114.295 123.425 ;
        RECT 110.870 122.485 111.120 122.945 ;
        RECT 111.290 122.655 111.540 122.985 ;
        RECT 111.755 122.655 112.435 122.985 ;
        RECT 112.605 123.085 113.680 123.255 ;
        RECT 114.125 123.115 114.685 123.285 ;
        RECT 114.990 123.165 115.450 123.455 ;
        RECT 115.620 123.375 116.840 123.545 ;
        RECT 112.605 122.745 112.775 123.085 ;
        RECT 113.010 122.485 113.340 122.915 ;
        RECT 113.510 122.745 113.680 123.085 ;
        RECT 113.975 122.485 114.345 122.945 ;
        RECT 114.515 122.655 114.685 123.115 ;
        RECT 115.620 122.995 115.790 123.375 ;
        RECT 117.010 123.205 117.180 123.825 ;
        RECT 119.050 123.665 119.460 124.215 ;
        RECT 114.920 122.655 115.790 122.995 ;
        RECT 116.380 123.035 117.180 123.205 ;
        RECT 115.960 122.485 116.210 122.945 ;
        RECT 116.380 122.745 116.550 123.035 ;
        RECT 116.730 122.485 117.060 122.865 ;
        RECT 117.355 122.485 117.525 123.545 ;
        RECT 117.735 123.495 119.460 123.665 ;
        RECT 120.125 123.635 120.375 124.235 ;
        RECT 120.625 124.215 120.855 125.035 ;
        RECT 121.105 124.215 121.335 125.035 ;
        RECT 121.505 124.235 121.835 124.865 ;
        RECT 120.545 123.795 120.875 124.045 ;
        RECT 121.085 123.795 121.415 124.045 ;
        RECT 121.585 123.635 121.835 124.235 ;
        RECT 122.005 124.215 122.215 125.035 ;
        RECT 122.445 124.265 124.115 125.035 ;
        RECT 124.285 124.285 125.495 125.035 ;
        RECT 122.445 123.745 123.195 124.265 ;
        RECT 117.735 122.655 118.025 123.495 ;
        RECT 118.195 122.485 118.365 123.325 ;
        RECT 118.575 122.655 118.825 123.495 ;
        RECT 119.035 122.485 119.205 123.325 ;
        RECT 119.745 122.485 119.955 123.625 ;
        RECT 120.125 122.655 120.455 123.635 ;
        RECT 120.625 122.485 120.855 123.625 ;
        RECT 121.105 122.485 121.335 123.625 ;
        RECT 121.505 122.655 121.835 123.635 ;
        RECT 122.005 122.485 122.215 123.625 ;
        RECT 123.365 123.575 124.115 124.095 ;
        RECT 122.445 122.485 124.115 123.575 ;
        RECT 124.285 123.575 124.805 124.115 ;
        RECT 124.975 123.745 125.495 124.285 ;
        RECT 124.285 122.485 125.495 123.575 ;
        RECT 5.520 122.315 125.580 122.485 ;
        RECT 5.605 121.225 6.815 122.315 ;
        RECT 7.295 121.475 7.465 122.315 ;
        RECT 7.675 121.305 7.925 122.145 ;
        RECT 8.135 121.475 8.305 122.315 ;
        RECT 8.475 121.305 8.765 122.145 ;
        RECT 5.605 120.515 6.125 121.055 ;
        RECT 6.295 120.685 6.815 121.225 ;
        RECT 7.040 121.135 8.765 121.305 ;
        RECT 8.975 121.255 9.145 122.315 ;
        RECT 9.440 121.935 9.770 122.315 ;
        RECT 9.950 121.765 10.120 122.055 ;
        RECT 10.290 121.855 10.540 122.315 ;
        RECT 9.320 121.595 10.120 121.765 ;
        RECT 10.710 121.805 11.580 122.145 ;
        RECT 7.040 120.585 7.450 121.135 ;
        RECT 9.320 120.975 9.490 121.595 ;
        RECT 10.710 121.425 10.880 121.805 ;
        RECT 11.815 121.685 11.985 122.145 ;
        RECT 12.155 121.855 12.525 122.315 ;
        RECT 12.820 121.715 12.990 122.055 ;
        RECT 13.160 121.885 13.490 122.315 ;
        RECT 13.725 121.715 13.895 122.055 ;
        RECT 9.660 121.255 10.880 121.425 ;
        RECT 11.050 121.345 11.510 121.635 ;
        RECT 11.815 121.515 12.375 121.685 ;
        RECT 12.820 121.545 13.895 121.715 ;
        RECT 14.065 121.815 14.745 122.145 ;
        RECT 14.960 121.815 15.210 122.145 ;
        RECT 15.380 121.855 15.630 122.315 ;
        RECT 12.205 121.375 12.375 121.515 ;
        RECT 11.050 121.335 12.015 121.345 ;
        RECT 10.710 121.165 10.880 121.255 ;
        RECT 11.340 121.175 12.015 121.335 ;
        RECT 9.320 120.965 9.665 120.975 ;
        RECT 7.635 120.755 9.665 120.965 ;
        RECT 5.605 119.765 6.815 120.515 ;
        RECT 7.040 120.415 8.805 120.585 ;
        RECT 7.295 119.765 7.465 120.235 ;
        RECT 7.635 119.935 7.965 120.415 ;
        RECT 8.135 119.765 8.305 120.235 ;
        RECT 8.475 119.935 8.805 120.415 ;
        RECT 8.975 119.765 9.145 120.575 ;
        RECT 9.340 120.500 9.665 120.755 ;
        RECT 9.345 120.145 9.665 120.500 ;
        RECT 9.835 120.715 10.375 121.085 ;
        RECT 10.710 120.995 11.115 121.165 ;
        RECT 9.835 120.315 10.075 120.715 ;
        RECT 10.555 120.545 10.775 120.825 ;
        RECT 10.245 120.375 10.775 120.545 ;
        RECT 10.245 120.145 10.415 120.375 ;
        RECT 10.945 120.215 11.115 120.995 ;
        RECT 11.285 120.385 11.635 121.005 ;
        RECT 11.805 120.385 12.015 121.175 ;
        RECT 12.205 121.205 13.705 121.375 ;
        RECT 12.205 120.515 12.375 121.205 ;
        RECT 14.065 121.035 14.235 121.815 ;
        RECT 15.040 121.685 15.210 121.815 ;
        RECT 12.545 120.865 14.235 121.035 ;
        RECT 14.405 121.255 14.870 121.645 ;
        RECT 15.040 121.515 15.435 121.685 ;
        RECT 12.545 120.685 12.715 120.865 ;
        RECT 9.345 119.975 10.415 120.145 ;
        RECT 10.585 119.765 10.775 120.205 ;
        RECT 10.945 119.935 11.895 120.215 ;
        RECT 12.205 120.125 12.465 120.515 ;
        RECT 12.885 120.445 13.675 120.695 ;
        RECT 12.115 119.955 12.465 120.125 ;
        RECT 12.675 119.765 13.005 120.225 ;
        RECT 13.880 120.155 14.050 120.865 ;
        RECT 14.405 120.665 14.575 121.255 ;
        RECT 14.220 120.445 14.575 120.665 ;
        RECT 14.745 120.445 15.095 121.065 ;
        RECT 15.265 120.155 15.435 121.515 ;
        RECT 15.800 121.345 16.125 122.130 ;
        RECT 15.605 120.295 16.065 121.345 ;
        RECT 13.880 119.985 14.735 120.155 ;
        RECT 14.940 119.985 15.435 120.155 ;
        RECT 15.605 119.765 15.935 120.125 ;
        RECT 16.295 120.025 16.465 122.145 ;
        RECT 16.635 121.815 16.965 122.315 ;
        RECT 17.135 121.645 17.390 122.145 ;
        RECT 16.640 121.475 17.390 121.645 ;
        RECT 16.640 120.485 16.870 121.475 ;
        RECT 17.040 120.655 17.390 121.305 ;
        RECT 18.485 121.150 18.775 122.315 ;
        RECT 18.945 121.225 20.615 122.315 ;
        RECT 18.945 120.535 19.695 121.055 ;
        RECT 19.865 120.705 20.615 121.225 ;
        RECT 21.245 121.240 21.515 122.145 ;
        RECT 21.685 121.555 22.015 122.315 ;
        RECT 22.195 121.385 22.365 122.145 ;
        RECT 16.640 120.315 17.390 120.485 ;
        RECT 16.635 119.765 16.965 120.145 ;
        RECT 17.135 120.025 17.390 120.315 ;
        RECT 18.485 119.765 18.775 120.490 ;
        RECT 18.945 119.765 20.615 120.535 ;
        RECT 21.245 120.440 21.415 121.240 ;
        RECT 21.700 121.215 22.365 121.385 ;
        RECT 23.545 121.240 23.815 122.145 ;
        RECT 23.985 121.555 24.315 122.315 ;
        RECT 24.495 121.385 24.665 122.145 ;
        RECT 21.700 121.070 21.870 121.215 ;
        RECT 21.585 120.740 21.870 121.070 ;
        RECT 21.700 120.485 21.870 120.740 ;
        RECT 22.105 120.665 22.435 121.035 ;
        RECT 21.245 119.935 21.505 120.440 ;
        RECT 21.700 120.315 22.365 120.485 ;
        RECT 21.685 119.765 22.015 120.145 ;
        RECT 22.195 119.935 22.365 120.315 ;
        RECT 23.545 120.440 23.715 121.240 ;
        RECT 24.000 121.215 24.665 121.385 ;
        RECT 24.000 121.070 24.170 121.215 ;
        RECT 24.985 121.175 25.195 122.315 ;
        RECT 23.885 120.740 24.170 121.070 ;
        RECT 25.365 121.165 25.695 122.145 ;
        RECT 25.865 121.175 26.095 122.315 ;
        RECT 26.305 121.225 27.515 122.315 ;
        RECT 24.000 120.485 24.170 120.740 ;
        RECT 24.405 120.665 24.735 121.035 ;
        RECT 23.545 119.935 23.805 120.440 ;
        RECT 24.000 120.315 24.665 120.485 ;
        RECT 23.985 119.765 24.315 120.145 ;
        RECT 24.495 119.935 24.665 120.315 ;
        RECT 24.985 119.765 25.195 120.585 ;
        RECT 25.365 120.565 25.615 121.165 ;
        RECT 25.785 120.755 26.115 121.005 ;
        RECT 25.365 119.935 25.695 120.565 ;
        RECT 25.865 119.765 26.095 120.585 ;
        RECT 26.305 120.515 26.825 121.055 ;
        RECT 26.995 120.685 27.515 121.225 ;
        RECT 27.685 121.240 27.955 122.145 ;
        RECT 28.125 121.555 28.455 122.315 ;
        RECT 28.635 121.385 28.805 122.145 ;
        RECT 29.065 121.880 34.410 122.315 ;
        RECT 26.305 119.765 27.515 120.515 ;
        RECT 27.685 120.440 27.855 121.240 ;
        RECT 28.140 121.215 28.805 121.385 ;
        RECT 28.140 121.070 28.310 121.215 ;
        RECT 28.025 120.740 28.310 121.070 ;
        RECT 28.140 120.485 28.310 120.740 ;
        RECT 28.545 120.665 28.875 121.035 ;
        RECT 27.685 119.935 27.945 120.440 ;
        RECT 28.140 120.315 28.805 120.485 ;
        RECT 28.125 119.765 28.455 120.145 ;
        RECT 28.635 119.935 28.805 120.315 ;
        RECT 30.650 120.310 30.990 121.140 ;
        RECT 32.470 120.630 32.820 121.880 ;
        RECT 34.585 121.240 34.855 122.145 ;
        RECT 35.025 121.555 35.355 122.315 ;
        RECT 35.535 121.385 35.705 122.145 ;
        RECT 34.585 120.440 34.755 121.240 ;
        RECT 35.040 121.215 35.705 121.385 ;
        RECT 35.965 121.225 39.475 122.315 ;
        RECT 35.040 121.070 35.210 121.215 ;
        RECT 34.925 120.740 35.210 121.070 ;
        RECT 35.040 120.485 35.210 120.740 ;
        RECT 35.445 120.665 35.775 121.035 ;
        RECT 35.965 120.535 37.615 121.055 ;
        RECT 37.785 120.705 39.475 121.225 ;
        RECT 40.565 121.240 40.835 122.145 ;
        RECT 41.005 121.555 41.335 122.315 ;
        RECT 41.515 121.385 41.685 122.145 ;
        RECT 29.065 119.765 34.410 120.310 ;
        RECT 34.585 119.935 34.845 120.440 ;
        RECT 35.040 120.315 35.705 120.485 ;
        RECT 35.025 119.765 35.355 120.145 ;
        RECT 35.535 119.935 35.705 120.315 ;
        RECT 35.965 119.765 39.475 120.535 ;
        RECT 40.565 120.440 40.735 121.240 ;
        RECT 41.020 121.215 41.685 121.385 ;
        RECT 41.945 121.225 43.615 122.315 ;
        RECT 41.020 121.070 41.190 121.215 ;
        RECT 40.905 120.740 41.190 121.070 ;
        RECT 41.020 120.485 41.190 120.740 ;
        RECT 41.425 120.665 41.755 121.035 ;
        RECT 41.945 120.535 42.695 121.055 ;
        RECT 42.865 120.705 43.615 121.225 ;
        RECT 44.245 121.150 44.535 122.315 ;
        RECT 45.625 121.240 45.895 122.145 ;
        RECT 46.065 121.555 46.395 122.315 ;
        RECT 46.575 121.385 46.745 122.145 ;
        RECT 47.005 121.880 52.350 122.315 ;
        RECT 40.565 119.935 40.825 120.440 ;
        RECT 41.020 120.315 41.685 120.485 ;
        RECT 41.005 119.765 41.335 120.145 ;
        RECT 41.515 119.935 41.685 120.315 ;
        RECT 41.945 119.765 43.615 120.535 ;
        RECT 44.245 119.765 44.535 120.490 ;
        RECT 45.625 120.440 45.795 121.240 ;
        RECT 46.080 121.215 46.745 121.385 ;
        RECT 46.080 121.070 46.250 121.215 ;
        RECT 45.965 120.740 46.250 121.070 ;
        RECT 46.080 120.485 46.250 120.740 ;
        RECT 46.485 120.665 46.815 121.035 ;
        RECT 45.625 119.935 45.885 120.440 ;
        RECT 46.080 120.315 46.745 120.485 ;
        RECT 46.065 119.765 46.395 120.145 ;
        RECT 46.575 119.935 46.745 120.315 ;
        RECT 48.590 120.310 48.930 121.140 ;
        RECT 50.410 120.630 50.760 121.880 ;
        RECT 52.675 121.165 53.005 122.315 ;
        RECT 53.175 121.295 53.345 122.145 ;
        RECT 53.515 121.515 53.845 122.315 ;
        RECT 54.015 121.295 54.185 122.145 ;
        RECT 54.365 121.515 54.605 122.315 ;
        RECT 54.775 121.335 55.105 122.145 ;
        RECT 53.175 121.125 54.185 121.295 ;
        RECT 54.390 121.165 55.105 121.335 ;
        RECT 55.285 121.225 57.875 122.315 ;
        RECT 53.175 120.585 53.670 121.125 ;
        RECT 54.390 120.925 54.560 121.165 ;
        RECT 54.060 120.755 54.560 120.925 ;
        RECT 54.730 120.755 55.110 120.995 ;
        RECT 54.390 120.585 54.560 120.755 ;
        RECT 47.005 119.765 52.350 120.310 ;
        RECT 52.675 119.765 53.005 120.565 ;
        RECT 53.175 120.415 54.185 120.585 ;
        RECT 54.390 120.415 55.025 120.585 ;
        RECT 53.175 119.935 53.345 120.415 ;
        RECT 53.515 119.765 53.845 120.245 ;
        RECT 54.015 119.935 54.185 120.415 ;
        RECT 54.435 119.765 54.675 120.245 ;
        RECT 54.855 119.935 55.025 120.415 ;
        RECT 55.285 120.535 56.495 121.055 ;
        RECT 56.665 120.705 57.875 121.225 ;
        RECT 58.545 121.175 58.775 122.315 ;
        RECT 58.945 121.165 59.275 122.145 ;
        RECT 59.445 121.175 59.655 122.315 ;
        RECT 59.885 121.880 65.230 122.315 ;
        RECT 58.525 120.755 58.855 121.005 ;
        RECT 55.285 119.765 57.875 120.535 ;
        RECT 58.545 119.765 58.775 120.585 ;
        RECT 59.025 120.565 59.275 121.165 ;
        RECT 58.945 119.935 59.275 120.565 ;
        RECT 59.445 119.765 59.655 120.585 ;
        RECT 61.470 120.310 61.810 121.140 ;
        RECT 63.290 120.630 63.640 121.880 ;
        RECT 65.405 121.225 67.075 122.315 ;
        RECT 65.405 120.535 66.155 121.055 ;
        RECT 66.325 120.705 67.075 121.225 ;
        RECT 67.705 121.240 67.975 122.145 ;
        RECT 68.145 121.555 68.475 122.315 ;
        RECT 68.655 121.385 68.825 122.145 ;
        RECT 59.885 119.765 65.230 120.310 ;
        RECT 65.405 119.765 67.075 120.535 ;
        RECT 67.705 120.440 67.875 121.240 ;
        RECT 68.160 121.215 68.825 121.385 ;
        RECT 68.160 121.070 68.330 121.215 ;
        RECT 70.005 121.150 70.295 122.315 ;
        RECT 70.525 121.175 70.735 122.315 ;
        RECT 70.905 121.165 71.235 122.145 ;
        RECT 71.405 121.175 71.635 122.315 ;
        RECT 72.915 121.165 73.245 122.315 ;
        RECT 73.415 121.295 73.585 122.145 ;
        RECT 73.755 121.515 74.085 122.315 ;
        RECT 74.255 121.295 74.425 122.145 ;
        RECT 74.605 121.515 74.845 122.315 ;
        RECT 75.015 121.335 75.345 122.145 ;
        RECT 68.045 120.740 68.330 121.070 ;
        RECT 68.160 120.485 68.330 120.740 ;
        RECT 68.565 120.665 68.895 121.035 ;
        RECT 67.705 119.935 67.965 120.440 ;
        RECT 68.160 120.315 68.825 120.485 ;
        RECT 68.145 119.765 68.475 120.145 ;
        RECT 68.655 119.935 68.825 120.315 ;
        RECT 70.005 119.765 70.295 120.490 ;
        RECT 70.525 119.765 70.735 120.585 ;
        RECT 70.905 120.565 71.155 121.165 ;
        RECT 73.415 121.125 74.425 121.295 ;
        RECT 74.630 121.165 75.345 121.335 ;
        RECT 75.525 121.240 75.795 122.145 ;
        RECT 75.965 121.555 76.295 122.315 ;
        RECT 76.475 121.385 76.645 122.145 ;
        RECT 71.325 120.755 71.655 121.005 ;
        RECT 73.415 120.585 73.910 121.125 ;
        RECT 74.630 120.925 74.800 121.165 ;
        RECT 74.300 120.755 74.800 120.925 ;
        RECT 74.970 120.755 75.350 120.995 ;
        RECT 74.630 120.585 74.800 120.755 ;
        RECT 70.905 119.935 71.235 120.565 ;
        RECT 71.405 119.765 71.635 120.585 ;
        RECT 72.915 119.765 73.245 120.565 ;
        RECT 73.415 120.415 74.425 120.585 ;
        RECT 74.630 120.415 75.265 120.585 ;
        RECT 73.415 119.935 73.585 120.415 ;
        RECT 73.755 119.765 74.085 120.245 ;
        RECT 74.255 119.935 74.425 120.415 ;
        RECT 74.675 119.765 74.915 120.245 ;
        RECT 75.095 119.935 75.265 120.415 ;
        RECT 75.525 120.440 75.695 121.240 ;
        RECT 75.980 121.215 76.645 121.385 ;
        RECT 76.905 121.225 78.575 122.315 ;
        RECT 75.980 121.070 76.150 121.215 ;
        RECT 75.865 120.740 76.150 121.070 ;
        RECT 75.980 120.485 76.150 120.740 ;
        RECT 76.385 120.665 76.715 121.035 ;
        RECT 76.905 120.535 77.655 121.055 ;
        RECT 77.825 120.705 78.575 121.225 ;
        RECT 78.745 121.240 79.015 122.145 ;
        RECT 79.185 121.555 79.515 122.315 ;
        RECT 79.695 121.385 79.865 122.145 ;
        RECT 75.525 119.935 75.785 120.440 ;
        RECT 75.980 120.315 76.645 120.485 ;
        RECT 75.965 119.765 76.295 120.145 ;
        RECT 76.475 119.935 76.645 120.315 ;
        RECT 76.905 119.765 78.575 120.535 ;
        RECT 78.745 120.440 78.915 121.240 ;
        RECT 79.200 121.215 79.865 121.385 ;
        RECT 80.125 121.225 83.635 122.315 ;
        RECT 79.200 121.070 79.370 121.215 ;
        RECT 79.085 120.740 79.370 121.070 ;
        RECT 79.200 120.485 79.370 120.740 ;
        RECT 79.605 120.665 79.935 121.035 ;
        RECT 80.125 120.535 81.775 121.055 ;
        RECT 81.945 120.705 83.635 121.225 ;
        RECT 84.355 121.385 84.525 122.145 ;
        RECT 84.705 121.555 85.035 122.315 ;
        RECT 84.355 121.215 85.020 121.385 ;
        RECT 85.205 121.240 85.475 122.145 ;
        RECT 84.850 121.070 85.020 121.215 ;
        RECT 84.285 120.665 84.615 121.035 ;
        RECT 84.850 120.740 85.135 121.070 ;
        RECT 78.745 119.935 79.005 120.440 ;
        RECT 79.200 120.315 79.865 120.485 ;
        RECT 79.185 119.765 79.515 120.145 ;
        RECT 79.695 119.935 79.865 120.315 ;
        RECT 80.125 119.765 83.635 120.535 ;
        RECT 84.850 120.485 85.020 120.740 ;
        RECT 84.355 120.315 85.020 120.485 ;
        RECT 85.305 120.440 85.475 121.240 ;
        RECT 85.645 121.225 89.155 122.315 ;
        RECT 84.355 119.935 84.525 120.315 ;
        RECT 84.705 119.765 85.035 120.145 ;
        RECT 85.215 119.935 85.475 120.440 ;
        RECT 85.645 120.535 87.295 121.055 ;
        RECT 87.465 120.705 89.155 121.225 ;
        RECT 89.325 121.240 89.595 122.145 ;
        RECT 89.765 121.555 90.095 122.315 ;
        RECT 90.275 121.385 90.445 122.145 ;
        RECT 85.645 119.765 89.155 120.535 ;
        RECT 89.325 120.440 89.495 121.240 ;
        RECT 89.780 121.215 90.445 121.385 ;
        RECT 90.705 121.225 91.915 122.315 ;
        RECT 89.780 121.070 89.950 121.215 ;
        RECT 89.665 120.740 89.950 121.070 ;
        RECT 89.780 120.485 89.950 120.740 ;
        RECT 90.185 120.665 90.515 121.035 ;
        RECT 90.705 120.515 91.225 121.055 ;
        RECT 91.395 120.685 91.915 121.225 ;
        RECT 92.175 121.385 92.345 122.145 ;
        RECT 92.525 121.555 92.855 122.315 ;
        RECT 92.175 121.215 92.840 121.385 ;
        RECT 93.025 121.240 93.295 122.145 ;
        RECT 92.670 121.070 92.840 121.215 ;
        RECT 92.105 120.665 92.435 121.035 ;
        RECT 92.670 120.740 92.955 121.070 ;
        RECT 89.325 119.935 89.585 120.440 ;
        RECT 89.780 120.315 90.445 120.485 ;
        RECT 89.765 119.765 90.095 120.145 ;
        RECT 90.275 119.935 90.445 120.315 ;
        RECT 90.705 119.765 91.915 120.515 ;
        RECT 92.670 120.485 92.840 120.740 ;
        RECT 92.175 120.315 92.840 120.485 ;
        RECT 93.125 120.440 93.295 121.240 ;
        RECT 93.525 121.175 93.735 122.315 ;
        RECT 93.905 121.165 94.235 122.145 ;
        RECT 94.405 121.175 94.635 122.315 ;
        RECT 92.175 119.935 92.345 120.315 ;
        RECT 92.525 119.765 92.855 120.145 ;
        RECT 93.035 119.935 93.295 120.440 ;
        RECT 93.525 119.765 93.735 120.585 ;
        RECT 93.905 120.565 94.155 121.165 ;
        RECT 95.765 121.150 96.055 122.315 ;
        RECT 96.225 121.880 101.570 122.315 ;
        RECT 94.325 120.755 94.655 121.005 ;
        RECT 93.905 119.935 94.235 120.565 ;
        RECT 94.405 119.765 94.635 120.585 ;
        RECT 95.765 119.765 96.055 120.490 ;
        RECT 97.810 120.310 98.150 121.140 ;
        RECT 99.630 120.630 99.980 121.880 ;
        RECT 102.295 121.385 102.465 122.145 ;
        RECT 102.645 121.555 102.975 122.315 ;
        RECT 102.295 121.215 102.960 121.385 ;
        RECT 103.145 121.240 103.415 122.145 ;
        RECT 102.790 121.070 102.960 121.215 ;
        RECT 102.225 120.665 102.555 121.035 ;
        RECT 102.790 120.740 103.075 121.070 ;
        RECT 102.790 120.485 102.960 120.740 ;
        RECT 102.295 120.315 102.960 120.485 ;
        RECT 103.245 120.440 103.415 121.240 ;
        RECT 103.585 121.225 105.255 122.315 ;
        RECT 96.225 119.765 101.570 120.310 ;
        RECT 102.295 119.935 102.465 120.315 ;
        RECT 102.645 119.765 102.975 120.145 ;
        RECT 103.155 119.935 103.415 120.440 ;
        RECT 103.585 120.535 104.335 121.055 ;
        RECT 104.505 120.705 105.255 121.225 ;
        RECT 105.975 121.385 106.145 122.145 ;
        RECT 106.325 121.555 106.655 122.315 ;
        RECT 105.975 121.215 106.640 121.385 ;
        RECT 106.825 121.240 107.095 122.145 ;
        RECT 106.470 121.070 106.640 121.215 ;
        RECT 105.905 120.665 106.235 121.035 ;
        RECT 106.470 120.740 106.755 121.070 ;
        RECT 103.585 119.765 105.255 120.535 ;
        RECT 106.470 120.485 106.640 120.740 ;
        RECT 105.975 120.315 106.640 120.485 ;
        RECT 106.925 120.440 107.095 121.240 ;
        RECT 107.355 121.385 107.525 122.145 ;
        RECT 107.705 121.555 108.035 122.315 ;
        RECT 107.355 121.215 108.020 121.385 ;
        RECT 108.205 121.240 108.475 122.145 ;
        RECT 107.850 121.070 108.020 121.215 ;
        RECT 107.285 120.665 107.615 121.035 ;
        RECT 107.850 120.740 108.135 121.070 ;
        RECT 107.850 120.485 108.020 120.740 ;
        RECT 105.975 119.935 106.145 120.315 ;
        RECT 106.325 119.765 106.655 120.145 ;
        RECT 106.835 119.935 107.095 120.440 ;
        RECT 107.355 120.315 108.020 120.485 ;
        RECT 108.305 120.440 108.475 121.240 ;
        RECT 109.655 121.385 109.825 122.145 ;
        RECT 110.005 121.555 110.335 122.315 ;
        RECT 109.655 121.215 110.320 121.385 ;
        RECT 110.505 121.240 110.775 122.145 ;
        RECT 110.950 121.645 111.205 122.145 ;
        RECT 111.375 121.815 111.705 122.315 ;
        RECT 110.950 121.475 111.700 121.645 ;
        RECT 110.150 121.070 110.320 121.215 ;
        RECT 109.585 120.665 109.915 121.035 ;
        RECT 110.150 120.740 110.435 121.070 ;
        RECT 110.150 120.485 110.320 120.740 ;
        RECT 107.355 119.935 107.525 120.315 ;
        RECT 107.705 119.765 108.035 120.145 ;
        RECT 108.215 119.935 108.475 120.440 ;
        RECT 109.655 120.315 110.320 120.485 ;
        RECT 110.605 120.440 110.775 121.240 ;
        RECT 110.950 120.655 111.300 121.305 ;
        RECT 111.470 120.485 111.700 121.475 ;
        RECT 109.655 119.935 109.825 120.315 ;
        RECT 110.005 119.765 110.335 120.145 ;
        RECT 110.515 119.935 110.775 120.440 ;
        RECT 110.950 120.315 111.700 120.485 ;
        RECT 110.950 120.025 111.205 120.315 ;
        RECT 111.375 119.765 111.705 120.145 ;
        RECT 111.875 120.025 112.045 122.145 ;
        RECT 112.215 121.345 112.540 122.130 ;
        RECT 112.710 121.855 112.960 122.315 ;
        RECT 113.130 121.815 113.380 122.145 ;
        RECT 113.595 121.815 114.275 122.145 ;
        RECT 113.130 121.685 113.300 121.815 ;
        RECT 112.905 121.515 113.300 121.685 ;
        RECT 112.275 120.295 112.735 121.345 ;
        RECT 112.905 120.155 113.075 121.515 ;
        RECT 113.470 121.255 113.935 121.645 ;
        RECT 113.245 120.445 113.595 121.065 ;
        RECT 113.765 120.665 113.935 121.255 ;
        RECT 114.105 121.035 114.275 121.815 ;
        RECT 114.445 121.715 114.615 122.055 ;
        RECT 114.850 121.885 115.180 122.315 ;
        RECT 115.350 121.715 115.520 122.055 ;
        RECT 115.815 121.855 116.185 122.315 ;
        RECT 114.445 121.545 115.520 121.715 ;
        RECT 116.355 121.685 116.525 122.145 ;
        RECT 116.760 121.805 117.630 122.145 ;
        RECT 117.800 121.855 118.050 122.315 ;
        RECT 115.965 121.515 116.525 121.685 ;
        RECT 115.965 121.375 116.135 121.515 ;
        RECT 114.635 121.205 116.135 121.375 ;
        RECT 116.830 121.345 117.290 121.635 ;
        RECT 114.105 120.865 115.795 121.035 ;
        RECT 113.765 120.445 114.120 120.665 ;
        RECT 114.290 120.155 114.460 120.865 ;
        RECT 114.665 120.445 115.455 120.695 ;
        RECT 115.625 120.685 115.795 120.865 ;
        RECT 115.965 120.515 116.135 121.205 ;
        RECT 112.405 119.765 112.735 120.125 ;
        RECT 112.905 119.985 113.400 120.155 ;
        RECT 113.605 119.985 114.460 120.155 ;
        RECT 115.335 119.765 115.665 120.225 ;
        RECT 115.875 120.125 116.135 120.515 ;
        RECT 116.325 121.335 117.290 121.345 ;
        RECT 117.460 121.425 117.630 121.805 ;
        RECT 118.220 121.765 118.390 122.055 ;
        RECT 118.570 121.935 118.900 122.315 ;
        RECT 118.220 121.595 119.020 121.765 ;
        RECT 116.325 121.175 117.000 121.335 ;
        RECT 117.460 121.255 118.680 121.425 ;
        RECT 116.325 120.385 116.535 121.175 ;
        RECT 117.460 121.165 117.630 121.255 ;
        RECT 116.705 120.385 117.055 121.005 ;
        RECT 117.225 120.995 117.630 121.165 ;
        RECT 117.225 120.215 117.395 120.995 ;
        RECT 117.565 120.545 117.785 120.825 ;
        RECT 117.965 120.715 118.505 121.085 ;
        RECT 118.850 120.975 119.020 121.595 ;
        RECT 119.195 121.255 119.365 122.315 ;
        RECT 119.575 121.305 119.865 122.145 ;
        RECT 120.035 121.475 120.205 122.315 ;
        RECT 120.415 121.305 120.665 122.145 ;
        RECT 120.875 121.475 121.045 122.315 ;
        RECT 119.575 121.135 121.300 121.305 ;
        RECT 121.525 121.150 121.815 122.315 ;
        RECT 121.985 121.225 123.655 122.315 ;
        RECT 117.565 120.375 118.095 120.545 ;
        RECT 115.875 119.955 116.225 120.125 ;
        RECT 116.445 119.935 117.395 120.215 ;
        RECT 117.565 119.765 117.755 120.205 ;
        RECT 117.925 120.145 118.095 120.375 ;
        RECT 118.265 120.315 118.505 120.715 ;
        RECT 118.675 120.965 119.020 120.975 ;
        RECT 118.675 120.755 120.705 120.965 ;
        RECT 118.675 120.500 119.000 120.755 ;
        RECT 120.890 120.585 121.300 121.135 ;
        RECT 118.675 120.145 118.995 120.500 ;
        RECT 117.925 119.975 118.995 120.145 ;
        RECT 119.195 119.765 119.365 120.575 ;
        RECT 119.535 120.415 121.300 120.585 ;
        RECT 121.985 120.535 122.735 121.055 ;
        RECT 122.905 120.705 123.655 121.225 ;
        RECT 124.285 121.225 125.495 122.315 ;
        RECT 124.285 120.685 124.805 121.225 ;
        RECT 119.535 119.935 119.865 120.415 ;
        RECT 120.035 119.765 120.205 120.235 ;
        RECT 120.375 119.935 120.705 120.415 ;
        RECT 120.875 119.765 121.045 120.235 ;
        RECT 121.525 119.765 121.815 120.490 ;
        RECT 121.985 119.765 123.655 120.535 ;
        RECT 124.975 120.515 125.495 121.055 ;
        RECT 124.285 119.765 125.495 120.515 ;
        RECT 5.520 119.595 125.580 119.765 ;
        RECT 5.605 118.845 6.815 119.595 ;
        RECT 7.075 119.045 7.245 119.425 ;
        RECT 7.425 119.215 7.755 119.595 ;
        RECT 7.075 118.875 7.740 119.045 ;
        RECT 7.935 118.920 8.195 119.425 ;
        RECT 5.605 118.305 6.125 118.845 ;
        RECT 6.295 118.135 6.815 118.675 ;
        RECT 7.005 118.325 7.345 118.695 ;
        RECT 7.570 118.620 7.740 118.875 ;
        RECT 7.570 118.290 7.845 118.620 ;
        RECT 7.570 118.145 7.740 118.290 ;
        RECT 5.605 117.045 6.815 118.135 ;
        RECT 7.065 117.975 7.740 118.145 ;
        RECT 8.015 118.120 8.195 118.920 ;
        RECT 8.365 118.825 10.035 119.595 ;
        RECT 10.295 119.045 10.465 119.425 ;
        RECT 10.645 119.215 10.975 119.595 ;
        RECT 10.295 118.875 10.960 119.045 ;
        RECT 11.155 118.920 11.415 119.425 ;
        RECT 8.365 118.305 9.115 118.825 ;
        RECT 9.285 118.135 10.035 118.655 ;
        RECT 10.225 118.325 10.555 118.695 ;
        RECT 10.790 118.620 10.960 118.875 ;
        RECT 10.790 118.290 11.075 118.620 ;
        RECT 10.790 118.145 10.960 118.290 ;
        RECT 7.065 117.215 7.245 117.975 ;
        RECT 7.425 117.045 7.755 117.805 ;
        RECT 7.925 117.215 8.195 118.120 ;
        RECT 8.365 117.045 10.035 118.135 ;
        RECT 10.295 117.975 10.960 118.145 ;
        RECT 11.245 118.120 11.415 118.920 ;
        RECT 11.675 119.045 11.845 119.425 ;
        RECT 12.025 119.215 12.355 119.595 ;
        RECT 11.675 118.875 12.340 119.045 ;
        RECT 12.535 118.920 12.795 119.425 ;
        RECT 11.605 118.325 11.935 118.695 ;
        RECT 12.170 118.620 12.340 118.875 ;
        RECT 12.170 118.290 12.455 118.620 ;
        RECT 12.170 118.145 12.340 118.290 ;
        RECT 10.295 117.215 10.465 117.975 ;
        RECT 10.645 117.045 10.975 117.805 ;
        RECT 11.145 117.215 11.415 118.120 ;
        RECT 11.675 117.975 12.340 118.145 ;
        RECT 12.625 118.120 12.795 118.920 ;
        RECT 13.025 118.775 13.235 119.595 ;
        RECT 13.405 118.795 13.735 119.425 ;
        RECT 13.405 118.195 13.655 118.795 ;
        RECT 13.905 118.775 14.135 119.595 ;
        RECT 14.345 119.050 19.690 119.595 ;
        RECT 19.865 119.050 25.210 119.595 ;
        RECT 25.385 119.050 30.730 119.595 ;
        RECT 13.825 118.355 14.155 118.605 ;
        RECT 15.930 118.220 16.270 119.050 ;
        RECT 11.675 117.215 11.845 117.975 ;
        RECT 12.025 117.045 12.355 117.805 ;
        RECT 12.525 117.215 12.795 118.120 ;
        RECT 13.025 117.045 13.235 118.185 ;
        RECT 13.405 117.215 13.735 118.195 ;
        RECT 13.905 117.045 14.135 118.185 ;
        RECT 17.750 117.480 18.100 118.730 ;
        RECT 21.450 118.220 21.790 119.050 ;
        RECT 23.270 117.480 23.620 118.730 ;
        RECT 26.970 118.220 27.310 119.050 ;
        RECT 31.365 118.870 31.655 119.595 ;
        RECT 31.825 119.050 37.170 119.595 ;
        RECT 37.345 119.050 42.690 119.595 ;
        RECT 42.865 119.050 48.210 119.595 ;
        RECT 48.385 119.050 53.730 119.595 ;
        RECT 28.790 117.480 29.140 118.730 ;
        RECT 33.410 118.220 33.750 119.050 ;
        RECT 14.345 117.045 19.690 117.480 ;
        RECT 19.865 117.045 25.210 117.480 ;
        RECT 25.385 117.045 30.730 117.480 ;
        RECT 31.365 117.045 31.655 118.210 ;
        RECT 35.230 117.480 35.580 118.730 ;
        RECT 38.930 118.220 39.270 119.050 ;
        RECT 40.750 117.480 41.100 118.730 ;
        RECT 44.450 118.220 44.790 119.050 ;
        RECT 46.270 117.480 46.620 118.730 ;
        RECT 49.970 118.220 50.310 119.050 ;
        RECT 53.905 118.825 56.495 119.595 ;
        RECT 57.125 118.870 57.415 119.595 ;
        RECT 57.585 119.050 62.930 119.595 ;
        RECT 63.105 119.050 68.450 119.595 ;
        RECT 68.625 119.050 73.970 119.595 ;
        RECT 74.145 119.050 79.490 119.595 ;
        RECT 51.790 117.480 52.140 118.730 ;
        RECT 53.905 118.305 55.115 118.825 ;
        RECT 55.285 118.135 56.495 118.655 ;
        RECT 59.170 118.220 59.510 119.050 ;
        RECT 31.825 117.045 37.170 117.480 ;
        RECT 37.345 117.045 42.690 117.480 ;
        RECT 42.865 117.045 48.210 117.480 ;
        RECT 48.385 117.045 53.730 117.480 ;
        RECT 53.905 117.045 56.495 118.135 ;
        RECT 57.125 117.045 57.415 118.210 ;
        RECT 60.990 117.480 61.340 118.730 ;
        RECT 64.690 118.220 65.030 119.050 ;
        RECT 66.510 117.480 66.860 118.730 ;
        RECT 70.210 118.220 70.550 119.050 ;
        RECT 72.030 117.480 72.380 118.730 ;
        RECT 75.730 118.220 76.070 119.050 ;
        RECT 79.665 118.825 82.255 119.595 ;
        RECT 82.885 118.870 83.175 119.595 ;
        RECT 83.345 118.825 86.855 119.595 ;
        RECT 87.025 118.845 88.235 119.595 ;
        RECT 77.550 117.480 77.900 118.730 ;
        RECT 79.665 118.305 80.875 118.825 ;
        RECT 81.045 118.135 82.255 118.655 ;
        RECT 83.345 118.305 84.995 118.825 ;
        RECT 57.585 117.045 62.930 117.480 ;
        RECT 63.105 117.045 68.450 117.480 ;
        RECT 68.625 117.045 73.970 117.480 ;
        RECT 74.145 117.045 79.490 117.480 ;
        RECT 79.665 117.045 82.255 118.135 ;
        RECT 82.885 117.045 83.175 118.210 ;
        RECT 85.165 118.135 86.855 118.655 ;
        RECT 87.025 118.305 87.545 118.845 ;
        RECT 88.465 118.775 88.675 119.595 ;
        RECT 88.845 118.795 89.175 119.425 ;
        RECT 87.715 118.135 88.235 118.675 ;
        RECT 88.845 118.195 89.095 118.795 ;
        RECT 89.345 118.775 89.575 119.595 ;
        RECT 89.785 119.050 95.130 119.595 ;
        RECT 95.305 119.050 100.650 119.595 ;
        RECT 100.825 119.050 106.170 119.595 ;
        RECT 89.265 118.355 89.595 118.605 ;
        RECT 91.370 118.220 91.710 119.050 ;
        RECT 83.345 117.045 86.855 118.135 ;
        RECT 87.025 117.045 88.235 118.135 ;
        RECT 88.465 117.045 88.675 118.185 ;
        RECT 88.845 117.215 89.175 118.195 ;
        RECT 89.345 117.045 89.575 118.185 ;
        RECT 93.190 117.480 93.540 118.730 ;
        RECT 96.890 118.220 97.230 119.050 ;
        RECT 98.710 117.480 99.060 118.730 ;
        RECT 102.410 118.220 102.750 119.050 ;
        RECT 106.345 118.825 108.015 119.595 ;
        RECT 108.645 118.870 108.935 119.595 ;
        RECT 109.105 119.050 114.450 119.595 ;
        RECT 114.625 119.050 119.970 119.595 ;
        RECT 104.230 117.480 104.580 118.730 ;
        RECT 106.345 118.305 107.095 118.825 ;
        RECT 107.265 118.135 108.015 118.655 ;
        RECT 110.690 118.220 111.030 119.050 ;
        RECT 89.785 117.045 95.130 117.480 ;
        RECT 95.305 117.045 100.650 117.480 ;
        RECT 100.825 117.045 106.170 117.480 ;
        RECT 106.345 117.045 108.015 118.135 ;
        RECT 108.645 117.045 108.935 118.210 ;
        RECT 112.510 117.480 112.860 118.730 ;
        RECT 116.210 118.220 116.550 119.050 ;
        RECT 120.145 118.825 123.655 119.595 ;
        RECT 124.285 118.845 125.495 119.595 ;
        RECT 118.030 117.480 118.380 118.730 ;
        RECT 120.145 118.305 121.795 118.825 ;
        RECT 121.965 118.135 123.655 118.655 ;
        RECT 109.105 117.045 114.450 117.480 ;
        RECT 114.625 117.045 119.970 117.480 ;
        RECT 120.145 117.045 123.655 118.135 ;
        RECT 124.285 118.135 124.805 118.675 ;
        RECT 124.975 118.305 125.495 118.845 ;
        RECT 124.285 117.045 125.495 118.135 ;
        RECT 5.520 116.875 125.580 117.045 ;
        RECT 5.605 115.785 6.815 116.875 ;
        RECT 6.985 116.440 12.330 116.875 ;
        RECT 5.605 115.075 6.125 115.615 ;
        RECT 6.295 115.245 6.815 115.785 ;
        RECT 5.605 114.325 6.815 115.075 ;
        RECT 8.570 114.870 8.910 115.700 ;
        RECT 10.390 115.190 10.740 116.440 ;
        RECT 12.505 115.785 15.095 116.875 ;
        RECT 12.505 115.095 13.715 115.615 ;
        RECT 13.885 115.265 15.095 115.785 ;
        RECT 15.265 115.800 15.535 116.705 ;
        RECT 15.705 116.115 16.035 116.875 ;
        RECT 16.215 115.945 16.385 116.705 ;
        RECT 6.985 114.325 12.330 114.870 ;
        RECT 12.505 114.325 15.095 115.095 ;
        RECT 15.265 115.000 15.435 115.800 ;
        RECT 15.720 115.775 16.385 115.945 ;
        RECT 16.645 115.785 18.315 116.875 ;
        RECT 15.720 115.630 15.890 115.775 ;
        RECT 15.605 115.300 15.890 115.630 ;
        RECT 15.720 115.045 15.890 115.300 ;
        RECT 16.125 115.225 16.455 115.595 ;
        RECT 16.645 115.095 17.395 115.615 ;
        RECT 17.565 115.265 18.315 115.785 ;
        RECT 18.485 115.710 18.775 116.875 ;
        RECT 18.945 116.440 24.290 116.875 ;
        RECT 24.465 116.440 29.810 116.875 ;
        RECT 29.985 116.440 35.330 116.875 ;
        RECT 35.505 116.440 40.850 116.875 ;
        RECT 15.265 114.495 15.525 115.000 ;
        RECT 15.720 114.875 16.385 115.045 ;
        RECT 15.705 114.325 16.035 114.705 ;
        RECT 16.215 114.495 16.385 114.875 ;
        RECT 16.645 114.325 18.315 115.095 ;
        RECT 18.485 114.325 18.775 115.050 ;
        RECT 20.530 114.870 20.870 115.700 ;
        RECT 22.350 115.190 22.700 116.440 ;
        RECT 26.050 114.870 26.390 115.700 ;
        RECT 27.870 115.190 28.220 116.440 ;
        RECT 31.570 114.870 31.910 115.700 ;
        RECT 33.390 115.190 33.740 116.440 ;
        RECT 37.090 114.870 37.430 115.700 ;
        RECT 38.910 115.190 39.260 116.440 ;
        RECT 41.025 115.785 43.615 116.875 ;
        RECT 41.025 115.095 42.235 115.615 ;
        RECT 42.405 115.265 43.615 115.785 ;
        RECT 44.245 115.710 44.535 116.875 ;
        RECT 44.705 115.785 47.295 116.875 ;
        RECT 44.705 115.095 45.915 115.615 ;
        RECT 46.085 115.265 47.295 115.785 ;
        RECT 47.965 115.735 48.195 116.875 ;
        RECT 48.365 115.725 48.695 116.705 ;
        RECT 48.865 115.735 49.075 116.875 ;
        RECT 49.305 116.440 54.650 116.875 ;
        RECT 47.945 115.315 48.275 115.565 ;
        RECT 18.945 114.325 24.290 114.870 ;
        RECT 24.465 114.325 29.810 114.870 ;
        RECT 29.985 114.325 35.330 114.870 ;
        RECT 35.505 114.325 40.850 114.870 ;
        RECT 41.025 114.325 43.615 115.095 ;
        RECT 44.245 114.325 44.535 115.050 ;
        RECT 44.705 114.325 47.295 115.095 ;
        RECT 47.965 114.325 48.195 115.145 ;
        RECT 48.445 115.125 48.695 115.725 ;
        RECT 48.365 114.495 48.695 115.125 ;
        RECT 48.865 114.325 49.075 115.145 ;
        RECT 50.890 114.870 51.230 115.700 ;
        RECT 52.710 115.190 53.060 116.440 ;
        RECT 55.835 115.945 56.005 116.705 ;
        RECT 56.185 116.115 56.515 116.875 ;
        RECT 55.835 115.775 56.500 115.945 ;
        RECT 56.685 115.800 56.955 116.705 ;
        RECT 56.330 115.630 56.500 115.775 ;
        RECT 55.765 115.225 56.095 115.595 ;
        RECT 56.330 115.300 56.615 115.630 ;
        RECT 56.330 115.045 56.500 115.300 ;
        RECT 55.835 114.875 56.500 115.045 ;
        RECT 56.785 115.000 56.955 115.800 ;
        RECT 57.125 115.785 60.635 116.875 ;
        RECT 49.305 114.325 54.650 114.870 ;
        RECT 55.835 114.495 56.005 114.875 ;
        RECT 56.185 114.325 56.515 114.705 ;
        RECT 56.695 114.495 56.955 115.000 ;
        RECT 57.125 115.095 58.775 115.615 ;
        RECT 58.945 115.265 60.635 115.785 ;
        RECT 60.845 115.735 61.075 116.875 ;
        RECT 61.245 115.725 61.575 116.705 ;
        RECT 61.745 115.735 61.955 116.875 ;
        RECT 62.185 116.440 67.530 116.875 ;
        RECT 60.825 115.315 61.155 115.565 ;
        RECT 57.125 114.325 60.635 115.095 ;
        RECT 60.845 114.325 61.075 115.145 ;
        RECT 61.325 115.125 61.575 115.725 ;
        RECT 61.245 114.495 61.575 115.125 ;
        RECT 61.745 114.325 61.955 115.145 ;
        RECT 63.770 114.870 64.110 115.700 ;
        RECT 65.590 115.190 65.940 116.440 ;
        RECT 67.705 115.785 69.375 116.875 ;
        RECT 67.705 115.095 68.455 115.615 ;
        RECT 68.625 115.265 69.375 115.785 ;
        RECT 70.005 115.710 70.295 116.875 ;
        RECT 70.465 116.440 75.810 116.875 ;
        RECT 75.985 116.440 81.330 116.875 ;
        RECT 62.185 114.325 67.530 114.870 ;
        RECT 67.705 114.325 69.375 115.095 ;
        RECT 70.005 114.325 70.295 115.050 ;
        RECT 72.050 114.870 72.390 115.700 ;
        RECT 73.870 115.190 74.220 116.440 ;
        RECT 77.570 114.870 77.910 115.700 ;
        RECT 79.390 115.190 79.740 116.440 ;
        RECT 81.505 115.785 83.175 116.875 ;
        RECT 81.505 115.095 82.255 115.615 ;
        RECT 82.425 115.265 83.175 115.785 ;
        RECT 83.720 115.895 83.975 116.565 ;
        RECT 84.155 116.075 84.440 116.875 ;
        RECT 84.620 116.155 84.950 116.665 ;
        RECT 70.465 114.325 75.810 114.870 ;
        RECT 75.985 114.325 81.330 114.870 ;
        RECT 81.505 114.325 83.175 115.095 ;
        RECT 83.720 115.035 83.900 115.895 ;
        RECT 84.620 115.565 84.870 116.155 ;
        RECT 85.220 116.005 85.390 116.615 ;
        RECT 85.560 116.185 85.890 116.875 ;
        RECT 86.120 116.325 86.360 116.615 ;
        RECT 86.560 116.495 86.980 116.875 ;
        RECT 87.160 116.405 87.790 116.655 ;
        RECT 88.260 116.495 88.590 116.875 ;
        RECT 87.160 116.325 87.330 116.405 ;
        RECT 88.760 116.325 88.930 116.615 ;
        RECT 89.110 116.495 89.490 116.875 ;
        RECT 89.730 116.490 90.560 116.660 ;
        RECT 86.120 116.155 87.330 116.325 ;
        RECT 84.070 115.235 84.870 115.565 ;
        RECT 83.720 114.835 83.975 115.035 ;
        RECT 83.635 114.665 83.975 114.835 ;
        RECT 83.720 114.505 83.975 114.665 ;
        RECT 84.155 114.325 84.440 114.785 ;
        RECT 84.620 114.585 84.870 115.235 ;
        RECT 85.070 115.985 85.390 116.005 ;
        RECT 85.070 115.815 86.990 115.985 ;
        RECT 85.070 114.920 85.260 115.815 ;
        RECT 87.160 115.645 87.330 116.155 ;
        RECT 87.500 115.895 88.020 116.205 ;
        RECT 85.430 115.475 87.330 115.645 ;
        RECT 85.430 115.415 85.760 115.475 ;
        RECT 85.910 115.245 86.240 115.305 ;
        RECT 85.580 114.975 86.240 115.245 ;
        RECT 85.070 114.590 85.390 114.920 ;
        RECT 85.570 114.325 86.230 114.805 ;
        RECT 86.430 114.715 86.600 115.475 ;
        RECT 87.500 115.305 87.680 115.715 ;
        RECT 86.770 115.135 87.100 115.255 ;
        RECT 87.850 115.135 88.020 115.895 ;
        RECT 86.770 114.965 88.020 115.135 ;
        RECT 88.190 116.075 89.560 116.325 ;
        RECT 88.190 115.305 88.380 116.075 ;
        RECT 89.310 115.815 89.560 116.075 ;
        RECT 88.550 115.645 88.800 115.805 ;
        RECT 89.730 115.645 89.900 116.490 ;
        RECT 90.795 116.205 90.965 116.705 ;
        RECT 91.135 116.375 91.465 116.875 ;
        RECT 90.070 115.815 90.570 116.195 ;
        RECT 90.795 116.035 91.490 116.205 ;
        RECT 88.550 115.475 89.900 115.645 ;
        RECT 89.480 115.435 89.900 115.475 ;
        RECT 88.190 114.965 88.610 115.305 ;
        RECT 88.900 114.975 89.310 115.305 ;
        RECT 86.430 114.545 87.280 114.715 ;
        RECT 87.840 114.325 88.160 114.785 ;
        RECT 88.360 114.535 88.610 114.965 ;
        RECT 88.900 114.325 89.310 114.765 ;
        RECT 89.480 114.705 89.650 115.435 ;
        RECT 89.820 114.885 90.170 115.255 ;
        RECT 90.350 114.945 90.570 115.815 ;
        RECT 90.740 115.245 91.150 115.865 ;
        RECT 91.320 115.065 91.490 116.035 ;
        RECT 90.795 114.875 91.490 115.065 ;
        RECT 89.480 114.505 90.495 114.705 ;
        RECT 90.795 114.545 90.965 114.875 ;
        RECT 91.135 114.325 91.465 114.705 ;
        RECT 91.680 114.585 91.905 116.705 ;
        RECT 92.075 116.375 92.405 116.875 ;
        RECT 92.575 116.205 92.745 116.705 ;
        RECT 92.080 116.035 92.745 116.205 ;
        RECT 92.080 115.045 92.310 116.035 ;
        RECT 92.480 115.215 92.830 115.865 ;
        RECT 93.005 115.785 95.595 116.875 ;
        RECT 93.005 115.095 94.215 115.615 ;
        RECT 94.385 115.265 95.595 115.785 ;
        RECT 95.765 115.710 96.055 116.875 ;
        RECT 96.235 115.895 96.565 116.705 ;
        RECT 96.735 116.075 96.975 116.875 ;
        RECT 96.235 115.725 96.950 115.895 ;
        RECT 96.230 115.315 96.610 115.555 ;
        RECT 96.780 115.485 96.950 115.725 ;
        RECT 97.155 115.855 97.325 116.705 ;
        RECT 97.495 116.075 97.825 116.875 ;
        RECT 97.995 115.855 98.165 116.705 ;
        RECT 97.155 115.685 98.165 115.855 ;
        RECT 98.335 115.725 98.665 116.875 ;
        RECT 99.505 115.735 99.715 116.875 ;
        RECT 99.885 115.725 100.215 116.705 ;
        RECT 100.385 115.735 100.615 116.875 ;
        RECT 100.825 115.785 103.415 116.875 ;
        RECT 97.670 115.515 98.165 115.685 ;
        RECT 96.780 115.315 97.280 115.485 ;
        RECT 97.665 115.345 98.165 115.515 ;
        RECT 96.780 115.145 96.950 115.315 ;
        RECT 97.670 115.145 98.165 115.345 ;
        RECT 92.080 114.875 92.745 115.045 ;
        RECT 92.075 114.325 92.405 114.705 ;
        RECT 92.575 114.585 92.745 114.875 ;
        RECT 93.005 114.325 95.595 115.095 ;
        RECT 95.765 114.325 96.055 115.050 ;
        RECT 96.315 114.975 96.950 115.145 ;
        RECT 97.155 114.975 98.165 115.145 ;
        RECT 96.315 114.495 96.485 114.975 ;
        RECT 96.665 114.325 96.905 114.805 ;
        RECT 97.155 114.495 97.325 114.975 ;
        RECT 97.495 114.325 97.825 114.805 ;
        RECT 97.995 114.495 98.165 114.975 ;
        RECT 98.335 114.325 98.665 115.125 ;
        RECT 99.505 114.325 99.715 115.145 ;
        RECT 99.885 115.125 100.135 115.725 ;
        RECT 100.305 115.315 100.635 115.565 ;
        RECT 99.885 114.495 100.215 115.125 ;
        RECT 100.385 114.325 100.615 115.145 ;
        RECT 100.825 115.095 102.035 115.615 ;
        RECT 102.205 115.265 103.415 115.785 ;
        RECT 103.675 115.945 103.845 116.705 ;
        RECT 104.025 116.115 104.355 116.875 ;
        RECT 103.675 115.775 104.340 115.945 ;
        RECT 104.525 115.800 104.795 116.705 ;
        RECT 104.965 116.440 110.310 116.875 ;
        RECT 104.170 115.630 104.340 115.775 ;
        RECT 103.605 115.225 103.935 115.595 ;
        RECT 104.170 115.300 104.455 115.630 ;
        RECT 100.825 114.325 103.415 115.095 ;
        RECT 104.170 115.045 104.340 115.300 ;
        RECT 103.675 114.875 104.340 115.045 ;
        RECT 104.625 115.000 104.795 115.800 ;
        RECT 103.675 114.495 103.845 114.875 ;
        RECT 104.025 114.325 104.355 114.705 ;
        RECT 104.535 114.495 104.795 115.000 ;
        RECT 106.550 114.870 106.890 115.700 ;
        RECT 108.370 115.190 108.720 116.440 ;
        RECT 110.485 115.785 111.695 116.875 ;
        RECT 111.955 116.205 112.125 116.705 ;
        RECT 112.295 116.375 112.625 116.875 ;
        RECT 111.955 116.035 112.620 116.205 ;
        RECT 110.485 115.075 111.005 115.615 ;
        RECT 111.175 115.245 111.695 115.785 ;
        RECT 111.870 115.215 112.220 115.865 ;
        RECT 104.965 114.325 110.310 114.870 ;
        RECT 110.485 114.325 111.695 115.075 ;
        RECT 112.390 115.045 112.620 116.035 ;
        RECT 111.955 114.875 112.620 115.045 ;
        RECT 111.955 114.585 112.125 114.875 ;
        RECT 112.295 114.325 112.625 114.705 ;
        RECT 112.795 114.585 113.020 116.705 ;
        RECT 113.235 116.375 113.565 116.875 ;
        RECT 113.735 116.205 113.905 116.705 ;
        RECT 114.140 116.490 114.970 116.660 ;
        RECT 115.210 116.495 115.590 116.875 ;
        RECT 113.210 116.035 113.905 116.205 ;
        RECT 113.210 115.065 113.380 116.035 ;
        RECT 113.550 115.245 113.960 115.865 ;
        RECT 114.130 115.815 114.630 116.195 ;
        RECT 113.210 114.875 113.905 115.065 ;
        RECT 114.130 114.945 114.350 115.815 ;
        RECT 114.800 115.645 114.970 116.490 ;
        RECT 115.770 116.325 115.940 116.615 ;
        RECT 116.110 116.495 116.440 116.875 ;
        RECT 116.910 116.405 117.540 116.655 ;
        RECT 117.720 116.495 118.140 116.875 ;
        RECT 117.370 116.325 117.540 116.405 ;
        RECT 118.340 116.325 118.580 116.615 ;
        RECT 115.140 116.075 116.510 116.325 ;
        RECT 115.140 115.815 115.390 116.075 ;
        RECT 115.900 115.645 116.150 115.805 ;
        RECT 114.800 115.475 116.150 115.645 ;
        RECT 114.800 115.435 115.220 115.475 ;
        RECT 114.530 114.885 114.880 115.255 ;
        RECT 113.235 114.325 113.565 114.705 ;
        RECT 113.735 114.545 113.905 114.875 ;
        RECT 115.050 114.705 115.220 115.435 ;
        RECT 116.320 115.305 116.510 116.075 ;
        RECT 115.390 114.975 115.800 115.305 ;
        RECT 116.090 114.965 116.510 115.305 ;
        RECT 116.680 115.895 117.200 116.205 ;
        RECT 117.370 116.155 118.580 116.325 ;
        RECT 118.810 116.185 119.140 116.875 ;
        RECT 116.680 115.135 116.850 115.895 ;
        RECT 117.020 115.305 117.200 115.715 ;
        RECT 117.370 115.645 117.540 116.155 ;
        RECT 119.310 116.005 119.480 116.615 ;
        RECT 119.750 116.155 120.080 116.665 ;
        RECT 119.310 115.985 119.630 116.005 ;
        RECT 117.710 115.815 119.630 115.985 ;
        RECT 117.370 115.475 119.270 115.645 ;
        RECT 117.600 115.135 117.930 115.255 ;
        RECT 116.680 114.965 117.930 115.135 ;
        RECT 114.205 114.505 115.220 114.705 ;
        RECT 115.390 114.325 115.800 114.765 ;
        RECT 116.090 114.535 116.340 114.965 ;
        RECT 116.540 114.325 116.860 114.785 ;
        RECT 118.100 114.715 118.270 115.475 ;
        RECT 118.940 115.415 119.270 115.475 ;
        RECT 118.460 115.245 118.790 115.305 ;
        RECT 118.460 114.975 119.120 115.245 ;
        RECT 119.440 114.920 119.630 115.815 ;
        RECT 117.420 114.545 118.270 114.715 ;
        RECT 118.470 114.325 119.130 114.805 ;
        RECT 119.310 114.590 119.630 114.920 ;
        RECT 119.830 115.565 120.080 116.155 ;
        RECT 120.260 116.075 120.545 116.875 ;
        RECT 120.725 115.895 120.980 116.565 ;
        RECT 119.830 115.235 120.630 115.565 ;
        RECT 119.830 114.585 120.080 115.235 ;
        RECT 120.800 115.035 120.980 115.895 ;
        RECT 121.525 115.710 121.815 116.875 ;
        RECT 121.985 115.785 123.655 116.875 ;
        RECT 121.985 115.095 122.735 115.615 ;
        RECT 122.905 115.265 123.655 115.785 ;
        RECT 124.285 115.785 125.495 116.875 ;
        RECT 124.285 115.245 124.805 115.785 ;
        RECT 120.725 114.835 120.980 115.035 ;
        RECT 120.260 114.325 120.545 114.785 ;
        RECT 120.725 114.665 121.065 114.835 ;
        RECT 120.725 114.505 120.980 114.665 ;
        RECT 121.525 114.325 121.815 115.050 ;
        RECT 121.985 114.325 123.655 115.095 ;
        RECT 124.975 115.075 125.495 115.615 ;
        RECT 124.285 114.325 125.495 115.075 ;
        RECT 5.520 114.155 125.580 114.325 ;
        RECT 5.605 113.405 6.815 114.155 ;
        RECT 5.605 112.865 6.125 113.405 ;
        RECT 6.985 113.385 10.495 114.155 ;
        RECT 11.675 113.605 11.845 113.895 ;
        RECT 12.015 113.775 12.345 114.155 ;
        RECT 11.675 113.435 12.340 113.605 ;
        RECT 6.295 112.695 6.815 113.235 ;
        RECT 6.985 112.865 8.635 113.385 ;
        RECT 8.805 112.695 10.495 113.215 ;
        RECT 5.605 111.605 6.815 112.695 ;
        RECT 6.985 111.605 10.495 112.695 ;
        RECT 11.590 112.615 11.940 113.265 ;
        RECT 12.110 112.445 12.340 113.435 ;
        RECT 11.675 112.275 12.340 112.445 ;
        RECT 11.675 111.775 11.845 112.275 ;
        RECT 12.015 111.605 12.345 112.105 ;
        RECT 12.515 111.775 12.740 113.895 ;
        RECT 12.955 113.775 13.285 114.155 ;
        RECT 13.455 113.605 13.625 113.935 ;
        RECT 13.925 113.775 14.940 113.975 ;
        RECT 12.930 113.415 13.625 113.605 ;
        RECT 12.930 112.445 13.100 113.415 ;
        RECT 13.270 112.615 13.680 113.235 ;
        RECT 13.850 112.665 14.070 113.535 ;
        RECT 14.250 113.225 14.600 113.595 ;
        RECT 14.770 113.045 14.940 113.775 ;
        RECT 15.110 113.715 15.520 114.155 ;
        RECT 15.810 113.515 16.060 113.945 ;
        RECT 16.260 113.695 16.580 114.155 ;
        RECT 17.140 113.765 17.990 113.935 ;
        RECT 15.110 113.175 15.520 113.505 ;
        RECT 15.810 113.175 16.230 113.515 ;
        RECT 14.520 113.005 14.940 113.045 ;
        RECT 14.520 112.835 15.870 113.005 ;
        RECT 12.930 112.275 13.625 112.445 ;
        RECT 13.850 112.285 14.350 112.665 ;
        RECT 12.955 111.605 13.285 112.105 ;
        RECT 13.455 111.775 13.625 112.275 ;
        RECT 14.520 111.990 14.690 112.835 ;
        RECT 15.620 112.675 15.870 112.835 ;
        RECT 14.860 112.405 15.110 112.665 ;
        RECT 16.040 112.405 16.230 113.175 ;
        RECT 14.860 112.155 16.230 112.405 ;
        RECT 16.400 113.345 17.650 113.515 ;
        RECT 16.400 112.585 16.570 113.345 ;
        RECT 17.320 113.225 17.650 113.345 ;
        RECT 16.740 112.765 16.920 113.175 ;
        RECT 17.820 113.005 17.990 113.765 ;
        RECT 18.190 113.675 18.850 114.155 ;
        RECT 19.030 113.560 19.350 113.890 ;
        RECT 18.180 113.235 18.840 113.505 ;
        RECT 18.180 113.175 18.510 113.235 ;
        RECT 18.660 113.005 18.990 113.065 ;
        RECT 17.090 112.835 18.990 113.005 ;
        RECT 16.400 112.275 16.920 112.585 ;
        RECT 17.090 112.325 17.260 112.835 ;
        RECT 19.160 112.665 19.350 113.560 ;
        RECT 17.430 112.495 19.350 112.665 ;
        RECT 19.030 112.475 19.350 112.495 ;
        RECT 19.550 113.245 19.800 113.895 ;
        RECT 19.980 113.695 20.265 114.155 ;
        RECT 20.445 113.445 20.700 113.975 ;
        RECT 19.550 112.915 20.350 113.245 ;
        RECT 17.090 112.155 18.300 112.325 ;
        RECT 13.860 111.820 14.690 111.990 ;
        RECT 14.930 111.605 15.310 111.985 ;
        RECT 15.490 111.865 15.660 112.155 ;
        RECT 17.090 112.075 17.260 112.155 ;
        RECT 15.830 111.605 16.160 111.985 ;
        RECT 16.630 111.825 17.260 112.075 ;
        RECT 17.440 111.605 17.860 111.985 ;
        RECT 18.060 111.865 18.300 112.155 ;
        RECT 18.530 111.605 18.860 112.295 ;
        RECT 19.030 111.865 19.200 112.475 ;
        RECT 19.550 112.325 19.800 112.915 ;
        RECT 20.520 112.585 20.700 113.445 ;
        RECT 21.795 113.605 21.965 113.895 ;
        RECT 22.135 113.775 22.465 114.155 ;
        RECT 21.795 113.435 22.460 113.605 ;
        RECT 21.710 112.615 22.060 113.265 ;
        RECT 19.470 111.815 19.800 112.325 ;
        RECT 19.980 111.605 20.265 112.405 ;
        RECT 20.445 112.115 20.700 112.585 ;
        RECT 22.230 112.445 22.460 113.435 ;
        RECT 21.795 112.275 22.460 112.445 ;
        RECT 20.445 111.945 20.785 112.115 ;
        RECT 20.445 111.915 20.700 111.945 ;
        RECT 21.795 111.775 21.965 112.275 ;
        RECT 22.135 111.605 22.465 112.105 ;
        RECT 22.635 111.775 22.860 113.895 ;
        RECT 23.075 113.775 23.405 114.155 ;
        RECT 23.575 113.605 23.745 113.935 ;
        RECT 24.045 113.775 25.060 113.975 ;
        RECT 23.050 113.415 23.745 113.605 ;
        RECT 23.050 112.445 23.220 113.415 ;
        RECT 23.390 112.615 23.800 113.235 ;
        RECT 23.970 112.665 24.190 113.535 ;
        RECT 24.370 113.225 24.720 113.595 ;
        RECT 24.890 113.045 25.060 113.775 ;
        RECT 25.230 113.715 25.640 114.155 ;
        RECT 25.930 113.515 26.180 113.945 ;
        RECT 26.380 113.695 26.700 114.155 ;
        RECT 27.260 113.765 28.110 113.935 ;
        RECT 25.230 113.175 25.640 113.505 ;
        RECT 25.930 113.175 26.350 113.515 ;
        RECT 24.640 113.005 25.060 113.045 ;
        RECT 24.640 112.835 25.990 113.005 ;
        RECT 23.050 112.275 23.745 112.445 ;
        RECT 23.970 112.285 24.470 112.665 ;
        RECT 23.075 111.605 23.405 112.105 ;
        RECT 23.575 111.775 23.745 112.275 ;
        RECT 24.640 111.990 24.810 112.835 ;
        RECT 25.740 112.675 25.990 112.835 ;
        RECT 24.980 112.405 25.230 112.665 ;
        RECT 26.160 112.405 26.350 113.175 ;
        RECT 24.980 112.155 26.350 112.405 ;
        RECT 26.520 113.345 27.770 113.515 ;
        RECT 26.520 112.585 26.690 113.345 ;
        RECT 27.440 113.225 27.770 113.345 ;
        RECT 26.860 112.765 27.040 113.175 ;
        RECT 27.940 113.005 28.110 113.765 ;
        RECT 28.310 113.675 28.970 114.155 ;
        RECT 29.150 113.560 29.470 113.890 ;
        RECT 28.300 113.235 28.960 113.505 ;
        RECT 28.300 113.175 28.630 113.235 ;
        RECT 28.780 113.005 29.110 113.065 ;
        RECT 27.210 112.835 29.110 113.005 ;
        RECT 26.520 112.275 27.040 112.585 ;
        RECT 27.210 112.325 27.380 112.835 ;
        RECT 29.280 112.665 29.470 113.560 ;
        RECT 27.550 112.495 29.470 112.665 ;
        RECT 29.150 112.475 29.470 112.495 ;
        RECT 29.670 113.245 29.920 113.895 ;
        RECT 30.100 113.695 30.385 114.155 ;
        RECT 30.565 113.445 30.820 113.975 ;
        RECT 29.670 112.915 30.470 113.245 ;
        RECT 27.210 112.155 28.420 112.325 ;
        RECT 23.980 111.820 24.810 111.990 ;
        RECT 25.050 111.605 25.430 111.985 ;
        RECT 25.610 111.865 25.780 112.155 ;
        RECT 27.210 112.075 27.380 112.155 ;
        RECT 25.950 111.605 26.280 111.985 ;
        RECT 26.750 111.825 27.380 112.075 ;
        RECT 27.560 111.605 27.980 111.985 ;
        RECT 28.180 111.865 28.420 112.155 ;
        RECT 28.650 111.605 28.980 112.295 ;
        RECT 29.150 111.865 29.320 112.475 ;
        RECT 29.670 112.325 29.920 112.915 ;
        RECT 30.640 112.585 30.820 113.445 ;
        RECT 31.365 113.430 31.655 114.155 ;
        RECT 31.830 113.415 32.085 113.985 ;
        RECT 32.255 113.755 32.585 114.155 ;
        RECT 33.010 113.620 33.540 113.985 ;
        RECT 33.010 113.585 33.185 113.620 ;
        RECT 32.255 113.415 33.185 113.585 ;
        RECT 30.565 112.455 30.820 112.585 ;
        RECT 29.590 111.815 29.920 112.325 ;
        RECT 30.100 111.605 30.385 112.405 ;
        RECT 30.565 112.285 30.905 112.455 ;
        RECT 30.565 111.915 30.820 112.285 ;
        RECT 31.365 111.605 31.655 112.770 ;
        RECT 31.830 112.745 32.000 113.415 ;
        RECT 32.255 113.245 32.425 113.415 ;
        RECT 32.170 112.915 32.425 113.245 ;
        RECT 32.650 112.915 32.845 113.245 ;
        RECT 31.830 111.775 32.165 112.745 ;
        RECT 32.335 111.605 32.505 112.745 ;
        RECT 32.675 111.945 32.845 112.915 ;
        RECT 33.015 112.285 33.185 113.415 ;
        RECT 33.355 112.625 33.525 113.425 ;
        RECT 33.730 113.135 34.005 113.985 ;
        RECT 33.725 112.965 34.005 113.135 ;
        RECT 33.730 112.825 34.005 112.965 ;
        RECT 34.175 112.625 34.365 113.985 ;
        RECT 34.545 113.620 35.055 114.155 ;
        RECT 35.275 113.345 35.520 113.950 ;
        RECT 35.965 113.480 36.225 113.985 ;
        RECT 36.405 113.775 36.735 114.155 ;
        RECT 36.915 113.605 37.085 113.985 ;
        RECT 34.565 113.175 35.795 113.345 ;
        RECT 33.355 112.455 34.365 112.625 ;
        RECT 34.535 112.610 35.285 112.800 ;
        RECT 33.015 112.115 34.140 112.285 ;
        RECT 34.535 111.945 34.705 112.610 ;
        RECT 35.455 112.365 35.795 113.175 ;
        RECT 32.675 111.775 34.705 111.945 ;
        RECT 34.875 111.605 35.045 112.365 ;
        RECT 35.280 111.955 35.795 112.365 ;
        RECT 35.965 112.680 36.135 113.480 ;
        RECT 36.420 113.435 37.085 113.605 ;
        RECT 36.420 113.180 36.590 113.435 ;
        RECT 37.345 113.405 38.555 114.155 ;
        RECT 38.815 113.605 38.985 113.985 ;
        RECT 39.165 113.775 39.495 114.155 ;
        RECT 38.815 113.435 39.480 113.605 ;
        RECT 39.675 113.480 39.935 113.985 ;
        RECT 36.305 112.850 36.590 113.180 ;
        RECT 36.825 112.885 37.155 113.255 ;
        RECT 37.345 112.865 37.865 113.405 ;
        RECT 36.420 112.705 36.590 112.850 ;
        RECT 35.965 111.775 36.235 112.680 ;
        RECT 36.420 112.535 37.085 112.705 ;
        RECT 38.035 112.695 38.555 113.235 ;
        RECT 38.745 112.885 39.075 113.255 ;
        RECT 39.310 113.180 39.480 113.435 ;
        RECT 39.310 112.850 39.595 113.180 ;
        RECT 39.310 112.705 39.480 112.850 ;
        RECT 36.405 111.605 36.735 112.365 ;
        RECT 36.915 111.775 37.085 112.535 ;
        RECT 37.345 111.605 38.555 112.695 ;
        RECT 38.815 112.535 39.480 112.705 ;
        RECT 39.765 112.680 39.935 113.480 ;
        RECT 40.165 113.335 40.375 114.155 ;
        RECT 40.545 113.355 40.875 113.985 ;
        RECT 40.545 112.755 40.795 113.355 ;
        RECT 41.045 113.335 41.275 114.155 ;
        RECT 41.960 113.630 42.255 114.155 ;
        RECT 42.425 113.515 42.650 113.960 ;
        RECT 42.820 113.685 43.150 114.155 ;
        RECT 42.425 113.345 43.155 113.515 ;
        RECT 43.700 113.475 43.955 113.975 ;
        RECT 44.135 113.695 44.420 114.155 ;
        RECT 40.965 112.915 41.295 113.165 ;
        RECT 41.485 112.950 42.705 113.175 ;
        RECT 42.875 112.780 43.155 113.345 ;
        RECT 43.615 113.445 43.955 113.475 ;
        RECT 43.615 113.305 43.880 113.445 ;
        RECT 38.815 111.775 38.985 112.535 ;
        RECT 39.165 111.605 39.495 112.365 ;
        RECT 39.665 111.775 39.935 112.680 ;
        RECT 40.165 111.605 40.375 112.745 ;
        RECT 40.545 111.775 40.875 112.755 ;
        RECT 41.045 111.605 41.275 112.745 ;
        RECT 41.555 112.610 43.155 112.780 ;
        RECT 41.555 111.805 41.810 112.610 ;
        RECT 41.980 111.605 42.240 112.440 ;
        RECT 42.410 111.805 42.670 112.610 ;
        RECT 43.700 112.585 43.880 113.305 ;
        RECT 44.600 113.245 44.850 113.895 ;
        RECT 44.050 112.915 44.850 113.245 ;
        RECT 42.840 111.605 43.095 112.440 ;
        RECT 43.700 111.915 43.955 112.585 ;
        RECT 44.135 111.605 44.420 112.405 ;
        RECT 44.600 112.325 44.850 112.915 ;
        RECT 45.050 113.560 45.370 113.890 ;
        RECT 45.550 113.675 46.210 114.155 ;
        RECT 46.410 113.765 47.260 113.935 ;
        RECT 45.050 112.665 45.240 113.560 ;
        RECT 45.560 113.235 46.220 113.505 ;
        RECT 45.890 113.175 46.220 113.235 ;
        RECT 45.410 113.005 45.740 113.065 ;
        RECT 46.410 113.005 46.580 113.765 ;
        RECT 47.820 113.695 48.140 114.155 ;
        RECT 48.340 113.515 48.590 113.945 ;
        RECT 48.880 113.715 49.290 114.155 ;
        RECT 49.460 113.775 50.475 113.975 ;
        RECT 46.750 113.345 48.000 113.515 ;
        RECT 46.750 113.225 47.080 113.345 ;
        RECT 45.410 112.835 47.310 113.005 ;
        RECT 45.050 112.495 46.970 112.665 ;
        RECT 45.050 112.475 45.370 112.495 ;
        RECT 44.600 111.815 44.930 112.325 ;
        RECT 45.200 111.865 45.370 112.475 ;
        RECT 47.140 112.325 47.310 112.835 ;
        RECT 47.480 112.765 47.660 113.175 ;
        RECT 47.830 112.585 48.000 113.345 ;
        RECT 45.540 111.605 45.870 112.295 ;
        RECT 46.100 112.155 47.310 112.325 ;
        RECT 47.480 112.275 48.000 112.585 ;
        RECT 48.170 113.175 48.590 113.515 ;
        RECT 48.880 113.175 49.290 113.505 ;
        RECT 48.170 112.405 48.360 113.175 ;
        RECT 49.460 113.045 49.630 113.775 ;
        RECT 50.775 113.605 50.945 113.935 ;
        RECT 51.115 113.775 51.445 114.155 ;
        RECT 49.800 113.225 50.150 113.595 ;
        RECT 49.460 113.005 49.880 113.045 ;
        RECT 48.530 112.835 49.880 113.005 ;
        RECT 48.530 112.675 48.780 112.835 ;
        RECT 49.290 112.405 49.540 112.665 ;
        RECT 48.170 112.155 49.540 112.405 ;
        RECT 46.100 111.865 46.340 112.155 ;
        RECT 47.140 112.075 47.310 112.155 ;
        RECT 46.540 111.605 46.960 111.985 ;
        RECT 47.140 111.825 47.770 112.075 ;
        RECT 48.240 111.605 48.570 111.985 ;
        RECT 48.740 111.865 48.910 112.155 ;
        RECT 49.710 111.990 49.880 112.835 ;
        RECT 50.330 112.665 50.550 113.535 ;
        RECT 50.775 113.415 51.470 113.605 ;
        RECT 50.050 112.285 50.550 112.665 ;
        RECT 50.720 112.615 51.130 113.235 ;
        RECT 51.300 112.445 51.470 113.415 ;
        RECT 50.775 112.275 51.470 112.445 ;
        RECT 49.090 111.605 49.470 111.985 ;
        RECT 49.710 111.820 50.540 111.990 ;
        RECT 50.775 111.775 50.945 112.275 ;
        RECT 51.115 111.605 51.445 112.105 ;
        RECT 51.660 111.775 51.885 113.895 ;
        RECT 52.055 113.775 52.385 114.155 ;
        RECT 52.555 113.605 52.725 113.895 ;
        RECT 52.060 113.435 52.725 113.605 ;
        RECT 52.060 112.445 52.290 113.435 ;
        RECT 53.260 113.345 53.505 113.950 ;
        RECT 53.725 113.620 54.235 114.155 ;
        RECT 52.460 112.615 52.810 113.265 ;
        RECT 52.985 113.175 54.215 113.345 ;
        RECT 52.060 112.275 52.725 112.445 ;
        RECT 52.055 111.605 52.385 112.105 ;
        RECT 52.555 111.775 52.725 112.275 ;
        RECT 52.985 112.365 53.325 113.175 ;
        RECT 53.495 112.610 54.245 112.800 ;
        RECT 52.985 111.955 53.500 112.365 ;
        RECT 53.735 111.605 53.905 112.365 ;
        RECT 54.075 111.945 54.245 112.610 ;
        RECT 54.415 112.625 54.605 113.985 ;
        RECT 54.775 113.135 55.050 113.985 ;
        RECT 55.240 113.620 55.770 113.985 ;
        RECT 56.195 113.755 56.525 114.155 ;
        RECT 55.595 113.585 55.770 113.620 ;
        RECT 54.775 112.965 55.055 113.135 ;
        RECT 54.775 112.825 55.050 112.965 ;
        RECT 55.255 112.625 55.425 113.425 ;
        RECT 54.415 112.455 55.425 112.625 ;
        RECT 55.595 113.415 56.525 113.585 ;
        RECT 56.695 113.415 56.950 113.985 ;
        RECT 57.125 113.430 57.415 114.155 ;
        RECT 57.960 113.445 58.215 113.975 ;
        RECT 58.395 113.695 58.680 114.155 ;
        RECT 55.595 112.285 55.765 113.415 ;
        RECT 56.355 113.245 56.525 113.415 ;
        RECT 54.640 112.115 55.765 112.285 ;
        RECT 55.935 112.915 56.130 113.245 ;
        RECT 56.355 112.915 56.610 113.245 ;
        RECT 55.935 111.945 56.105 112.915 ;
        RECT 56.780 112.745 56.950 113.415 ;
        RECT 54.075 111.775 56.105 111.945 ;
        RECT 56.275 111.605 56.445 112.745 ;
        RECT 56.615 111.775 56.950 112.745 ;
        RECT 57.125 111.605 57.415 112.770 ;
        RECT 57.960 112.585 58.140 113.445 ;
        RECT 58.860 113.245 59.110 113.895 ;
        RECT 58.310 112.915 59.110 113.245 ;
        RECT 57.960 112.115 58.215 112.585 ;
        RECT 57.875 111.945 58.215 112.115 ;
        RECT 57.960 111.915 58.215 111.945 ;
        RECT 58.395 111.605 58.680 112.405 ;
        RECT 58.860 112.325 59.110 112.915 ;
        RECT 59.310 113.560 59.630 113.890 ;
        RECT 59.810 113.675 60.470 114.155 ;
        RECT 60.670 113.765 61.520 113.935 ;
        RECT 59.310 112.665 59.500 113.560 ;
        RECT 59.820 113.235 60.480 113.505 ;
        RECT 60.150 113.175 60.480 113.235 ;
        RECT 59.670 113.005 60.000 113.065 ;
        RECT 60.670 113.005 60.840 113.765 ;
        RECT 62.080 113.695 62.400 114.155 ;
        RECT 62.600 113.515 62.850 113.945 ;
        RECT 63.140 113.715 63.550 114.155 ;
        RECT 63.720 113.775 64.735 113.975 ;
        RECT 61.010 113.345 62.260 113.515 ;
        RECT 61.010 113.225 61.340 113.345 ;
        RECT 59.670 112.835 61.570 113.005 ;
        RECT 59.310 112.495 61.230 112.665 ;
        RECT 59.310 112.475 59.630 112.495 ;
        RECT 58.860 111.815 59.190 112.325 ;
        RECT 59.460 111.865 59.630 112.475 ;
        RECT 61.400 112.325 61.570 112.835 ;
        RECT 61.740 112.765 61.920 113.175 ;
        RECT 62.090 112.585 62.260 113.345 ;
        RECT 59.800 111.605 60.130 112.295 ;
        RECT 60.360 112.155 61.570 112.325 ;
        RECT 61.740 112.275 62.260 112.585 ;
        RECT 62.430 113.175 62.850 113.515 ;
        RECT 63.140 113.175 63.550 113.505 ;
        RECT 62.430 112.405 62.620 113.175 ;
        RECT 63.720 113.045 63.890 113.775 ;
        RECT 65.035 113.605 65.205 113.935 ;
        RECT 65.375 113.775 65.705 114.155 ;
        RECT 64.060 113.225 64.410 113.595 ;
        RECT 63.720 113.005 64.140 113.045 ;
        RECT 62.790 112.835 64.140 113.005 ;
        RECT 62.790 112.675 63.040 112.835 ;
        RECT 63.550 112.405 63.800 112.665 ;
        RECT 62.430 112.155 63.800 112.405 ;
        RECT 60.360 111.865 60.600 112.155 ;
        RECT 61.400 112.075 61.570 112.155 ;
        RECT 60.800 111.605 61.220 111.985 ;
        RECT 61.400 111.825 62.030 112.075 ;
        RECT 62.500 111.605 62.830 111.985 ;
        RECT 63.000 111.865 63.170 112.155 ;
        RECT 63.970 111.990 64.140 112.835 ;
        RECT 64.590 112.665 64.810 113.535 ;
        RECT 65.035 113.415 65.730 113.605 ;
        RECT 64.310 112.285 64.810 112.665 ;
        RECT 64.980 112.615 65.390 113.235 ;
        RECT 65.560 112.445 65.730 113.415 ;
        RECT 65.035 112.275 65.730 112.445 ;
        RECT 63.350 111.605 63.730 111.985 ;
        RECT 63.970 111.820 64.800 111.990 ;
        RECT 65.035 111.775 65.205 112.275 ;
        RECT 65.375 111.605 65.705 112.105 ;
        RECT 65.920 111.775 66.145 113.895 ;
        RECT 66.315 113.775 66.645 114.155 ;
        RECT 66.815 113.605 66.985 113.895 ;
        RECT 66.320 113.435 66.985 113.605 ;
        RECT 66.320 112.445 66.550 113.435 ;
        RECT 67.245 113.385 69.835 114.155 ;
        RECT 70.095 113.605 70.265 113.895 ;
        RECT 70.435 113.775 70.765 114.155 ;
        RECT 70.095 113.435 70.760 113.605 ;
        RECT 66.720 112.615 67.070 113.265 ;
        RECT 67.245 112.865 68.455 113.385 ;
        RECT 68.625 112.695 69.835 113.215 ;
        RECT 66.320 112.275 66.985 112.445 ;
        RECT 66.315 111.605 66.645 112.105 ;
        RECT 66.815 111.775 66.985 112.275 ;
        RECT 67.245 111.605 69.835 112.695 ;
        RECT 70.010 112.615 70.360 113.265 ;
        RECT 70.530 112.445 70.760 113.435 ;
        RECT 70.095 112.275 70.760 112.445 ;
        RECT 70.095 111.775 70.265 112.275 ;
        RECT 70.435 111.605 70.765 112.105 ;
        RECT 70.935 111.775 71.160 113.895 ;
        RECT 71.375 113.775 71.705 114.155 ;
        RECT 71.875 113.605 72.045 113.935 ;
        RECT 72.345 113.775 73.360 113.975 ;
        RECT 71.350 113.415 72.045 113.605 ;
        RECT 71.350 112.445 71.520 113.415 ;
        RECT 71.690 112.615 72.100 113.235 ;
        RECT 72.270 112.665 72.490 113.535 ;
        RECT 72.670 113.225 73.020 113.595 ;
        RECT 73.190 113.045 73.360 113.775 ;
        RECT 73.530 113.715 73.940 114.155 ;
        RECT 74.230 113.515 74.480 113.945 ;
        RECT 74.680 113.695 75.000 114.155 ;
        RECT 75.560 113.765 76.410 113.935 ;
        RECT 73.530 113.175 73.940 113.505 ;
        RECT 74.230 113.175 74.650 113.515 ;
        RECT 72.940 113.005 73.360 113.045 ;
        RECT 72.940 112.835 74.290 113.005 ;
        RECT 71.350 112.275 72.045 112.445 ;
        RECT 72.270 112.285 72.770 112.665 ;
        RECT 71.375 111.605 71.705 112.105 ;
        RECT 71.875 111.775 72.045 112.275 ;
        RECT 72.940 111.990 73.110 112.835 ;
        RECT 74.040 112.675 74.290 112.835 ;
        RECT 73.280 112.405 73.530 112.665 ;
        RECT 74.460 112.405 74.650 113.175 ;
        RECT 73.280 112.155 74.650 112.405 ;
        RECT 74.820 113.345 76.070 113.515 ;
        RECT 74.820 112.585 74.990 113.345 ;
        RECT 75.740 113.225 76.070 113.345 ;
        RECT 75.160 112.765 75.340 113.175 ;
        RECT 76.240 113.005 76.410 113.765 ;
        RECT 76.610 113.675 77.270 114.155 ;
        RECT 77.450 113.560 77.770 113.890 ;
        RECT 76.600 113.235 77.260 113.505 ;
        RECT 76.600 113.175 76.930 113.235 ;
        RECT 77.080 113.005 77.410 113.065 ;
        RECT 75.510 112.835 77.410 113.005 ;
        RECT 74.820 112.275 75.340 112.585 ;
        RECT 75.510 112.325 75.680 112.835 ;
        RECT 77.580 112.665 77.770 113.560 ;
        RECT 75.850 112.495 77.770 112.665 ;
        RECT 77.450 112.475 77.770 112.495 ;
        RECT 77.970 113.245 78.220 113.895 ;
        RECT 78.400 113.695 78.685 114.155 ;
        RECT 78.865 113.445 79.120 113.975 ;
        RECT 77.970 112.915 78.770 113.245 ;
        RECT 75.510 112.155 76.720 112.325 ;
        RECT 72.280 111.820 73.110 111.990 ;
        RECT 73.350 111.605 73.730 111.985 ;
        RECT 73.910 111.865 74.080 112.155 ;
        RECT 75.510 112.075 75.680 112.155 ;
        RECT 74.250 111.605 74.580 111.985 ;
        RECT 75.050 111.825 75.680 112.075 ;
        RECT 75.860 111.605 76.280 111.985 ;
        RECT 76.480 111.865 76.720 112.155 ;
        RECT 76.950 111.605 77.280 112.295 ;
        RECT 77.450 111.865 77.620 112.475 ;
        RECT 77.970 112.325 78.220 112.915 ;
        RECT 78.940 112.585 79.120 113.445 ;
        RECT 79.665 113.385 82.255 114.155 ;
        RECT 82.885 113.430 83.175 114.155 ;
        RECT 79.665 112.865 80.875 113.385 ;
        RECT 83.385 113.335 83.615 114.155 ;
        RECT 83.785 113.355 84.115 113.985 ;
        RECT 81.045 112.695 82.255 113.215 ;
        RECT 83.365 112.915 83.695 113.165 ;
        RECT 77.890 111.815 78.220 112.325 ;
        RECT 78.400 111.605 78.685 112.405 ;
        RECT 78.865 112.115 79.120 112.585 ;
        RECT 78.865 111.945 79.205 112.115 ;
        RECT 78.865 111.915 79.120 111.945 ;
        RECT 79.665 111.605 82.255 112.695 ;
        RECT 82.885 111.605 83.175 112.770 ;
        RECT 83.865 112.755 84.115 113.355 ;
        RECT 84.285 113.335 84.495 114.155 ;
        RECT 85.000 113.345 85.245 113.950 ;
        RECT 85.465 113.620 85.975 114.155 ;
        RECT 83.385 111.605 83.615 112.745 ;
        RECT 83.785 111.775 84.115 112.755 ;
        RECT 84.725 113.175 85.955 113.345 ;
        RECT 84.285 111.605 84.495 112.745 ;
        RECT 84.725 112.365 85.065 113.175 ;
        RECT 85.235 112.610 85.985 112.800 ;
        RECT 84.725 111.955 85.240 112.365 ;
        RECT 85.475 111.605 85.645 112.365 ;
        RECT 85.815 111.945 85.985 112.610 ;
        RECT 86.155 112.625 86.345 113.985 ;
        RECT 86.515 113.135 86.790 113.985 ;
        RECT 86.980 113.620 87.510 113.985 ;
        RECT 87.935 113.755 88.265 114.155 ;
        RECT 87.335 113.585 87.510 113.620 ;
        RECT 86.515 112.965 86.795 113.135 ;
        RECT 86.515 112.825 86.790 112.965 ;
        RECT 86.995 112.625 87.165 113.425 ;
        RECT 86.155 112.455 87.165 112.625 ;
        RECT 87.335 113.415 88.265 113.585 ;
        RECT 88.435 113.415 88.690 113.985 ;
        RECT 88.955 113.605 89.125 113.985 ;
        RECT 89.305 113.775 89.635 114.155 ;
        RECT 88.955 113.435 89.620 113.605 ;
        RECT 89.815 113.480 90.075 113.985 ;
        RECT 87.335 112.285 87.505 113.415 ;
        RECT 88.095 113.245 88.265 113.415 ;
        RECT 86.380 112.115 87.505 112.285 ;
        RECT 87.675 112.915 87.870 113.245 ;
        RECT 88.095 112.915 88.350 113.245 ;
        RECT 87.675 111.945 87.845 112.915 ;
        RECT 88.520 112.745 88.690 113.415 ;
        RECT 88.885 112.885 89.215 113.255 ;
        RECT 89.450 113.180 89.620 113.435 ;
        RECT 85.815 111.775 87.845 111.945 ;
        RECT 88.015 111.605 88.185 112.745 ;
        RECT 88.355 111.775 88.690 112.745 ;
        RECT 89.450 112.850 89.735 113.180 ;
        RECT 89.450 112.705 89.620 112.850 ;
        RECT 88.955 112.535 89.620 112.705 ;
        RECT 89.905 112.680 90.075 113.480 ;
        RECT 90.245 113.385 91.915 114.155 ;
        RECT 92.635 113.605 92.805 113.985 ;
        RECT 92.985 113.775 93.315 114.155 ;
        RECT 92.635 113.435 93.300 113.605 ;
        RECT 93.495 113.480 93.755 113.985 ;
        RECT 90.245 112.865 90.995 113.385 ;
        RECT 91.165 112.695 91.915 113.215 ;
        RECT 92.565 112.885 92.895 113.255 ;
        RECT 93.130 113.180 93.300 113.435 ;
        RECT 93.130 112.850 93.415 113.180 ;
        RECT 93.130 112.705 93.300 112.850 ;
        RECT 88.955 111.775 89.125 112.535 ;
        RECT 89.305 111.605 89.635 112.365 ;
        RECT 89.805 111.775 90.075 112.680 ;
        RECT 90.245 111.605 91.915 112.695 ;
        RECT 92.635 112.535 93.300 112.705 ;
        RECT 93.585 112.680 93.755 113.480 ;
        RECT 94.015 113.605 94.185 113.895 ;
        RECT 94.355 113.775 94.685 114.155 ;
        RECT 94.015 113.435 94.680 113.605 ;
        RECT 92.635 111.775 92.805 112.535 ;
        RECT 92.985 111.605 93.315 112.365 ;
        RECT 93.485 111.775 93.755 112.680 ;
        RECT 93.930 112.615 94.280 113.265 ;
        RECT 94.450 112.445 94.680 113.435 ;
        RECT 94.015 112.275 94.680 112.445 ;
        RECT 94.015 111.775 94.185 112.275 ;
        RECT 94.355 111.605 94.685 112.105 ;
        RECT 94.855 111.775 95.080 113.895 ;
        RECT 95.295 113.775 95.625 114.155 ;
        RECT 95.795 113.605 95.965 113.935 ;
        RECT 96.265 113.775 97.280 113.975 ;
        RECT 95.270 113.415 95.965 113.605 ;
        RECT 95.270 112.445 95.440 113.415 ;
        RECT 95.610 112.615 96.020 113.235 ;
        RECT 96.190 112.665 96.410 113.535 ;
        RECT 96.590 113.225 96.940 113.595 ;
        RECT 97.110 113.045 97.280 113.775 ;
        RECT 97.450 113.715 97.860 114.155 ;
        RECT 98.150 113.515 98.400 113.945 ;
        RECT 98.600 113.695 98.920 114.155 ;
        RECT 99.480 113.765 100.330 113.935 ;
        RECT 97.450 113.175 97.860 113.505 ;
        RECT 98.150 113.175 98.570 113.515 ;
        RECT 96.860 113.005 97.280 113.045 ;
        RECT 96.860 112.835 98.210 113.005 ;
        RECT 95.270 112.275 95.965 112.445 ;
        RECT 96.190 112.285 96.690 112.665 ;
        RECT 95.295 111.605 95.625 112.105 ;
        RECT 95.795 111.775 95.965 112.275 ;
        RECT 96.860 111.990 97.030 112.835 ;
        RECT 97.960 112.675 98.210 112.835 ;
        RECT 97.200 112.405 97.450 112.665 ;
        RECT 98.380 112.405 98.570 113.175 ;
        RECT 97.200 112.155 98.570 112.405 ;
        RECT 98.740 113.345 99.990 113.515 ;
        RECT 98.740 112.585 98.910 113.345 ;
        RECT 99.660 113.225 99.990 113.345 ;
        RECT 99.080 112.765 99.260 113.175 ;
        RECT 100.160 113.005 100.330 113.765 ;
        RECT 100.530 113.675 101.190 114.155 ;
        RECT 101.370 113.560 101.690 113.890 ;
        RECT 100.520 113.235 101.180 113.505 ;
        RECT 100.520 113.175 100.850 113.235 ;
        RECT 101.000 113.005 101.330 113.065 ;
        RECT 99.430 112.835 101.330 113.005 ;
        RECT 98.740 112.275 99.260 112.585 ;
        RECT 99.430 112.325 99.600 112.835 ;
        RECT 101.500 112.665 101.690 113.560 ;
        RECT 99.770 112.495 101.690 112.665 ;
        RECT 101.370 112.475 101.690 112.495 ;
        RECT 101.890 113.245 102.140 113.895 ;
        RECT 102.320 113.695 102.605 114.155 ;
        RECT 102.785 113.445 103.040 113.975 ;
        RECT 101.890 112.915 102.690 113.245 ;
        RECT 99.430 112.155 100.640 112.325 ;
        RECT 96.200 111.820 97.030 111.990 ;
        RECT 97.270 111.605 97.650 111.985 ;
        RECT 97.830 111.865 98.000 112.155 ;
        RECT 99.430 112.075 99.600 112.155 ;
        RECT 98.170 111.605 98.500 111.985 ;
        RECT 98.970 111.825 99.600 112.075 ;
        RECT 99.780 111.605 100.200 111.985 ;
        RECT 100.400 111.865 100.640 112.155 ;
        RECT 100.870 111.605 101.200 112.295 ;
        RECT 101.370 111.865 101.540 112.475 ;
        RECT 101.890 112.325 102.140 112.915 ;
        RECT 102.860 112.795 103.040 113.445 ;
        RECT 103.590 113.415 103.845 113.985 ;
        RECT 104.015 113.755 104.345 114.155 ;
        RECT 104.770 113.620 105.300 113.985 ;
        RECT 104.770 113.585 104.945 113.620 ;
        RECT 104.015 113.415 104.945 113.585 ;
        RECT 102.860 112.625 103.125 112.795 ;
        RECT 103.590 112.745 103.760 113.415 ;
        RECT 104.015 113.245 104.185 113.415 ;
        RECT 103.930 112.915 104.185 113.245 ;
        RECT 104.410 112.915 104.605 113.245 ;
        RECT 102.860 112.585 103.040 112.625 ;
        RECT 101.810 111.815 102.140 112.325 ;
        RECT 102.320 111.605 102.605 112.405 ;
        RECT 102.785 111.915 103.040 112.585 ;
        RECT 103.590 111.775 103.925 112.745 ;
        RECT 104.095 111.605 104.265 112.745 ;
        RECT 104.435 111.945 104.605 112.915 ;
        RECT 104.775 112.285 104.945 113.415 ;
        RECT 105.115 112.625 105.285 113.425 ;
        RECT 105.490 113.135 105.765 113.985 ;
        RECT 105.485 112.965 105.765 113.135 ;
        RECT 105.490 112.825 105.765 112.965 ;
        RECT 105.935 112.625 106.125 113.985 ;
        RECT 106.305 113.620 106.815 114.155 ;
        RECT 107.035 113.345 107.280 113.950 ;
        RECT 108.645 113.430 108.935 114.155 ;
        RECT 109.105 113.385 110.775 114.155 ;
        RECT 111.035 113.605 111.205 113.895 ;
        RECT 111.375 113.775 111.705 114.155 ;
        RECT 111.035 113.435 111.700 113.605 ;
        RECT 106.325 113.175 107.555 113.345 ;
        RECT 105.115 112.455 106.125 112.625 ;
        RECT 106.295 112.610 107.045 112.800 ;
        RECT 104.775 112.115 105.900 112.285 ;
        RECT 106.295 111.945 106.465 112.610 ;
        RECT 107.215 112.365 107.555 113.175 ;
        RECT 109.105 112.865 109.855 113.385 ;
        RECT 104.435 111.775 106.465 111.945 ;
        RECT 106.635 111.605 106.805 112.365 ;
        RECT 107.040 111.955 107.555 112.365 ;
        RECT 108.645 111.605 108.935 112.770 ;
        RECT 110.025 112.695 110.775 113.215 ;
        RECT 109.105 111.605 110.775 112.695 ;
        RECT 110.950 112.615 111.300 113.265 ;
        RECT 111.470 112.445 111.700 113.435 ;
        RECT 111.035 112.275 111.700 112.445 ;
        RECT 111.035 111.775 111.205 112.275 ;
        RECT 111.375 111.605 111.705 112.105 ;
        RECT 111.875 111.775 112.100 113.895 ;
        RECT 112.315 113.775 112.645 114.155 ;
        RECT 112.815 113.605 112.985 113.935 ;
        RECT 113.285 113.775 114.300 113.975 ;
        RECT 112.290 113.415 112.985 113.605 ;
        RECT 112.290 112.445 112.460 113.415 ;
        RECT 112.630 112.615 113.040 113.235 ;
        RECT 113.210 112.665 113.430 113.535 ;
        RECT 113.610 113.225 113.960 113.595 ;
        RECT 114.130 113.045 114.300 113.775 ;
        RECT 114.470 113.715 114.880 114.155 ;
        RECT 115.170 113.515 115.420 113.945 ;
        RECT 115.620 113.695 115.940 114.155 ;
        RECT 116.500 113.765 117.350 113.935 ;
        RECT 114.470 113.175 114.880 113.505 ;
        RECT 115.170 113.175 115.590 113.515 ;
        RECT 113.880 113.005 114.300 113.045 ;
        RECT 113.880 112.835 115.230 113.005 ;
        RECT 112.290 112.275 112.985 112.445 ;
        RECT 113.210 112.285 113.710 112.665 ;
        RECT 112.315 111.605 112.645 112.105 ;
        RECT 112.815 111.775 112.985 112.275 ;
        RECT 113.880 111.990 114.050 112.835 ;
        RECT 114.980 112.675 115.230 112.835 ;
        RECT 114.220 112.405 114.470 112.665 ;
        RECT 115.400 112.405 115.590 113.175 ;
        RECT 114.220 112.155 115.590 112.405 ;
        RECT 115.760 113.345 117.010 113.515 ;
        RECT 115.760 112.585 115.930 113.345 ;
        RECT 116.680 113.225 117.010 113.345 ;
        RECT 116.100 112.765 116.280 113.175 ;
        RECT 117.180 113.005 117.350 113.765 ;
        RECT 117.550 113.675 118.210 114.155 ;
        RECT 118.390 113.560 118.710 113.890 ;
        RECT 117.540 113.235 118.200 113.505 ;
        RECT 117.540 113.175 117.870 113.235 ;
        RECT 118.020 113.005 118.350 113.065 ;
        RECT 116.450 112.835 118.350 113.005 ;
        RECT 115.760 112.275 116.280 112.585 ;
        RECT 116.450 112.325 116.620 112.835 ;
        RECT 118.520 112.665 118.710 113.560 ;
        RECT 116.790 112.495 118.710 112.665 ;
        RECT 118.390 112.475 118.710 112.495 ;
        RECT 118.910 113.245 119.160 113.895 ;
        RECT 119.340 113.695 119.625 114.155 ;
        RECT 119.805 113.445 120.060 113.975 ;
        RECT 118.910 112.915 119.710 113.245 ;
        RECT 116.450 112.155 117.660 112.325 ;
        RECT 113.220 111.820 114.050 111.990 ;
        RECT 114.290 111.605 114.670 111.985 ;
        RECT 114.850 111.865 115.020 112.155 ;
        RECT 116.450 112.075 116.620 112.155 ;
        RECT 115.190 111.605 115.520 111.985 ;
        RECT 115.990 111.825 116.620 112.075 ;
        RECT 116.800 111.605 117.220 111.985 ;
        RECT 117.420 111.865 117.660 112.155 ;
        RECT 117.890 111.605 118.220 112.295 ;
        RECT 118.390 111.865 118.560 112.475 ;
        RECT 118.910 112.325 119.160 112.915 ;
        RECT 119.880 112.585 120.060 113.445 ;
        RECT 120.605 113.385 124.115 114.155 ;
        RECT 124.285 113.405 125.495 114.155 ;
        RECT 120.605 112.865 122.255 113.385 ;
        RECT 122.425 112.695 124.115 113.215 ;
        RECT 118.830 111.815 119.160 112.325 ;
        RECT 119.340 111.605 119.625 112.405 ;
        RECT 119.805 112.115 120.060 112.585 ;
        RECT 119.805 111.945 120.145 112.115 ;
        RECT 119.805 111.915 120.060 111.945 ;
        RECT 120.605 111.605 124.115 112.695 ;
        RECT 124.285 112.695 124.805 113.235 ;
        RECT 124.975 112.865 125.495 113.405 ;
        RECT 124.285 111.605 125.495 112.695 ;
        RECT 5.520 111.435 125.580 111.605 ;
        RECT 5.605 110.345 6.815 111.435 ;
        RECT 6.985 111.000 12.330 111.435 ;
        RECT 5.605 109.635 6.125 110.175 ;
        RECT 6.295 109.805 6.815 110.345 ;
        RECT 5.605 108.885 6.815 109.635 ;
        RECT 8.570 109.430 8.910 110.260 ;
        RECT 10.390 109.750 10.740 111.000 ;
        RECT 12.505 110.345 16.015 111.435 ;
        RECT 12.505 109.655 14.155 110.175 ;
        RECT 14.325 109.825 16.015 110.345 ;
        RECT 16.225 110.295 16.455 111.435 ;
        RECT 16.625 110.285 16.955 111.265 ;
        RECT 17.125 110.295 17.335 111.435 ;
        RECT 16.205 109.875 16.535 110.125 ;
        RECT 6.985 108.885 12.330 109.430 ;
        RECT 12.505 108.885 16.015 109.655 ;
        RECT 16.225 108.885 16.455 109.705 ;
        RECT 16.705 109.685 16.955 110.285 ;
        RECT 18.485 110.270 18.775 111.435 ;
        RECT 18.950 110.295 19.285 111.265 ;
        RECT 19.455 110.295 19.625 111.435 ;
        RECT 19.795 111.095 21.825 111.265 ;
        RECT 16.625 109.055 16.955 109.685 ;
        RECT 17.125 108.885 17.335 109.705 ;
        RECT 18.950 109.625 19.120 110.295 ;
        RECT 19.795 110.125 19.965 111.095 ;
        RECT 19.290 109.795 19.545 110.125 ;
        RECT 19.770 109.795 19.965 110.125 ;
        RECT 20.135 110.755 21.260 110.925 ;
        RECT 19.375 109.625 19.545 109.795 ;
        RECT 20.135 109.625 20.305 110.755 ;
        RECT 18.485 108.885 18.775 109.610 ;
        RECT 18.950 109.055 19.205 109.625 ;
        RECT 19.375 109.455 20.305 109.625 ;
        RECT 20.475 110.415 21.485 110.585 ;
        RECT 20.475 109.615 20.645 110.415 ;
        RECT 20.130 109.420 20.305 109.455 ;
        RECT 19.375 108.885 19.705 109.285 ;
        RECT 20.130 109.055 20.660 109.420 ;
        RECT 20.850 109.395 21.125 110.215 ;
        RECT 20.845 109.225 21.125 109.395 ;
        RECT 20.850 109.055 21.125 109.225 ;
        RECT 21.295 109.055 21.485 110.415 ;
        RECT 21.655 110.430 21.825 111.095 ;
        RECT 21.995 110.675 22.165 111.435 ;
        RECT 22.400 110.675 22.915 111.085 ;
        RECT 21.655 110.240 22.405 110.430 ;
        RECT 22.575 109.865 22.915 110.675 ;
        RECT 21.685 109.695 22.915 109.865 ;
        RECT 23.545 110.360 23.815 111.265 ;
        RECT 23.985 110.675 24.315 111.435 ;
        RECT 24.495 110.505 24.665 111.265 ;
        RECT 25.015 110.690 25.285 111.435 ;
        RECT 25.915 111.430 32.190 111.435 ;
        RECT 25.455 110.520 25.745 111.260 ;
        RECT 25.915 110.705 26.170 111.430 ;
        RECT 26.355 110.535 26.615 111.260 ;
        RECT 26.785 110.705 27.030 111.430 ;
        RECT 27.215 110.535 27.475 111.260 ;
        RECT 27.645 110.705 27.890 111.430 ;
        RECT 28.075 110.535 28.335 111.260 ;
        RECT 28.505 110.705 28.750 111.430 ;
        RECT 28.920 110.535 29.180 111.260 ;
        RECT 29.350 110.705 29.610 111.430 ;
        RECT 29.780 110.535 30.040 111.260 ;
        RECT 30.210 110.705 30.470 111.430 ;
        RECT 30.640 110.535 30.900 111.260 ;
        RECT 31.070 110.705 31.330 111.430 ;
        RECT 31.500 110.535 31.760 111.260 ;
        RECT 31.930 110.635 32.190 111.430 ;
        RECT 26.355 110.520 31.760 110.535 ;
        RECT 21.665 108.885 22.175 109.420 ;
        RECT 22.395 109.090 22.640 109.695 ;
        RECT 23.545 109.560 23.715 110.360 ;
        RECT 24.000 110.335 24.665 110.505 ;
        RECT 24.000 110.190 24.170 110.335 ;
        RECT 23.885 109.860 24.170 110.190 ;
        RECT 25.015 110.295 31.760 110.520 ;
        RECT 24.000 109.605 24.170 109.860 ;
        RECT 24.405 109.785 24.735 110.155 ;
        RECT 25.015 109.705 26.180 110.295 ;
        RECT 32.360 110.125 32.610 111.260 ;
        RECT 32.790 110.625 33.050 111.435 ;
        RECT 33.225 110.125 33.470 111.265 ;
        RECT 33.650 110.625 33.945 111.435 ;
        RECT 34.215 110.765 34.385 111.265 ;
        RECT 34.555 110.935 34.885 111.435 ;
        RECT 34.215 110.595 34.880 110.765 ;
        RECT 26.350 109.875 33.470 110.125 ;
        RECT 23.545 109.055 23.805 109.560 ;
        RECT 24.000 109.435 24.665 109.605 ;
        RECT 25.015 109.535 31.760 109.705 ;
        RECT 23.985 108.885 24.315 109.265 ;
        RECT 24.495 109.055 24.665 109.435 ;
        RECT 25.015 108.885 25.315 109.365 ;
        RECT 25.485 109.080 25.745 109.535 ;
        RECT 25.915 108.885 26.175 109.365 ;
        RECT 26.355 109.080 26.615 109.535 ;
        RECT 26.785 108.885 27.035 109.365 ;
        RECT 27.215 109.080 27.475 109.535 ;
        RECT 27.645 108.885 27.895 109.365 ;
        RECT 28.075 109.080 28.335 109.535 ;
        RECT 28.505 108.885 28.750 109.365 ;
        RECT 28.920 109.080 29.195 109.535 ;
        RECT 29.365 108.885 29.610 109.365 ;
        RECT 29.780 109.080 30.040 109.535 ;
        RECT 30.210 108.885 30.470 109.365 ;
        RECT 30.640 109.080 30.900 109.535 ;
        RECT 31.070 108.885 31.330 109.365 ;
        RECT 31.500 109.080 31.760 109.535 ;
        RECT 31.930 108.885 32.190 109.445 ;
        RECT 32.360 109.065 32.610 109.875 ;
        RECT 32.790 108.885 33.050 109.410 ;
        RECT 33.220 109.065 33.470 109.875 ;
        RECT 33.640 109.565 33.955 110.125 ;
        RECT 34.130 109.775 34.480 110.425 ;
        RECT 34.650 109.605 34.880 110.595 ;
        RECT 34.215 109.435 34.880 109.605 ;
        RECT 33.650 108.885 33.955 109.395 ;
        RECT 34.215 109.145 34.385 109.435 ;
        RECT 34.555 108.885 34.885 109.265 ;
        RECT 35.055 109.145 35.280 111.265 ;
        RECT 35.495 110.935 35.825 111.435 ;
        RECT 35.995 110.765 36.165 111.265 ;
        RECT 36.400 111.050 37.230 111.220 ;
        RECT 37.470 111.055 37.850 111.435 ;
        RECT 35.470 110.595 36.165 110.765 ;
        RECT 35.470 109.625 35.640 110.595 ;
        RECT 35.810 109.805 36.220 110.425 ;
        RECT 36.390 110.375 36.890 110.755 ;
        RECT 35.470 109.435 36.165 109.625 ;
        RECT 36.390 109.505 36.610 110.375 ;
        RECT 37.060 110.205 37.230 111.050 ;
        RECT 38.030 110.885 38.200 111.175 ;
        RECT 38.370 111.055 38.700 111.435 ;
        RECT 39.170 110.965 39.800 111.215 ;
        RECT 39.980 111.055 40.400 111.435 ;
        RECT 39.630 110.885 39.800 110.965 ;
        RECT 40.600 110.885 40.840 111.175 ;
        RECT 37.400 110.635 38.770 110.885 ;
        RECT 37.400 110.375 37.650 110.635 ;
        RECT 38.160 110.205 38.410 110.365 ;
        RECT 37.060 110.035 38.410 110.205 ;
        RECT 37.060 109.995 37.480 110.035 ;
        RECT 36.790 109.445 37.140 109.815 ;
        RECT 35.495 108.885 35.825 109.265 ;
        RECT 35.995 109.105 36.165 109.435 ;
        RECT 37.310 109.265 37.480 109.995 ;
        RECT 38.580 109.865 38.770 110.635 ;
        RECT 37.650 109.535 38.060 109.865 ;
        RECT 38.350 109.525 38.770 109.865 ;
        RECT 38.940 110.455 39.460 110.765 ;
        RECT 39.630 110.715 40.840 110.885 ;
        RECT 41.070 110.745 41.400 111.435 ;
        RECT 38.940 109.695 39.110 110.455 ;
        RECT 39.280 109.865 39.460 110.275 ;
        RECT 39.630 110.205 39.800 110.715 ;
        RECT 41.570 110.565 41.740 111.175 ;
        RECT 42.010 110.715 42.340 111.225 ;
        RECT 41.570 110.545 41.890 110.565 ;
        RECT 39.970 110.375 41.890 110.545 ;
        RECT 39.630 110.035 41.530 110.205 ;
        RECT 39.860 109.695 40.190 109.815 ;
        RECT 38.940 109.525 40.190 109.695 ;
        RECT 36.465 109.065 37.480 109.265 ;
        RECT 37.650 108.885 38.060 109.325 ;
        RECT 38.350 109.095 38.600 109.525 ;
        RECT 38.800 108.885 39.120 109.345 ;
        RECT 40.360 109.275 40.530 110.035 ;
        RECT 41.200 109.975 41.530 110.035 ;
        RECT 40.720 109.805 41.050 109.865 ;
        RECT 40.720 109.535 41.380 109.805 ;
        RECT 41.700 109.480 41.890 110.375 ;
        RECT 39.680 109.105 40.530 109.275 ;
        RECT 40.730 108.885 41.390 109.365 ;
        RECT 41.570 109.150 41.890 109.480 ;
        RECT 42.090 110.125 42.340 110.715 ;
        RECT 42.520 110.635 42.805 111.435 ;
        RECT 42.985 110.455 43.240 111.125 ;
        RECT 42.090 109.795 42.890 110.125 ;
        RECT 42.090 109.145 42.340 109.795 ;
        RECT 43.060 109.595 43.240 110.455 ;
        RECT 44.245 110.270 44.535 111.435 ;
        RECT 44.795 110.690 45.065 111.435 ;
        RECT 45.695 111.430 51.970 111.435 ;
        RECT 45.235 110.520 45.525 111.260 ;
        RECT 45.695 110.705 45.950 111.430 ;
        RECT 46.135 110.535 46.395 111.260 ;
        RECT 46.565 110.705 46.810 111.430 ;
        RECT 46.995 110.535 47.255 111.260 ;
        RECT 47.425 110.705 47.670 111.430 ;
        RECT 47.855 110.535 48.115 111.260 ;
        RECT 48.285 110.705 48.530 111.430 ;
        RECT 48.700 110.535 48.960 111.260 ;
        RECT 49.130 110.705 49.390 111.430 ;
        RECT 49.560 110.535 49.820 111.260 ;
        RECT 49.990 110.705 50.250 111.430 ;
        RECT 50.420 110.535 50.680 111.260 ;
        RECT 50.850 110.705 51.110 111.430 ;
        RECT 51.280 110.535 51.540 111.260 ;
        RECT 51.710 110.635 51.970 111.430 ;
        RECT 46.135 110.520 51.540 110.535 ;
        RECT 44.795 110.295 51.540 110.520 ;
        RECT 44.795 109.705 45.960 110.295 ;
        RECT 52.140 110.125 52.390 111.260 ;
        RECT 52.570 110.625 52.830 111.435 ;
        RECT 53.005 110.125 53.250 111.265 ;
        RECT 53.430 110.625 53.725 111.435 ;
        RECT 54.455 110.765 54.625 111.265 ;
        RECT 54.795 110.935 55.125 111.435 ;
        RECT 54.455 110.595 55.120 110.765 ;
        RECT 46.130 109.875 53.250 110.125 ;
        RECT 42.985 109.395 43.240 109.595 ;
        RECT 42.520 108.885 42.805 109.345 ;
        RECT 42.985 109.225 43.325 109.395 ;
        RECT 42.985 109.065 43.240 109.225 ;
        RECT 44.245 108.885 44.535 109.610 ;
        RECT 44.795 109.535 51.540 109.705 ;
        RECT 44.795 108.885 45.095 109.365 ;
        RECT 45.265 109.080 45.525 109.535 ;
        RECT 45.695 108.885 45.955 109.365 ;
        RECT 46.135 109.080 46.395 109.535 ;
        RECT 46.565 108.885 46.815 109.365 ;
        RECT 46.995 109.080 47.255 109.535 ;
        RECT 47.425 108.885 47.675 109.365 ;
        RECT 47.855 109.080 48.115 109.535 ;
        RECT 48.285 108.885 48.530 109.365 ;
        RECT 48.700 109.080 48.975 109.535 ;
        RECT 49.145 108.885 49.390 109.365 ;
        RECT 49.560 109.080 49.820 109.535 ;
        RECT 49.990 108.885 50.250 109.365 ;
        RECT 50.420 109.080 50.680 109.535 ;
        RECT 50.850 108.885 51.110 109.365 ;
        RECT 51.280 109.080 51.540 109.535 ;
        RECT 51.710 108.885 51.970 109.445 ;
        RECT 52.140 109.065 52.390 109.875 ;
        RECT 52.570 108.885 52.830 109.410 ;
        RECT 53.000 109.065 53.250 109.875 ;
        RECT 53.420 109.565 53.735 110.125 ;
        RECT 54.370 109.775 54.720 110.425 ;
        RECT 54.890 109.605 55.120 110.595 ;
        RECT 54.455 109.435 55.120 109.605 ;
        RECT 53.430 108.885 53.735 109.395 ;
        RECT 54.455 109.145 54.625 109.435 ;
        RECT 54.795 108.885 55.125 109.265 ;
        RECT 55.295 109.145 55.520 111.265 ;
        RECT 55.735 110.935 56.065 111.435 ;
        RECT 56.235 110.765 56.405 111.265 ;
        RECT 56.640 111.050 57.470 111.220 ;
        RECT 57.710 111.055 58.090 111.435 ;
        RECT 55.710 110.595 56.405 110.765 ;
        RECT 55.710 109.625 55.880 110.595 ;
        RECT 56.050 109.805 56.460 110.425 ;
        RECT 56.630 110.375 57.130 110.755 ;
        RECT 55.710 109.435 56.405 109.625 ;
        RECT 56.630 109.505 56.850 110.375 ;
        RECT 57.300 110.205 57.470 111.050 ;
        RECT 58.270 110.885 58.440 111.175 ;
        RECT 58.610 111.055 58.940 111.435 ;
        RECT 59.410 110.965 60.040 111.215 ;
        RECT 60.220 111.055 60.640 111.435 ;
        RECT 59.870 110.885 60.040 110.965 ;
        RECT 60.840 110.885 61.080 111.175 ;
        RECT 57.640 110.635 59.010 110.885 ;
        RECT 57.640 110.375 57.890 110.635 ;
        RECT 58.400 110.205 58.650 110.365 ;
        RECT 57.300 110.035 58.650 110.205 ;
        RECT 57.300 109.995 57.720 110.035 ;
        RECT 57.030 109.445 57.380 109.815 ;
        RECT 55.735 108.885 56.065 109.265 ;
        RECT 56.235 109.105 56.405 109.435 ;
        RECT 57.550 109.265 57.720 109.995 ;
        RECT 58.820 109.865 59.010 110.635 ;
        RECT 57.890 109.535 58.300 109.865 ;
        RECT 58.590 109.525 59.010 109.865 ;
        RECT 59.180 110.455 59.700 110.765 ;
        RECT 59.870 110.715 61.080 110.885 ;
        RECT 61.310 110.745 61.640 111.435 ;
        RECT 59.180 109.695 59.350 110.455 ;
        RECT 59.520 109.865 59.700 110.275 ;
        RECT 59.870 110.205 60.040 110.715 ;
        RECT 61.810 110.565 61.980 111.175 ;
        RECT 62.250 110.715 62.580 111.225 ;
        RECT 61.810 110.545 62.130 110.565 ;
        RECT 60.210 110.375 62.130 110.545 ;
        RECT 59.870 110.035 61.770 110.205 ;
        RECT 60.100 109.695 60.430 109.815 ;
        RECT 59.180 109.525 60.430 109.695 ;
        RECT 56.705 109.065 57.720 109.265 ;
        RECT 57.890 108.885 58.300 109.325 ;
        RECT 58.590 109.095 58.840 109.525 ;
        RECT 59.040 108.885 59.360 109.345 ;
        RECT 60.600 109.275 60.770 110.035 ;
        RECT 61.440 109.975 61.770 110.035 ;
        RECT 60.960 109.805 61.290 109.865 ;
        RECT 60.960 109.535 61.620 109.805 ;
        RECT 61.940 109.480 62.130 110.375 ;
        RECT 59.920 109.105 60.770 109.275 ;
        RECT 60.970 108.885 61.630 109.365 ;
        RECT 61.810 109.150 62.130 109.480 ;
        RECT 62.330 110.125 62.580 110.715 ;
        RECT 62.760 110.635 63.045 111.435 ;
        RECT 63.225 110.455 63.480 111.125 ;
        RECT 62.330 109.795 63.130 110.125 ;
        RECT 62.330 109.145 62.580 109.795 ;
        RECT 63.300 109.595 63.480 110.455 ;
        RECT 64.085 110.295 64.295 111.435 ;
        RECT 64.465 110.285 64.795 111.265 ;
        RECT 64.965 110.295 65.195 111.435 ;
        RECT 65.405 110.345 67.995 111.435 ;
        RECT 63.225 109.395 63.480 109.595 ;
        RECT 62.760 108.885 63.045 109.345 ;
        RECT 63.225 109.225 63.565 109.395 ;
        RECT 63.225 109.065 63.480 109.225 ;
        RECT 64.085 108.885 64.295 109.705 ;
        RECT 64.465 109.685 64.715 110.285 ;
        RECT 64.885 109.875 65.215 110.125 ;
        RECT 64.465 109.055 64.795 109.685 ;
        RECT 64.965 108.885 65.195 109.705 ;
        RECT 65.405 109.655 66.615 110.175 ;
        RECT 66.785 109.825 67.995 110.345 ;
        RECT 68.715 110.505 68.885 111.265 ;
        RECT 69.065 110.675 69.395 111.435 ;
        RECT 68.715 110.335 69.380 110.505 ;
        RECT 69.565 110.360 69.835 111.265 ;
        RECT 69.210 110.190 69.380 110.335 ;
        RECT 68.645 109.785 68.975 110.155 ;
        RECT 69.210 109.860 69.495 110.190 ;
        RECT 65.405 108.885 67.995 109.655 ;
        RECT 69.210 109.605 69.380 109.860 ;
        RECT 68.715 109.435 69.380 109.605 ;
        RECT 69.665 109.560 69.835 110.360 ;
        RECT 70.005 110.270 70.295 111.435 ;
        RECT 70.555 110.765 70.725 111.265 ;
        RECT 70.895 110.935 71.225 111.435 ;
        RECT 70.555 110.595 71.220 110.765 ;
        RECT 70.470 109.775 70.820 110.425 ;
        RECT 68.715 109.055 68.885 109.435 ;
        RECT 69.065 108.885 69.395 109.265 ;
        RECT 69.575 109.055 69.835 109.560 ;
        RECT 70.005 108.885 70.295 109.610 ;
        RECT 70.990 109.605 71.220 110.595 ;
        RECT 70.555 109.435 71.220 109.605 ;
        RECT 70.555 109.145 70.725 109.435 ;
        RECT 70.895 108.885 71.225 109.265 ;
        RECT 71.395 109.145 71.620 111.265 ;
        RECT 71.835 110.935 72.165 111.435 ;
        RECT 72.335 110.765 72.505 111.265 ;
        RECT 72.740 111.050 73.570 111.220 ;
        RECT 73.810 111.055 74.190 111.435 ;
        RECT 71.810 110.595 72.505 110.765 ;
        RECT 71.810 109.625 71.980 110.595 ;
        RECT 72.150 109.805 72.560 110.425 ;
        RECT 72.730 110.375 73.230 110.755 ;
        RECT 71.810 109.435 72.505 109.625 ;
        RECT 72.730 109.505 72.950 110.375 ;
        RECT 73.400 110.205 73.570 111.050 ;
        RECT 74.370 110.885 74.540 111.175 ;
        RECT 74.710 111.055 75.040 111.435 ;
        RECT 75.510 110.965 76.140 111.215 ;
        RECT 76.320 111.055 76.740 111.435 ;
        RECT 75.970 110.885 76.140 110.965 ;
        RECT 76.940 110.885 77.180 111.175 ;
        RECT 73.740 110.635 75.110 110.885 ;
        RECT 73.740 110.375 73.990 110.635 ;
        RECT 74.500 110.205 74.750 110.365 ;
        RECT 73.400 110.035 74.750 110.205 ;
        RECT 73.400 109.995 73.820 110.035 ;
        RECT 73.130 109.445 73.480 109.815 ;
        RECT 71.835 108.885 72.165 109.265 ;
        RECT 72.335 109.105 72.505 109.435 ;
        RECT 73.650 109.265 73.820 109.995 ;
        RECT 74.920 109.865 75.110 110.635 ;
        RECT 73.990 109.535 74.400 109.865 ;
        RECT 74.690 109.525 75.110 109.865 ;
        RECT 75.280 110.455 75.800 110.765 ;
        RECT 75.970 110.715 77.180 110.885 ;
        RECT 77.410 110.745 77.740 111.435 ;
        RECT 75.280 109.695 75.450 110.455 ;
        RECT 75.620 109.865 75.800 110.275 ;
        RECT 75.970 110.205 76.140 110.715 ;
        RECT 77.910 110.565 78.080 111.175 ;
        RECT 78.350 110.715 78.680 111.225 ;
        RECT 77.910 110.545 78.230 110.565 ;
        RECT 76.310 110.375 78.230 110.545 ;
        RECT 75.970 110.035 77.870 110.205 ;
        RECT 76.200 109.695 76.530 109.815 ;
        RECT 75.280 109.525 76.530 109.695 ;
        RECT 72.805 109.065 73.820 109.265 ;
        RECT 73.990 108.885 74.400 109.325 ;
        RECT 74.690 109.095 74.940 109.525 ;
        RECT 75.140 108.885 75.460 109.345 ;
        RECT 76.700 109.275 76.870 110.035 ;
        RECT 77.540 109.975 77.870 110.035 ;
        RECT 77.060 109.805 77.390 109.865 ;
        RECT 77.060 109.535 77.720 109.805 ;
        RECT 78.040 109.480 78.230 110.375 ;
        RECT 76.020 109.105 76.870 109.275 ;
        RECT 77.070 108.885 77.730 109.365 ;
        RECT 77.910 109.150 78.230 109.480 ;
        RECT 78.430 110.125 78.680 110.715 ;
        RECT 78.860 110.635 79.145 111.435 ;
        RECT 79.325 110.455 79.580 111.125 ;
        RECT 80.215 110.765 80.385 111.265 ;
        RECT 80.555 110.935 80.885 111.435 ;
        RECT 80.215 110.595 80.880 110.765 ;
        RECT 78.430 109.795 79.230 110.125 ;
        RECT 78.430 109.145 78.680 109.795 ;
        RECT 79.400 109.595 79.580 110.455 ;
        RECT 80.130 109.775 80.480 110.425 ;
        RECT 80.650 109.605 80.880 110.595 ;
        RECT 79.325 109.395 79.580 109.595 ;
        RECT 80.215 109.435 80.880 109.605 ;
        RECT 78.860 108.885 79.145 109.345 ;
        RECT 79.325 109.225 79.665 109.395 ;
        RECT 79.325 109.065 79.580 109.225 ;
        RECT 80.215 109.145 80.385 109.435 ;
        RECT 80.555 108.885 80.885 109.265 ;
        RECT 81.055 109.145 81.280 111.265 ;
        RECT 81.495 110.935 81.825 111.435 ;
        RECT 81.995 110.765 82.165 111.265 ;
        RECT 82.400 111.050 83.230 111.220 ;
        RECT 83.470 111.055 83.850 111.435 ;
        RECT 81.470 110.595 82.165 110.765 ;
        RECT 81.470 109.625 81.640 110.595 ;
        RECT 81.810 109.805 82.220 110.425 ;
        RECT 82.390 110.375 82.890 110.755 ;
        RECT 81.470 109.435 82.165 109.625 ;
        RECT 82.390 109.505 82.610 110.375 ;
        RECT 83.060 110.205 83.230 111.050 ;
        RECT 84.030 110.885 84.200 111.175 ;
        RECT 84.370 111.055 84.700 111.435 ;
        RECT 85.170 110.965 85.800 111.215 ;
        RECT 85.980 111.055 86.400 111.435 ;
        RECT 85.630 110.885 85.800 110.965 ;
        RECT 86.600 110.885 86.840 111.175 ;
        RECT 83.400 110.635 84.770 110.885 ;
        RECT 83.400 110.375 83.650 110.635 ;
        RECT 84.160 110.205 84.410 110.365 ;
        RECT 83.060 110.035 84.410 110.205 ;
        RECT 83.060 109.995 83.480 110.035 ;
        RECT 82.790 109.445 83.140 109.815 ;
        RECT 81.495 108.885 81.825 109.265 ;
        RECT 81.995 109.105 82.165 109.435 ;
        RECT 83.310 109.265 83.480 109.995 ;
        RECT 84.580 109.865 84.770 110.635 ;
        RECT 83.650 109.535 84.060 109.865 ;
        RECT 84.350 109.525 84.770 109.865 ;
        RECT 84.940 110.455 85.460 110.765 ;
        RECT 85.630 110.715 86.840 110.885 ;
        RECT 87.070 110.745 87.400 111.435 ;
        RECT 84.940 109.695 85.110 110.455 ;
        RECT 85.280 109.865 85.460 110.275 ;
        RECT 85.630 110.205 85.800 110.715 ;
        RECT 87.570 110.565 87.740 111.175 ;
        RECT 88.010 110.715 88.340 111.225 ;
        RECT 87.570 110.545 87.890 110.565 ;
        RECT 85.970 110.375 87.890 110.545 ;
        RECT 85.630 110.035 87.530 110.205 ;
        RECT 85.860 109.695 86.190 109.815 ;
        RECT 84.940 109.525 86.190 109.695 ;
        RECT 82.465 109.065 83.480 109.265 ;
        RECT 83.650 108.885 84.060 109.325 ;
        RECT 84.350 109.095 84.600 109.525 ;
        RECT 84.800 108.885 85.120 109.345 ;
        RECT 86.360 109.275 86.530 110.035 ;
        RECT 87.200 109.975 87.530 110.035 ;
        RECT 86.720 109.805 87.050 109.865 ;
        RECT 86.720 109.535 87.380 109.805 ;
        RECT 87.700 109.480 87.890 110.375 ;
        RECT 85.680 109.105 86.530 109.275 ;
        RECT 86.730 108.885 87.390 109.365 ;
        RECT 87.570 109.150 87.890 109.480 ;
        RECT 88.090 110.125 88.340 110.715 ;
        RECT 88.520 110.635 88.805 111.435 ;
        RECT 88.985 110.755 89.240 111.125 ;
        RECT 88.985 110.585 89.325 110.755 ;
        RECT 88.985 110.455 89.240 110.585 ;
        RECT 88.090 109.795 88.890 110.125 ;
        RECT 88.090 109.145 88.340 109.795 ;
        RECT 89.060 109.595 89.240 110.455 ;
        RECT 89.795 110.295 90.125 111.435 ;
        RECT 88.520 108.885 88.805 109.345 ;
        RECT 88.985 109.065 89.240 109.595 ;
        RECT 89.785 109.545 90.125 110.125 ;
        RECT 90.295 110.095 90.655 111.265 ;
        RECT 90.855 110.265 91.185 111.435 ;
        RECT 91.385 110.095 91.715 111.265 ;
        RECT 91.915 110.265 92.245 111.435 ;
        RECT 92.545 110.345 95.135 111.435 ;
        RECT 90.295 109.815 91.715 110.095 ;
        RECT 90.295 109.480 90.655 109.815 ;
        RECT 92.545 109.655 93.755 110.175 ;
        RECT 93.925 109.825 95.135 110.345 ;
        RECT 95.765 110.270 96.055 111.435 ;
        RECT 96.230 110.295 96.565 111.265 ;
        RECT 96.735 110.295 96.905 111.435 ;
        RECT 97.075 111.095 99.105 111.265 ;
        RECT 89.795 108.885 90.125 109.375 ;
        RECT 90.295 109.055 90.915 109.480 ;
        RECT 91.375 108.885 91.705 109.575 ;
        RECT 92.545 108.885 95.135 109.655 ;
        RECT 96.230 109.625 96.400 110.295 ;
        RECT 97.075 110.125 97.245 111.095 ;
        RECT 96.570 109.795 96.825 110.125 ;
        RECT 97.050 109.795 97.245 110.125 ;
        RECT 97.415 110.755 98.540 110.925 ;
        RECT 96.655 109.625 96.825 109.795 ;
        RECT 97.415 109.625 97.585 110.755 ;
        RECT 95.765 108.885 96.055 109.610 ;
        RECT 96.230 109.055 96.485 109.625 ;
        RECT 96.655 109.455 97.585 109.625 ;
        RECT 97.755 110.415 98.765 110.585 ;
        RECT 97.755 109.615 97.925 110.415 ;
        RECT 97.410 109.420 97.585 109.455 ;
        RECT 96.655 108.885 96.985 109.285 ;
        RECT 97.410 109.055 97.940 109.420 ;
        RECT 98.130 109.395 98.405 110.215 ;
        RECT 98.125 109.225 98.405 109.395 ;
        RECT 98.130 109.055 98.405 109.225 ;
        RECT 98.575 109.055 98.765 110.415 ;
        RECT 98.935 110.430 99.105 111.095 ;
        RECT 99.275 110.675 99.445 111.435 ;
        RECT 99.680 110.675 100.195 111.085 ;
        RECT 98.935 110.240 99.685 110.430 ;
        RECT 99.855 109.865 100.195 110.675 ;
        RECT 100.365 110.345 103.875 111.435 ;
        RECT 104.135 110.765 104.305 111.265 ;
        RECT 104.475 110.935 104.805 111.435 ;
        RECT 104.135 110.595 104.800 110.765 ;
        RECT 98.965 109.695 100.195 109.865 ;
        RECT 98.945 108.885 99.455 109.420 ;
        RECT 99.675 109.090 99.920 109.695 ;
        RECT 100.365 109.655 102.015 110.175 ;
        RECT 102.185 109.825 103.875 110.345 ;
        RECT 104.050 109.775 104.400 110.425 ;
        RECT 100.365 108.885 103.875 109.655 ;
        RECT 104.570 109.605 104.800 110.595 ;
        RECT 104.135 109.435 104.800 109.605 ;
        RECT 104.135 109.145 104.305 109.435 ;
        RECT 104.475 108.885 104.805 109.265 ;
        RECT 104.975 109.145 105.200 111.265 ;
        RECT 105.415 110.935 105.745 111.435 ;
        RECT 105.915 110.765 106.085 111.265 ;
        RECT 106.320 111.050 107.150 111.220 ;
        RECT 107.390 111.055 107.770 111.435 ;
        RECT 105.390 110.595 106.085 110.765 ;
        RECT 105.390 109.625 105.560 110.595 ;
        RECT 105.730 109.805 106.140 110.425 ;
        RECT 106.310 110.375 106.810 110.755 ;
        RECT 105.390 109.435 106.085 109.625 ;
        RECT 106.310 109.505 106.530 110.375 ;
        RECT 106.980 110.205 107.150 111.050 ;
        RECT 107.950 110.885 108.120 111.175 ;
        RECT 108.290 111.055 108.620 111.435 ;
        RECT 109.090 110.965 109.720 111.215 ;
        RECT 109.900 111.055 110.320 111.435 ;
        RECT 109.550 110.885 109.720 110.965 ;
        RECT 110.520 110.885 110.760 111.175 ;
        RECT 107.320 110.635 108.690 110.885 ;
        RECT 107.320 110.375 107.570 110.635 ;
        RECT 108.080 110.205 108.330 110.365 ;
        RECT 106.980 110.035 108.330 110.205 ;
        RECT 106.980 109.995 107.400 110.035 ;
        RECT 106.710 109.445 107.060 109.815 ;
        RECT 105.415 108.885 105.745 109.265 ;
        RECT 105.915 109.105 106.085 109.435 ;
        RECT 107.230 109.265 107.400 109.995 ;
        RECT 108.500 109.865 108.690 110.635 ;
        RECT 107.570 109.535 107.980 109.865 ;
        RECT 108.270 109.525 108.690 109.865 ;
        RECT 108.860 110.455 109.380 110.765 ;
        RECT 109.550 110.715 110.760 110.885 ;
        RECT 110.990 110.745 111.320 111.435 ;
        RECT 108.860 109.695 109.030 110.455 ;
        RECT 109.200 109.865 109.380 110.275 ;
        RECT 109.550 110.205 109.720 110.715 ;
        RECT 111.490 110.565 111.660 111.175 ;
        RECT 111.930 110.715 112.260 111.225 ;
        RECT 111.490 110.545 111.810 110.565 ;
        RECT 109.890 110.375 111.810 110.545 ;
        RECT 109.550 110.035 111.450 110.205 ;
        RECT 109.780 109.695 110.110 109.815 ;
        RECT 108.860 109.525 110.110 109.695 ;
        RECT 106.385 109.065 107.400 109.265 ;
        RECT 107.570 108.885 107.980 109.325 ;
        RECT 108.270 109.095 108.520 109.525 ;
        RECT 108.720 108.885 109.040 109.345 ;
        RECT 110.280 109.275 110.450 110.035 ;
        RECT 111.120 109.975 111.450 110.035 ;
        RECT 110.640 109.805 110.970 109.865 ;
        RECT 110.640 109.535 111.300 109.805 ;
        RECT 111.620 109.480 111.810 110.375 ;
        RECT 109.600 109.105 110.450 109.275 ;
        RECT 110.650 108.885 111.310 109.365 ;
        RECT 111.490 109.150 111.810 109.480 ;
        RECT 112.010 110.125 112.260 110.715 ;
        RECT 112.440 110.635 112.725 111.435 ;
        RECT 112.905 110.455 113.160 111.125 ;
        RECT 112.010 109.795 112.810 110.125 ;
        RECT 112.980 110.075 113.160 110.455 ;
        RECT 113.710 110.295 114.045 111.265 ;
        RECT 114.215 110.295 114.385 111.435 ;
        RECT 114.555 111.095 116.585 111.265 ;
        RECT 112.980 109.905 113.245 110.075 ;
        RECT 112.010 109.145 112.260 109.795 ;
        RECT 112.980 109.595 113.160 109.905 ;
        RECT 112.440 108.885 112.725 109.345 ;
        RECT 112.905 109.065 113.160 109.595 ;
        RECT 113.710 109.625 113.880 110.295 ;
        RECT 114.555 110.125 114.725 111.095 ;
        RECT 114.050 109.795 114.305 110.125 ;
        RECT 114.530 109.795 114.725 110.125 ;
        RECT 114.895 110.755 116.020 110.925 ;
        RECT 114.135 109.625 114.305 109.795 ;
        RECT 114.895 109.625 115.065 110.755 ;
        RECT 113.710 109.055 113.965 109.625 ;
        RECT 114.135 109.455 115.065 109.625 ;
        RECT 115.235 110.415 116.245 110.585 ;
        RECT 115.235 109.615 115.405 110.415 ;
        RECT 114.890 109.420 115.065 109.455 ;
        RECT 114.135 108.885 114.465 109.285 ;
        RECT 114.890 109.055 115.420 109.420 ;
        RECT 115.610 109.395 115.885 110.215 ;
        RECT 115.605 109.225 115.885 109.395 ;
        RECT 115.610 109.055 115.885 109.225 ;
        RECT 116.055 109.055 116.245 110.415 ;
        RECT 116.415 110.430 116.585 111.095 ;
        RECT 116.755 110.675 116.925 111.435 ;
        RECT 117.160 110.675 117.675 111.085 ;
        RECT 116.415 110.240 117.165 110.430 ;
        RECT 117.335 109.865 117.675 110.675 ;
        RECT 117.905 110.295 118.115 111.435 ;
        RECT 116.445 109.695 117.675 109.865 ;
        RECT 118.285 110.285 118.615 111.265 ;
        RECT 118.785 110.295 119.015 111.435 ;
        RECT 119.225 110.360 119.495 111.265 ;
        RECT 119.665 110.675 119.995 111.435 ;
        RECT 120.175 110.505 120.345 111.265 ;
        RECT 116.425 108.885 116.935 109.420 ;
        RECT 117.155 109.090 117.400 109.695 ;
        RECT 117.905 108.885 118.115 109.705 ;
        RECT 118.285 109.685 118.535 110.285 ;
        RECT 118.705 109.875 119.035 110.125 ;
        RECT 118.285 109.055 118.615 109.685 ;
        RECT 118.785 108.885 119.015 109.705 ;
        RECT 119.225 109.560 119.395 110.360 ;
        RECT 119.680 110.335 120.345 110.505 ;
        RECT 119.680 110.190 119.850 110.335 ;
        RECT 121.525 110.270 121.815 111.435 ;
        RECT 122.025 110.295 122.255 111.435 ;
        RECT 122.425 110.285 122.755 111.265 ;
        RECT 122.925 110.295 123.135 111.435 ;
        RECT 124.285 110.345 125.495 111.435 ;
        RECT 119.565 109.860 119.850 110.190 ;
        RECT 119.680 109.605 119.850 109.860 ;
        RECT 120.085 109.785 120.415 110.155 ;
        RECT 122.005 109.875 122.335 110.125 ;
        RECT 119.225 109.055 119.485 109.560 ;
        RECT 119.680 109.435 120.345 109.605 ;
        RECT 119.665 108.885 119.995 109.265 ;
        RECT 120.175 109.055 120.345 109.435 ;
        RECT 121.525 108.885 121.815 109.610 ;
        RECT 122.025 108.885 122.255 109.705 ;
        RECT 122.505 109.685 122.755 110.285 ;
        RECT 124.285 109.805 124.805 110.345 ;
        RECT 122.425 109.055 122.755 109.685 ;
        RECT 122.925 108.885 123.135 109.705 ;
        RECT 124.975 109.635 125.495 110.175 ;
        RECT 124.285 108.885 125.495 109.635 ;
        RECT 5.520 108.715 125.580 108.885 ;
        RECT 5.605 107.965 6.815 108.715 ;
        RECT 5.605 107.425 6.125 107.965 ;
        RECT 6.985 107.945 10.495 108.715 ;
        RECT 10.665 107.965 11.875 108.715 ;
        RECT 12.045 108.040 12.305 108.545 ;
        RECT 12.485 108.335 12.815 108.715 ;
        RECT 12.995 108.165 13.165 108.545 ;
        RECT 6.295 107.255 6.815 107.795 ;
        RECT 6.985 107.425 8.635 107.945 ;
        RECT 8.805 107.255 10.495 107.775 ;
        RECT 10.665 107.425 11.185 107.965 ;
        RECT 11.355 107.255 11.875 107.795 ;
        RECT 5.605 106.165 6.815 107.255 ;
        RECT 6.985 106.165 10.495 107.255 ;
        RECT 10.665 106.165 11.875 107.255 ;
        RECT 12.045 107.240 12.215 108.040 ;
        RECT 12.500 107.995 13.165 108.165 ;
        RECT 13.425 108.040 13.685 108.545 ;
        RECT 13.865 108.335 14.195 108.715 ;
        RECT 14.375 108.165 14.545 108.545 ;
        RECT 12.500 107.740 12.670 107.995 ;
        RECT 12.385 107.410 12.670 107.740 ;
        RECT 12.905 107.445 13.235 107.815 ;
        RECT 12.500 107.265 12.670 107.410 ;
        RECT 12.045 106.335 12.315 107.240 ;
        RECT 12.500 107.095 13.165 107.265 ;
        RECT 12.485 106.165 12.815 106.925 ;
        RECT 12.995 106.335 13.165 107.095 ;
        RECT 13.425 107.240 13.595 108.040 ;
        RECT 13.880 107.995 14.545 108.165 ;
        RECT 13.880 107.740 14.050 107.995 ;
        RECT 15.325 107.895 15.535 108.715 ;
        RECT 15.705 107.915 16.035 108.545 ;
        RECT 13.765 107.410 14.050 107.740 ;
        RECT 14.285 107.445 14.615 107.815 ;
        RECT 13.880 107.265 14.050 107.410 ;
        RECT 15.705 107.315 15.955 107.915 ;
        RECT 16.205 107.895 16.435 108.715 ;
        RECT 16.650 107.975 16.905 108.545 ;
        RECT 17.075 108.315 17.405 108.715 ;
        RECT 17.830 108.180 18.360 108.545 ;
        RECT 17.830 108.145 18.005 108.180 ;
        RECT 17.075 107.975 18.005 108.145 ;
        RECT 16.125 107.475 16.455 107.725 ;
        RECT 13.425 106.335 13.695 107.240 ;
        RECT 13.880 107.095 14.545 107.265 ;
        RECT 13.865 106.165 14.195 106.925 ;
        RECT 14.375 106.335 14.545 107.095 ;
        RECT 15.325 106.165 15.535 107.305 ;
        RECT 15.705 106.335 16.035 107.315 ;
        RECT 16.650 107.305 16.820 107.975 ;
        RECT 17.075 107.805 17.245 107.975 ;
        RECT 16.990 107.475 17.245 107.805 ;
        RECT 17.470 107.475 17.665 107.805 ;
        RECT 16.205 106.165 16.435 107.305 ;
        RECT 16.650 106.335 16.985 107.305 ;
        RECT 17.155 106.165 17.325 107.305 ;
        RECT 17.495 106.505 17.665 107.475 ;
        RECT 17.835 106.845 18.005 107.975 ;
        RECT 18.175 107.185 18.345 107.985 ;
        RECT 18.550 107.695 18.825 108.545 ;
        RECT 18.545 107.525 18.825 107.695 ;
        RECT 18.550 107.385 18.825 107.525 ;
        RECT 18.995 107.185 19.185 108.545 ;
        RECT 19.365 108.180 19.875 108.715 ;
        RECT 20.095 107.905 20.340 108.510 ;
        RECT 20.785 107.945 23.375 108.715 ;
        RECT 23.635 108.165 23.805 108.545 ;
        RECT 23.985 108.335 24.315 108.715 ;
        RECT 23.635 107.995 24.300 108.165 ;
        RECT 24.495 108.040 24.755 108.545 ;
        RECT 19.385 107.735 20.615 107.905 ;
        RECT 18.175 107.015 19.185 107.185 ;
        RECT 19.355 107.170 20.105 107.360 ;
        RECT 17.835 106.675 18.960 106.845 ;
        RECT 19.355 106.505 19.525 107.170 ;
        RECT 20.275 106.925 20.615 107.735 ;
        RECT 20.785 107.425 21.995 107.945 ;
        RECT 22.165 107.255 23.375 107.775 ;
        RECT 23.565 107.445 23.895 107.815 ;
        RECT 24.130 107.740 24.300 107.995 ;
        RECT 24.130 107.410 24.415 107.740 ;
        RECT 24.130 107.265 24.300 107.410 ;
        RECT 17.495 106.335 19.525 106.505 ;
        RECT 19.695 106.165 19.865 106.925 ;
        RECT 20.100 106.515 20.615 106.925 ;
        RECT 20.785 106.165 23.375 107.255 ;
        RECT 23.635 107.095 24.300 107.265 ;
        RECT 24.585 107.240 24.755 108.040 ;
        RECT 23.635 106.335 23.805 107.095 ;
        RECT 23.985 106.165 24.315 106.925 ;
        RECT 24.485 106.335 24.755 107.240 ;
        RECT 24.925 108.215 25.225 108.545 ;
        RECT 25.395 108.235 25.670 108.715 ;
        RECT 24.925 107.305 25.095 108.215 ;
        RECT 25.850 108.065 26.145 108.455 ;
        RECT 26.315 108.235 26.570 108.715 ;
        RECT 26.745 108.065 27.005 108.455 ;
        RECT 27.175 108.235 27.455 108.715 ;
        RECT 25.265 107.475 25.615 108.045 ;
        RECT 25.850 107.895 27.500 108.065 ;
        RECT 28.205 107.895 28.415 108.715 ;
        RECT 28.585 107.915 28.915 108.545 ;
        RECT 25.785 107.555 26.925 107.725 ;
        RECT 25.785 107.305 25.955 107.555 ;
        RECT 27.095 107.385 27.500 107.895 ;
        RECT 24.925 107.135 25.955 107.305 ;
        RECT 26.745 107.215 27.500 107.385 ;
        RECT 28.585 107.315 28.835 107.915 ;
        RECT 29.085 107.895 29.315 108.715 ;
        RECT 29.565 107.895 29.795 108.715 ;
        RECT 29.965 107.915 30.295 108.545 ;
        RECT 29.005 107.475 29.335 107.725 ;
        RECT 29.545 107.475 29.875 107.725 ;
        RECT 30.045 107.315 30.295 107.915 ;
        RECT 30.465 107.895 30.675 108.715 ;
        RECT 31.365 107.990 31.655 108.715 ;
        RECT 31.825 107.945 33.495 108.715 ;
        RECT 31.825 107.425 32.575 107.945 ;
        RECT 33.940 107.905 34.185 108.510 ;
        RECT 34.405 108.180 34.915 108.715 ;
        RECT 24.925 106.335 25.235 107.135 ;
        RECT 26.745 106.965 27.005 107.215 ;
        RECT 25.405 106.165 25.715 106.965 ;
        RECT 25.885 106.795 27.005 106.965 ;
        RECT 25.885 106.335 26.145 106.795 ;
        RECT 26.315 106.165 26.570 106.625 ;
        RECT 26.745 106.335 27.005 106.795 ;
        RECT 27.175 106.165 27.460 107.035 ;
        RECT 28.205 106.165 28.415 107.305 ;
        RECT 28.585 106.335 28.915 107.315 ;
        RECT 29.085 106.165 29.315 107.305 ;
        RECT 29.565 106.165 29.795 107.305 ;
        RECT 29.965 106.335 30.295 107.315 ;
        RECT 30.465 106.165 30.675 107.305 ;
        RECT 31.365 106.165 31.655 107.330 ;
        RECT 32.745 107.255 33.495 107.775 ;
        RECT 31.825 106.165 33.495 107.255 ;
        RECT 33.665 107.735 34.895 107.905 ;
        RECT 33.665 106.925 34.005 107.735 ;
        RECT 34.175 107.170 34.925 107.360 ;
        RECT 33.665 106.515 34.180 106.925 ;
        RECT 34.415 106.165 34.585 106.925 ;
        RECT 34.755 106.505 34.925 107.170 ;
        RECT 35.095 107.185 35.285 108.545 ;
        RECT 35.455 107.695 35.730 108.545 ;
        RECT 35.920 108.180 36.450 108.545 ;
        RECT 36.875 108.315 37.205 108.715 ;
        RECT 36.275 108.145 36.450 108.180 ;
        RECT 35.455 107.525 35.735 107.695 ;
        RECT 35.455 107.385 35.730 107.525 ;
        RECT 35.935 107.185 36.105 107.985 ;
        RECT 35.095 107.015 36.105 107.185 ;
        RECT 36.275 107.975 37.205 108.145 ;
        RECT 37.375 107.975 37.630 108.545 ;
        RECT 38.355 108.165 38.525 108.455 ;
        RECT 38.695 108.335 39.025 108.715 ;
        RECT 38.355 107.995 39.020 108.165 ;
        RECT 36.275 106.845 36.445 107.975 ;
        RECT 37.035 107.805 37.205 107.975 ;
        RECT 35.320 106.675 36.445 106.845 ;
        RECT 36.615 107.475 36.810 107.805 ;
        RECT 37.035 107.475 37.290 107.805 ;
        RECT 36.615 106.505 36.785 107.475 ;
        RECT 37.460 107.305 37.630 107.975 ;
        RECT 34.755 106.335 36.785 106.505 ;
        RECT 36.955 106.165 37.125 107.305 ;
        RECT 37.295 106.335 37.630 107.305 ;
        RECT 38.270 107.175 38.620 107.825 ;
        RECT 38.790 107.005 39.020 107.995 ;
        RECT 38.355 106.835 39.020 107.005 ;
        RECT 38.355 106.335 38.525 106.835 ;
        RECT 38.695 106.165 39.025 106.665 ;
        RECT 39.195 106.335 39.420 108.455 ;
        RECT 39.635 108.335 39.965 108.715 ;
        RECT 40.135 108.165 40.305 108.495 ;
        RECT 40.605 108.335 41.620 108.535 ;
        RECT 39.610 107.975 40.305 108.165 ;
        RECT 39.610 107.005 39.780 107.975 ;
        RECT 39.950 107.175 40.360 107.795 ;
        RECT 40.530 107.225 40.750 108.095 ;
        RECT 40.930 107.785 41.280 108.155 ;
        RECT 41.450 107.605 41.620 108.335 ;
        RECT 41.790 108.275 42.200 108.715 ;
        RECT 42.490 108.075 42.740 108.505 ;
        RECT 42.940 108.255 43.260 108.715 ;
        RECT 43.820 108.325 44.670 108.495 ;
        RECT 41.790 107.735 42.200 108.065 ;
        RECT 42.490 107.735 42.910 108.075 ;
        RECT 41.200 107.565 41.620 107.605 ;
        RECT 41.200 107.395 42.550 107.565 ;
        RECT 39.610 106.835 40.305 107.005 ;
        RECT 40.530 106.845 41.030 107.225 ;
        RECT 39.635 106.165 39.965 106.665 ;
        RECT 40.135 106.335 40.305 106.835 ;
        RECT 41.200 106.550 41.370 107.395 ;
        RECT 42.300 107.235 42.550 107.395 ;
        RECT 41.540 106.965 41.790 107.225 ;
        RECT 42.720 106.965 42.910 107.735 ;
        RECT 41.540 106.715 42.910 106.965 ;
        RECT 43.080 107.905 44.330 108.075 ;
        RECT 43.080 107.145 43.250 107.905 ;
        RECT 44.000 107.785 44.330 107.905 ;
        RECT 43.420 107.325 43.600 107.735 ;
        RECT 44.500 107.565 44.670 108.325 ;
        RECT 44.870 108.235 45.530 108.715 ;
        RECT 45.710 108.120 46.030 108.450 ;
        RECT 44.860 107.795 45.520 108.065 ;
        RECT 44.860 107.735 45.190 107.795 ;
        RECT 45.340 107.565 45.670 107.625 ;
        RECT 43.770 107.395 45.670 107.565 ;
        RECT 43.080 106.835 43.600 107.145 ;
        RECT 43.770 106.885 43.940 107.395 ;
        RECT 45.840 107.225 46.030 108.120 ;
        RECT 44.110 107.055 46.030 107.225 ;
        RECT 45.710 107.035 46.030 107.055 ;
        RECT 46.230 107.805 46.480 108.455 ;
        RECT 46.660 108.255 46.945 108.715 ;
        RECT 47.125 108.005 47.380 108.535 ;
        RECT 46.230 107.475 47.030 107.805 ;
        RECT 43.770 106.715 44.980 106.885 ;
        RECT 40.540 106.380 41.370 106.550 ;
        RECT 41.610 106.165 41.990 106.545 ;
        RECT 42.170 106.425 42.340 106.715 ;
        RECT 43.770 106.635 43.940 106.715 ;
        RECT 42.510 106.165 42.840 106.545 ;
        RECT 43.310 106.385 43.940 106.635 ;
        RECT 44.120 106.165 44.540 106.545 ;
        RECT 44.740 106.425 44.980 106.715 ;
        RECT 45.210 106.165 45.540 106.855 ;
        RECT 45.710 106.425 45.880 107.035 ;
        RECT 46.230 106.885 46.480 107.475 ;
        RECT 47.200 107.145 47.380 108.005 ;
        RECT 47.985 107.895 48.195 108.715 ;
        RECT 48.365 107.915 48.695 108.545 ;
        RECT 48.365 107.315 48.615 107.915 ;
        RECT 48.865 107.895 49.095 108.715 ;
        RECT 49.395 108.165 49.565 108.545 ;
        RECT 49.745 108.335 50.075 108.715 ;
        RECT 49.395 107.995 50.060 108.165 ;
        RECT 50.255 108.040 50.515 108.545 ;
        RECT 48.785 107.475 49.115 107.725 ;
        RECT 49.325 107.445 49.655 107.815 ;
        RECT 49.890 107.740 50.060 107.995 ;
        RECT 49.890 107.410 50.175 107.740 ;
        RECT 46.150 106.375 46.480 106.885 ;
        RECT 46.660 106.165 46.945 106.965 ;
        RECT 47.125 106.675 47.380 107.145 ;
        RECT 47.125 106.505 47.465 106.675 ;
        RECT 47.125 106.475 47.380 106.505 ;
        RECT 47.985 106.165 48.195 107.305 ;
        RECT 48.365 106.335 48.695 107.315 ;
        RECT 48.865 106.165 49.095 107.305 ;
        RECT 49.890 107.265 50.060 107.410 ;
        RECT 49.395 107.095 50.060 107.265 ;
        RECT 50.345 107.240 50.515 108.040 ;
        RECT 49.395 106.335 49.565 107.095 ;
        RECT 49.745 106.165 50.075 106.925 ;
        RECT 50.245 106.335 50.515 107.240 ;
        RECT 50.690 107.975 50.945 108.545 ;
        RECT 51.115 108.315 51.445 108.715 ;
        RECT 51.870 108.180 52.400 108.545 ;
        RECT 51.870 108.145 52.045 108.180 ;
        RECT 51.115 107.975 52.045 108.145 ;
        RECT 50.690 107.305 50.860 107.975 ;
        RECT 51.115 107.805 51.285 107.975 ;
        RECT 51.030 107.475 51.285 107.805 ;
        RECT 51.510 107.475 51.705 107.805 ;
        RECT 50.690 106.335 51.025 107.305 ;
        RECT 51.195 106.165 51.365 107.305 ;
        RECT 51.535 106.505 51.705 107.475 ;
        RECT 51.875 106.845 52.045 107.975 ;
        RECT 52.215 107.185 52.385 107.985 ;
        RECT 52.590 107.695 52.865 108.545 ;
        RECT 52.585 107.525 52.865 107.695 ;
        RECT 52.590 107.385 52.865 107.525 ;
        RECT 53.035 107.185 53.225 108.545 ;
        RECT 53.405 108.180 53.915 108.715 ;
        RECT 54.135 107.905 54.380 108.510 ;
        RECT 55.285 108.040 55.545 108.545 ;
        RECT 55.725 108.335 56.055 108.715 ;
        RECT 56.235 108.165 56.405 108.545 ;
        RECT 53.425 107.735 54.655 107.905 ;
        RECT 52.215 107.015 53.225 107.185 ;
        RECT 53.395 107.170 54.145 107.360 ;
        RECT 51.875 106.675 53.000 106.845 ;
        RECT 53.395 106.505 53.565 107.170 ;
        RECT 54.315 106.925 54.655 107.735 ;
        RECT 51.535 106.335 53.565 106.505 ;
        RECT 53.735 106.165 53.905 106.925 ;
        RECT 54.140 106.515 54.655 106.925 ;
        RECT 55.285 107.240 55.455 108.040 ;
        RECT 55.740 107.995 56.405 108.165 ;
        RECT 55.740 107.740 55.910 107.995 ;
        RECT 57.125 107.990 57.415 108.715 ;
        RECT 57.590 107.975 57.845 108.545 ;
        RECT 58.015 108.315 58.345 108.715 ;
        RECT 58.770 108.180 59.300 108.545 ;
        RECT 59.490 108.375 59.765 108.545 ;
        RECT 59.485 108.205 59.765 108.375 ;
        RECT 58.770 108.145 58.945 108.180 ;
        RECT 58.015 107.975 58.945 108.145 ;
        RECT 55.625 107.410 55.910 107.740 ;
        RECT 56.145 107.445 56.475 107.815 ;
        RECT 55.740 107.265 55.910 107.410 ;
        RECT 55.285 106.335 55.555 107.240 ;
        RECT 55.740 107.095 56.405 107.265 ;
        RECT 55.725 106.165 56.055 106.925 ;
        RECT 56.235 106.335 56.405 107.095 ;
        RECT 57.125 106.165 57.415 107.330 ;
        RECT 57.590 107.305 57.760 107.975 ;
        RECT 58.015 107.805 58.185 107.975 ;
        RECT 57.930 107.475 58.185 107.805 ;
        RECT 58.410 107.475 58.605 107.805 ;
        RECT 57.590 106.335 57.925 107.305 ;
        RECT 58.095 106.165 58.265 107.305 ;
        RECT 58.435 106.505 58.605 107.475 ;
        RECT 58.775 106.845 58.945 107.975 ;
        RECT 59.115 107.185 59.285 107.985 ;
        RECT 59.490 107.385 59.765 108.205 ;
        RECT 59.935 107.185 60.125 108.545 ;
        RECT 60.305 108.180 60.815 108.715 ;
        RECT 61.035 107.905 61.280 108.510 ;
        RECT 61.725 108.170 67.070 108.715 ;
        RECT 60.325 107.735 61.555 107.905 ;
        RECT 59.115 107.015 60.125 107.185 ;
        RECT 60.295 107.170 61.045 107.360 ;
        RECT 58.775 106.675 59.900 106.845 ;
        RECT 60.295 106.505 60.465 107.170 ;
        RECT 61.215 106.925 61.555 107.735 ;
        RECT 63.310 107.340 63.650 108.170 ;
        RECT 67.245 107.945 68.915 108.715 ;
        RECT 69.635 108.165 69.805 108.545 ;
        RECT 69.985 108.335 70.315 108.715 ;
        RECT 69.635 107.995 70.300 108.165 ;
        RECT 70.495 108.040 70.755 108.545 ;
        RECT 58.435 106.335 60.465 106.505 ;
        RECT 60.635 106.165 60.805 106.925 ;
        RECT 61.040 106.515 61.555 106.925 ;
        RECT 65.130 106.600 65.480 107.850 ;
        RECT 67.245 107.425 67.995 107.945 ;
        RECT 68.165 107.255 68.915 107.775 ;
        RECT 69.565 107.445 69.895 107.815 ;
        RECT 70.130 107.740 70.300 107.995 ;
        RECT 70.130 107.410 70.415 107.740 ;
        RECT 70.130 107.265 70.300 107.410 ;
        RECT 61.725 106.165 67.070 106.600 ;
        RECT 67.245 106.165 68.915 107.255 ;
        RECT 69.635 107.095 70.300 107.265 ;
        RECT 70.585 107.240 70.755 108.040 ;
        RECT 71.885 107.895 72.115 108.715 ;
        RECT 72.285 107.915 72.615 108.545 ;
        RECT 71.865 107.475 72.195 107.725 ;
        RECT 72.365 107.315 72.615 107.915 ;
        RECT 72.785 107.895 72.995 108.715 ;
        RECT 74.150 107.975 74.405 108.545 ;
        RECT 74.575 108.315 74.905 108.715 ;
        RECT 75.330 108.180 75.860 108.545 ;
        RECT 75.330 108.145 75.505 108.180 ;
        RECT 74.575 107.975 75.505 108.145 ;
        RECT 76.050 108.035 76.325 108.545 ;
        RECT 69.635 106.335 69.805 107.095 ;
        RECT 69.985 106.165 70.315 106.925 ;
        RECT 70.485 106.335 70.755 107.240 ;
        RECT 71.885 106.165 72.115 107.305 ;
        RECT 72.285 106.335 72.615 107.315 ;
        RECT 74.150 107.305 74.320 107.975 ;
        RECT 74.575 107.805 74.745 107.975 ;
        RECT 74.490 107.475 74.745 107.805 ;
        RECT 74.970 107.475 75.165 107.805 ;
        RECT 72.785 106.165 72.995 107.305 ;
        RECT 74.150 106.335 74.485 107.305 ;
        RECT 74.655 106.165 74.825 107.305 ;
        RECT 74.995 106.505 75.165 107.475 ;
        RECT 75.335 106.845 75.505 107.975 ;
        RECT 75.675 107.185 75.845 107.985 ;
        RECT 76.045 107.865 76.325 108.035 ;
        RECT 76.050 107.385 76.325 107.865 ;
        RECT 76.495 107.185 76.685 108.545 ;
        RECT 76.865 108.180 77.375 108.715 ;
        RECT 77.595 107.905 77.840 108.510 ;
        RECT 76.885 107.735 78.115 107.905 ;
        RECT 78.345 107.895 78.555 108.715 ;
        RECT 78.725 107.915 79.055 108.545 ;
        RECT 75.675 107.015 76.685 107.185 ;
        RECT 76.855 107.170 77.605 107.360 ;
        RECT 75.335 106.675 76.460 106.845 ;
        RECT 76.855 106.505 77.025 107.170 ;
        RECT 77.775 106.925 78.115 107.735 ;
        RECT 78.725 107.315 78.975 107.915 ;
        RECT 79.225 107.895 79.455 108.715 ;
        RECT 79.755 108.165 79.925 108.545 ;
        RECT 80.105 108.335 80.435 108.715 ;
        RECT 79.755 107.995 80.420 108.165 ;
        RECT 80.615 108.040 80.875 108.545 ;
        RECT 79.145 107.475 79.475 107.725 ;
        RECT 79.685 107.445 80.015 107.815 ;
        RECT 80.250 107.740 80.420 107.995 ;
        RECT 80.250 107.410 80.535 107.740 ;
        RECT 74.995 106.335 77.025 106.505 ;
        RECT 77.195 106.165 77.365 106.925 ;
        RECT 77.600 106.515 78.115 106.925 ;
        RECT 78.345 106.165 78.555 107.305 ;
        RECT 78.725 106.335 79.055 107.315 ;
        RECT 79.225 106.165 79.455 107.305 ;
        RECT 80.250 107.265 80.420 107.410 ;
        RECT 79.755 107.095 80.420 107.265 ;
        RECT 80.705 107.240 80.875 108.040 ;
        RECT 81.045 107.945 82.715 108.715 ;
        RECT 82.885 107.990 83.175 108.715 ;
        RECT 83.345 108.205 83.650 108.715 ;
        RECT 81.045 107.425 81.795 107.945 ;
        RECT 81.965 107.255 82.715 107.775 ;
        RECT 83.345 107.475 83.660 108.035 ;
        RECT 83.830 107.725 84.080 108.535 ;
        RECT 84.250 108.190 84.510 108.715 ;
        RECT 84.690 107.725 84.940 108.535 ;
        RECT 85.110 108.155 85.370 108.715 ;
        RECT 85.540 108.065 85.800 108.520 ;
        RECT 85.970 108.235 86.230 108.715 ;
        RECT 86.400 108.065 86.660 108.520 ;
        RECT 86.830 108.235 87.090 108.715 ;
        RECT 87.260 108.065 87.520 108.520 ;
        RECT 87.690 108.235 87.935 108.715 ;
        RECT 88.105 108.065 88.380 108.520 ;
        RECT 88.550 108.235 88.795 108.715 ;
        RECT 88.965 108.065 89.225 108.520 ;
        RECT 89.405 108.235 89.655 108.715 ;
        RECT 89.825 108.065 90.085 108.520 ;
        RECT 90.265 108.235 90.515 108.715 ;
        RECT 90.685 108.065 90.945 108.520 ;
        RECT 91.125 108.235 91.385 108.715 ;
        RECT 91.555 108.065 91.815 108.520 ;
        RECT 91.985 108.235 92.285 108.715 ;
        RECT 85.540 107.895 92.285 108.065 ;
        RECT 83.830 107.475 90.950 107.725 ;
        RECT 79.755 106.335 79.925 107.095 ;
        RECT 80.105 106.165 80.435 106.925 ;
        RECT 80.605 106.335 80.875 107.240 ;
        RECT 81.045 106.165 82.715 107.255 ;
        RECT 82.885 106.165 83.175 107.330 ;
        RECT 83.355 106.165 83.650 106.975 ;
        RECT 83.830 106.335 84.075 107.475 ;
        RECT 84.250 106.165 84.510 106.975 ;
        RECT 84.690 106.340 84.940 107.475 ;
        RECT 91.120 107.305 92.285 107.895 ;
        RECT 92.545 107.945 95.135 108.715 ;
        RECT 95.855 108.165 96.025 108.455 ;
        RECT 96.195 108.335 96.525 108.715 ;
        RECT 95.855 107.995 96.520 108.165 ;
        RECT 92.545 107.425 93.755 107.945 ;
        RECT 85.540 107.080 92.285 107.305 ;
        RECT 93.925 107.255 95.135 107.775 ;
        RECT 85.540 107.065 90.945 107.080 ;
        RECT 85.110 106.170 85.370 106.965 ;
        RECT 85.540 106.340 85.800 107.065 ;
        RECT 85.970 106.170 86.230 106.895 ;
        RECT 86.400 106.340 86.660 107.065 ;
        RECT 86.830 106.170 87.090 106.895 ;
        RECT 87.260 106.340 87.520 107.065 ;
        RECT 87.690 106.170 87.950 106.895 ;
        RECT 88.120 106.340 88.380 107.065 ;
        RECT 88.550 106.170 88.795 106.895 ;
        RECT 88.965 106.340 89.225 107.065 ;
        RECT 89.410 106.170 89.655 106.895 ;
        RECT 89.825 106.340 90.085 107.065 ;
        RECT 90.270 106.170 90.515 106.895 ;
        RECT 90.685 106.340 90.945 107.065 ;
        RECT 91.130 106.170 91.385 106.895 ;
        RECT 91.555 106.340 91.845 107.080 ;
        RECT 85.110 106.165 91.385 106.170 ;
        RECT 92.015 106.165 92.285 106.910 ;
        RECT 92.545 106.165 95.135 107.255 ;
        RECT 95.770 107.175 96.120 107.825 ;
        RECT 96.290 107.005 96.520 107.995 ;
        RECT 95.855 106.835 96.520 107.005 ;
        RECT 95.855 106.335 96.025 106.835 ;
        RECT 96.195 106.165 96.525 106.665 ;
        RECT 96.695 106.335 96.920 108.455 ;
        RECT 97.135 108.335 97.465 108.715 ;
        RECT 97.635 108.165 97.805 108.495 ;
        RECT 98.105 108.335 99.120 108.535 ;
        RECT 97.110 107.975 97.805 108.165 ;
        RECT 97.110 107.005 97.280 107.975 ;
        RECT 97.450 107.175 97.860 107.795 ;
        RECT 98.030 107.225 98.250 108.095 ;
        RECT 98.430 107.785 98.780 108.155 ;
        RECT 98.950 107.605 99.120 108.335 ;
        RECT 99.290 108.275 99.700 108.715 ;
        RECT 99.990 108.075 100.240 108.505 ;
        RECT 100.440 108.255 100.760 108.715 ;
        RECT 101.320 108.325 102.170 108.495 ;
        RECT 99.290 107.735 99.700 108.065 ;
        RECT 99.990 107.735 100.410 108.075 ;
        RECT 98.700 107.565 99.120 107.605 ;
        RECT 98.700 107.395 100.050 107.565 ;
        RECT 97.110 106.835 97.805 107.005 ;
        RECT 98.030 106.845 98.530 107.225 ;
        RECT 97.135 106.165 97.465 106.665 ;
        RECT 97.635 106.335 97.805 106.835 ;
        RECT 98.700 106.550 98.870 107.395 ;
        RECT 99.800 107.235 100.050 107.395 ;
        RECT 99.040 106.965 99.290 107.225 ;
        RECT 100.220 106.965 100.410 107.735 ;
        RECT 99.040 106.715 100.410 106.965 ;
        RECT 100.580 107.905 101.830 108.075 ;
        RECT 100.580 107.145 100.750 107.905 ;
        RECT 101.500 107.785 101.830 107.905 ;
        RECT 100.920 107.325 101.100 107.735 ;
        RECT 102.000 107.565 102.170 108.325 ;
        RECT 102.370 108.235 103.030 108.715 ;
        RECT 103.210 108.120 103.530 108.450 ;
        RECT 102.360 107.795 103.020 108.065 ;
        RECT 102.360 107.735 102.690 107.795 ;
        RECT 102.840 107.565 103.170 107.625 ;
        RECT 101.270 107.395 103.170 107.565 ;
        RECT 100.580 106.835 101.100 107.145 ;
        RECT 101.270 106.885 101.440 107.395 ;
        RECT 103.340 107.225 103.530 108.120 ;
        RECT 101.610 107.055 103.530 107.225 ;
        RECT 103.210 107.035 103.530 107.055 ;
        RECT 103.730 107.805 103.980 108.455 ;
        RECT 104.160 108.255 104.445 108.715 ;
        RECT 104.625 108.005 104.880 108.535 ;
        RECT 103.730 107.475 104.530 107.805 ;
        RECT 101.270 106.715 102.480 106.885 ;
        RECT 98.040 106.380 98.870 106.550 ;
        RECT 99.110 106.165 99.490 106.545 ;
        RECT 99.670 106.425 99.840 106.715 ;
        RECT 101.270 106.635 101.440 106.715 ;
        RECT 100.010 106.165 100.340 106.545 ;
        RECT 100.810 106.385 101.440 106.635 ;
        RECT 101.620 106.165 102.040 106.545 ;
        RECT 102.240 106.425 102.480 106.715 ;
        RECT 102.710 106.165 103.040 106.855 ;
        RECT 103.210 106.425 103.380 107.035 ;
        RECT 103.730 106.885 103.980 107.475 ;
        RECT 104.700 107.145 104.880 108.005 ;
        RECT 105.485 107.895 105.695 108.715 ;
        RECT 105.865 107.915 106.195 108.545 ;
        RECT 105.865 107.315 106.115 107.915 ;
        RECT 106.365 107.895 106.595 108.715 ;
        RECT 106.805 107.945 108.475 108.715 ;
        RECT 108.645 107.990 108.935 108.715 ;
        RECT 106.285 107.475 106.615 107.725 ;
        RECT 106.805 107.425 107.555 107.945 ;
        RECT 109.165 107.895 109.375 108.715 ;
        RECT 109.545 107.915 109.875 108.545 ;
        RECT 103.650 106.375 103.980 106.885 ;
        RECT 104.160 106.165 104.445 106.965 ;
        RECT 104.625 106.675 104.880 107.145 ;
        RECT 104.625 106.505 104.965 106.675 ;
        RECT 104.625 106.475 104.880 106.505 ;
        RECT 105.485 106.165 105.695 107.305 ;
        RECT 105.865 106.335 106.195 107.315 ;
        RECT 106.365 106.165 106.595 107.305 ;
        RECT 107.725 107.255 108.475 107.775 ;
        RECT 106.805 106.165 108.475 107.255 ;
        RECT 108.645 106.165 108.935 107.330 ;
        RECT 109.545 107.315 109.795 107.915 ;
        RECT 110.045 107.895 110.275 108.715 ;
        RECT 110.485 107.965 111.695 108.715 ;
        RECT 111.865 108.040 112.125 108.545 ;
        RECT 112.305 108.335 112.635 108.715 ;
        RECT 112.815 108.165 112.985 108.545 ;
        RECT 109.965 107.475 110.295 107.725 ;
        RECT 110.485 107.425 111.005 107.965 ;
        RECT 109.165 106.165 109.375 107.305 ;
        RECT 109.545 106.335 109.875 107.315 ;
        RECT 110.045 106.165 110.275 107.305 ;
        RECT 111.175 107.255 111.695 107.795 ;
        RECT 110.485 106.165 111.695 107.255 ;
        RECT 111.865 107.240 112.035 108.040 ;
        RECT 112.320 107.995 112.985 108.165 ;
        RECT 112.320 107.740 112.490 107.995 ;
        RECT 113.245 107.945 114.915 108.715 ;
        RECT 112.205 107.410 112.490 107.740 ;
        RECT 112.725 107.445 113.055 107.815 ;
        RECT 113.245 107.425 113.995 107.945 ;
        RECT 115.820 107.905 116.065 108.510 ;
        RECT 116.285 108.180 116.795 108.715 ;
        RECT 112.320 107.265 112.490 107.410 ;
        RECT 111.865 106.335 112.135 107.240 ;
        RECT 112.320 107.095 112.985 107.265 ;
        RECT 114.165 107.255 114.915 107.775 ;
        RECT 112.305 106.165 112.635 106.925 ;
        RECT 112.815 106.335 112.985 107.095 ;
        RECT 113.245 106.165 114.915 107.255 ;
        RECT 115.545 107.735 116.775 107.905 ;
        RECT 115.545 106.925 115.885 107.735 ;
        RECT 116.055 107.170 116.805 107.360 ;
        RECT 115.545 106.515 116.060 106.925 ;
        RECT 116.295 106.165 116.465 106.925 ;
        RECT 116.635 106.505 116.805 107.170 ;
        RECT 116.975 107.185 117.165 108.545 ;
        RECT 117.335 107.695 117.610 108.545 ;
        RECT 117.800 108.180 118.330 108.545 ;
        RECT 118.755 108.315 119.085 108.715 ;
        RECT 118.155 108.145 118.330 108.180 ;
        RECT 117.335 107.525 117.615 107.695 ;
        RECT 117.335 107.385 117.610 107.525 ;
        RECT 117.815 107.185 117.985 107.985 ;
        RECT 116.975 107.015 117.985 107.185 ;
        RECT 118.155 107.975 119.085 108.145 ;
        RECT 119.255 107.975 119.510 108.545 ;
        RECT 118.155 106.845 118.325 107.975 ;
        RECT 118.915 107.805 119.085 107.975 ;
        RECT 117.200 106.675 118.325 106.845 ;
        RECT 118.495 107.475 118.690 107.805 ;
        RECT 118.915 107.475 119.170 107.805 ;
        RECT 118.495 106.505 118.665 107.475 ;
        RECT 119.340 107.305 119.510 107.975 ;
        RECT 119.685 107.945 123.195 108.715 ;
        RECT 124.285 107.965 125.495 108.715 ;
        RECT 119.685 107.425 121.335 107.945 ;
        RECT 116.635 106.335 118.665 106.505 ;
        RECT 118.835 106.165 119.005 107.305 ;
        RECT 119.175 106.335 119.510 107.305 ;
        RECT 121.505 107.255 123.195 107.775 ;
        RECT 119.685 106.165 123.195 107.255 ;
        RECT 124.285 107.255 124.805 107.795 ;
        RECT 124.975 107.425 125.495 107.965 ;
        RECT 124.285 106.165 125.495 107.255 ;
        RECT 5.520 105.995 125.580 106.165 ;
        RECT 5.605 104.905 6.815 105.995 ;
        RECT 6.985 104.905 8.195 105.995 ;
        RECT 8.455 105.325 8.625 105.825 ;
        RECT 8.795 105.495 9.125 105.995 ;
        RECT 8.455 105.155 9.120 105.325 ;
        RECT 5.605 104.195 6.125 104.735 ;
        RECT 6.295 104.365 6.815 104.905 ;
        RECT 6.985 104.195 7.505 104.735 ;
        RECT 7.675 104.365 8.195 104.905 ;
        RECT 8.370 104.335 8.720 104.985 ;
        RECT 5.605 103.445 6.815 104.195 ;
        RECT 6.985 103.445 8.195 104.195 ;
        RECT 8.890 104.165 9.120 105.155 ;
        RECT 8.455 103.995 9.120 104.165 ;
        RECT 8.455 103.705 8.625 103.995 ;
        RECT 8.795 103.445 9.125 103.825 ;
        RECT 9.295 103.705 9.520 105.825 ;
        RECT 9.735 105.495 10.065 105.995 ;
        RECT 10.235 105.325 10.405 105.825 ;
        RECT 10.640 105.610 11.470 105.780 ;
        RECT 11.710 105.615 12.090 105.995 ;
        RECT 9.710 105.155 10.405 105.325 ;
        RECT 9.710 104.185 9.880 105.155 ;
        RECT 10.050 104.365 10.460 104.985 ;
        RECT 10.630 104.935 11.130 105.315 ;
        RECT 9.710 103.995 10.405 104.185 ;
        RECT 10.630 104.065 10.850 104.935 ;
        RECT 11.300 104.765 11.470 105.610 ;
        RECT 12.270 105.445 12.440 105.735 ;
        RECT 12.610 105.615 12.940 105.995 ;
        RECT 13.410 105.525 14.040 105.775 ;
        RECT 14.220 105.615 14.640 105.995 ;
        RECT 13.870 105.445 14.040 105.525 ;
        RECT 14.840 105.445 15.080 105.735 ;
        RECT 11.640 105.195 13.010 105.445 ;
        RECT 11.640 104.935 11.890 105.195 ;
        RECT 12.400 104.765 12.650 104.925 ;
        RECT 11.300 104.595 12.650 104.765 ;
        RECT 11.300 104.555 11.720 104.595 ;
        RECT 11.030 104.005 11.380 104.375 ;
        RECT 9.735 103.445 10.065 103.825 ;
        RECT 10.235 103.665 10.405 103.995 ;
        RECT 11.550 103.825 11.720 104.555 ;
        RECT 12.820 104.425 13.010 105.195 ;
        RECT 11.890 104.095 12.300 104.425 ;
        RECT 12.590 104.085 13.010 104.425 ;
        RECT 13.180 105.015 13.700 105.325 ;
        RECT 13.870 105.275 15.080 105.445 ;
        RECT 15.310 105.305 15.640 105.995 ;
        RECT 13.180 104.255 13.350 105.015 ;
        RECT 13.520 104.425 13.700 104.835 ;
        RECT 13.870 104.765 14.040 105.275 ;
        RECT 15.810 105.125 15.980 105.735 ;
        RECT 16.250 105.275 16.580 105.785 ;
        RECT 15.810 105.105 16.130 105.125 ;
        RECT 14.210 104.935 16.130 105.105 ;
        RECT 13.870 104.595 15.770 104.765 ;
        RECT 14.100 104.255 14.430 104.375 ;
        RECT 13.180 104.085 14.430 104.255 ;
        RECT 10.705 103.625 11.720 103.825 ;
        RECT 11.890 103.445 12.300 103.885 ;
        RECT 12.590 103.655 12.840 104.085 ;
        RECT 13.040 103.445 13.360 103.905 ;
        RECT 14.600 103.835 14.770 104.595 ;
        RECT 15.440 104.535 15.770 104.595 ;
        RECT 14.960 104.365 15.290 104.425 ;
        RECT 14.960 104.095 15.620 104.365 ;
        RECT 15.940 104.040 16.130 104.935 ;
        RECT 13.920 103.665 14.770 103.835 ;
        RECT 14.970 103.445 15.630 103.925 ;
        RECT 15.810 103.710 16.130 104.040 ;
        RECT 16.330 104.685 16.580 105.275 ;
        RECT 16.760 105.195 17.045 105.995 ;
        RECT 17.225 105.015 17.480 105.685 ;
        RECT 16.330 104.355 17.130 104.685 ;
        RECT 16.330 103.705 16.580 104.355 ;
        RECT 17.300 104.155 17.480 105.015 ;
        RECT 18.485 104.830 18.775 105.995 ;
        RECT 18.950 104.855 19.285 105.825 ;
        RECT 19.455 104.855 19.625 105.995 ;
        RECT 19.795 105.655 21.825 105.825 ;
        RECT 18.950 104.185 19.120 104.855 ;
        RECT 19.795 104.685 19.965 105.655 ;
        RECT 19.290 104.355 19.545 104.685 ;
        RECT 19.770 104.355 19.965 104.685 ;
        RECT 20.135 105.315 21.260 105.485 ;
        RECT 19.375 104.185 19.545 104.355 ;
        RECT 20.135 104.185 20.305 105.315 ;
        RECT 17.225 103.955 17.480 104.155 ;
        RECT 16.760 103.445 17.045 103.905 ;
        RECT 17.225 103.785 17.565 103.955 ;
        RECT 17.225 103.625 17.480 103.785 ;
        RECT 18.485 103.445 18.775 104.170 ;
        RECT 18.950 103.615 19.205 104.185 ;
        RECT 19.375 104.015 20.305 104.185 ;
        RECT 20.475 104.975 21.485 105.145 ;
        RECT 20.475 104.175 20.645 104.975 ;
        RECT 20.130 103.980 20.305 104.015 ;
        RECT 19.375 103.445 19.705 103.845 ;
        RECT 20.130 103.615 20.660 103.980 ;
        RECT 20.850 103.955 21.125 104.775 ;
        RECT 20.845 103.785 21.125 103.955 ;
        RECT 20.850 103.615 21.125 103.785 ;
        RECT 21.295 103.615 21.485 104.975 ;
        RECT 21.655 104.990 21.825 105.655 ;
        RECT 21.995 105.235 22.165 105.995 ;
        RECT 22.400 105.235 22.915 105.645 ;
        RECT 21.655 104.800 22.405 104.990 ;
        RECT 22.575 104.425 22.915 105.235 ;
        RECT 23.085 104.905 24.755 105.995 ;
        RECT 25.015 105.325 25.185 105.825 ;
        RECT 25.355 105.495 25.685 105.995 ;
        RECT 25.015 105.155 25.680 105.325 ;
        RECT 21.685 104.255 22.915 104.425 ;
        RECT 21.665 103.445 22.175 103.980 ;
        RECT 22.395 103.650 22.640 104.255 ;
        RECT 23.085 104.215 23.835 104.735 ;
        RECT 24.005 104.385 24.755 104.905 ;
        RECT 24.930 104.335 25.280 104.985 ;
        RECT 23.085 103.445 24.755 104.215 ;
        RECT 25.450 104.165 25.680 105.155 ;
        RECT 25.015 103.995 25.680 104.165 ;
        RECT 25.015 103.705 25.185 103.995 ;
        RECT 25.355 103.445 25.685 103.825 ;
        RECT 25.855 103.705 26.080 105.825 ;
        RECT 26.295 105.495 26.625 105.995 ;
        RECT 26.795 105.325 26.965 105.825 ;
        RECT 27.200 105.610 28.030 105.780 ;
        RECT 28.270 105.615 28.650 105.995 ;
        RECT 26.270 105.155 26.965 105.325 ;
        RECT 26.270 104.185 26.440 105.155 ;
        RECT 26.610 104.365 27.020 104.985 ;
        RECT 27.190 104.935 27.690 105.315 ;
        RECT 26.270 103.995 26.965 104.185 ;
        RECT 27.190 104.065 27.410 104.935 ;
        RECT 27.860 104.765 28.030 105.610 ;
        RECT 28.830 105.445 29.000 105.735 ;
        RECT 29.170 105.615 29.500 105.995 ;
        RECT 29.970 105.525 30.600 105.775 ;
        RECT 30.780 105.615 31.200 105.995 ;
        RECT 30.430 105.445 30.600 105.525 ;
        RECT 31.400 105.445 31.640 105.735 ;
        RECT 28.200 105.195 29.570 105.445 ;
        RECT 28.200 104.935 28.450 105.195 ;
        RECT 28.960 104.765 29.210 104.925 ;
        RECT 27.860 104.595 29.210 104.765 ;
        RECT 27.860 104.555 28.280 104.595 ;
        RECT 27.590 104.005 27.940 104.375 ;
        RECT 26.295 103.445 26.625 103.825 ;
        RECT 26.795 103.665 26.965 103.995 ;
        RECT 28.110 103.825 28.280 104.555 ;
        RECT 29.380 104.425 29.570 105.195 ;
        RECT 28.450 104.095 28.860 104.425 ;
        RECT 29.150 104.085 29.570 104.425 ;
        RECT 29.740 105.015 30.260 105.325 ;
        RECT 30.430 105.275 31.640 105.445 ;
        RECT 31.870 105.305 32.200 105.995 ;
        RECT 29.740 104.255 29.910 105.015 ;
        RECT 30.080 104.425 30.260 104.835 ;
        RECT 30.430 104.765 30.600 105.275 ;
        RECT 32.370 105.125 32.540 105.735 ;
        RECT 32.810 105.275 33.140 105.785 ;
        RECT 32.370 105.105 32.690 105.125 ;
        RECT 30.770 104.935 32.690 105.105 ;
        RECT 30.430 104.595 32.330 104.765 ;
        RECT 30.660 104.255 30.990 104.375 ;
        RECT 29.740 104.085 30.990 104.255 ;
        RECT 27.265 103.625 28.280 103.825 ;
        RECT 28.450 103.445 28.860 103.885 ;
        RECT 29.150 103.655 29.400 104.085 ;
        RECT 29.600 103.445 29.920 103.905 ;
        RECT 31.160 103.835 31.330 104.595 ;
        RECT 32.000 104.535 32.330 104.595 ;
        RECT 31.520 104.365 31.850 104.425 ;
        RECT 31.520 104.095 32.180 104.365 ;
        RECT 32.500 104.040 32.690 104.935 ;
        RECT 30.480 103.665 31.330 103.835 ;
        RECT 31.530 103.445 32.190 103.925 ;
        RECT 32.370 103.710 32.690 104.040 ;
        RECT 32.890 104.685 33.140 105.275 ;
        RECT 33.320 105.195 33.605 105.995 ;
        RECT 33.785 105.015 34.040 105.685 ;
        RECT 34.585 105.560 39.930 105.995 ;
        RECT 32.890 104.355 33.690 104.685 ;
        RECT 32.890 103.705 33.140 104.355 ;
        RECT 33.860 104.155 34.040 105.015 ;
        RECT 33.785 103.955 34.040 104.155 ;
        RECT 36.170 103.990 36.510 104.820 ;
        RECT 37.990 104.310 38.340 105.560 ;
        RECT 40.105 104.905 43.615 105.995 ;
        RECT 40.105 104.215 41.755 104.735 ;
        RECT 41.925 104.385 43.615 104.905 ;
        RECT 44.245 104.830 44.535 105.995 ;
        RECT 44.710 104.855 45.045 105.825 ;
        RECT 45.215 104.855 45.385 105.995 ;
        RECT 45.555 105.655 47.585 105.825 ;
        RECT 33.320 103.445 33.605 103.905 ;
        RECT 33.785 103.785 34.125 103.955 ;
        RECT 33.785 103.625 34.040 103.785 ;
        RECT 34.585 103.445 39.930 103.990 ;
        RECT 40.105 103.445 43.615 104.215 ;
        RECT 44.710 104.185 44.880 104.855 ;
        RECT 45.555 104.685 45.725 105.655 ;
        RECT 45.050 104.355 45.305 104.685 ;
        RECT 45.530 104.355 45.725 104.685 ;
        RECT 45.895 105.315 47.020 105.485 ;
        RECT 45.135 104.185 45.305 104.355 ;
        RECT 45.895 104.185 46.065 105.315 ;
        RECT 44.245 103.445 44.535 104.170 ;
        RECT 44.710 103.615 44.965 104.185 ;
        RECT 45.135 104.015 46.065 104.185 ;
        RECT 46.235 104.975 47.245 105.145 ;
        RECT 46.235 104.175 46.405 104.975 ;
        RECT 46.610 104.635 46.885 104.775 ;
        RECT 46.605 104.465 46.885 104.635 ;
        RECT 45.890 103.980 46.065 104.015 ;
        RECT 45.135 103.445 45.465 103.845 ;
        RECT 45.890 103.615 46.420 103.980 ;
        RECT 46.610 103.615 46.885 104.465 ;
        RECT 47.055 103.615 47.245 104.975 ;
        RECT 47.415 104.990 47.585 105.655 ;
        RECT 47.755 105.235 47.925 105.995 ;
        RECT 48.160 105.235 48.675 105.645 ;
        RECT 48.845 105.560 54.190 105.995 ;
        RECT 47.415 104.800 48.165 104.990 ;
        RECT 48.335 104.425 48.675 105.235 ;
        RECT 47.445 104.255 48.675 104.425 ;
        RECT 47.425 103.445 47.935 103.980 ;
        RECT 48.155 103.650 48.400 104.255 ;
        RECT 50.430 103.990 50.770 104.820 ;
        RECT 52.250 104.310 52.600 105.560 ;
        RECT 54.365 104.905 56.035 105.995 ;
        RECT 56.865 105.325 57.145 105.995 ;
        RECT 57.315 105.105 57.615 105.655 ;
        RECT 57.815 105.275 58.145 105.995 ;
        RECT 58.335 105.275 58.795 105.825 ;
        RECT 54.365 104.215 55.115 104.735 ;
        RECT 55.285 104.385 56.035 104.905 ;
        RECT 56.680 104.685 56.945 105.045 ;
        RECT 57.315 104.935 58.255 105.105 ;
        RECT 58.085 104.685 58.255 104.935 ;
        RECT 56.680 104.435 57.355 104.685 ;
        RECT 57.575 104.435 57.915 104.685 ;
        RECT 58.085 104.355 58.375 104.685 ;
        RECT 58.085 104.265 58.255 104.355 ;
        RECT 48.845 103.445 54.190 103.990 ;
        RECT 54.365 103.445 56.035 104.215 ;
        RECT 56.865 104.075 58.255 104.265 ;
        RECT 56.865 103.715 57.195 104.075 ;
        RECT 58.545 103.905 58.795 105.275 ;
        RECT 57.815 103.445 58.065 103.905 ;
        RECT 58.235 103.615 58.795 103.905 ;
        RECT 58.965 105.275 59.425 105.825 ;
        RECT 59.615 105.275 59.945 105.995 ;
        RECT 58.965 103.905 59.215 105.275 ;
        RECT 60.145 105.105 60.445 105.655 ;
        RECT 60.615 105.325 60.895 105.995 ;
        RECT 61.265 105.560 66.610 105.995 ;
        RECT 59.505 104.935 60.445 105.105 ;
        RECT 59.505 104.685 59.675 104.935 ;
        RECT 60.815 104.685 61.080 105.045 ;
        RECT 59.385 104.355 59.675 104.685 ;
        RECT 59.845 104.435 60.185 104.685 ;
        RECT 60.405 104.435 61.080 104.685 ;
        RECT 59.505 104.265 59.675 104.355 ;
        RECT 59.505 104.075 60.895 104.265 ;
        RECT 58.965 103.615 59.525 103.905 ;
        RECT 59.695 103.445 59.945 103.905 ;
        RECT 60.565 103.715 60.895 104.075 ;
        RECT 62.850 103.990 63.190 104.820 ;
        RECT 64.670 104.310 65.020 105.560 ;
        RECT 66.785 104.905 69.375 105.995 ;
        RECT 66.785 104.215 67.995 104.735 ;
        RECT 68.165 104.385 69.375 104.905 ;
        RECT 70.005 104.830 70.295 105.995 ;
        RECT 71.390 104.855 71.725 105.825 ;
        RECT 71.895 104.855 72.065 105.995 ;
        RECT 72.235 105.655 74.265 105.825 ;
        RECT 61.265 103.445 66.610 103.990 ;
        RECT 66.785 103.445 69.375 104.215 ;
        RECT 71.390 104.185 71.560 104.855 ;
        RECT 72.235 104.685 72.405 105.655 ;
        RECT 71.730 104.355 71.985 104.685 ;
        RECT 72.210 104.355 72.405 104.685 ;
        RECT 72.575 105.315 73.700 105.485 ;
        RECT 71.815 104.185 71.985 104.355 ;
        RECT 72.575 104.185 72.745 105.315 ;
        RECT 70.005 103.445 70.295 104.170 ;
        RECT 71.390 103.615 71.645 104.185 ;
        RECT 71.815 104.015 72.745 104.185 ;
        RECT 72.915 104.975 73.925 105.145 ;
        RECT 72.915 104.175 73.085 104.975 ;
        RECT 73.290 104.295 73.565 104.775 ;
        RECT 73.285 104.125 73.565 104.295 ;
        RECT 72.570 103.980 72.745 104.015 ;
        RECT 71.815 103.445 72.145 103.845 ;
        RECT 72.570 103.615 73.100 103.980 ;
        RECT 73.290 103.615 73.565 104.125 ;
        RECT 73.735 103.615 73.925 104.975 ;
        RECT 74.095 104.990 74.265 105.655 ;
        RECT 74.435 105.235 74.605 105.995 ;
        RECT 74.840 105.235 75.355 105.645 ;
        RECT 75.525 105.560 80.870 105.995 ;
        RECT 74.095 104.800 74.845 104.990 ;
        RECT 75.015 104.425 75.355 105.235 ;
        RECT 74.125 104.255 75.355 104.425 ;
        RECT 74.105 103.445 74.615 103.980 ;
        RECT 74.835 103.650 75.080 104.255 ;
        RECT 77.110 103.990 77.450 104.820 ;
        RECT 78.930 104.310 79.280 105.560 ;
        RECT 81.045 104.905 82.715 105.995 ;
        RECT 81.045 104.215 81.795 104.735 ;
        RECT 81.965 104.385 82.715 104.905 ;
        RECT 83.350 104.855 83.685 105.825 ;
        RECT 83.855 104.855 84.025 105.995 ;
        RECT 84.195 105.655 86.225 105.825 ;
        RECT 75.525 103.445 80.870 103.990 ;
        RECT 81.045 103.445 82.715 104.215 ;
        RECT 83.350 104.185 83.520 104.855 ;
        RECT 84.195 104.685 84.365 105.655 ;
        RECT 83.690 104.355 83.945 104.685 ;
        RECT 84.170 104.355 84.365 104.685 ;
        RECT 84.535 105.315 85.660 105.485 ;
        RECT 83.775 104.185 83.945 104.355 ;
        RECT 84.535 104.185 84.705 105.315 ;
        RECT 83.350 103.615 83.605 104.185 ;
        RECT 83.775 104.015 84.705 104.185 ;
        RECT 84.875 104.975 85.885 105.145 ;
        RECT 84.875 104.175 85.045 104.975 ;
        RECT 85.250 104.635 85.525 104.775 ;
        RECT 85.245 104.465 85.525 104.635 ;
        RECT 84.530 103.980 84.705 104.015 ;
        RECT 83.775 103.445 84.105 103.845 ;
        RECT 84.530 103.615 85.060 103.980 ;
        RECT 85.250 103.615 85.525 104.465 ;
        RECT 85.695 103.615 85.885 104.975 ;
        RECT 86.055 104.990 86.225 105.655 ;
        RECT 86.395 105.235 86.565 105.995 ;
        RECT 86.800 105.235 87.315 105.645 ;
        RECT 86.055 104.800 86.805 104.990 ;
        RECT 86.975 104.425 87.315 105.235 ;
        RECT 87.485 104.905 89.155 105.995 ;
        RECT 86.085 104.255 87.315 104.425 ;
        RECT 86.065 103.445 86.575 103.980 ;
        RECT 86.795 103.650 87.040 104.255 ;
        RECT 87.485 104.215 88.235 104.735 ;
        RECT 88.405 104.385 89.155 104.905 ;
        RECT 89.325 105.275 89.785 105.825 ;
        RECT 89.975 105.275 90.305 105.995 ;
        RECT 87.485 103.445 89.155 104.215 ;
        RECT 89.325 103.905 89.575 105.275 ;
        RECT 90.505 105.105 90.805 105.655 ;
        RECT 90.975 105.325 91.255 105.995 ;
        RECT 89.865 104.935 90.805 105.105 ;
        RECT 91.625 105.275 92.085 105.825 ;
        RECT 92.275 105.275 92.605 105.995 ;
        RECT 89.865 104.685 90.035 104.935 ;
        RECT 91.175 104.685 91.440 105.045 ;
        RECT 89.745 104.355 90.035 104.685 ;
        RECT 90.205 104.435 90.545 104.685 ;
        RECT 90.765 104.435 91.440 104.685 ;
        RECT 89.865 104.265 90.035 104.355 ;
        RECT 89.865 104.075 91.255 104.265 ;
        RECT 89.325 103.615 89.885 103.905 ;
        RECT 90.055 103.445 90.305 103.905 ;
        RECT 90.925 103.715 91.255 104.075 ;
        RECT 91.625 103.905 91.875 105.275 ;
        RECT 92.805 105.105 93.105 105.655 ;
        RECT 93.275 105.325 93.555 105.995 ;
        RECT 92.165 104.935 93.105 105.105 ;
        RECT 92.165 104.685 92.335 104.935 ;
        RECT 93.475 104.685 93.740 105.045 ;
        RECT 93.925 104.905 95.595 105.995 ;
        RECT 92.045 104.355 92.335 104.685 ;
        RECT 92.505 104.435 92.845 104.685 ;
        RECT 93.065 104.435 93.740 104.685 ;
        RECT 92.165 104.265 92.335 104.355 ;
        RECT 92.165 104.075 93.555 104.265 ;
        RECT 91.625 103.615 92.185 103.905 ;
        RECT 92.355 103.445 92.605 103.905 ;
        RECT 93.225 103.715 93.555 104.075 ;
        RECT 93.925 104.215 94.675 104.735 ;
        RECT 94.845 104.385 95.595 104.905 ;
        RECT 95.765 104.830 96.055 105.995 ;
        RECT 96.315 105.065 96.485 105.825 ;
        RECT 96.665 105.235 96.995 105.995 ;
        RECT 96.315 104.895 96.980 105.065 ;
        RECT 97.165 104.920 97.435 105.825 ;
        RECT 96.810 104.750 96.980 104.895 ;
        RECT 96.245 104.345 96.575 104.715 ;
        RECT 96.810 104.420 97.095 104.750 ;
        RECT 93.925 103.445 95.595 104.215 ;
        RECT 95.765 103.445 96.055 104.170 ;
        RECT 96.810 104.165 96.980 104.420 ;
        RECT 96.315 103.995 96.980 104.165 ;
        RECT 97.265 104.120 97.435 104.920 ;
        RECT 96.315 103.615 96.485 103.995 ;
        RECT 96.665 103.445 96.995 103.825 ;
        RECT 97.175 103.615 97.435 104.120 ;
        RECT 97.610 104.855 97.945 105.825 ;
        RECT 98.115 104.855 98.285 105.995 ;
        RECT 98.455 105.655 100.485 105.825 ;
        RECT 97.610 104.185 97.780 104.855 ;
        RECT 98.455 104.685 98.625 105.655 ;
        RECT 97.950 104.355 98.205 104.685 ;
        RECT 98.430 104.355 98.625 104.685 ;
        RECT 98.795 105.315 99.920 105.485 ;
        RECT 98.035 104.185 98.205 104.355 ;
        RECT 98.795 104.185 98.965 105.315 ;
        RECT 97.610 103.615 97.865 104.185 ;
        RECT 98.035 104.015 98.965 104.185 ;
        RECT 99.135 104.975 100.145 105.145 ;
        RECT 99.135 104.175 99.305 104.975 ;
        RECT 98.790 103.980 98.965 104.015 ;
        RECT 98.035 103.445 98.365 103.845 ;
        RECT 98.790 103.615 99.320 103.980 ;
        RECT 99.510 103.955 99.785 104.775 ;
        RECT 99.505 103.785 99.785 103.955 ;
        RECT 99.510 103.615 99.785 103.785 ;
        RECT 99.955 103.615 100.145 104.975 ;
        RECT 100.315 104.990 100.485 105.655 ;
        RECT 100.655 105.235 100.825 105.995 ;
        RECT 101.060 105.235 101.575 105.645 ;
        RECT 100.315 104.800 101.065 104.990 ;
        RECT 101.235 104.425 101.575 105.235 ;
        RECT 101.745 104.905 102.955 105.995 ;
        RECT 103.135 105.185 103.430 105.995 ;
        RECT 100.345 104.255 101.575 104.425 ;
        RECT 100.325 103.445 100.835 103.980 ;
        RECT 101.055 103.650 101.300 104.255 ;
        RECT 101.745 104.195 102.265 104.735 ;
        RECT 102.435 104.365 102.955 104.905 ;
        RECT 103.610 104.685 103.855 105.825 ;
        RECT 104.030 105.185 104.290 105.995 ;
        RECT 104.890 105.990 111.165 105.995 ;
        RECT 104.470 104.685 104.720 105.820 ;
        RECT 104.890 105.195 105.150 105.990 ;
        RECT 105.320 105.095 105.580 105.820 ;
        RECT 105.750 105.265 106.010 105.990 ;
        RECT 106.180 105.095 106.440 105.820 ;
        RECT 106.610 105.265 106.870 105.990 ;
        RECT 107.040 105.095 107.300 105.820 ;
        RECT 107.470 105.265 107.730 105.990 ;
        RECT 107.900 105.095 108.160 105.820 ;
        RECT 108.330 105.265 108.575 105.990 ;
        RECT 108.745 105.095 109.005 105.820 ;
        RECT 109.190 105.265 109.435 105.990 ;
        RECT 109.605 105.095 109.865 105.820 ;
        RECT 110.050 105.265 110.295 105.990 ;
        RECT 110.465 105.095 110.725 105.820 ;
        RECT 110.910 105.265 111.165 105.990 ;
        RECT 105.320 105.080 110.725 105.095 ;
        RECT 111.335 105.080 111.625 105.820 ;
        RECT 111.795 105.250 112.065 105.995 ;
        RECT 112.325 105.560 117.670 105.995 ;
        RECT 105.320 104.855 112.065 105.080 ;
        RECT 101.745 103.445 102.955 104.195 ;
        RECT 103.125 104.125 103.440 104.685 ;
        RECT 103.610 104.435 110.730 104.685 ;
        RECT 103.125 103.445 103.430 103.955 ;
        RECT 103.610 103.625 103.860 104.435 ;
        RECT 104.030 103.445 104.290 103.970 ;
        RECT 104.470 103.625 104.720 104.435 ;
        RECT 110.900 104.265 112.065 104.855 ;
        RECT 105.320 104.095 112.065 104.265 ;
        RECT 104.890 103.445 105.150 104.005 ;
        RECT 105.320 103.640 105.580 104.095 ;
        RECT 105.750 103.445 106.010 103.925 ;
        RECT 106.180 103.640 106.440 104.095 ;
        RECT 106.610 103.445 106.870 103.925 ;
        RECT 107.040 103.640 107.300 104.095 ;
        RECT 107.470 103.445 107.715 103.925 ;
        RECT 107.885 103.640 108.160 104.095 ;
        RECT 108.330 103.445 108.575 103.925 ;
        RECT 108.745 103.640 109.005 104.095 ;
        RECT 109.185 103.445 109.435 103.925 ;
        RECT 109.605 103.640 109.865 104.095 ;
        RECT 110.045 103.445 110.295 103.925 ;
        RECT 110.465 103.640 110.725 104.095 ;
        RECT 110.905 103.445 111.165 103.925 ;
        RECT 111.335 103.640 111.595 104.095 ;
        RECT 113.910 103.990 114.250 104.820 ;
        RECT 115.730 104.310 116.080 105.560 ;
        RECT 117.845 104.905 121.355 105.995 ;
        RECT 117.845 104.215 119.495 104.735 ;
        RECT 119.665 104.385 121.355 104.905 ;
        RECT 121.525 104.830 121.815 105.995 ;
        RECT 121.985 104.905 123.655 105.995 ;
        RECT 121.985 104.215 122.735 104.735 ;
        RECT 122.905 104.385 123.655 104.905 ;
        RECT 124.285 104.905 125.495 105.995 ;
        RECT 124.285 104.365 124.805 104.905 ;
        RECT 111.765 103.445 112.065 103.925 ;
        RECT 112.325 103.445 117.670 103.990 ;
        RECT 117.845 103.445 121.355 104.215 ;
        RECT 121.525 103.445 121.815 104.170 ;
        RECT 121.985 103.445 123.655 104.215 ;
        RECT 124.975 104.195 125.495 104.735 ;
        RECT 124.285 103.445 125.495 104.195 ;
        RECT 5.520 103.275 125.580 103.445 ;
        RECT 5.605 102.525 6.815 103.275 ;
        RECT 5.605 101.985 6.125 102.525 ;
        RECT 6.985 102.505 9.575 103.275 ;
        RECT 10.295 102.725 10.465 103.015 ;
        RECT 10.635 102.895 10.965 103.275 ;
        RECT 10.295 102.555 10.960 102.725 ;
        RECT 6.295 101.815 6.815 102.355 ;
        RECT 6.985 101.985 8.195 102.505 ;
        RECT 8.365 101.815 9.575 102.335 ;
        RECT 5.605 100.725 6.815 101.815 ;
        RECT 6.985 100.725 9.575 101.815 ;
        RECT 10.210 101.735 10.560 102.385 ;
        RECT 10.730 101.565 10.960 102.555 ;
        RECT 10.295 101.395 10.960 101.565 ;
        RECT 10.295 100.895 10.465 101.395 ;
        RECT 10.635 100.725 10.965 101.225 ;
        RECT 11.135 100.895 11.360 103.015 ;
        RECT 11.575 102.895 11.905 103.275 ;
        RECT 12.075 102.725 12.245 103.055 ;
        RECT 12.545 102.895 13.560 103.095 ;
        RECT 11.550 102.535 12.245 102.725 ;
        RECT 11.550 101.565 11.720 102.535 ;
        RECT 11.890 101.735 12.300 102.355 ;
        RECT 12.470 101.785 12.690 102.655 ;
        RECT 12.870 102.345 13.220 102.715 ;
        RECT 13.390 102.165 13.560 102.895 ;
        RECT 13.730 102.835 14.140 103.275 ;
        RECT 14.430 102.635 14.680 103.065 ;
        RECT 14.880 102.815 15.200 103.275 ;
        RECT 15.760 102.885 16.610 103.055 ;
        RECT 13.730 102.295 14.140 102.625 ;
        RECT 14.430 102.295 14.850 102.635 ;
        RECT 13.140 102.125 13.560 102.165 ;
        RECT 13.140 101.955 14.490 102.125 ;
        RECT 11.550 101.395 12.245 101.565 ;
        RECT 12.470 101.405 12.970 101.785 ;
        RECT 11.575 100.725 11.905 101.225 ;
        RECT 12.075 100.895 12.245 101.395 ;
        RECT 13.140 101.110 13.310 101.955 ;
        RECT 14.240 101.795 14.490 101.955 ;
        RECT 13.480 101.525 13.730 101.785 ;
        RECT 14.660 101.525 14.850 102.295 ;
        RECT 13.480 101.275 14.850 101.525 ;
        RECT 15.020 102.465 16.270 102.635 ;
        RECT 15.020 101.705 15.190 102.465 ;
        RECT 15.940 102.345 16.270 102.465 ;
        RECT 15.360 101.885 15.540 102.295 ;
        RECT 16.440 102.125 16.610 102.885 ;
        RECT 16.810 102.795 17.470 103.275 ;
        RECT 17.650 102.680 17.970 103.010 ;
        RECT 16.800 102.355 17.460 102.625 ;
        RECT 16.800 102.295 17.130 102.355 ;
        RECT 17.280 102.125 17.610 102.185 ;
        RECT 15.710 101.955 17.610 102.125 ;
        RECT 15.020 101.395 15.540 101.705 ;
        RECT 15.710 101.445 15.880 101.955 ;
        RECT 17.780 101.785 17.970 102.680 ;
        RECT 16.050 101.615 17.970 101.785 ;
        RECT 17.650 101.595 17.970 101.615 ;
        RECT 18.170 102.365 18.420 103.015 ;
        RECT 18.600 102.815 18.885 103.275 ;
        RECT 19.065 102.935 19.320 103.095 ;
        RECT 19.065 102.765 19.405 102.935 ;
        RECT 19.065 102.565 19.320 102.765 ;
        RECT 18.170 102.035 18.970 102.365 ;
        RECT 15.710 101.275 16.920 101.445 ;
        RECT 12.480 100.940 13.310 101.110 ;
        RECT 13.550 100.725 13.930 101.105 ;
        RECT 14.110 100.985 14.280 101.275 ;
        RECT 15.710 101.195 15.880 101.275 ;
        RECT 14.450 100.725 14.780 101.105 ;
        RECT 15.250 100.945 15.880 101.195 ;
        RECT 16.060 100.725 16.480 101.105 ;
        RECT 16.680 100.985 16.920 101.275 ;
        RECT 17.150 100.725 17.480 101.415 ;
        RECT 17.650 100.985 17.820 101.595 ;
        RECT 18.170 101.445 18.420 102.035 ;
        RECT 19.140 101.705 19.320 102.565 ;
        RECT 19.865 102.505 23.375 103.275 ;
        RECT 23.545 102.525 24.755 103.275 ;
        RECT 24.930 102.535 25.185 103.105 ;
        RECT 25.355 102.875 25.685 103.275 ;
        RECT 26.110 102.740 26.640 103.105 ;
        RECT 26.830 102.935 27.105 103.105 ;
        RECT 26.825 102.765 27.105 102.935 ;
        RECT 26.110 102.705 26.285 102.740 ;
        RECT 25.355 102.535 26.285 102.705 ;
        RECT 19.865 101.985 21.515 102.505 ;
        RECT 21.685 101.815 23.375 102.335 ;
        RECT 23.545 101.985 24.065 102.525 ;
        RECT 24.235 101.815 24.755 102.355 ;
        RECT 18.090 100.935 18.420 101.445 ;
        RECT 18.600 100.725 18.885 101.525 ;
        RECT 19.065 101.035 19.320 101.705 ;
        RECT 19.865 100.725 23.375 101.815 ;
        RECT 23.545 100.725 24.755 101.815 ;
        RECT 24.930 101.865 25.100 102.535 ;
        RECT 25.355 102.365 25.525 102.535 ;
        RECT 25.270 102.035 25.525 102.365 ;
        RECT 25.750 102.035 25.945 102.365 ;
        RECT 24.930 100.895 25.265 101.865 ;
        RECT 25.435 100.725 25.605 101.865 ;
        RECT 25.775 101.065 25.945 102.035 ;
        RECT 26.115 101.405 26.285 102.535 ;
        RECT 26.455 101.745 26.625 102.545 ;
        RECT 26.830 101.945 27.105 102.765 ;
        RECT 27.275 101.745 27.465 103.105 ;
        RECT 27.645 102.740 28.155 103.275 ;
        RECT 28.375 102.465 28.620 103.070 ;
        RECT 29.065 102.505 30.735 103.275 ;
        RECT 31.365 102.550 31.655 103.275 ;
        RECT 31.825 102.730 37.170 103.275 ;
        RECT 37.345 102.730 42.690 103.275 ;
        RECT 27.665 102.295 28.895 102.465 ;
        RECT 26.455 101.575 27.465 101.745 ;
        RECT 27.635 101.730 28.385 101.920 ;
        RECT 26.115 101.235 27.240 101.405 ;
        RECT 27.635 101.065 27.805 101.730 ;
        RECT 28.555 101.485 28.895 102.295 ;
        RECT 29.065 101.985 29.815 102.505 ;
        RECT 29.985 101.815 30.735 102.335 ;
        RECT 33.410 101.900 33.750 102.730 ;
        RECT 25.775 100.895 27.805 101.065 ;
        RECT 27.975 100.725 28.145 101.485 ;
        RECT 28.380 101.075 28.895 101.485 ;
        RECT 29.065 100.725 30.735 101.815 ;
        RECT 31.365 100.725 31.655 101.890 ;
        RECT 35.230 101.160 35.580 102.410 ;
        RECT 38.930 101.900 39.270 102.730 ;
        RECT 42.865 102.505 46.375 103.275 ;
        RECT 46.545 102.525 47.755 103.275 ;
        RECT 40.750 101.160 41.100 102.410 ;
        RECT 42.865 101.985 44.515 102.505 ;
        RECT 44.685 101.815 46.375 102.335 ;
        RECT 46.545 101.985 47.065 102.525 ;
        RECT 47.965 102.455 48.195 103.275 ;
        RECT 48.365 102.475 48.695 103.105 ;
        RECT 47.235 101.815 47.755 102.355 ;
        RECT 47.945 102.035 48.275 102.285 ;
        RECT 48.445 101.875 48.695 102.475 ;
        RECT 48.865 102.455 49.075 103.275 ;
        RECT 49.305 102.730 54.650 103.275 ;
        RECT 50.890 101.900 51.230 102.730 ;
        RECT 55.025 102.645 55.355 103.005 ;
        RECT 55.975 102.815 56.225 103.275 ;
        RECT 56.395 102.815 56.955 103.105 ;
        RECT 55.025 102.455 56.415 102.645 ;
        RECT 31.825 100.725 37.170 101.160 ;
        RECT 37.345 100.725 42.690 101.160 ;
        RECT 42.865 100.725 46.375 101.815 ;
        RECT 46.545 100.725 47.755 101.815 ;
        RECT 47.965 100.725 48.195 101.865 ;
        RECT 48.365 100.895 48.695 101.875 ;
        RECT 48.865 100.725 49.075 101.865 ;
        RECT 52.710 101.160 53.060 102.410 ;
        RECT 56.245 102.365 56.415 102.455 ;
        RECT 54.840 102.035 55.515 102.285 ;
        RECT 55.735 102.035 56.075 102.285 ;
        RECT 56.245 102.035 56.535 102.365 ;
        RECT 54.840 101.675 55.105 102.035 ;
        RECT 56.245 101.785 56.415 102.035 ;
        RECT 55.475 101.615 56.415 101.785 ;
        RECT 49.305 100.725 54.650 101.160 ;
        RECT 55.025 100.725 55.305 101.395 ;
        RECT 55.475 101.065 55.775 101.615 ;
        RECT 56.705 101.445 56.955 102.815 ;
        RECT 57.125 102.550 57.415 103.275 ;
        RECT 57.585 102.815 58.145 103.105 ;
        RECT 58.315 102.815 58.565 103.275 ;
        RECT 55.975 100.725 56.305 101.445 ;
        RECT 56.495 100.895 56.955 101.445 ;
        RECT 57.125 100.725 57.415 101.890 ;
        RECT 57.585 101.445 57.835 102.815 ;
        RECT 59.185 102.645 59.515 103.005 ;
        RECT 58.125 102.455 59.515 102.645 ;
        RECT 59.885 102.505 61.555 103.275 ;
        RECT 62.245 102.795 62.525 103.275 ;
        RECT 62.695 102.625 62.955 103.015 ;
        RECT 63.130 102.795 63.385 103.275 ;
        RECT 63.555 102.625 63.850 103.015 ;
        RECT 64.030 102.795 64.305 103.275 ;
        RECT 64.475 102.775 64.775 103.105 ;
        RECT 58.125 102.365 58.295 102.455 ;
        RECT 58.005 102.035 58.295 102.365 ;
        RECT 58.465 102.035 58.805 102.285 ;
        RECT 59.025 102.035 59.700 102.285 ;
        RECT 58.125 101.785 58.295 102.035 ;
        RECT 58.125 101.615 59.065 101.785 ;
        RECT 59.435 101.675 59.700 102.035 ;
        RECT 59.885 101.985 60.635 102.505 ;
        RECT 62.200 102.455 63.850 102.625 ;
        RECT 60.805 101.815 61.555 102.335 ;
        RECT 57.585 100.895 58.045 101.445 ;
        RECT 58.235 100.725 58.565 101.445 ;
        RECT 58.765 101.065 59.065 101.615 ;
        RECT 59.235 100.725 59.515 101.395 ;
        RECT 59.885 100.725 61.555 101.815 ;
        RECT 62.200 101.945 62.605 102.455 ;
        RECT 62.775 102.115 63.915 102.285 ;
        RECT 62.200 101.775 62.955 101.945 ;
        RECT 62.240 100.725 62.525 101.595 ;
        RECT 62.695 101.525 62.955 101.775 ;
        RECT 63.745 101.865 63.915 102.115 ;
        RECT 64.085 102.035 64.435 102.605 ;
        RECT 64.605 101.865 64.775 102.775 ;
        RECT 64.945 102.730 70.290 103.275 ;
        RECT 70.465 102.730 75.810 103.275 ;
        RECT 75.985 102.730 81.330 103.275 ;
        RECT 66.530 101.900 66.870 102.730 ;
        RECT 63.745 101.695 64.775 101.865 ;
        RECT 62.695 101.355 63.815 101.525 ;
        RECT 62.695 100.895 62.955 101.355 ;
        RECT 63.130 100.725 63.385 101.185 ;
        RECT 63.555 100.895 63.815 101.355 ;
        RECT 63.985 100.725 64.295 101.525 ;
        RECT 64.465 100.895 64.775 101.695 ;
        RECT 68.350 101.160 68.700 102.410 ;
        RECT 72.050 101.900 72.390 102.730 ;
        RECT 73.870 101.160 74.220 102.410 ;
        RECT 77.570 101.900 77.910 102.730 ;
        RECT 81.505 102.525 82.715 103.275 ;
        RECT 82.885 102.550 83.175 103.275 ;
        RECT 79.390 101.160 79.740 102.410 ;
        RECT 81.505 101.985 82.025 102.525 ;
        RECT 83.345 102.505 85.935 103.275 ;
        RECT 86.115 102.775 86.445 103.275 ;
        RECT 86.645 102.705 86.815 103.055 ;
        RECT 87.015 102.875 87.345 103.275 ;
        RECT 87.515 102.705 87.685 103.055 ;
        RECT 87.855 102.875 88.235 103.275 ;
        RECT 82.195 101.815 82.715 102.355 ;
        RECT 83.345 101.985 84.555 102.505 ;
        RECT 64.945 100.725 70.290 101.160 ;
        RECT 70.465 100.725 75.810 101.160 ;
        RECT 75.985 100.725 81.330 101.160 ;
        RECT 81.505 100.725 82.715 101.815 ;
        RECT 82.885 100.725 83.175 101.890 ;
        RECT 84.725 101.815 85.935 102.335 ;
        RECT 86.110 102.035 86.460 102.605 ;
        RECT 86.645 102.535 88.255 102.705 ;
        RECT 88.425 102.600 88.695 102.945 ;
        RECT 88.875 102.775 89.205 103.275 ;
        RECT 89.405 102.705 89.575 103.055 ;
        RECT 89.775 102.875 90.105 103.275 ;
        RECT 90.275 102.705 90.445 103.055 ;
        RECT 90.615 102.875 90.995 103.275 ;
        RECT 88.085 102.365 88.255 102.535 ;
        RECT 83.345 100.725 85.935 101.815 ;
        RECT 86.110 101.575 86.430 101.865 ;
        RECT 86.630 101.745 87.340 102.365 ;
        RECT 87.510 102.035 87.915 102.365 ;
        RECT 88.085 102.035 88.355 102.365 ;
        RECT 88.085 101.865 88.255 102.035 ;
        RECT 88.525 101.865 88.695 102.600 ;
        RECT 88.870 102.035 89.220 102.605 ;
        RECT 89.405 102.535 91.015 102.705 ;
        RECT 91.185 102.600 91.455 102.945 ;
        RECT 90.845 102.365 91.015 102.535 ;
        RECT 87.530 101.695 88.255 101.865 ;
        RECT 87.530 101.575 87.700 101.695 ;
        RECT 86.110 101.405 87.700 101.575 ;
        RECT 86.110 100.945 87.765 101.235 ;
        RECT 87.935 100.725 88.215 101.525 ;
        RECT 88.425 100.895 88.695 101.865 ;
        RECT 88.870 101.575 89.190 101.865 ;
        RECT 89.390 101.745 90.100 102.365 ;
        RECT 90.270 102.035 90.675 102.365 ;
        RECT 90.845 102.035 91.115 102.365 ;
        RECT 90.845 101.865 91.015 102.035 ;
        RECT 91.285 101.865 91.455 102.600 ;
        RECT 90.290 101.695 91.015 101.865 ;
        RECT 90.290 101.575 90.460 101.695 ;
        RECT 88.870 101.405 90.460 101.575 ;
        RECT 88.870 100.945 90.525 101.235 ;
        RECT 90.695 100.725 90.975 101.525 ;
        RECT 91.185 100.895 91.455 101.865 ;
        RECT 92.085 102.815 92.645 103.105 ;
        RECT 92.815 102.815 93.065 103.275 ;
        RECT 92.085 101.445 92.335 102.815 ;
        RECT 93.685 102.645 94.015 103.005 ;
        RECT 92.625 102.455 94.015 102.645 ;
        RECT 94.385 102.815 94.945 103.105 ;
        RECT 95.115 102.815 95.365 103.275 ;
        RECT 92.625 102.365 92.795 102.455 ;
        RECT 92.505 102.035 92.795 102.365 ;
        RECT 92.965 102.035 93.305 102.285 ;
        RECT 93.525 102.035 94.200 102.285 ;
        RECT 92.625 101.785 92.795 102.035 ;
        RECT 92.625 101.615 93.565 101.785 ;
        RECT 93.935 101.675 94.200 102.035 ;
        RECT 92.085 100.895 92.545 101.445 ;
        RECT 92.735 100.725 93.065 101.445 ;
        RECT 93.265 101.065 93.565 101.615 ;
        RECT 94.385 101.445 94.635 102.815 ;
        RECT 95.985 102.645 96.315 103.005 ;
        RECT 96.685 102.730 102.030 103.275 ;
        RECT 102.205 102.730 107.550 103.275 ;
        RECT 94.925 102.455 96.315 102.645 ;
        RECT 94.925 102.365 95.095 102.455 ;
        RECT 94.805 102.035 95.095 102.365 ;
        RECT 95.265 102.035 95.605 102.285 ;
        RECT 95.825 102.035 96.500 102.285 ;
        RECT 94.925 101.785 95.095 102.035 ;
        RECT 94.925 101.615 95.865 101.785 ;
        RECT 96.235 101.675 96.500 102.035 ;
        RECT 98.270 101.900 98.610 102.730 ;
        RECT 93.735 100.725 94.015 101.395 ;
        RECT 94.385 100.895 94.845 101.445 ;
        RECT 95.035 100.725 95.365 101.445 ;
        RECT 95.565 101.065 95.865 101.615 ;
        RECT 96.035 100.725 96.315 101.395 ;
        RECT 100.090 101.160 100.440 102.410 ;
        RECT 103.790 101.900 104.130 102.730 ;
        RECT 108.645 102.550 108.935 103.275 ;
        RECT 109.105 102.525 110.315 103.275 ;
        RECT 105.610 101.160 105.960 102.410 ;
        RECT 109.105 101.985 109.625 102.525 ;
        RECT 110.545 102.455 110.755 103.275 ;
        RECT 110.925 102.475 111.255 103.105 ;
        RECT 96.685 100.725 102.030 101.160 ;
        RECT 102.205 100.725 107.550 101.160 ;
        RECT 108.645 100.725 108.935 101.890 ;
        RECT 109.795 101.815 110.315 102.355 ;
        RECT 110.925 101.875 111.175 102.475 ;
        RECT 111.425 102.455 111.655 103.275 ;
        RECT 111.865 102.730 117.210 103.275 ;
        RECT 117.385 102.730 122.730 103.275 ;
        RECT 111.345 102.035 111.675 102.285 ;
        RECT 113.450 101.900 113.790 102.730 ;
        RECT 109.105 100.725 110.315 101.815 ;
        RECT 110.545 100.725 110.755 101.865 ;
        RECT 110.925 100.895 111.255 101.875 ;
        RECT 111.425 100.725 111.655 101.865 ;
        RECT 115.270 101.160 115.620 102.410 ;
        RECT 118.970 101.900 119.310 102.730 ;
        RECT 122.905 102.525 124.115 103.275 ;
        RECT 124.285 102.525 125.495 103.275 ;
        RECT 120.790 101.160 121.140 102.410 ;
        RECT 122.905 101.985 123.425 102.525 ;
        RECT 123.595 101.815 124.115 102.355 ;
        RECT 111.865 100.725 117.210 101.160 ;
        RECT 117.385 100.725 122.730 101.160 ;
        RECT 122.905 100.725 124.115 101.815 ;
        RECT 124.285 101.815 124.805 102.355 ;
        RECT 124.975 101.985 125.495 102.525 ;
        RECT 124.285 100.725 125.495 101.815 ;
        RECT 5.520 100.555 125.580 100.725 ;
        RECT 5.605 99.465 6.815 100.555 ;
        RECT 6.985 100.120 12.330 100.555 ;
        RECT 5.605 98.755 6.125 99.295 ;
        RECT 6.295 98.925 6.815 99.465 ;
        RECT 5.605 98.005 6.815 98.755 ;
        RECT 8.570 98.550 8.910 99.380 ;
        RECT 10.390 98.870 10.740 100.120 ;
        RECT 12.505 99.465 14.175 100.555 ;
        RECT 12.505 98.775 13.255 99.295 ;
        RECT 13.425 98.945 14.175 99.465 ;
        RECT 14.405 99.415 14.615 100.555 ;
        RECT 14.785 99.405 15.115 100.385 ;
        RECT 15.285 99.415 15.515 100.555 ;
        RECT 15.725 99.465 18.315 100.555 ;
        RECT 6.985 98.005 12.330 98.550 ;
        RECT 12.505 98.005 14.175 98.775 ;
        RECT 14.405 98.005 14.615 98.825 ;
        RECT 14.785 98.805 15.035 99.405 ;
        RECT 15.205 98.995 15.535 99.245 ;
        RECT 14.785 98.175 15.115 98.805 ;
        RECT 15.285 98.005 15.515 98.825 ;
        RECT 15.725 98.775 16.935 99.295 ;
        RECT 17.105 98.945 18.315 99.465 ;
        RECT 18.485 99.390 18.775 100.555 ;
        RECT 18.945 99.465 20.615 100.555 ;
        RECT 21.445 99.885 21.725 100.555 ;
        RECT 21.895 99.665 22.195 100.215 ;
        RECT 22.395 99.835 22.725 100.555 ;
        RECT 22.915 99.835 23.375 100.385 ;
        RECT 23.745 99.885 24.025 100.555 ;
        RECT 18.945 98.775 19.695 99.295 ;
        RECT 19.865 98.945 20.615 99.465 ;
        RECT 21.260 99.245 21.525 99.605 ;
        RECT 21.895 99.495 22.835 99.665 ;
        RECT 22.665 99.245 22.835 99.495 ;
        RECT 21.260 98.995 21.935 99.245 ;
        RECT 22.155 98.995 22.495 99.245 ;
        RECT 22.665 98.915 22.955 99.245 ;
        RECT 22.665 98.825 22.835 98.915 ;
        RECT 15.725 98.005 18.315 98.775 ;
        RECT 18.485 98.005 18.775 98.730 ;
        RECT 18.945 98.005 20.615 98.775 ;
        RECT 21.445 98.635 22.835 98.825 ;
        RECT 21.445 98.275 21.775 98.635 ;
        RECT 23.125 98.465 23.375 99.835 ;
        RECT 24.195 99.665 24.495 100.215 ;
        RECT 24.695 99.835 25.025 100.555 ;
        RECT 25.215 99.835 25.675 100.385 ;
        RECT 23.560 99.245 23.825 99.605 ;
        RECT 24.195 99.495 25.135 99.665 ;
        RECT 24.965 99.245 25.135 99.495 ;
        RECT 23.560 98.995 24.235 99.245 ;
        RECT 24.455 98.995 24.795 99.245 ;
        RECT 24.965 98.915 25.255 99.245 ;
        RECT 24.965 98.825 25.135 98.915 ;
        RECT 22.395 98.005 22.645 98.465 ;
        RECT 22.815 98.175 23.375 98.465 ;
        RECT 23.745 98.635 25.135 98.825 ;
        RECT 23.745 98.275 24.075 98.635 ;
        RECT 25.425 98.465 25.675 99.835 ;
        RECT 24.695 98.005 24.945 98.465 ;
        RECT 25.115 98.175 25.675 98.465 ;
        RECT 25.845 99.835 26.305 100.385 ;
        RECT 26.495 99.835 26.825 100.555 ;
        RECT 25.845 98.465 26.095 99.835 ;
        RECT 27.025 99.665 27.325 100.215 ;
        RECT 27.495 99.885 27.775 100.555 ;
        RECT 28.345 99.885 28.625 100.555 ;
        RECT 26.385 99.495 27.325 99.665 ;
        RECT 28.795 99.665 29.095 100.215 ;
        RECT 29.295 99.835 29.625 100.555 ;
        RECT 29.815 99.835 30.275 100.385 ;
        RECT 26.385 99.245 26.555 99.495 ;
        RECT 27.695 99.245 27.960 99.605 ;
        RECT 26.265 98.915 26.555 99.245 ;
        RECT 26.725 98.995 27.065 99.245 ;
        RECT 27.285 98.995 27.960 99.245 ;
        RECT 28.160 99.245 28.425 99.605 ;
        RECT 28.795 99.495 29.735 99.665 ;
        RECT 29.565 99.245 29.735 99.495 ;
        RECT 28.160 98.995 28.835 99.245 ;
        RECT 29.055 98.995 29.395 99.245 ;
        RECT 26.385 98.825 26.555 98.915 ;
        RECT 29.565 98.915 29.855 99.245 ;
        RECT 29.565 98.825 29.735 98.915 ;
        RECT 26.385 98.635 27.775 98.825 ;
        RECT 25.845 98.175 26.405 98.465 ;
        RECT 26.575 98.005 26.825 98.465 ;
        RECT 27.445 98.275 27.775 98.635 ;
        RECT 28.345 98.635 29.735 98.825 ;
        RECT 28.345 98.275 28.675 98.635 ;
        RECT 30.025 98.465 30.275 99.835 ;
        RECT 29.295 98.005 29.545 98.465 ;
        RECT 29.715 98.175 30.275 98.465 ;
        RECT 30.445 99.835 30.905 100.385 ;
        RECT 31.095 99.835 31.425 100.555 ;
        RECT 30.445 98.465 30.695 99.835 ;
        RECT 31.625 99.665 31.925 100.215 ;
        RECT 32.095 99.885 32.375 100.555 ;
        RECT 30.985 99.495 31.925 99.665 ;
        RECT 30.985 99.245 31.155 99.495 ;
        RECT 32.295 99.245 32.560 99.605 ;
        RECT 32.745 99.465 36.255 100.555 ;
        RECT 36.625 99.885 36.905 100.555 ;
        RECT 37.075 99.665 37.375 100.215 ;
        RECT 37.575 99.835 37.905 100.555 ;
        RECT 38.095 99.835 38.555 100.385 ;
        RECT 30.865 98.915 31.155 99.245 ;
        RECT 31.325 98.995 31.665 99.245 ;
        RECT 31.885 98.995 32.560 99.245 ;
        RECT 30.985 98.825 31.155 98.915 ;
        RECT 30.985 98.635 32.375 98.825 ;
        RECT 30.445 98.175 31.005 98.465 ;
        RECT 31.175 98.005 31.425 98.465 ;
        RECT 32.045 98.275 32.375 98.635 ;
        RECT 32.745 98.775 34.395 99.295 ;
        RECT 34.565 98.945 36.255 99.465 ;
        RECT 36.440 99.245 36.705 99.605 ;
        RECT 37.075 99.495 38.015 99.665 ;
        RECT 37.845 99.245 38.015 99.495 ;
        RECT 36.440 98.995 37.115 99.245 ;
        RECT 37.335 98.995 37.675 99.245 ;
        RECT 37.845 98.915 38.135 99.245 ;
        RECT 37.845 98.825 38.015 98.915 ;
        RECT 32.745 98.005 36.255 98.775 ;
        RECT 36.625 98.635 38.015 98.825 ;
        RECT 36.625 98.275 36.955 98.635 ;
        RECT 38.305 98.465 38.555 99.835 ;
        RECT 38.815 99.625 38.985 100.385 ;
        RECT 39.165 99.795 39.495 100.555 ;
        RECT 38.815 99.455 39.480 99.625 ;
        RECT 39.665 99.480 39.935 100.385 ;
        RECT 39.310 99.310 39.480 99.455 ;
        RECT 38.745 98.905 39.075 99.275 ;
        RECT 39.310 98.980 39.595 99.310 ;
        RECT 39.310 98.725 39.480 98.980 ;
        RECT 37.575 98.005 37.825 98.465 ;
        RECT 37.995 98.175 38.555 98.465 ;
        RECT 38.815 98.555 39.480 98.725 ;
        RECT 39.765 98.680 39.935 99.480 ;
        RECT 40.105 99.465 43.615 100.555 ;
        RECT 38.815 98.175 38.985 98.555 ;
        RECT 39.165 98.005 39.495 98.385 ;
        RECT 39.675 98.175 39.935 98.680 ;
        RECT 40.105 98.775 41.755 99.295 ;
        RECT 41.925 98.945 43.615 99.465 ;
        RECT 44.245 99.390 44.535 100.555 ;
        RECT 44.795 99.885 44.965 100.385 ;
        RECT 45.135 100.055 45.465 100.555 ;
        RECT 44.795 99.715 45.460 99.885 ;
        RECT 44.710 98.895 45.060 99.545 ;
        RECT 40.105 98.005 43.615 98.775 ;
        RECT 44.245 98.005 44.535 98.730 ;
        RECT 45.230 98.725 45.460 99.715 ;
        RECT 44.795 98.555 45.460 98.725 ;
        RECT 44.795 98.265 44.965 98.555 ;
        RECT 45.135 98.005 45.465 98.385 ;
        RECT 45.635 98.265 45.860 100.385 ;
        RECT 46.075 100.055 46.405 100.555 ;
        RECT 46.575 99.885 46.745 100.385 ;
        RECT 46.980 100.170 47.810 100.340 ;
        RECT 48.050 100.175 48.430 100.555 ;
        RECT 46.050 99.715 46.745 99.885 ;
        RECT 46.050 98.745 46.220 99.715 ;
        RECT 46.390 98.925 46.800 99.545 ;
        RECT 46.970 99.495 47.470 99.875 ;
        RECT 46.050 98.555 46.745 98.745 ;
        RECT 46.970 98.625 47.190 99.495 ;
        RECT 47.640 99.325 47.810 100.170 ;
        RECT 48.610 100.005 48.780 100.295 ;
        RECT 48.950 100.175 49.280 100.555 ;
        RECT 49.750 100.085 50.380 100.335 ;
        RECT 50.560 100.175 50.980 100.555 ;
        RECT 50.210 100.005 50.380 100.085 ;
        RECT 51.180 100.005 51.420 100.295 ;
        RECT 47.980 99.755 49.350 100.005 ;
        RECT 47.980 99.495 48.230 99.755 ;
        RECT 48.740 99.325 48.990 99.485 ;
        RECT 47.640 99.155 48.990 99.325 ;
        RECT 47.640 99.115 48.060 99.155 ;
        RECT 47.370 98.565 47.720 98.935 ;
        RECT 46.075 98.005 46.405 98.385 ;
        RECT 46.575 98.225 46.745 98.555 ;
        RECT 47.890 98.385 48.060 99.115 ;
        RECT 49.160 98.985 49.350 99.755 ;
        RECT 48.230 98.655 48.640 98.985 ;
        RECT 48.930 98.645 49.350 98.985 ;
        RECT 49.520 99.575 50.040 99.885 ;
        RECT 50.210 99.835 51.420 100.005 ;
        RECT 51.650 99.865 51.980 100.555 ;
        RECT 49.520 98.815 49.690 99.575 ;
        RECT 49.860 98.985 50.040 99.395 ;
        RECT 50.210 99.325 50.380 99.835 ;
        RECT 52.150 99.685 52.320 100.295 ;
        RECT 52.590 99.835 52.920 100.345 ;
        RECT 52.150 99.665 52.470 99.685 ;
        RECT 50.550 99.495 52.470 99.665 ;
        RECT 50.210 99.155 52.110 99.325 ;
        RECT 50.440 98.815 50.770 98.935 ;
        RECT 49.520 98.645 50.770 98.815 ;
        RECT 47.045 98.185 48.060 98.385 ;
        RECT 48.230 98.005 48.640 98.445 ;
        RECT 48.930 98.215 49.180 98.645 ;
        RECT 49.380 98.005 49.700 98.465 ;
        RECT 50.940 98.395 51.110 99.155 ;
        RECT 51.780 99.095 52.110 99.155 ;
        RECT 51.300 98.925 51.630 98.985 ;
        RECT 51.300 98.655 51.960 98.925 ;
        RECT 52.280 98.600 52.470 99.495 ;
        RECT 50.260 98.225 51.110 98.395 ;
        RECT 51.310 98.005 51.970 98.485 ;
        RECT 52.150 98.270 52.470 98.600 ;
        RECT 52.670 99.245 52.920 99.835 ;
        RECT 53.100 99.755 53.385 100.555 ;
        RECT 53.565 99.575 53.820 100.245 ;
        RECT 52.670 98.915 53.470 99.245 ;
        RECT 52.670 98.265 52.920 98.915 ;
        RECT 53.640 98.715 53.820 99.575 ;
        RECT 54.365 99.465 55.575 100.555 ;
        RECT 55.750 100.045 57.405 100.335 ;
        RECT 53.565 98.515 53.820 98.715 ;
        RECT 54.365 98.755 54.885 99.295 ;
        RECT 55.055 98.925 55.575 99.465 ;
        RECT 55.750 99.705 57.340 99.875 ;
        RECT 57.575 99.755 57.855 100.555 ;
        RECT 55.750 99.415 56.070 99.705 ;
        RECT 57.170 99.585 57.340 99.705 ;
        RECT 56.265 99.365 56.980 99.535 ;
        RECT 57.170 99.415 57.895 99.585 ;
        RECT 58.065 99.415 58.335 100.385 ;
        RECT 58.505 100.120 63.850 100.555 ;
        RECT 53.100 98.005 53.385 98.465 ;
        RECT 53.565 98.345 53.905 98.515 ;
        RECT 53.565 98.185 53.820 98.345 ;
        RECT 54.365 98.005 55.575 98.755 ;
        RECT 55.750 98.675 56.100 99.245 ;
        RECT 56.270 98.915 56.980 99.365 ;
        RECT 57.725 99.245 57.895 99.415 ;
        RECT 57.150 98.915 57.555 99.245 ;
        RECT 57.725 98.915 57.995 99.245 ;
        RECT 57.725 98.745 57.895 98.915 ;
        RECT 56.285 98.575 57.895 98.745 ;
        RECT 58.165 98.680 58.335 99.415 ;
        RECT 55.755 98.005 56.085 98.505 ;
        RECT 56.285 98.225 56.455 98.575 ;
        RECT 56.655 98.005 56.985 98.405 ;
        RECT 57.155 98.225 57.325 98.575 ;
        RECT 57.495 98.005 57.875 98.405 ;
        RECT 58.065 98.335 58.335 98.680 ;
        RECT 60.090 98.550 60.430 99.380 ;
        RECT 61.910 98.870 62.260 100.120 ;
        RECT 64.025 99.465 66.615 100.555 ;
        RECT 64.025 98.775 65.235 99.295 ;
        RECT 65.405 98.945 66.615 99.465 ;
        RECT 67.245 99.585 67.555 100.385 ;
        RECT 67.725 99.755 68.035 100.555 ;
        RECT 68.205 99.925 68.465 100.385 ;
        RECT 68.635 100.095 68.890 100.555 ;
        RECT 69.065 99.925 69.325 100.385 ;
        RECT 68.205 99.755 69.325 99.925 ;
        RECT 67.245 99.415 68.275 99.585 ;
        RECT 58.505 98.005 63.850 98.550 ;
        RECT 64.025 98.005 66.615 98.775 ;
        RECT 67.245 98.505 67.415 99.415 ;
        RECT 67.585 98.675 67.935 99.245 ;
        RECT 68.105 99.165 68.275 99.415 ;
        RECT 69.065 99.505 69.325 99.755 ;
        RECT 69.495 99.685 69.780 100.555 ;
        RECT 69.065 99.335 69.820 99.505 ;
        RECT 70.005 99.390 70.295 100.555 ;
        RECT 70.985 99.415 71.195 100.555 ;
        RECT 71.365 99.405 71.695 100.385 ;
        RECT 71.865 99.415 72.095 100.555 ;
        RECT 72.305 99.480 72.575 100.385 ;
        RECT 72.745 99.795 73.075 100.555 ;
        RECT 73.255 99.625 73.425 100.385 ;
        RECT 68.105 98.995 69.245 99.165 ;
        RECT 69.415 98.825 69.820 99.335 ;
        RECT 68.170 98.655 69.820 98.825 ;
        RECT 67.245 98.175 67.545 98.505 ;
        RECT 67.715 98.005 67.990 98.485 ;
        RECT 68.170 98.265 68.465 98.655 ;
        RECT 68.635 98.005 68.890 98.485 ;
        RECT 69.065 98.265 69.325 98.655 ;
        RECT 69.495 98.005 69.775 98.485 ;
        RECT 70.005 98.005 70.295 98.730 ;
        RECT 70.985 98.005 71.195 98.825 ;
        RECT 71.365 98.805 71.615 99.405 ;
        RECT 71.785 98.995 72.115 99.245 ;
        RECT 71.365 98.175 71.695 98.805 ;
        RECT 71.865 98.005 72.095 98.825 ;
        RECT 72.305 98.680 72.475 99.480 ;
        RECT 72.760 99.455 73.425 99.625 ;
        RECT 73.685 99.465 77.195 100.555 ;
        RECT 72.760 99.310 72.930 99.455 ;
        RECT 72.645 98.980 72.930 99.310 ;
        RECT 72.760 98.725 72.930 98.980 ;
        RECT 73.165 98.905 73.495 99.275 ;
        RECT 73.685 98.775 75.335 99.295 ;
        RECT 75.505 98.945 77.195 99.465 ;
        RECT 77.570 99.585 77.900 100.385 ;
        RECT 78.070 99.755 78.400 100.555 ;
        RECT 78.700 99.585 79.030 100.385 ;
        RECT 79.675 99.755 79.925 100.555 ;
        RECT 77.570 99.415 80.005 99.585 ;
        RECT 80.195 99.415 80.365 100.555 ;
        RECT 80.535 99.415 80.875 100.385 ;
        RECT 81.250 99.585 81.580 100.385 ;
        RECT 81.750 99.755 82.080 100.555 ;
        RECT 82.380 99.585 82.710 100.385 ;
        RECT 83.355 99.755 83.605 100.555 ;
        RECT 81.250 99.415 83.685 99.585 ;
        RECT 83.875 99.415 84.045 100.555 ;
        RECT 84.215 99.415 84.555 100.385 ;
        RECT 84.930 99.585 85.260 100.385 ;
        RECT 85.430 99.755 85.760 100.555 ;
        RECT 86.060 99.585 86.390 100.385 ;
        RECT 87.035 99.755 87.285 100.555 ;
        RECT 84.930 99.415 87.365 99.585 ;
        RECT 87.555 99.415 87.725 100.555 ;
        RECT 87.895 99.415 88.235 100.385 ;
        RECT 88.405 99.465 91.915 100.555 ;
        RECT 92.085 99.465 93.295 100.555 ;
        RECT 77.365 98.995 77.715 99.245 ;
        RECT 77.900 98.785 78.070 99.415 ;
        RECT 78.240 98.995 78.570 99.195 ;
        RECT 78.740 98.995 79.070 99.195 ;
        RECT 79.240 98.995 79.660 99.195 ;
        RECT 79.835 99.165 80.005 99.415 ;
        RECT 79.835 98.995 80.530 99.165 ;
        RECT 72.305 98.175 72.565 98.680 ;
        RECT 72.760 98.555 73.425 98.725 ;
        RECT 72.745 98.005 73.075 98.385 ;
        RECT 73.255 98.175 73.425 98.555 ;
        RECT 73.685 98.005 77.195 98.775 ;
        RECT 77.570 98.175 78.070 98.785 ;
        RECT 78.700 98.655 79.925 98.825 ;
        RECT 80.700 98.805 80.875 99.415 ;
        RECT 81.045 98.995 81.395 99.245 ;
        RECT 78.700 98.175 79.030 98.655 ;
        RECT 79.200 98.005 79.425 98.465 ;
        RECT 79.595 98.175 79.925 98.655 ;
        RECT 80.115 98.005 80.365 98.805 ;
        RECT 80.535 98.175 80.875 98.805 ;
        RECT 81.580 98.785 81.750 99.415 ;
        RECT 81.920 98.995 82.250 99.195 ;
        RECT 82.420 98.995 82.750 99.195 ;
        RECT 82.920 98.995 83.340 99.195 ;
        RECT 83.515 99.165 83.685 99.415 ;
        RECT 83.515 98.995 84.210 99.165 ;
        RECT 81.250 98.175 81.750 98.785 ;
        RECT 82.380 98.655 83.605 98.825 ;
        RECT 84.380 98.805 84.555 99.415 ;
        RECT 84.725 98.995 85.075 99.245 ;
        RECT 82.380 98.175 82.710 98.655 ;
        RECT 82.880 98.005 83.105 98.465 ;
        RECT 83.275 98.175 83.605 98.655 ;
        RECT 83.795 98.005 84.045 98.805 ;
        RECT 84.215 98.175 84.555 98.805 ;
        RECT 85.260 98.785 85.430 99.415 ;
        RECT 85.600 98.995 85.930 99.195 ;
        RECT 86.100 98.995 86.430 99.195 ;
        RECT 86.600 98.995 87.020 99.195 ;
        RECT 87.195 99.165 87.365 99.415 ;
        RECT 87.195 98.995 87.890 99.165 ;
        RECT 84.930 98.175 85.430 98.785 ;
        RECT 86.060 98.655 87.285 98.825 ;
        RECT 88.060 98.805 88.235 99.415 ;
        RECT 86.060 98.175 86.390 98.655 ;
        RECT 86.560 98.005 86.785 98.465 ;
        RECT 86.955 98.175 87.285 98.655 ;
        RECT 87.475 98.005 87.725 98.805 ;
        RECT 87.895 98.175 88.235 98.805 ;
        RECT 88.405 98.775 90.055 99.295 ;
        RECT 90.225 98.945 91.915 99.465 ;
        RECT 88.405 98.005 91.915 98.775 ;
        RECT 92.085 98.755 92.605 99.295 ;
        RECT 92.775 98.925 93.295 99.465 ;
        RECT 93.465 99.835 93.925 100.385 ;
        RECT 94.115 99.835 94.445 100.555 ;
        RECT 92.085 98.005 93.295 98.755 ;
        RECT 93.465 98.465 93.715 99.835 ;
        RECT 94.645 99.665 94.945 100.215 ;
        RECT 95.115 99.885 95.395 100.555 ;
        RECT 94.005 99.495 94.945 99.665 ;
        RECT 94.005 99.245 94.175 99.495 ;
        RECT 95.315 99.245 95.580 99.605 ;
        RECT 95.765 99.390 96.055 100.555 ;
        RECT 97.145 99.480 97.415 100.385 ;
        RECT 97.585 99.795 97.915 100.555 ;
        RECT 98.095 99.625 98.265 100.385 ;
        RECT 93.885 98.915 94.175 99.245 ;
        RECT 94.345 98.995 94.685 99.245 ;
        RECT 94.905 98.995 95.580 99.245 ;
        RECT 94.005 98.825 94.175 98.915 ;
        RECT 94.005 98.635 95.395 98.825 ;
        RECT 93.465 98.175 94.025 98.465 ;
        RECT 94.195 98.005 94.445 98.465 ;
        RECT 95.065 98.275 95.395 98.635 ;
        RECT 95.765 98.005 96.055 98.730 ;
        RECT 97.145 98.680 97.315 99.480 ;
        RECT 97.600 99.455 98.265 99.625 ;
        RECT 98.525 99.465 100.195 100.555 ;
        RECT 97.600 99.310 97.770 99.455 ;
        RECT 97.485 98.980 97.770 99.310 ;
        RECT 97.600 98.725 97.770 98.980 ;
        RECT 98.005 98.905 98.335 99.275 ;
        RECT 98.525 98.775 99.275 99.295 ;
        RECT 99.445 98.945 100.195 99.465 ;
        RECT 100.885 99.415 101.095 100.555 ;
        RECT 101.265 99.405 101.595 100.385 ;
        RECT 101.765 99.415 101.995 100.555 ;
        RECT 102.205 99.465 104.795 100.555 ;
        RECT 105.515 99.885 105.685 100.385 ;
        RECT 105.855 100.055 106.185 100.555 ;
        RECT 105.515 99.715 106.180 99.885 ;
        RECT 97.145 98.175 97.405 98.680 ;
        RECT 97.600 98.555 98.265 98.725 ;
        RECT 97.585 98.005 97.915 98.385 ;
        RECT 98.095 98.175 98.265 98.555 ;
        RECT 98.525 98.005 100.195 98.775 ;
        RECT 100.885 98.005 101.095 98.825 ;
        RECT 101.265 98.805 101.515 99.405 ;
        RECT 101.685 98.995 102.015 99.245 ;
        RECT 101.265 98.175 101.595 98.805 ;
        RECT 101.765 98.005 101.995 98.825 ;
        RECT 102.205 98.775 103.415 99.295 ;
        RECT 103.585 98.945 104.795 99.465 ;
        RECT 105.430 98.895 105.780 99.545 ;
        RECT 102.205 98.005 104.795 98.775 ;
        RECT 105.950 98.725 106.180 99.715 ;
        RECT 105.515 98.555 106.180 98.725 ;
        RECT 105.515 98.265 105.685 98.555 ;
        RECT 105.855 98.005 106.185 98.385 ;
        RECT 106.355 98.265 106.580 100.385 ;
        RECT 106.795 100.055 107.125 100.555 ;
        RECT 107.295 99.885 107.465 100.385 ;
        RECT 107.700 100.170 108.530 100.340 ;
        RECT 108.770 100.175 109.150 100.555 ;
        RECT 106.770 99.715 107.465 99.885 ;
        RECT 106.770 98.745 106.940 99.715 ;
        RECT 107.110 98.925 107.520 99.545 ;
        RECT 107.690 99.495 108.190 99.875 ;
        RECT 106.770 98.555 107.465 98.745 ;
        RECT 107.690 98.625 107.910 99.495 ;
        RECT 108.360 99.325 108.530 100.170 ;
        RECT 109.330 100.005 109.500 100.295 ;
        RECT 109.670 100.175 110.000 100.555 ;
        RECT 110.470 100.085 111.100 100.335 ;
        RECT 111.280 100.175 111.700 100.555 ;
        RECT 110.930 100.005 111.100 100.085 ;
        RECT 111.900 100.005 112.140 100.295 ;
        RECT 108.700 99.755 110.070 100.005 ;
        RECT 108.700 99.495 108.950 99.755 ;
        RECT 109.460 99.325 109.710 99.485 ;
        RECT 108.360 99.155 109.710 99.325 ;
        RECT 108.360 99.115 108.780 99.155 ;
        RECT 108.090 98.565 108.440 98.935 ;
        RECT 106.795 98.005 107.125 98.385 ;
        RECT 107.295 98.225 107.465 98.555 ;
        RECT 108.610 98.385 108.780 99.115 ;
        RECT 109.880 98.985 110.070 99.755 ;
        RECT 108.950 98.655 109.360 98.985 ;
        RECT 109.650 98.645 110.070 98.985 ;
        RECT 110.240 99.575 110.760 99.885 ;
        RECT 110.930 99.835 112.140 100.005 ;
        RECT 112.370 99.865 112.700 100.555 ;
        RECT 110.240 98.815 110.410 99.575 ;
        RECT 110.580 98.985 110.760 99.395 ;
        RECT 110.930 99.325 111.100 99.835 ;
        RECT 112.870 99.685 113.040 100.295 ;
        RECT 113.310 99.835 113.640 100.345 ;
        RECT 112.870 99.665 113.190 99.685 ;
        RECT 111.270 99.495 113.190 99.665 ;
        RECT 110.930 99.155 112.830 99.325 ;
        RECT 111.160 98.815 111.490 98.935 ;
        RECT 110.240 98.645 111.490 98.815 ;
        RECT 107.765 98.185 108.780 98.385 ;
        RECT 108.950 98.005 109.360 98.445 ;
        RECT 109.650 98.215 109.900 98.645 ;
        RECT 110.100 98.005 110.420 98.465 ;
        RECT 111.660 98.395 111.830 99.155 ;
        RECT 112.500 99.095 112.830 99.155 ;
        RECT 112.020 98.925 112.350 98.985 ;
        RECT 112.020 98.655 112.680 98.925 ;
        RECT 113.000 98.600 113.190 99.495 ;
        RECT 110.980 98.225 111.830 98.395 ;
        RECT 112.030 98.005 112.690 98.485 ;
        RECT 112.870 98.270 113.190 98.600 ;
        RECT 113.390 99.245 113.640 99.835 ;
        RECT 113.820 99.755 114.105 100.555 ;
        RECT 114.285 99.575 114.540 100.245 ;
        RECT 113.390 98.915 114.190 99.245 ;
        RECT 113.390 98.265 113.640 98.915 ;
        RECT 114.360 98.715 114.540 99.575 ;
        RECT 115.085 99.795 115.600 100.205 ;
        RECT 115.835 99.795 116.005 100.555 ;
        RECT 116.175 100.215 118.205 100.385 ;
        RECT 115.085 98.985 115.425 99.795 ;
        RECT 116.175 99.550 116.345 100.215 ;
        RECT 116.740 99.875 117.865 100.045 ;
        RECT 115.595 99.360 116.345 99.550 ;
        RECT 116.515 99.535 117.525 99.705 ;
        RECT 115.085 98.815 116.315 98.985 ;
        RECT 114.285 98.515 114.540 98.715 ;
        RECT 113.820 98.005 114.105 98.465 ;
        RECT 114.285 98.345 114.625 98.515 ;
        RECT 114.285 98.185 114.540 98.345 ;
        RECT 115.360 98.210 115.605 98.815 ;
        RECT 115.825 98.005 116.335 98.540 ;
        RECT 116.515 98.175 116.705 99.535 ;
        RECT 116.875 98.515 117.150 99.335 ;
        RECT 117.355 98.735 117.525 99.535 ;
        RECT 117.695 98.745 117.865 99.875 ;
        RECT 118.035 99.245 118.205 100.215 ;
        RECT 118.375 99.415 118.545 100.555 ;
        RECT 118.715 99.415 119.050 100.385 ;
        RECT 118.035 98.915 118.230 99.245 ;
        RECT 118.455 98.915 118.710 99.245 ;
        RECT 118.455 98.745 118.625 98.915 ;
        RECT 118.880 98.745 119.050 99.415 ;
        RECT 117.695 98.575 118.625 98.745 ;
        RECT 117.695 98.540 117.870 98.575 ;
        RECT 116.875 98.345 117.155 98.515 ;
        RECT 116.875 98.175 117.150 98.345 ;
        RECT 117.340 98.175 117.870 98.540 ;
        RECT 118.295 98.005 118.625 98.405 ;
        RECT 118.795 98.175 119.050 98.745 ;
        RECT 119.225 99.480 119.495 100.385 ;
        RECT 119.665 99.795 119.995 100.555 ;
        RECT 120.175 99.625 120.345 100.385 ;
        RECT 119.225 98.680 119.395 99.480 ;
        RECT 119.680 99.455 120.345 99.625 ;
        RECT 119.680 99.310 119.850 99.455 ;
        RECT 121.525 99.390 121.815 100.555 ;
        RECT 122.025 99.415 122.255 100.555 ;
        RECT 122.425 99.405 122.755 100.385 ;
        RECT 122.925 99.415 123.135 100.555 ;
        RECT 124.285 99.465 125.495 100.555 ;
        RECT 119.565 98.980 119.850 99.310 ;
        RECT 119.680 98.725 119.850 98.980 ;
        RECT 120.085 98.905 120.415 99.275 ;
        RECT 122.005 98.995 122.335 99.245 ;
        RECT 119.225 98.175 119.485 98.680 ;
        RECT 119.680 98.555 120.345 98.725 ;
        RECT 119.665 98.005 119.995 98.385 ;
        RECT 120.175 98.175 120.345 98.555 ;
        RECT 121.525 98.005 121.815 98.730 ;
        RECT 122.025 98.005 122.255 98.825 ;
        RECT 122.505 98.805 122.755 99.405 ;
        RECT 124.285 98.925 124.805 99.465 ;
        RECT 122.425 98.175 122.755 98.805 ;
        RECT 122.925 98.005 123.135 98.825 ;
        RECT 124.975 98.755 125.495 99.295 ;
        RECT 124.285 98.005 125.495 98.755 ;
        RECT 5.520 97.835 125.580 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 6.985 97.290 12.330 97.835 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 8.570 96.460 8.910 97.290 ;
        RECT 13.425 97.160 13.685 97.665 ;
        RECT 13.865 97.455 14.195 97.835 ;
        RECT 14.375 97.285 14.545 97.665 ;
        RECT 14.805 97.290 20.150 97.835 ;
        RECT 20.325 97.290 25.670 97.835 ;
        RECT 25.845 97.290 31.190 97.835 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 10.390 95.720 10.740 96.970 ;
        RECT 13.425 96.360 13.595 97.160 ;
        RECT 13.880 97.115 14.545 97.285 ;
        RECT 13.880 96.860 14.050 97.115 ;
        RECT 13.765 96.530 14.050 96.860 ;
        RECT 14.285 96.565 14.615 96.935 ;
        RECT 13.880 96.385 14.050 96.530 ;
        RECT 16.390 96.460 16.730 97.290 ;
        RECT 6.985 95.285 12.330 95.720 ;
        RECT 13.425 95.455 13.695 96.360 ;
        RECT 13.880 96.215 14.545 96.385 ;
        RECT 13.865 95.285 14.195 96.045 ;
        RECT 14.375 95.455 14.545 96.215 ;
        RECT 18.210 95.720 18.560 96.970 ;
        RECT 21.910 96.460 22.250 97.290 ;
        RECT 23.730 95.720 24.080 96.970 ;
        RECT 27.430 96.460 27.770 97.290 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 32.805 97.015 33.015 97.835 ;
        RECT 33.185 97.035 33.515 97.665 ;
        RECT 29.250 95.720 29.600 96.970 ;
        RECT 14.805 95.285 20.150 95.720 ;
        RECT 20.325 95.285 25.670 95.720 ;
        RECT 25.845 95.285 31.190 95.720 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 33.185 96.435 33.435 97.035 ;
        RECT 33.685 97.015 33.915 97.835 ;
        RECT 34.125 97.065 36.715 97.835 ;
        RECT 37.435 97.285 37.605 97.575 ;
        RECT 37.775 97.455 38.105 97.835 ;
        RECT 37.435 97.115 38.100 97.285 ;
        RECT 33.605 96.595 33.935 96.845 ;
        RECT 34.125 96.545 35.335 97.065 ;
        RECT 32.805 95.285 33.015 96.425 ;
        RECT 33.185 95.455 33.515 96.435 ;
        RECT 33.685 95.285 33.915 96.425 ;
        RECT 35.505 96.375 36.715 96.895 ;
        RECT 34.125 95.285 36.715 96.375 ;
        RECT 37.350 96.295 37.700 96.945 ;
        RECT 37.870 96.125 38.100 97.115 ;
        RECT 37.435 95.955 38.100 96.125 ;
        RECT 37.435 95.455 37.605 95.955 ;
        RECT 37.775 95.285 38.105 95.785 ;
        RECT 38.275 95.455 38.500 97.575 ;
        RECT 38.715 97.455 39.045 97.835 ;
        RECT 39.215 97.285 39.385 97.615 ;
        RECT 39.685 97.455 40.700 97.655 ;
        RECT 38.690 97.095 39.385 97.285 ;
        RECT 38.690 96.125 38.860 97.095 ;
        RECT 39.030 96.295 39.440 96.915 ;
        RECT 39.610 96.345 39.830 97.215 ;
        RECT 40.010 96.905 40.360 97.275 ;
        RECT 40.530 96.725 40.700 97.455 ;
        RECT 40.870 97.395 41.280 97.835 ;
        RECT 41.570 97.195 41.820 97.625 ;
        RECT 42.020 97.375 42.340 97.835 ;
        RECT 42.900 97.445 43.750 97.615 ;
        RECT 40.870 96.855 41.280 97.185 ;
        RECT 41.570 96.855 41.990 97.195 ;
        RECT 40.280 96.685 40.700 96.725 ;
        RECT 40.280 96.515 41.630 96.685 ;
        RECT 38.690 95.955 39.385 96.125 ;
        RECT 39.610 95.965 40.110 96.345 ;
        RECT 38.715 95.285 39.045 95.785 ;
        RECT 39.215 95.455 39.385 95.955 ;
        RECT 40.280 95.670 40.450 96.515 ;
        RECT 41.380 96.355 41.630 96.515 ;
        RECT 40.620 96.085 40.870 96.345 ;
        RECT 41.800 96.085 41.990 96.855 ;
        RECT 40.620 95.835 41.990 96.085 ;
        RECT 42.160 97.025 43.410 97.195 ;
        RECT 42.160 96.265 42.330 97.025 ;
        RECT 43.080 96.905 43.410 97.025 ;
        RECT 42.500 96.445 42.680 96.855 ;
        RECT 43.580 96.685 43.750 97.445 ;
        RECT 43.950 97.355 44.610 97.835 ;
        RECT 44.790 97.240 45.110 97.570 ;
        RECT 43.940 96.915 44.600 97.185 ;
        RECT 43.940 96.855 44.270 96.915 ;
        RECT 44.420 96.685 44.750 96.745 ;
        RECT 42.850 96.515 44.750 96.685 ;
        RECT 42.160 95.955 42.680 96.265 ;
        RECT 42.850 96.005 43.020 96.515 ;
        RECT 44.920 96.345 45.110 97.240 ;
        RECT 43.190 96.175 45.110 96.345 ;
        RECT 44.790 96.155 45.110 96.175 ;
        RECT 45.310 96.925 45.560 97.575 ;
        RECT 45.740 97.375 46.025 97.835 ;
        RECT 46.205 97.125 46.460 97.655 ;
        RECT 45.310 96.595 46.110 96.925 ;
        RECT 42.850 95.835 44.060 96.005 ;
        RECT 39.620 95.500 40.450 95.670 ;
        RECT 40.690 95.285 41.070 95.665 ;
        RECT 41.250 95.545 41.420 95.835 ;
        RECT 42.850 95.755 43.020 95.835 ;
        RECT 41.590 95.285 41.920 95.665 ;
        RECT 42.390 95.505 43.020 95.755 ;
        RECT 43.200 95.285 43.620 95.665 ;
        RECT 43.820 95.545 44.060 95.835 ;
        RECT 44.290 95.285 44.620 95.975 ;
        RECT 44.790 95.545 44.960 96.155 ;
        RECT 45.310 96.005 45.560 96.595 ;
        RECT 46.280 96.265 46.460 97.125 ;
        RECT 45.230 95.495 45.560 96.005 ;
        RECT 45.740 95.285 46.025 96.085 ;
        RECT 46.205 95.795 46.460 96.265 ;
        RECT 47.005 97.160 47.265 97.665 ;
        RECT 47.445 97.455 47.775 97.835 ;
        RECT 47.955 97.285 48.125 97.665 ;
        RECT 47.005 96.360 47.175 97.160 ;
        RECT 47.460 97.115 48.125 97.285 ;
        RECT 47.460 96.860 47.630 97.115 ;
        RECT 48.390 97.095 48.645 97.665 ;
        RECT 48.815 97.435 49.145 97.835 ;
        RECT 49.570 97.300 50.100 97.665 ;
        RECT 49.570 97.265 49.745 97.300 ;
        RECT 48.815 97.095 49.745 97.265 ;
        RECT 47.345 96.530 47.630 96.860 ;
        RECT 47.865 96.565 48.195 96.935 ;
        RECT 47.460 96.385 47.630 96.530 ;
        RECT 48.390 96.425 48.560 97.095 ;
        RECT 48.815 96.925 48.985 97.095 ;
        RECT 48.730 96.595 48.985 96.925 ;
        RECT 49.210 96.595 49.405 96.925 ;
        RECT 46.205 95.625 46.545 95.795 ;
        RECT 46.205 95.595 46.460 95.625 ;
        RECT 47.005 95.455 47.275 96.360 ;
        RECT 47.460 96.215 48.125 96.385 ;
        RECT 47.445 95.285 47.775 96.045 ;
        RECT 47.955 95.455 48.125 96.215 ;
        RECT 48.390 95.455 48.725 96.425 ;
        RECT 48.895 95.285 49.065 96.425 ;
        RECT 49.235 95.625 49.405 96.595 ;
        RECT 49.575 95.965 49.745 97.095 ;
        RECT 49.915 96.305 50.085 97.105 ;
        RECT 50.290 96.815 50.565 97.665 ;
        RECT 50.285 96.645 50.565 96.815 ;
        RECT 50.290 96.505 50.565 96.645 ;
        RECT 50.735 96.305 50.925 97.665 ;
        RECT 51.105 97.300 51.615 97.835 ;
        RECT 51.835 97.025 52.080 97.630 ;
        RECT 53.445 97.035 53.785 97.665 ;
        RECT 53.955 97.035 54.205 97.835 ;
        RECT 54.395 97.185 54.725 97.665 ;
        RECT 54.895 97.375 55.120 97.835 ;
        RECT 55.290 97.185 55.620 97.665 ;
        RECT 51.125 96.855 52.355 97.025 ;
        RECT 49.915 96.135 50.925 96.305 ;
        RECT 51.095 96.290 51.845 96.480 ;
        RECT 49.575 95.795 50.700 95.965 ;
        RECT 51.095 95.625 51.265 96.290 ;
        RECT 52.015 96.045 52.355 96.855 ;
        RECT 49.235 95.455 51.265 95.625 ;
        RECT 51.435 95.285 51.605 96.045 ;
        RECT 51.840 95.635 52.355 96.045 ;
        RECT 53.445 96.425 53.620 97.035 ;
        RECT 54.395 97.015 55.620 97.185 ;
        RECT 56.250 97.055 56.750 97.665 ;
        RECT 57.125 97.110 57.415 97.835 ;
        RECT 57.790 97.055 58.290 97.665 ;
        RECT 53.790 96.675 54.485 96.845 ;
        RECT 54.315 96.425 54.485 96.675 ;
        RECT 54.660 96.645 55.080 96.845 ;
        RECT 55.250 96.645 55.580 96.845 ;
        RECT 55.750 96.645 56.080 96.845 ;
        RECT 56.250 96.425 56.420 97.055 ;
        RECT 56.605 96.595 56.955 96.845 ;
        RECT 57.585 96.595 57.935 96.845 ;
        RECT 53.445 95.455 53.785 96.425 ;
        RECT 53.955 95.285 54.125 96.425 ;
        RECT 54.315 96.255 56.750 96.425 ;
        RECT 54.395 95.285 54.645 96.085 ;
        RECT 55.290 95.455 55.620 96.255 ;
        RECT 55.920 95.285 56.250 96.085 ;
        RECT 56.420 95.455 56.750 96.255 ;
        RECT 57.125 95.285 57.415 96.450 ;
        RECT 58.120 96.425 58.290 97.055 ;
        RECT 58.920 97.185 59.250 97.665 ;
        RECT 59.420 97.375 59.645 97.835 ;
        RECT 59.815 97.185 60.145 97.665 ;
        RECT 58.920 97.015 60.145 97.185 ;
        RECT 60.335 97.035 60.585 97.835 ;
        RECT 60.755 97.035 61.095 97.665 ;
        RECT 58.460 96.645 58.790 96.845 ;
        RECT 58.960 96.645 59.290 96.845 ;
        RECT 59.460 96.645 59.880 96.845 ;
        RECT 60.055 96.675 60.750 96.845 ;
        RECT 60.055 96.425 60.225 96.675 ;
        RECT 60.920 96.425 61.095 97.035 ;
        RECT 61.265 97.065 62.935 97.835 ;
        RECT 63.305 97.205 63.635 97.565 ;
        RECT 64.255 97.375 64.505 97.835 ;
        RECT 64.675 97.375 65.235 97.665 ;
        RECT 61.265 96.545 62.015 97.065 ;
        RECT 63.305 97.015 64.695 97.205 ;
        RECT 64.525 96.925 64.695 97.015 ;
        RECT 57.790 96.255 60.225 96.425 ;
        RECT 57.790 95.455 58.120 96.255 ;
        RECT 58.290 95.285 58.620 96.085 ;
        RECT 58.920 95.455 59.250 96.255 ;
        RECT 59.895 95.285 60.145 96.085 ;
        RECT 60.415 95.285 60.585 96.425 ;
        RECT 60.755 95.455 61.095 96.425 ;
        RECT 62.185 96.375 62.935 96.895 ;
        RECT 61.265 95.285 62.935 96.375 ;
        RECT 63.120 96.595 63.795 96.845 ;
        RECT 64.015 96.595 64.355 96.845 ;
        RECT 64.525 96.595 64.815 96.925 ;
        RECT 63.120 96.235 63.385 96.595 ;
        RECT 64.525 96.345 64.695 96.595 ;
        RECT 63.755 96.175 64.695 96.345 ;
        RECT 63.305 95.285 63.585 95.955 ;
        RECT 63.755 95.625 64.055 96.175 ;
        RECT 64.985 96.005 65.235 97.375 ;
        RECT 65.955 97.285 66.125 97.575 ;
        RECT 66.295 97.455 66.625 97.835 ;
        RECT 65.955 97.115 66.620 97.285 ;
        RECT 65.870 96.295 66.220 96.945 ;
        RECT 66.390 96.125 66.620 97.115 ;
        RECT 64.255 95.285 64.585 96.005 ;
        RECT 64.775 95.455 65.235 96.005 ;
        RECT 65.955 95.955 66.620 96.125 ;
        RECT 65.955 95.455 66.125 95.955 ;
        RECT 66.295 95.285 66.625 95.785 ;
        RECT 66.795 95.455 67.020 97.575 ;
        RECT 67.235 97.455 67.565 97.835 ;
        RECT 67.735 97.285 67.905 97.615 ;
        RECT 68.205 97.455 69.220 97.655 ;
        RECT 67.210 97.095 67.905 97.285 ;
        RECT 67.210 96.125 67.380 97.095 ;
        RECT 67.550 96.295 67.960 96.915 ;
        RECT 68.130 96.345 68.350 97.215 ;
        RECT 68.530 96.905 68.880 97.275 ;
        RECT 69.050 96.725 69.220 97.455 ;
        RECT 69.390 97.395 69.800 97.835 ;
        RECT 70.090 97.195 70.340 97.625 ;
        RECT 70.540 97.375 70.860 97.835 ;
        RECT 71.420 97.445 72.270 97.615 ;
        RECT 69.390 96.855 69.800 97.185 ;
        RECT 70.090 96.855 70.510 97.195 ;
        RECT 68.800 96.685 69.220 96.725 ;
        RECT 68.800 96.515 70.150 96.685 ;
        RECT 67.210 95.955 67.905 96.125 ;
        RECT 68.130 95.965 68.630 96.345 ;
        RECT 67.235 95.285 67.565 95.785 ;
        RECT 67.735 95.455 67.905 95.955 ;
        RECT 68.800 95.670 68.970 96.515 ;
        RECT 69.900 96.355 70.150 96.515 ;
        RECT 69.140 96.085 69.390 96.345 ;
        RECT 70.320 96.085 70.510 96.855 ;
        RECT 69.140 95.835 70.510 96.085 ;
        RECT 70.680 97.025 71.930 97.195 ;
        RECT 70.680 96.265 70.850 97.025 ;
        RECT 71.600 96.905 71.930 97.025 ;
        RECT 71.020 96.445 71.200 96.855 ;
        RECT 72.100 96.685 72.270 97.445 ;
        RECT 72.470 97.355 73.130 97.835 ;
        RECT 73.310 97.240 73.630 97.570 ;
        RECT 72.460 96.915 73.120 97.185 ;
        RECT 72.460 96.855 72.790 96.915 ;
        RECT 72.940 96.685 73.270 96.745 ;
        RECT 71.370 96.515 73.270 96.685 ;
        RECT 70.680 95.955 71.200 96.265 ;
        RECT 71.370 96.005 71.540 96.515 ;
        RECT 73.440 96.345 73.630 97.240 ;
        RECT 71.710 96.175 73.630 96.345 ;
        RECT 73.310 96.155 73.630 96.175 ;
        RECT 73.830 96.925 74.080 97.575 ;
        RECT 74.260 97.375 74.545 97.835 ;
        RECT 74.725 97.155 74.980 97.655 ;
        RECT 74.725 97.125 75.065 97.155 ;
        RECT 74.800 96.985 75.065 97.125 ;
        RECT 75.730 97.055 76.230 97.665 ;
        RECT 73.830 96.595 74.630 96.925 ;
        RECT 71.370 95.835 72.580 96.005 ;
        RECT 68.140 95.500 68.970 95.670 ;
        RECT 69.210 95.285 69.590 95.665 ;
        RECT 69.770 95.545 69.940 95.835 ;
        RECT 71.370 95.755 71.540 95.835 ;
        RECT 70.110 95.285 70.440 95.665 ;
        RECT 70.910 95.505 71.540 95.755 ;
        RECT 71.720 95.285 72.140 95.665 ;
        RECT 72.340 95.545 72.580 95.835 ;
        RECT 72.810 95.285 73.140 95.975 ;
        RECT 73.310 95.545 73.480 96.155 ;
        RECT 73.830 96.005 74.080 96.595 ;
        RECT 74.800 96.265 74.980 96.985 ;
        RECT 75.525 96.595 75.875 96.845 ;
        RECT 76.060 96.425 76.230 97.055 ;
        RECT 76.860 97.185 77.190 97.665 ;
        RECT 77.360 97.375 77.585 97.835 ;
        RECT 77.755 97.185 78.085 97.665 ;
        RECT 76.860 97.015 78.085 97.185 ;
        RECT 78.275 97.035 78.525 97.835 ;
        RECT 78.695 97.035 79.035 97.665 ;
        RECT 76.400 96.645 76.730 96.845 ;
        RECT 76.900 96.645 77.230 96.845 ;
        RECT 77.400 96.645 77.820 96.845 ;
        RECT 77.995 96.675 78.690 96.845 ;
        RECT 77.995 96.425 78.165 96.675 ;
        RECT 78.860 96.425 79.035 97.035 ;
        RECT 79.205 97.065 82.715 97.835 ;
        RECT 82.885 97.110 83.175 97.835 ;
        RECT 83.345 97.160 83.615 97.505 ;
        RECT 83.805 97.435 84.185 97.835 ;
        RECT 84.355 97.265 84.525 97.615 ;
        RECT 84.695 97.435 85.025 97.835 ;
        RECT 85.225 97.265 85.395 97.615 ;
        RECT 85.595 97.335 85.925 97.835 ;
        RECT 86.105 97.290 91.450 97.835 ;
        RECT 79.205 96.545 80.855 97.065 ;
        RECT 73.750 95.495 74.080 96.005 ;
        RECT 74.260 95.285 74.545 96.085 ;
        RECT 74.725 95.595 74.980 96.265 ;
        RECT 75.730 96.255 78.165 96.425 ;
        RECT 75.730 95.455 76.060 96.255 ;
        RECT 76.230 95.285 76.560 96.085 ;
        RECT 76.860 95.455 77.190 96.255 ;
        RECT 77.835 95.285 78.085 96.085 ;
        RECT 78.355 95.285 78.525 96.425 ;
        RECT 78.695 95.455 79.035 96.425 ;
        RECT 81.025 96.375 82.715 96.895 ;
        RECT 79.205 95.285 82.715 96.375 ;
        RECT 82.885 95.285 83.175 96.450 ;
        RECT 83.345 96.425 83.515 97.160 ;
        RECT 83.785 97.095 85.395 97.265 ;
        RECT 83.785 96.925 83.955 97.095 ;
        RECT 83.685 96.595 83.955 96.925 ;
        RECT 84.125 96.595 84.530 96.925 ;
        RECT 83.785 96.425 83.955 96.595 ;
        RECT 83.345 95.455 83.615 96.425 ;
        RECT 83.785 96.255 84.510 96.425 ;
        RECT 84.700 96.305 85.410 96.925 ;
        RECT 85.580 96.595 85.930 97.165 ;
        RECT 87.690 96.460 88.030 97.290 ;
        RECT 91.625 97.085 92.835 97.835 ;
        RECT 93.005 97.160 93.275 97.505 ;
        RECT 93.465 97.435 93.845 97.835 ;
        RECT 94.015 97.265 94.185 97.615 ;
        RECT 94.355 97.435 94.685 97.835 ;
        RECT 94.885 97.265 95.055 97.615 ;
        RECT 95.255 97.335 95.585 97.835 ;
        RECT 84.340 96.135 84.510 96.255 ;
        RECT 85.610 96.135 85.930 96.425 ;
        RECT 83.825 95.285 84.105 96.085 ;
        RECT 84.340 95.965 85.930 96.135 ;
        RECT 84.275 95.505 85.930 95.795 ;
        RECT 89.510 95.720 89.860 96.970 ;
        RECT 91.625 96.545 92.145 97.085 ;
        RECT 92.315 96.375 92.835 96.915 ;
        RECT 86.105 95.285 91.450 95.720 ;
        RECT 91.625 95.285 92.835 96.375 ;
        RECT 93.005 96.425 93.175 97.160 ;
        RECT 93.445 97.095 95.055 97.265 ;
        RECT 95.855 97.285 96.025 97.575 ;
        RECT 96.195 97.455 96.525 97.835 ;
        RECT 93.445 96.925 93.615 97.095 ;
        RECT 93.345 96.595 93.615 96.925 ;
        RECT 93.785 96.595 94.190 96.925 ;
        RECT 93.445 96.425 93.615 96.595 ;
        RECT 93.005 95.455 93.275 96.425 ;
        RECT 93.445 96.255 94.170 96.425 ;
        RECT 94.360 96.305 95.070 96.925 ;
        RECT 95.240 96.595 95.590 97.165 ;
        RECT 95.855 97.115 96.520 97.285 ;
        RECT 94.000 96.135 94.170 96.255 ;
        RECT 95.270 96.135 95.590 96.425 ;
        RECT 95.770 96.295 96.120 96.945 ;
        RECT 93.485 95.285 93.765 96.085 ;
        RECT 94.000 95.965 95.590 96.135 ;
        RECT 96.290 96.125 96.520 97.115 ;
        RECT 95.855 95.955 96.520 96.125 ;
        RECT 93.935 95.505 95.590 95.795 ;
        RECT 95.855 95.455 96.025 95.955 ;
        RECT 96.195 95.285 96.525 95.785 ;
        RECT 96.695 95.455 96.920 97.575 ;
        RECT 97.135 97.455 97.465 97.835 ;
        RECT 97.635 97.285 97.805 97.615 ;
        RECT 98.105 97.455 99.120 97.655 ;
        RECT 97.110 97.095 97.805 97.285 ;
        RECT 97.110 96.125 97.280 97.095 ;
        RECT 97.450 96.295 97.860 96.915 ;
        RECT 98.030 96.345 98.250 97.215 ;
        RECT 98.430 96.905 98.780 97.275 ;
        RECT 98.950 96.725 99.120 97.455 ;
        RECT 99.290 97.395 99.700 97.835 ;
        RECT 99.990 97.195 100.240 97.625 ;
        RECT 100.440 97.375 100.760 97.835 ;
        RECT 101.320 97.445 102.170 97.615 ;
        RECT 99.290 96.855 99.700 97.185 ;
        RECT 99.990 96.855 100.410 97.195 ;
        RECT 98.700 96.685 99.120 96.725 ;
        RECT 98.700 96.515 100.050 96.685 ;
        RECT 97.110 95.955 97.805 96.125 ;
        RECT 98.030 95.965 98.530 96.345 ;
        RECT 97.135 95.285 97.465 95.785 ;
        RECT 97.635 95.455 97.805 95.955 ;
        RECT 98.700 95.670 98.870 96.515 ;
        RECT 99.800 96.355 100.050 96.515 ;
        RECT 99.040 96.085 99.290 96.345 ;
        RECT 100.220 96.085 100.410 96.855 ;
        RECT 99.040 95.835 100.410 96.085 ;
        RECT 100.580 97.025 101.830 97.195 ;
        RECT 100.580 96.265 100.750 97.025 ;
        RECT 101.500 96.905 101.830 97.025 ;
        RECT 100.920 96.445 101.100 96.855 ;
        RECT 102.000 96.685 102.170 97.445 ;
        RECT 102.370 97.355 103.030 97.835 ;
        RECT 103.210 97.240 103.530 97.570 ;
        RECT 102.360 96.915 103.020 97.185 ;
        RECT 102.360 96.855 102.690 96.915 ;
        RECT 102.840 96.685 103.170 96.745 ;
        RECT 101.270 96.515 103.170 96.685 ;
        RECT 100.580 95.955 101.100 96.265 ;
        RECT 101.270 96.005 101.440 96.515 ;
        RECT 103.340 96.345 103.530 97.240 ;
        RECT 101.610 96.175 103.530 96.345 ;
        RECT 103.210 96.155 103.530 96.175 ;
        RECT 103.730 96.925 103.980 97.575 ;
        RECT 104.160 97.375 104.445 97.835 ;
        RECT 104.625 97.125 104.880 97.655 ;
        RECT 103.730 96.595 104.530 96.925 ;
        RECT 101.270 95.835 102.480 96.005 ;
        RECT 98.040 95.500 98.870 95.670 ;
        RECT 99.110 95.285 99.490 95.665 ;
        RECT 99.670 95.545 99.840 95.835 ;
        RECT 101.270 95.755 101.440 95.835 ;
        RECT 100.010 95.285 100.340 95.665 ;
        RECT 100.810 95.505 101.440 95.755 ;
        RECT 101.620 95.285 102.040 95.665 ;
        RECT 102.240 95.545 102.480 95.835 ;
        RECT 102.710 95.285 103.040 95.975 ;
        RECT 103.210 95.545 103.380 96.155 ;
        RECT 103.730 96.005 103.980 96.595 ;
        RECT 104.700 96.265 104.880 97.125 ;
        RECT 103.650 95.495 103.980 96.005 ;
        RECT 104.160 95.285 104.445 96.085 ;
        RECT 104.625 95.795 104.880 96.265 ;
        RECT 105.425 97.375 105.985 97.665 ;
        RECT 106.155 97.375 106.405 97.835 ;
        RECT 105.425 96.005 105.675 97.375 ;
        RECT 107.025 97.205 107.355 97.565 ;
        RECT 105.965 97.015 107.355 97.205 ;
        RECT 108.645 97.110 108.935 97.835 ;
        RECT 109.110 97.095 109.365 97.665 ;
        RECT 109.535 97.435 109.865 97.835 ;
        RECT 110.290 97.300 110.820 97.665 ;
        RECT 111.010 97.495 111.285 97.665 ;
        RECT 111.005 97.325 111.285 97.495 ;
        RECT 110.290 97.265 110.465 97.300 ;
        RECT 109.535 97.095 110.465 97.265 ;
        RECT 105.965 96.925 106.135 97.015 ;
        RECT 105.845 96.595 106.135 96.925 ;
        RECT 106.305 96.595 106.645 96.845 ;
        RECT 106.865 96.595 107.540 96.845 ;
        RECT 105.965 96.345 106.135 96.595 ;
        RECT 105.965 96.175 106.905 96.345 ;
        RECT 107.275 96.235 107.540 96.595 ;
        RECT 104.625 95.625 104.965 95.795 ;
        RECT 104.625 95.595 104.880 95.625 ;
        RECT 105.425 95.455 105.885 96.005 ;
        RECT 106.075 95.285 106.405 96.005 ;
        RECT 106.605 95.625 106.905 96.175 ;
        RECT 107.075 95.285 107.355 95.955 ;
        RECT 108.645 95.285 108.935 96.450 ;
        RECT 109.110 96.425 109.280 97.095 ;
        RECT 109.535 96.925 109.705 97.095 ;
        RECT 109.450 96.595 109.705 96.925 ;
        RECT 109.930 96.595 110.125 96.925 ;
        RECT 109.110 95.455 109.445 96.425 ;
        RECT 109.615 95.285 109.785 96.425 ;
        RECT 109.955 95.625 110.125 96.595 ;
        RECT 110.295 95.965 110.465 97.095 ;
        RECT 110.635 96.305 110.805 97.105 ;
        RECT 111.010 96.505 111.285 97.325 ;
        RECT 111.455 96.305 111.645 97.665 ;
        RECT 111.825 97.300 112.335 97.835 ;
        RECT 112.555 97.025 112.800 97.630 ;
        RECT 113.795 97.285 113.965 97.575 ;
        RECT 114.135 97.455 114.465 97.835 ;
        RECT 113.795 97.115 114.460 97.285 ;
        RECT 111.845 96.855 113.075 97.025 ;
        RECT 110.635 96.135 111.645 96.305 ;
        RECT 111.815 96.290 112.565 96.480 ;
        RECT 110.295 95.795 111.420 95.965 ;
        RECT 111.815 95.625 111.985 96.290 ;
        RECT 112.735 96.045 113.075 96.855 ;
        RECT 113.710 96.295 114.060 96.945 ;
        RECT 114.230 96.125 114.460 97.115 ;
        RECT 109.955 95.455 111.985 95.625 ;
        RECT 112.155 95.285 112.325 96.045 ;
        RECT 112.560 95.635 113.075 96.045 ;
        RECT 113.795 95.955 114.460 96.125 ;
        RECT 113.795 95.455 113.965 95.955 ;
        RECT 114.135 95.285 114.465 95.785 ;
        RECT 114.635 95.455 114.860 97.575 ;
        RECT 115.075 97.455 115.405 97.835 ;
        RECT 115.575 97.285 115.745 97.615 ;
        RECT 116.045 97.455 117.060 97.655 ;
        RECT 115.050 97.095 115.745 97.285 ;
        RECT 115.050 96.125 115.220 97.095 ;
        RECT 115.390 96.295 115.800 96.915 ;
        RECT 115.970 96.345 116.190 97.215 ;
        RECT 116.370 96.905 116.720 97.275 ;
        RECT 116.890 96.725 117.060 97.455 ;
        RECT 117.230 97.395 117.640 97.835 ;
        RECT 117.930 97.195 118.180 97.625 ;
        RECT 118.380 97.375 118.700 97.835 ;
        RECT 119.260 97.445 120.110 97.615 ;
        RECT 117.230 96.855 117.640 97.185 ;
        RECT 117.930 96.855 118.350 97.195 ;
        RECT 116.640 96.685 117.060 96.725 ;
        RECT 116.640 96.515 117.990 96.685 ;
        RECT 115.050 95.955 115.745 96.125 ;
        RECT 115.970 95.965 116.470 96.345 ;
        RECT 115.075 95.285 115.405 95.785 ;
        RECT 115.575 95.455 115.745 95.955 ;
        RECT 116.640 95.670 116.810 96.515 ;
        RECT 117.740 96.355 117.990 96.515 ;
        RECT 116.980 96.085 117.230 96.345 ;
        RECT 118.160 96.085 118.350 96.855 ;
        RECT 116.980 95.835 118.350 96.085 ;
        RECT 118.520 97.025 119.770 97.195 ;
        RECT 118.520 96.265 118.690 97.025 ;
        RECT 119.440 96.905 119.770 97.025 ;
        RECT 118.860 96.445 119.040 96.855 ;
        RECT 119.940 96.685 120.110 97.445 ;
        RECT 120.310 97.355 120.970 97.835 ;
        RECT 121.150 97.240 121.470 97.570 ;
        RECT 120.300 96.915 120.960 97.185 ;
        RECT 120.300 96.855 120.630 96.915 ;
        RECT 120.780 96.685 121.110 96.745 ;
        RECT 119.210 96.515 121.110 96.685 ;
        RECT 118.520 95.955 119.040 96.265 ;
        RECT 119.210 96.005 119.380 96.515 ;
        RECT 121.280 96.345 121.470 97.240 ;
        RECT 119.550 96.175 121.470 96.345 ;
        RECT 121.150 96.155 121.470 96.175 ;
        RECT 121.670 96.925 121.920 97.575 ;
        RECT 122.100 97.375 122.385 97.835 ;
        RECT 122.565 97.125 122.820 97.655 ;
        RECT 121.670 96.595 122.470 96.925 ;
        RECT 119.210 95.835 120.420 96.005 ;
        RECT 115.980 95.500 116.810 95.670 ;
        RECT 117.050 95.285 117.430 95.665 ;
        RECT 117.610 95.545 117.780 95.835 ;
        RECT 119.210 95.755 119.380 95.835 ;
        RECT 117.950 95.285 118.280 95.665 ;
        RECT 118.750 95.505 119.380 95.755 ;
        RECT 119.560 95.285 119.980 95.665 ;
        RECT 120.180 95.545 120.420 95.835 ;
        RECT 120.650 95.285 120.980 95.975 ;
        RECT 121.150 95.545 121.320 96.155 ;
        RECT 121.670 96.005 121.920 96.595 ;
        RECT 122.640 96.265 122.820 97.125 ;
        RECT 124.285 97.085 125.495 97.835 ;
        RECT 121.590 95.495 121.920 96.005 ;
        RECT 122.100 95.285 122.385 96.085 ;
        RECT 122.565 95.795 122.820 96.265 ;
        RECT 124.285 96.375 124.805 96.915 ;
        RECT 124.975 96.545 125.495 97.085 ;
        RECT 122.565 95.625 122.905 95.795 ;
        RECT 122.565 95.595 122.820 95.625 ;
        RECT 124.285 95.285 125.495 96.375 ;
        RECT 5.520 95.115 125.580 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 6.985 94.025 8.655 95.115 ;
        RECT 8.915 94.445 9.085 94.945 ;
        RECT 9.255 94.615 9.585 95.115 ;
        RECT 8.915 94.275 9.580 94.445 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 6.985 93.335 7.735 93.855 ;
        RECT 7.905 93.505 8.655 94.025 ;
        RECT 8.830 93.455 9.180 94.105 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 6.985 92.565 8.655 93.335 ;
        RECT 9.350 93.285 9.580 94.275 ;
        RECT 8.915 93.115 9.580 93.285 ;
        RECT 8.915 92.825 9.085 93.115 ;
        RECT 9.255 92.565 9.585 92.945 ;
        RECT 9.755 92.825 9.980 94.945 ;
        RECT 10.195 94.615 10.525 95.115 ;
        RECT 10.695 94.445 10.865 94.945 ;
        RECT 11.100 94.730 11.930 94.900 ;
        RECT 12.170 94.735 12.550 95.115 ;
        RECT 10.170 94.275 10.865 94.445 ;
        RECT 10.170 93.305 10.340 94.275 ;
        RECT 10.510 93.485 10.920 94.105 ;
        RECT 11.090 94.055 11.590 94.435 ;
        RECT 10.170 93.115 10.865 93.305 ;
        RECT 11.090 93.185 11.310 94.055 ;
        RECT 11.760 93.885 11.930 94.730 ;
        RECT 12.730 94.565 12.900 94.855 ;
        RECT 13.070 94.735 13.400 95.115 ;
        RECT 13.870 94.645 14.500 94.895 ;
        RECT 14.680 94.735 15.100 95.115 ;
        RECT 14.330 94.565 14.500 94.645 ;
        RECT 15.300 94.565 15.540 94.855 ;
        RECT 12.100 94.315 13.470 94.565 ;
        RECT 12.100 94.055 12.350 94.315 ;
        RECT 12.860 93.885 13.110 94.045 ;
        RECT 11.760 93.715 13.110 93.885 ;
        RECT 11.760 93.675 12.180 93.715 ;
        RECT 11.490 93.125 11.840 93.495 ;
        RECT 10.195 92.565 10.525 92.945 ;
        RECT 10.695 92.785 10.865 93.115 ;
        RECT 12.010 92.945 12.180 93.675 ;
        RECT 13.280 93.545 13.470 94.315 ;
        RECT 12.350 93.215 12.760 93.545 ;
        RECT 13.050 93.205 13.470 93.545 ;
        RECT 13.640 94.135 14.160 94.445 ;
        RECT 14.330 94.395 15.540 94.565 ;
        RECT 15.770 94.425 16.100 95.115 ;
        RECT 13.640 93.375 13.810 94.135 ;
        RECT 13.980 93.545 14.160 93.955 ;
        RECT 14.330 93.885 14.500 94.395 ;
        RECT 16.270 94.245 16.440 94.855 ;
        RECT 16.710 94.395 17.040 94.905 ;
        RECT 16.270 94.225 16.590 94.245 ;
        RECT 14.670 94.055 16.590 94.225 ;
        RECT 14.330 93.715 16.230 93.885 ;
        RECT 14.560 93.375 14.890 93.495 ;
        RECT 13.640 93.205 14.890 93.375 ;
        RECT 11.165 92.745 12.180 92.945 ;
        RECT 12.350 92.565 12.760 93.005 ;
        RECT 13.050 92.775 13.300 93.205 ;
        RECT 13.500 92.565 13.820 93.025 ;
        RECT 15.060 92.955 15.230 93.715 ;
        RECT 15.900 93.655 16.230 93.715 ;
        RECT 15.420 93.485 15.750 93.545 ;
        RECT 15.420 93.215 16.080 93.485 ;
        RECT 16.400 93.160 16.590 94.055 ;
        RECT 14.380 92.785 15.230 92.955 ;
        RECT 15.430 92.565 16.090 93.045 ;
        RECT 16.270 92.830 16.590 93.160 ;
        RECT 16.790 93.805 17.040 94.395 ;
        RECT 17.220 94.315 17.505 95.115 ;
        RECT 17.685 94.135 17.940 94.805 ;
        RECT 16.790 93.475 17.590 93.805 ;
        RECT 16.790 92.825 17.040 93.475 ;
        RECT 17.760 93.275 17.940 94.135 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 18.945 94.680 24.290 95.115 ;
        RECT 17.685 93.075 17.940 93.275 ;
        RECT 17.220 92.565 17.505 93.025 ;
        RECT 17.685 92.905 18.025 93.075 ;
        RECT 17.685 92.745 17.940 92.905 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 20.530 93.110 20.870 93.940 ;
        RECT 22.350 93.430 22.700 94.680 ;
        RECT 24.465 94.025 26.135 95.115 ;
        RECT 24.465 93.335 25.215 93.855 ;
        RECT 25.385 93.505 26.135 94.025 ;
        RECT 26.395 94.185 26.565 94.945 ;
        RECT 26.745 94.355 27.075 95.115 ;
        RECT 26.395 94.015 27.060 94.185 ;
        RECT 27.245 94.040 27.515 94.945 ;
        RECT 27.775 94.445 27.945 94.945 ;
        RECT 28.115 94.615 28.445 95.115 ;
        RECT 27.775 94.275 28.440 94.445 ;
        RECT 26.890 93.870 27.060 94.015 ;
        RECT 26.325 93.465 26.655 93.835 ;
        RECT 26.890 93.540 27.175 93.870 ;
        RECT 18.945 92.565 24.290 93.110 ;
        RECT 24.465 92.565 26.135 93.335 ;
        RECT 26.890 93.285 27.060 93.540 ;
        RECT 26.395 93.115 27.060 93.285 ;
        RECT 27.345 93.240 27.515 94.040 ;
        RECT 27.690 93.455 28.040 94.105 ;
        RECT 28.210 93.285 28.440 94.275 ;
        RECT 26.395 92.735 26.565 93.115 ;
        RECT 26.745 92.565 27.075 92.945 ;
        RECT 27.255 92.735 27.515 93.240 ;
        RECT 27.775 93.115 28.440 93.285 ;
        RECT 27.775 92.825 27.945 93.115 ;
        RECT 28.115 92.565 28.445 92.945 ;
        RECT 28.615 92.825 28.840 94.945 ;
        RECT 29.055 94.615 29.385 95.115 ;
        RECT 29.555 94.445 29.725 94.945 ;
        RECT 29.960 94.730 30.790 94.900 ;
        RECT 31.030 94.735 31.410 95.115 ;
        RECT 29.030 94.275 29.725 94.445 ;
        RECT 29.030 93.305 29.200 94.275 ;
        RECT 29.370 93.485 29.780 94.105 ;
        RECT 29.950 94.055 30.450 94.435 ;
        RECT 29.030 93.115 29.725 93.305 ;
        RECT 29.950 93.185 30.170 94.055 ;
        RECT 30.620 93.885 30.790 94.730 ;
        RECT 31.590 94.565 31.760 94.855 ;
        RECT 31.930 94.735 32.260 95.115 ;
        RECT 32.730 94.645 33.360 94.895 ;
        RECT 33.540 94.735 33.960 95.115 ;
        RECT 33.190 94.565 33.360 94.645 ;
        RECT 34.160 94.565 34.400 94.855 ;
        RECT 30.960 94.315 32.330 94.565 ;
        RECT 30.960 94.055 31.210 94.315 ;
        RECT 31.720 93.885 31.970 94.045 ;
        RECT 30.620 93.715 31.970 93.885 ;
        RECT 30.620 93.675 31.040 93.715 ;
        RECT 30.350 93.125 30.700 93.495 ;
        RECT 29.055 92.565 29.385 92.945 ;
        RECT 29.555 92.785 29.725 93.115 ;
        RECT 30.870 92.945 31.040 93.675 ;
        RECT 32.140 93.545 32.330 94.315 ;
        RECT 31.210 93.215 31.620 93.545 ;
        RECT 31.910 93.205 32.330 93.545 ;
        RECT 32.500 94.135 33.020 94.445 ;
        RECT 33.190 94.395 34.400 94.565 ;
        RECT 34.630 94.425 34.960 95.115 ;
        RECT 32.500 93.375 32.670 94.135 ;
        RECT 32.840 93.545 33.020 93.955 ;
        RECT 33.190 93.885 33.360 94.395 ;
        RECT 35.130 94.245 35.300 94.855 ;
        RECT 35.570 94.395 35.900 94.905 ;
        RECT 35.130 94.225 35.450 94.245 ;
        RECT 33.530 94.055 35.450 94.225 ;
        RECT 33.190 93.715 35.090 93.885 ;
        RECT 33.420 93.375 33.750 93.495 ;
        RECT 32.500 93.205 33.750 93.375 ;
        RECT 30.025 92.745 31.040 92.945 ;
        RECT 31.210 92.565 31.620 93.005 ;
        RECT 31.910 92.775 32.160 93.205 ;
        RECT 32.360 92.565 32.680 93.025 ;
        RECT 33.920 92.955 34.090 93.715 ;
        RECT 34.760 93.655 35.090 93.715 ;
        RECT 34.280 93.485 34.610 93.545 ;
        RECT 34.280 93.215 34.940 93.485 ;
        RECT 35.260 93.160 35.450 94.055 ;
        RECT 33.240 92.785 34.090 92.955 ;
        RECT 34.290 92.565 34.950 93.045 ;
        RECT 35.130 92.830 35.450 93.160 ;
        RECT 35.650 93.805 35.900 94.395 ;
        RECT 36.080 94.315 36.365 95.115 ;
        RECT 36.545 94.135 36.800 94.805 ;
        RECT 35.650 93.475 36.450 93.805 ;
        RECT 35.650 92.825 35.900 93.475 ;
        RECT 36.620 93.275 36.800 94.135 ;
        RECT 36.545 93.075 36.800 93.275 ;
        RECT 38.270 93.975 38.605 94.945 ;
        RECT 38.775 93.975 38.945 95.115 ;
        RECT 39.115 94.775 41.145 94.945 ;
        RECT 38.270 93.305 38.440 93.975 ;
        RECT 39.115 93.805 39.285 94.775 ;
        RECT 38.610 93.475 38.865 93.805 ;
        RECT 39.090 93.475 39.285 93.805 ;
        RECT 39.455 94.435 40.580 94.605 ;
        RECT 38.695 93.305 38.865 93.475 ;
        RECT 39.455 93.305 39.625 94.435 ;
        RECT 36.080 92.565 36.365 93.025 ;
        RECT 36.545 92.905 36.885 93.075 ;
        RECT 36.545 92.745 36.800 92.905 ;
        RECT 38.270 92.735 38.525 93.305 ;
        RECT 38.695 93.135 39.625 93.305 ;
        RECT 39.795 94.095 40.805 94.265 ;
        RECT 39.795 93.295 39.965 94.095 ;
        RECT 39.450 93.100 39.625 93.135 ;
        RECT 38.695 92.565 39.025 92.965 ;
        RECT 39.450 92.735 39.980 93.100 ;
        RECT 40.170 93.075 40.445 93.895 ;
        RECT 40.165 92.905 40.445 93.075 ;
        RECT 40.170 92.735 40.445 92.905 ;
        RECT 40.615 92.735 40.805 94.095 ;
        RECT 40.975 94.110 41.145 94.775 ;
        RECT 41.315 94.355 41.485 95.115 ;
        RECT 41.720 94.355 42.235 94.765 ;
        RECT 40.975 93.920 41.725 94.110 ;
        RECT 41.895 93.545 42.235 94.355 ;
        RECT 42.465 93.975 42.675 95.115 ;
        RECT 41.005 93.375 42.235 93.545 ;
        RECT 42.845 93.965 43.175 94.945 ;
        RECT 43.345 93.975 43.575 95.115 ;
        RECT 40.985 92.565 41.495 93.100 ;
        RECT 41.715 92.770 41.960 93.375 ;
        RECT 42.465 92.565 42.675 93.385 ;
        RECT 42.845 93.365 43.095 93.965 ;
        RECT 44.245 93.950 44.535 95.115 ;
        RECT 44.705 94.680 50.050 95.115 ;
        RECT 50.225 94.680 55.570 95.115 ;
        RECT 43.265 93.555 43.595 93.805 ;
        RECT 42.845 92.735 43.175 93.365 ;
        RECT 43.345 92.565 43.575 93.385 ;
        RECT 44.245 92.565 44.535 93.290 ;
        RECT 46.290 93.110 46.630 93.940 ;
        RECT 48.110 93.430 48.460 94.680 ;
        RECT 51.810 93.110 52.150 93.940 ;
        RECT 53.630 93.430 53.980 94.680 ;
        RECT 56.665 93.975 56.935 94.945 ;
        RECT 57.145 94.315 57.425 95.115 ;
        RECT 57.595 94.605 59.250 94.895 ;
        RECT 57.660 94.265 59.250 94.435 ;
        RECT 57.660 94.145 57.830 94.265 ;
        RECT 57.105 93.975 57.830 94.145 ;
        RECT 56.665 93.240 56.835 93.975 ;
        RECT 57.105 93.805 57.275 93.975 ;
        RECT 58.020 93.925 58.735 94.095 ;
        RECT 58.930 93.975 59.250 94.265 ;
        RECT 59.425 94.025 62.935 95.115 ;
        RECT 57.005 93.475 57.275 93.805 ;
        RECT 57.445 93.475 57.850 93.805 ;
        RECT 58.020 93.475 58.730 93.925 ;
        RECT 57.105 93.305 57.275 93.475 ;
        RECT 44.705 92.565 50.050 93.110 ;
        RECT 50.225 92.565 55.570 93.110 ;
        RECT 56.665 92.895 56.935 93.240 ;
        RECT 57.105 93.135 58.715 93.305 ;
        RECT 58.900 93.235 59.250 93.805 ;
        RECT 59.425 93.335 61.075 93.855 ;
        RECT 61.245 93.505 62.935 94.025 ;
        RECT 64.025 94.145 64.295 94.915 ;
        RECT 64.465 94.335 64.795 95.115 ;
        RECT 65.000 94.510 65.185 94.915 ;
        RECT 65.355 94.690 65.690 95.115 ;
        RECT 65.000 94.335 65.665 94.510 ;
        RECT 64.025 93.975 65.155 94.145 ;
        RECT 57.125 92.565 57.505 92.965 ;
        RECT 57.675 92.785 57.845 93.135 ;
        RECT 58.015 92.565 58.345 92.965 ;
        RECT 58.545 92.785 58.715 93.135 ;
        RECT 58.915 92.565 59.245 93.065 ;
        RECT 59.425 92.565 62.935 93.335 ;
        RECT 64.025 93.065 64.195 93.975 ;
        RECT 64.365 93.225 64.725 93.805 ;
        RECT 64.905 93.475 65.155 93.975 ;
        RECT 65.325 93.305 65.665 94.335 ;
        RECT 65.865 94.025 69.375 95.115 ;
        RECT 64.980 93.135 65.665 93.305 ;
        RECT 65.865 93.335 67.515 93.855 ;
        RECT 67.685 93.505 69.375 94.025 ;
        RECT 70.005 93.950 70.295 95.115 ;
        RECT 70.465 94.355 70.980 94.765 ;
        RECT 71.215 94.355 71.385 95.115 ;
        RECT 71.555 94.775 73.585 94.945 ;
        RECT 70.465 93.545 70.805 94.355 ;
        RECT 71.555 94.110 71.725 94.775 ;
        RECT 72.120 94.435 73.245 94.605 ;
        RECT 70.975 93.920 71.725 94.110 ;
        RECT 71.895 94.095 72.905 94.265 ;
        RECT 70.465 93.375 71.695 93.545 ;
        RECT 64.025 92.735 64.285 93.065 ;
        RECT 64.495 92.565 64.770 93.045 ;
        RECT 64.980 92.735 65.185 93.135 ;
        RECT 65.355 92.565 65.690 92.965 ;
        RECT 65.865 92.565 69.375 93.335 ;
        RECT 70.005 92.565 70.295 93.290 ;
        RECT 70.740 92.770 70.985 93.375 ;
        RECT 71.205 92.565 71.715 93.100 ;
        RECT 71.895 92.735 72.085 94.095 ;
        RECT 72.255 93.075 72.530 93.895 ;
        RECT 72.735 93.295 72.905 94.095 ;
        RECT 73.075 93.305 73.245 94.435 ;
        RECT 73.415 93.805 73.585 94.775 ;
        RECT 73.755 93.975 73.925 95.115 ;
        RECT 74.095 93.975 74.430 94.945 ;
        RECT 74.605 94.025 78.115 95.115 ;
        RECT 73.415 93.475 73.610 93.805 ;
        RECT 73.835 93.475 74.090 93.805 ;
        RECT 73.835 93.305 74.005 93.475 ;
        RECT 74.260 93.305 74.430 93.975 ;
        RECT 73.075 93.135 74.005 93.305 ;
        RECT 73.075 93.100 73.250 93.135 ;
        RECT 72.255 92.905 72.535 93.075 ;
        RECT 72.255 92.735 72.530 92.905 ;
        RECT 72.720 92.735 73.250 93.100 ;
        RECT 73.675 92.565 74.005 92.965 ;
        RECT 74.175 92.735 74.430 93.305 ;
        RECT 74.605 93.335 76.255 93.855 ;
        RECT 76.425 93.505 78.115 94.025 ;
        RECT 78.285 93.975 78.555 94.945 ;
        RECT 78.765 94.315 79.045 95.115 ;
        RECT 79.215 94.605 80.870 94.895 ;
        RECT 79.280 94.265 80.870 94.435 ;
        RECT 79.280 94.145 79.450 94.265 ;
        RECT 78.725 93.975 79.450 94.145 ;
        RECT 74.605 92.565 78.115 93.335 ;
        RECT 78.285 93.240 78.455 93.975 ;
        RECT 78.725 93.805 78.895 93.975 ;
        RECT 79.640 93.925 80.355 94.095 ;
        RECT 80.550 93.975 80.870 94.265 ;
        RECT 81.045 94.025 83.635 95.115 ;
        RECT 78.625 93.475 78.895 93.805 ;
        RECT 79.065 93.475 79.470 93.805 ;
        RECT 79.640 93.475 80.350 93.925 ;
        RECT 78.725 93.305 78.895 93.475 ;
        RECT 78.285 92.895 78.555 93.240 ;
        RECT 78.725 93.135 80.335 93.305 ;
        RECT 80.520 93.235 80.870 93.805 ;
        RECT 81.045 93.335 82.255 93.855 ;
        RECT 82.425 93.505 83.635 94.025 ;
        RECT 84.470 94.145 84.800 94.945 ;
        RECT 84.970 94.315 85.300 95.115 ;
        RECT 85.600 94.145 85.930 94.945 ;
        RECT 86.575 94.315 86.825 95.115 ;
        RECT 84.470 93.975 86.905 94.145 ;
        RECT 87.095 93.975 87.265 95.115 ;
        RECT 87.435 93.975 87.775 94.945 ;
        RECT 87.945 94.680 93.290 95.115 ;
        RECT 84.265 93.555 84.615 93.805 ;
        RECT 84.800 93.345 84.970 93.975 ;
        RECT 85.140 93.555 85.470 93.755 ;
        RECT 85.640 93.555 85.970 93.755 ;
        RECT 86.140 93.555 86.560 93.755 ;
        RECT 86.735 93.725 86.905 93.975 ;
        RECT 86.735 93.555 87.430 93.725 ;
        RECT 78.745 92.565 79.125 92.965 ;
        RECT 79.295 92.785 79.465 93.135 ;
        RECT 79.635 92.565 79.965 92.965 ;
        RECT 80.165 92.785 80.335 93.135 ;
        RECT 80.535 92.565 80.865 93.065 ;
        RECT 81.045 92.565 83.635 93.335 ;
        RECT 84.470 92.735 84.970 93.345 ;
        RECT 85.600 93.215 86.825 93.385 ;
        RECT 87.600 93.365 87.775 93.975 ;
        RECT 85.600 92.735 85.930 93.215 ;
        RECT 86.100 92.565 86.325 93.025 ;
        RECT 86.495 92.735 86.825 93.215 ;
        RECT 87.015 92.565 87.265 93.365 ;
        RECT 87.435 92.735 87.775 93.365 ;
        RECT 89.530 93.110 89.870 93.940 ;
        RECT 91.350 93.430 91.700 94.680 ;
        RECT 93.465 94.395 93.925 94.945 ;
        RECT 94.115 94.395 94.445 95.115 ;
        RECT 87.945 92.565 93.290 93.110 ;
        RECT 93.465 93.025 93.715 94.395 ;
        RECT 94.645 94.225 94.945 94.775 ;
        RECT 95.115 94.445 95.395 95.115 ;
        RECT 94.005 94.055 94.945 94.225 ;
        RECT 94.005 93.805 94.175 94.055 ;
        RECT 95.315 93.805 95.580 94.165 ;
        RECT 95.765 93.950 96.055 95.115 ;
        RECT 96.225 94.025 97.435 95.115 ;
        RECT 93.885 93.475 94.175 93.805 ;
        RECT 94.345 93.555 94.685 93.805 ;
        RECT 94.905 93.555 95.580 93.805 ;
        RECT 94.005 93.385 94.175 93.475 ;
        RECT 94.005 93.195 95.395 93.385 ;
        RECT 96.225 93.315 96.745 93.855 ;
        RECT 96.915 93.485 97.435 94.025 ;
        RECT 97.610 93.975 97.945 94.945 ;
        RECT 98.115 93.975 98.285 95.115 ;
        RECT 98.455 94.775 100.485 94.945 ;
        RECT 93.465 92.735 94.025 93.025 ;
        RECT 94.195 92.565 94.445 93.025 ;
        RECT 95.065 92.835 95.395 93.195 ;
        RECT 95.765 92.565 96.055 93.290 ;
        RECT 96.225 92.565 97.435 93.315 ;
        RECT 97.610 93.305 97.780 93.975 ;
        RECT 98.455 93.805 98.625 94.775 ;
        RECT 97.950 93.475 98.205 93.805 ;
        RECT 98.430 93.475 98.625 93.805 ;
        RECT 98.795 94.435 99.920 94.605 ;
        RECT 98.035 93.305 98.205 93.475 ;
        RECT 98.795 93.305 98.965 94.435 ;
        RECT 97.610 92.735 97.865 93.305 ;
        RECT 98.035 93.135 98.965 93.305 ;
        RECT 99.135 94.095 100.145 94.265 ;
        RECT 99.135 93.295 99.305 94.095 ;
        RECT 99.510 93.415 99.785 93.895 ;
        RECT 99.505 93.245 99.785 93.415 ;
        RECT 98.790 93.100 98.965 93.135 ;
        RECT 98.035 92.565 98.365 92.965 ;
        RECT 98.790 92.735 99.320 93.100 ;
        RECT 99.510 92.735 99.785 93.245 ;
        RECT 99.955 92.735 100.145 94.095 ;
        RECT 100.315 94.110 100.485 94.775 ;
        RECT 100.655 94.355 100.825 95.115 ;
        RECT 101.060 94.355 101.575 94.765 ;
        RECT 100.315 93.920 101.065 94.110 ;
        RECT 101.235 93.545 101.575 94.355 ;
        RECT 101.745 94.025 105.255 95.115 ;
        RECT 105.425 94.025 106.635 95.115 ;
        RECT 100.345 93.375 101.575 93.545 ;
        RECT 100.325 92.565 100.835 93.100 ;
        RECT 101.055 92.770 101.300 93.375 ;
        RECT 101.745 93.335 103.395 93.855 ;
        RECT 103.565 93.505 105.255 94.025 ;
        RECT 101.745 92.565 105.255 93.335 ;
        RECT 105.425 93.315 105.945 93.855 ;
        RECT 106.115 93.485 106.635 94.025 ;
        RECT 106.805 94.040 107.075 94.945 ;
        RECT 107.245 94.355 107.575 95.115 ;
        RECT 107.755 94.185 107.925 94.945 ;
        RECT 108.185 94.680 113.530 95.115 ;
        RECT 105.425 92.565 106.635 93.315 ;
        RECT 106.805 93.240 106.975 94.040 ;
        RECT 107.260 94.015 107.925 94.185 ;
        RECT 107.260 93.870 107.430 94.015 ;
        RECT 107.145 93.540 107.430 93.870 ;
        RECT 107.260 93.285 107.430 93.540 ;
        RECT 107.665 93.465 107.995 93.835 ;
        RECT 106.805 92.735 107.065 93.240 ;
        RECT 107.260 93.115 107.925 93.285 ;
        RECT 107.245 92.565 107.575 92.945 ;
        RECT 107.755 92.735 107.925 93.115 ;
        RECT 109.770 93.110 110.110 93.940 ;
        RECT 111.590 93.430 111.940 94.680 ;
        RECT 113.705 94.025 117.215 95.115 ;
        RECT 113.705 93.335 115.355 93.855 ;
        RECT 115.525 93.505 117.215 94.025 ;
        RECT 117.905 93.975 118.115 95.115 ;
        RECT 118.285 93.965 118.615 94.945 ;
        RECT 118.785 93.975 119.015 95.115 ;
        RECT 119.225 94.025 120.895 95.115 ;
        RECT 108.185 92.565 113.530 93.110 ;
        RECT 113.705 92.565 117.215 93.335 ;
        RECT 117.905 92.565 118.115 93.385 ;
        RECT 118.285 93.365 118.535 93.965 ;
        RECT 118.705 93.555 119.035 93.805 ;
        RECT 118.285 92.735 118.615 93.365 ;
        RECT 118.785 92.565 119.015 93.385 ;
        RECT 119.225 93.335 119.975 93.855 ;
        RECT 120.145 93.505 120.895 94.025 ;
        RECT 121.525 93.950 121.815 95.115 ;
        RECT 121.985 94.025 123.655 95.115 ;
        RECT 121.985 93.335 122.735 93.855 ;
        RECT 122.905 93.505 123.655 94.025 ;
        RECT 124.285 94.025 125.495 95.115 ;
        RECT 124.285 93.485 124.805 94.025 ;
        RECT 119.225 92.565 120.895 93.335 ;
        RECT 121.525 92.565 121.815 93.290 ;
        RECT 121.985 92.565 123.655 93.335 ;
        RECT 124.975 93.315 125.495 93.855 ;
        RECT 124.285 92.565 125.495 93.315 ;
        RECT 5.520 92.395 125.580 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 7.535 91.845 7.705 92.135 ;
        RECT 7.875 92.015 8.205 92.395 ;
        RECT 7.535 91.675 8.200 91.845 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 7.450 90.855 7.800 91.505 ;
        RECT 7.970 90.685 8.200 91.675 ;
        RECT 7.535 90.515 8.200 90.685 ;
        RECT 7.535 90.015 7.705 90.515 ;
        RECT 7.875 89.845 8.205 90.345 ;
        RECT 8.375 90.015 8.600 92.135 ;
        RECT 8.815 92.015 9.145 92.395 ;
        RECT 9.315 91.845 9.485 92.175 ;
        RECT 9.785 92.015 10.800 92.215 ;
        RECT 8.790 91.655 9.485 91.845 ;
        RECT 8.790 90.685 8.960 91.655 ;
        RECT 9.130 90.855 9.540 91.475 ;
        RECT 9.710 90.905 9.930 91.775 ;
        RECT 10.110 91.465 10.460 91.835 ;
        RECT 10.630 91.285 10.800 92.015 ;
        RECT 10.970 91.955 11.380 92.395 ;
        RECT 11.670 91.755 11.920 92.185 ;
        RECT 12.120 91.935 12.440 92.395 ;
        RECT 13.000 92.005 13.850 92.175 ;
        RECT 10.970 91.415 11.380 91.745 ;
        RECT 11.670 91.415 12.090 91.755 ;
        RECT 10.380 91.245 10.800 91.285 ;
        RECT 10.380 91.075 11.730 91.245 ;
        RECT 8.790 90.515 9.485 90.685 ;
        RECT 9.710 90.525 10.210 90.905 ;
        RECT 8.815 89.845 9.145 90.345 ;
        RECT 9.315 90.015 9.485 90.515 ;
        RECT 10.380 90.230 10.550 91.075 ;
        RECT 11.480 90.915 11.730 91.075 ;
        RECT 10.720 90.645 10.970 90.905 ;
        RECT 11.900 90.645 12.090 91.415 ;
        RECT 10.720 90.395 12.090 90.645 ;
        RECT 12.260 91.585 13.510 91.755 ;
        RECT 12.260 90.825 12.430 91.585 ;
        RECT 13.180 91.465 13.510 91.585 ;
        RECT 12.600 91.005 12.780 91.415 ;
        RECT 13.680 91.245 13.850 92.005 ;
        RECT 14.050 91.915 14.710 92.395 ;
        RECT 14.890 91.800 15.210 92.130 ;
        RECT 14.040 91.475 14.700 91.745 ;
        RECT 14.040 91.415 14.370 91.475 ;
        RECT 14.520 91.245 14.850 91.305 ;
        RECT 12.950 91.075 14.850 91.245 ;
        RECT 12.260 90.515 12.780 90.825 ;
        RECT 12.950 90.565 13.120 91.075 ;
        RECT 15.020 90.905 15.210 91.800 ;
        RECT 13.290 90.735 15.210 90.905 ;
        RECT 14.890 90.715 15.210 90.735 ;
        RECT 15.410 91.485 15.660 92.135 ;
        RECT 15.840 91.935 16.125 92.395 ;
        RECT 16.305 91.685 16.560 92.215 ;
        RECT 15.410 91.155 16.210 91.485 ;
        RECT 16.380 91.375 16.560 91.685 ;
        RECT 17.110 91.655 17.365 92.225 ;
        RECT 17.535 91.995 17.865 92.395 ;
        RECT 18.290 91.860 18.820 92.225 ;
        RECT 18.290 91.825 18.465 91.860 ;
        RECT 17.535 91.655 18.465 91.825 ;
        RECT 16.380 91.205 16.645 91.375 ;
        RECT 12.950 90.395 14.160 90.565 ;
        RECT 9.720 90.060 10.550 90.230 ;
        RECT 10.790 89.845 11.170 90.225 ;
        RECT 11.350 90.105 11.520 90.395 ;
        RECT 12.950 90.315 13.120 90.395 ;
        RECT 11.690 89.845 12.020 90.225 ;
        RECT 12.490 90.065 13.120 90.315 ;
        RECT 13.300 89.845 13.720 90.225 ;
        RECT 13.920 90.105 14.160 90.395 ;
        RECT 14.390 89.845 14.720 90.535 ;
        RECT 14.890 90.105 15.060 90.715 ;
        RECT 15.410 90.565 15.660 91.155 ;
        RECT 16.380 90.825 16.560 91.205 ;
        RECT 15.330 90.055 15.660 90.565 ;
        RECT 15.840 89.845 16.125 90.645 ;
        RECT 16.305 90.155 16.560 90.825 ;
        RECT 17.110 90.985 17.280 91.655 ;
        RECT 17.535 91.485 17.705 91.655 ;
        RECT 17.450 91.155 17.705 91.485 ;
        RECT 17.930 91.155 18.125 91.485 ;
        RECT 17.110 90.015 17.445 90.985 ;
        RECT 17.615 89.845 17.785 90.985 ;
        RECT 17.955 90.185 18.125 91.155 ;
        RECT 18.295 90.525 18.465 91.655 ;
        RECT 18.635 90.865 18.805 91.665 ;
        RECT 19.010 91.375 19.285 92.225 ;
        RECT 19.005 91.205 19.285 91.375 ;
        RECT 19.010 91.065 19.285 91.205 ;
        RECT 19.455 90.865 19.645 92.225 ;
        RECT 19.825 91.860 20.335 92.395 ;
        RECT 20.555 91.585 20.800 92.190 ;
        RECT 19.845 91.415 21.075 91.585 ;
        RECT 21.305 91.575 21.515 92.395 ;
        RECT 21.685 91.595 22.015 92.225 ;
        RECT 18.635 90.695 19.645 90.865 ;
        RECT 19.815 90.850 20.565 91.040 ;
        RECT 18.295 90.355 19.420 90.525 ;
        RECT 19.815 90.185 19.985 90.850 ;
        RECT 20.735 90.605 21.075 91.415 ;
        RECT 21.685 90.995 21.935 91.595 ;
        RECT 22.185 91.575 22.415 92.395 ;
        RECT 22.625 91.625 24.295 92.395 ;
        RECT 24.475 91.895 24.805 92.395 ;
        RECT 25.005 91.825 25.175 92.175 ;
        RECT 25.375 91.995 25.705 92.395 ;
        RECT 25.875 91.825 26.045 92.175 ;
        RECT 26.215 91.995 26.595 92.395 ;
        RECT 22.105 91.155 22.435 91.405 ;
        RECT 22.625 91.105 23.375 91.625 ;
        RECT 17.955 90.015 19.985 90.185 ;
        RECT 20.155 89.845 20.325 90.605 ;
        RECT 20.560 90.195 21.075 90.605 ;
        RECT 21.305 89.845 21.515 90.985 ;
        RECT 21.685 90.015 22.015 90.995 ;
        RECT 22.185 89.845 22.415 90.985 ;
        RECT 23.545 90.935 24.295 91.455 ;
        RECT 24.470 91.155 24.820 91.725 ;
        RECT 25.005 91.655 26.615 91.825 ;
        RECT 26.785 91.720 27.055 92.065 ;
        RECT 26.445 91.485 26.615 91.655 ;
        RECT 24.990 91.035 25.700 91.485 ;
        RECT 25.870 91.155 26.275 91.485 ;
        RECT 26.445 91.155 26.715 91.485 ;
        RECT 22.625 89.845 24.295 90.935 ;
        RECT 24.470 90.695 24.790 90.985 ;
        RECT 24.985 90.865 25.700 91.035 ;
        RECT 26.445 90.985 26.615 91.155 ;
        RECT 26.885 90.985 27.055 91.720 ;
        RECT 27.225 91.645 28.435 92.395 ;
        RECT 28.605 91.720 28.875 92.065 ;
        RECT 29.065 91.995 29.445 92.395 ;
        RECT 29.615 91.825 29.785 92.175 ;
        RECT 29.955 91.995 30.285 92.395 ;
        RECT 30.485 91.825 30.655 92.175 ;
        RECT 30.855 91.895 31.185 92.395 ;
        RECT 27.225 91.105 27.745 91.645 ;
        RECT 25.890 90.815 26.615 90.985 ;
        RECT 25.890 90.695 26.060 90.815 ;
        RECT 24.470 90.525 26.060 90.695 ;
        RECT 24.470 90.065 26.125 90.355 ;
        RECT 26.295 89.845 26.575 90.645 ;
        RECT 26.785 90.015 27.055 90.985 ;
        RECT 27.915 90.935 28.435 91.475 ;
        RECT 27.225 89.845 28.435 90.935 ;
        RECT 28.605 90.985 28.775 91.720 ;
        RECT 29.045 91.655 30.655 91.825 ;
        RECT 29.045 91.485 29.215 91.655 ;
        RECT 28.945 91.155 29.215 91.485 ;
        RECT 29.385 91.155 29.790 91.485 ;
        RECT 29.045 90.985 29.215 91.155 ;
        RECT 29.960 91.035 30.670 91.485 ;
        RECT 30.840 91.155 31.190 91.725 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 31.830 91.655 32.085 92.225 ;
        RECT 32.255 91.995 32.585 92.395 ;
        RECT 33.010 91.860 33.540 92.225 ;
        RECT 33.010 91.825 33.185 91.860 ;
        RECT 32.255 91.655 33.185 91.825 ;
        RECT 33.730 91.715 34.005 92.225 ;
        RECT 28.605 90.015 28.875 90.985 ;
        RECT 29.045 90.815 29.770 90.985 ;
        RECT 29.960 90.865 30.675 91.035 ;
        RECT 29.600 90.695 29.770 90.815 ;
        RECT 30.870 90.695 31.190 90.985 ;
        RECT 29.085 89.845 29.365 90.645 ;
        RECT 29.600 90.525 31.190 90.695 ;
        RECT 29.535 90.065 31.190 90.355 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 31.830 90.985 32.000 91.655 ;
        RECT 32.255 91.485 32.425 91.655 ;
        RECT 32.170 91.155 32.425 91.485 ;
        RECT 32.650 91.155 32.845 91.485 ;
        RECT 31.830 90.015 32.165 90.985 ;
        RECT 32.335 89.845 32.505 90.985 ;
        RECT 32.675 90.185 32.845 91.155 ;
        RECT 33.015 90.525 33.185 91.655 ;
        RECT 33.355 90.865 33.525 91.665 ;
        RECT 33.725 91.545 34.005 91.715 ;
        RECT 33.730 91.065 34.005 91.545 ;
        RECT 34.175 90.865 34.365 92.225 ;
        RECT 34.545 91.860 35.055 92.395 ;
        RECT 35.275 91.585 35.520 92.190 ;
        RECT 35.965 91.850 41.310 92.395 ;
        RECT 41.485 91.850 46.830 92.395 ;
        RECT 47.005 91.850 52.350 92.395 ;
        RECT 34.565 91.415 35.795 91.585 ;
        RECT 33.355 90.695 34.365 90.865 ;
        RECT 34.535 90.850 35.285 91.040 ;
        RECT 33.015 90.355 34.140 90.525 ;
        RECT 34.535 90.185 34.705 90.850 ;
        RECT 35.455 90.605 35.795 91.415 ;
        RECT 37.550 91.020 37.890 91.850 ;
        RECT 32.675 90.015 34.705 90.185 ;
        RECT 34.875 89.845 35.045 90.605 ;
        RECT 35.280 90.195 35.795 90.605 ;
        RECT 39.370 90.280 39.720 91.530 ;
        RECT 43.070 91.020 43.410 91.850 ;
        RECT 44.890 90.280 45.240 91.530 ;
        RECT 48.590 91.020 48.930 91.850 ;
        RECT 52.525 91.625 56.035 92.395 ;
        RECT 57.125 91.670 57.415 92.395 ;
        RECT 57.595 91.895 57.925 92.395 ;
        RECT 58.125 91.825 58.295 92.175 ;
        RECT 58.495 91.995 58.825 92.395 ;
        RECT 58.995 91.825 59.165 92.175 ;
        RECT 59.335 91.995 59.715 92.395 ;
        RECT 50.410 90.280 50.760 91.530 ;
        RECT 52.525 91.105 54.175 91.625 ;
        RECT 54.345 90.935 56.035 91.455 ;
        RECT 57.590 91.155 57.940 91.725 ;
        RECT 58.125 91.655 59.735 91.825 ;
        RECT 59.905 91.720 60.175 92.065 ;
        RECT 59.565 91.485 59.735 91.655 ;
        RECT 35.965 89.845 41.310 90.280 ;
        RECT 41.485 89.845 46.830 90.280 ;
        RECT 47.005 89.845 52.350 90.280 ;
        RECT 52.525 89.845 56.035 90.935 ;
        RECT 57.125 89.845 57.415 91.010 ;
        RECT 57.590 90.695 57.910 90.985 ;
        RECT 58.110 90.865 58.820 91.485 ;
        RECT 58.990 91.155 59.395 91.485 ;
        RECT 59.565 91.155 59.835 91.485 ;
        RECT 59.565 90.985 59.735 91.155 ;
        RECT 60.005 90.985 60.175 91.720 ;
        RECT 60.345 91.625 62.935 92.395 ;
        RECT 63.570 91.995 63.905 92.395 ;
        RECT 64.075 91.825 64.280 92.225 ;
        RECT 64.490 91.915 64.765 92.395 ;
        RECT 64.975 91.895 65.235 92.225 ;
        RECT 63.595 91.655 64.280 91.825 ;
        RECT 60.345 91.105 61.555 91.625 ;
        RECT 59.010 90.815 59.735 90.985 ;
        RECT 59.010 90.695 59.180 90.815 ;
        RECT 57.590 90.525 59.180 90.695 ;
        RECT 57.590 90.065 59.245 90.355 ;
        RECT 59.415 89.845 59.695 90.645 ;
        RECT 59.905 90.015 60.175 90.985 ;
        RECT 61.725 90.935 62.935 91.455 ;
        RECT 60.345 89.845 62.935 90.935 ;
        RECT 63.595 90.625 63.935 91.655 ;
        RECT 64.105 90.985 64.355 91.485 ;
        RECT 64.535 91.155 64.895 91.735 ;
        RECT 65.065 90.985 65.235 91.895 ;
        RECT 65.410 91.845 65.665 92.135 ;
        RECT 65.835 92.015 66.165 92.395 ;
        RECT 65.410 91.675 66.160 91.845 ;
        RECT 64.105 90.815 65.235 90.985 ;
        RECT 65.410 90.855 65.760 91.505 ;
        RECT 63.595 90.450 64.260 90.625 ;
        RECT 63.570 89.845 63.905 90.270 ;
        RECT 64.075 90.045 64.260 90.450 ;
        RECT 64.465 89.845 64.795 90.625 ;
        RECT 64.965 90.045 65.235 90.815 ;
        RECT 65.930 90.685 66.160 91.675 ;
        RECT 65.410 90.515 66.160 90.685 ;
        RECT 65.410 90.015 65.665 90.515 ;
        RECT 65.835 89.845 66.165 90.345 ;
        RECT 66.335 90.015 66.505 92.135 ;
        RECT 66.865 92.035 67.195 92.395 ;
        RECT 67.365 92.005 67.860 92.175 ;
        RECT 68.065 92.005 68.920 92.175 ;
        RECT 66.735 90.815 67.195 91.865 ;
        RECT 66.675 90.030 67.000 90.815 ;
        RECT 67.365 90.645 67.535 92.005 ;
        RECT 67.705 91.095 68.055 91.715 ;
        RECT 68.225 91.495 68.580 91.715 ;
        RECT 68.225 90.905 68.395 91.495 ;
        RECT 68.750 91.295 68.920 92.005 ;
        RECT 69.795 91.935 70.125 92.395 ;
        RECT 70.335 92.035 70.685 92.205 ;
        RECT 69.125 91.465 69.915 91.715 ;
        RECT 70.335 91.645 70.595 92.035 ;
        RECT 70.905 91.945 71.855 92.225 ;
        RECT 72.025 91.955 72.215 92.395 ;
        RECT 72.385 92.015 73.455 92.185 ;
        RECT 70.085 91.295 70.255 91.475 ;
        RECT 67.365 90.475 67.760 90.645 ;
        RECT 67.930 90.515 68.395 90.905 ;
        RECT 68.565 91.125 70.255 91.295 ;
        RECT 67.590 90.345 67.760 90.475 ;
        RECT 68.565 90.345 68.735 91.125 ;
        RECT 70.425 90.955 70.595 91.645 ;
        RECT 69.095 90.785 70.595 90.955 ;
        RECT 70.785 90.985 70.995 91.775 ;
        RECT 71.165 91.155 71.515 91.775 ;
        RECT 71.685 91.165 71.855 91.945 ;
        RECT 72.385 91.785 72.555 92.015 ;
        RECT 72.025 91.615 72.555 91.785 ;
        RECT 72.025 91.335 72.245 91.615 ;
        RECT 72.725 91.445 72.965 91.845 ;
        RECT 71.685 90.995 72.090 91.165 ;
        RECT 72.425 91.075 72.965 91.445 ;
        RECT 73.135 91.660 73.455 92.015 ;
        RECT 73.700 91.935 74.005 92.395 ;
        RECT 74.175 91.685 74.430 92.215 ;
        RECT 73.135 91.485 73.460 91.660 ;
        RECT 73.135 91.185 74.050 91.485 ;
        RECT 73.310 91.155 74.050 91.185 ;
        RECT 70.785 90.825 71.460 90.985 ;
        RECT 71.920 90.905 72.090 90.995 ;
        RECT 70.785 90.815 71.750 90.825 ;
        RECT 70.425 90.645 70.595 90.785 ;
        RECT 67.170 89.845 67.420 90.305 ;
        RECT 67.590 90.015 67.840 90.345 ;
        RECT 68.055 90.015 68.735 90.345 ;
        RECT 68.905 90.445 69.980 90.615 ;
        RECT 70.425 90.475 70.985 90.645 ;
        RECT 71.290 90.525 71.750 90.815 ;
        RECT 71.920 90.735 73.140 90.905 ;
        RECT 68.905 90.105 69.075 90.445 ;
        RECT 69.310 89.845 69.640 90.275 ;
        RECT 69.810 90.105 69.980 90.445 ;
        RECT 70.275 89.845 70.645 90.305 ;
        RECT 70.815 90.015 70.985 90.475 ;
        RECT 71.920 90.355 72.090 90.735 ;
        RECT 73.310 90.565 73.480 91.155 ;
        RECT 74.220 91.035 74.430 91.685 ;
        RECT 71.220 90.015 72.090 90.355 ;
        RECT 72.680 90.395 73.480 90.565 ;
        RECT 72.260 89.845 72.510 90.305 ;
        RECT 72.680 90.105 72.850 90.395 ;
        RECT 73.030 89.845 73.360 90.225 ;
        RECT 73.700 89.845 74.005 90.985 ;
        RECT 74.175 90.155 74.430 91.035 ;
        RECT 74.605 91.655 74.990 92.225 ;
        RECT 75.160 91.935 75.485 92.395 ;
        RECT 76.005 91.765 76.285 92.225 ;
        RECT 74.605 90.985 74.885 91.655 ;
        RECT 75.160 91.595 76.285 91.765 ;
        RECT 75.160 91.485 75.610 91.595 ;
        RECT 75.055 91.155 75.610 91.485 ;
        RECT 76.475 91.425 76.875 92.225 ;
        RECT 77.275 91.935 77.545 92.395 ;
        RECT 77.715 91.765 78.000 92.225 ;
        RECT 74.605 90.015 74.990 90.985 ;
        RECT 75.160 90.695 75.610 91.155 ;
        RECT 75.780 90.865 76.875 91.425 ;
        RECT 75.160 90.475 76.285 90.695 ;
        RECT 75.160 89.845 75.485 90.305 ;
        RECT 76.005 90.015 76.285 90.475 ;
        RECT 76.475 90.015 76.875 90.865 ;
        RECT 77.045 91.595 78.000 91.765 ;
        RECT 78.490 91.615 78.990 92.225 ;
        RECT 77.045 90.695 77.255 91.595 ;
        RECT 77.425 90.865 78.115 91.425 ;
        RECT 78.285 91.155 78.635 91.405 ;
        RECT 78.820 90.985 78.990 91.615 ;
        RECT 79.620 91.745 79.950 92.225 ;
        RECT 80.120 91.935 80.345 92.395 ;
        RECT 80.515 91.745 80.845 92.225 ;
        RECT 79.620 91.575 80.845 91.745 ;
        RECT 81.035 91.595 81.285 92.395 ;
        RECT 81.455 91.595 81.795 92.225 ;
        RECT 82.885 91.670 83.175 92.395 ;
        RECT 83.345 91.720 83.615 92.065 ;
        RECT 83.805 91.995 84.185 92.395 ;
        RECT 84.355 91.825 84.525 92.175 ;
        RECT 84.695 91.995 85.025 92.395 ;
        RECT 85.225 91.825 85.395 92.175 ;
        RECT 85.595 91.895 85.925 92.395 ;
        RECT 81.565 91.545 81.795 91.595 ;
        RECT 79.160 91.205 79.490 91.405 ;
        RECT 79.660 91.205 79.990 91.405 ;
        RECT 80.160 91.205 80.580 91.405 ;
        RECT 80.755 91.235 81.450 91.405 ;
        RECT 80.755 90.985 80.925 91.235 ;
        RECT 81.620 90.985 81.795 91.545 ;
        RECT 78.490 90.815 80.925 90.985 ;
        RECT 77.045 90.475 78.000 90.695 ;
        RECT 77.275 89.845 77.545 90.305 ;
        RECT 77.715 90.015 78.000 90.475 ;
        RECT 78.490 90.015 78.820 90.815 ;
        RECT 78.990 89.845 79.320 90.645 ;
        RECT 79.620 90.015 79.950 90.815 ;
        RECT 80.595 89.845 80.845 90.645 ;
        RECT 81.115 89.845 81.285 90.985 ;
        RECT 81.455 90.015 81.795 90.985 ;
        RECT 82.885 89.845 83.175 91.010 ;
        RECT 83.345 90.985 83.515 91.720 ;
        RECT 83.785 91.655 85.395 91.825 ;
        RECT 83.785 91.485 83.955 91.655 ;
        RECT 83.685 91.155 83.955 91.485 ;
        RECT 84.125 91.155 84.530 91.485 ;
        RECT 83.785 90.985 83.955 91.155 ;
        RECT 84.700 91.035 85.410 91.485 ;
        RECT 85.580 91.155 85.930 91.725 ;
        RECT 86.105 91.645 87.315 92.395 ;
        RECT 86.105 91.105 86.625 91.645 ;
        RECT 87.760 91.585 88.005 92.190 ;
        RECT 88.225 91.860 88.735 92.395 ;
        RECT 83.345 90.015 83.615 90.985 ;
        RECT 83.785 90.815 84.510 90.985 ;
        RECT 84.700 90.865 85.415 91.035 ;
        RECT 84.340 90.695 84.510 90.815 ;
        RECT 85.610 90.695 85.930 90.985 ;
        RECT 86.795 90.935 87.315 91.475 ;
        RECT 83.825 89.845 84.105 90.645 ;
        RECT 84.340 90.525 85.930 90.695 ;
        RECT 84.275 90.065 85.930 90.355 ;
        RECT 86.105 89.845 87.315 90.935 ;
        RECT 87.485 91.415 88.715 91.585 ;
        RECT 87.485 90.605 87.825 91.415 ;
        RECT 87.995 90.850 88.745 91.040 ;
        RECT 87.485 90.195 88.000 90.605 ;
        RECT 88.235 89.845 88.405 90.605 ;
        RECT 88.575 90.185 88.745 90.850 ;
        RECT 88.915 90.865 89.105 92.225 ;
        RECT 89.275 92.055 89.550 92.225 ;
        RECT 89.275 91.885 89.555 92.055 ;
        RECT 89.275 91.065 89.550 91.885 ;
        RECT 89.740 91.860 90.270 92.225 ;
        RECT 90.695 91.995 91.025 92.395 ;
        RECT 90.095 91.825 90.270 91.860 ;
        RECT 89.755 90.865 89.925 91.665 ;
        RECT 88.915 90.695 89.925 90.865 ;
        RECT 90.095 91.655 91.025 91.825 ;
        RECT 91.195 91.655 91.450 92.225 ;
        RECT 90.095 90.525 90.265 91.655 ;
        RECT 90.855 91.485 91.025 91.655 ;
        RECT 89.140 90.355 90.265 90.525 ;
        RECT 90.435 91.155 90.630 91.485 ;
        RECT 90.855 91.155 91.110 91.485 ;
        RECT 90.435 90.185 90.605 91.155 ;
        RECT 91.280 90.985 91.450 91.655 ;
        RECT 88.575 90.015 90.605 90.185 ;
        RECT 90.775 89.845 90.945 90.985 ;
        RECT 91.115 90.015 91.450 90.985 ;
        RECT 91.625 91.720 91.885 92.225 ;
        RECT 92.065 92.015 92.395 92.395 ;
        RECT 92.575 91.845 92.745 92.225 ;
        RECT 91.625 90.920 91.795 91.720 ;
        RECT 92.080 91.675 92.745 91.845 ;
        RECT 92.080 91.420 92.250 91.675 ;
        RECT 93.065 91.575 93.275 92.395 ;
        RECT 93.445 91.595 93.775 92.225 ;
        RECT 91.965 91.090 92.250 91.420 ;
        RECT 92.485 91.125 92.815 91.495 ;
        RECT 92.080 90.945 92.250 91.090 ;
        RECT 93.445 90.995 93.695 91.595 ;
        RECT 93.945 91.575 94.175 92.395 ;
        RECT 94.385 91.850 99.730 92.395 ;
        RECT 99.905 91.850 105.250 92.395 ;
        RECT 93.865 91.155 94.195 91.405 ;
        RECT 95.970 91.020 96.310 91.850 ;
        RECT 91.625 90.015 91.895 90.920 ;
        RECT 92.080 90.775 92.745 90.945 ;
        RECT 92.065 89.845 92.395 90.605 ;
        RECT 92.575 90.015 92.745 90.775 ;
        RECT 93.065 89.845 93.275 90.985 ;
        RECT 93.445 90.015 93.775 90.995 ;
        RECT 93.945 89.845 94.175 90.985 ;
        RECT 97.790 90.280 98.140 91.530 ;
        RECT 101.490 91.020 101.830 91.850 ;
        RECT 105.425 91.625 108.015 92.395 ;
        RECT 108.645 91.670 108.935 92.395 ;
        RECT 109.105 91.625 112.615 92.395 ;
        RECT 112.785 91.645 113.995 92.395 ;
        RECT 114.170 91.655 114.425 92.225 ;
        RECT 114.595 91.995 114.925 92.395 ;
        RECT 115.350 91.860 115.880 92.225 ;
        RECT 115.350 91.825 115.525 91.860 ;
        RECT 114.595 91.655 115.525 91.825 ;
        RECT 103.310 90.280 103.660 91.530 ;
        RECT 105.425 91.105 106.635 91.625 ;
        RECT 106.805 90.935 108.015 91.455 ;
        RECT 109.105 91.105 110.755 91.625 ;
        RECT 94.385 89.845 99.730 90.280 ;
        RECT 99.905 89.845 105.250 90.280 ;
        RECT 105.425 89.845 108.015 90.935 ;
        RECT 108.645 89.845 108.935 91.010 ;
        RECT 110.925 90.935 112.615 91.455 ;
        RECT 112.785 91.105 113.305 91.645 ;
        RECT 113.475 90.935 113.995 91.475 ;
        RECT 109.105 89.845 112.615 90.935 ;
        RECT 112.785 89.845 113.995 90.935 ;
        RECT 114.170 90.985 114.340 91.655 ;
        RECT 114.595 91.485 114.765 91.655 ;
        RECT 114.510 91.155 114.765 91.485 ;
        RECT 114.990 91.155 115.185 91.485 ;
        RECT 114.170 90.015 114.505 90.985 ;
        RECT 114.675 89.845 114.845 90.985 ;
        RECT 115.015 90.185 115.185 91.155 ;
        RECT 115.355 90.525 115.525 91.655 ;
        RECT 115.695 90.865 115.865 91.665 ;
        RECT 116.070 91.375 116.345 92.225 ;
        RECT 116.065 91.205 116.345 91.375 ;
        RECT 116.070 91.065 116.345 91.205 ;
        RECT 116.515 90.865 116.705 92.225 ;
        RECT 116.885 91.860 117.395 92.395 ;
        RECT 117.615 91.585 117.860 92.190 ;
        RECT 118.580 91.585 118.825 92.190 ;
        RECT 119.045 91.860 119.555 92.395 ;
        RECT 116.905 91.415 118.135 91.585 ;
        RECT 115.695 90.695 116.705 90.865 ;
        RECT 116.875 90.850 117.625 91.040 ;
        RECT 115.355 90.355 116.480 90.525 ;
        RECT 116.875 90.185 117.045 90.850 ;
        RECT 117.795 90.605 118.135 91.415 ;
        RECT 115.015 90.015 117.045 90.185 ;
        RECT 117.215 89.845 117.385 90.605 ;
        RECT 117.620 90.195 118.135 90.605 ;
        RECT 118.305 91.415 119.535 91.585 ;
        RECT 118.305 90.605 118.645 91.415 ;
        RECT 118.815 90.850 119.565 91.040 ;
        RECT 118.305 90.195 118.820 90.605 ;
        RECT 119.055 89.845 119.225 90.605 ;
        RECT 119.395 90.185 119.565 90.850 ;
        RECT 119.735 90.865 119.925 92.225 ;
        RECT 120.095 91.375 120.370 92.225 ;
        RECT 120.560 91.860 121.090 92.225 ;
        RECT 121.515 91.995 121.845 92.395 ;
        RECT 120.915 91.825 121.090 91.860 ;
        RECT 120.095 91.205 120.375 91.375 ;
        RECT 120.095 91.065 120.370 91.205 ;
        RECT 120.575 90.865 120.745 91.665 ;
        RECT 119.735 90.695 120.745 90.865 ;
        RECT 120.915 91.655 121.845 91.825 ;
        RECT 122.015 91.655 122.270 92.225 ;
        RECT 120.915 90.525 121.085 91.655 ;
        RECT 121.675 91.485 121.845 91.655 ;
        RECT 119.960 90.355 121.085 90.525 ;
        RECT 121.255 91.155 121.450 91.485 ;
        RECT 121.675 91.155 121.930 91.485 ;
        RECT 121.255 90.185 121.425 91.155 ;
        RECT 122.100 90.985 122.270 91.655 ;
        RECT 122.445 91.625 124.115 92.395 ;
        RECT 124.285 91.645 125.495 92.395 ;
        RECT 122.445 91.105 123.195 91.625 ;
        RECT 119.395 90.015 121.425 90.185 ;
        RECT 121.595 89.845 121.765 90.985 ;
        RECT 121.935 90.015 122.270 90.985 ;
        RECT 123.365 90.935 124.115 91.455 ;
        RECT 122.445 89.845 124.115 90.935 ;
        RECT 124.285 90.935 124.805 91.475 ;
        RECT 124.975 91.105 125.495 91.645 ;
        RECT 124.285 89.845 125.495 90.935 ;
        RECT 5.520 89.675 125.580 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 6.985 88.585 10.495 89.675 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 6.985 87.895 8.635 88.415 ;
        RECT 8.805 88.065 10.495 88.585 ;
        RECT 10.665 88.600 10.935 89.505 ;
        RECT 11.105 88.915 11.435 89.675 ;
        RECT 11.615 88.745 11.785 89.505 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 6.985 87.125 10.495 87.895 ;
        RECT 10.665 87.800 10.835 88.600 ;
        RECT 11.120 88.575 11.785 88.745 ;
        RECT 11.120 88.430 11.290 88.575 ;
        RECT 12.565 88.535 12.775 89.675 ;
        RECT 11.005 88.100 11.290 88.430 ;
        RECT 12.945 88.525 13.275 89.505 ;
        RECT 13.445 88.535 13.675 89.675 ;
        RECT 13.890 88.535 14.225 89.505 ;
        RECT 14.395 88.535 14.565 89.675 ;
        RECT 14.735 89.335 16.765 89.505 ;
        RECT 11.120 87.845 11.290 88.100 ;
        RECT 11.525 88.025 11.855 88.395 ;
        RECT 10.665 87.295 10.925 87.800 ;
        RECT 11.120 87.675 11.785 87.845 ;
        RECT 11.105 87.125 11.435 87.505 ;
        RECT 11.615 87.295 11.785 87.675 ;
        RECT 12.565 87.125 12.775 87.945 ;
        RECT 12.945 87.925 13.195 88.525 ;
        RECT 13.365 88.115 13.695 88.365 ;
        RECT 12.945 87.295 13.275 87.925 ;
        RECT 13.445 87.125 13.675 87.945 ;
        RECT 13.890 87.865 14.060 88.535 ;
        RECT 14.735 88.365 14.905 89.335 ;
        RECT 14.230 88.035 14.485 88.365 ;
        RECT 14.710 88.035 14.905 88.365 ;
        RECT 15.075 88.995 16.200 89.165 ;
        RECT 14.315 87.865 14.485 88.035 ;
        RECT 15.075 87.865 15.245 88.995 ;
        RECT 13.890 87.295 14.145 87.865 ;
        RECT 14.315 87.695 15.245 87.865 ;
        RECT 15.415 88.655 16.425 88.825 ;
        RECT 15.415 87.855 15.585 88.655 ;
        RECT 15.070 87.660 15.245 87.695 ;
        RECT 14.315 87.125 14.645 87.525 ;
        RECT 15.070 87.295 15.600 87.660 ;
        RECT 15.790 87.635 16.065 88.455 ;
        RECT 15.785 87.465 16.065 87.635 ;
        RECT 15.790 87.295 16.065 87.465 ;
        RECT 16.235 87.295 16.425 88.655 ;
        RECT 16.595 88.670 16.765 89.335 ;
        RECT 16.935 88.915 17.105 89.675 ;
        RECT 17.340 88.915 17.855 89.325 ;
        RECT 16.595 88.480 17.345 88.670 ;
        RECT 17.515 88.105 17.855 88.915 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 18.945 88.585 20.615 89.675 ;
        RECT 16.625 87.935 17.855 88.105 ;
        RECT 16.605 87.125 17.115 87.660 ;
        RECT 17.335 87.330 17.580 87.935 ;
        RECT 18.945 87.895 19.695 88.415 ;
        RECT 19.865 88.065 20.615 88.585 ;
        RECT 21.450 88.705 21.780 89.505 ;
        RECT 21.950 88.875 22.280 89.675 ;
        RECT 22.580 88.705 22.910 89.505 ;
        RECT 23.555 88.875 23.805 89.675 ;
        RECT 21.450 88.535 23.885 88.705 ;
        RECT 24.075 88.535 24.245 89.675 ;
        RECT 24.415 88.535 24.755 89.505 ;
        RECT 26.050 88.705 26.380 89.505 ;
        RECT 26.550 88.875 26.880 89.675 ;
        RECT 27.180 88.705 27.510 89.505 ;
        RECT 28.155 88.875 28.405 89.675 ;
        RECT 26.050 88.535 28.485 88.705 ;
        RECT 28.675 88.535 28.845 89.675 ;
        RECT 29.015 88.535 29.355 89.505 ;
        RECT 29.525 88.585 33.035 89.675 ;
        RECT 21.245 88.115 21.595 88.365 ;
        RECT 21.780 87.905 21.950 88.535 ;
        RECT 22.120 88.115 22.450 88.315 ;
        RECT 22.620 88.115 22.950 88.315 ;
        RECT 23.120 88.115 23.540 88.315 ;
        RECT 23.715 88.285 23.885 88.535 ;
        RECT 23.715 88.115 24.410 88.285 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 18.945 87.125 20.615 87.895 ;
        RECT 21.450 87.295 21.950 87.905 ;
        RECT 22.580 87.775 23.805 87.945 ;
        RECT 24.580 87.925 24.755 88.535 ;
        RECT 25.845 88.115 26.195 88.365 ;
        RECT 22.580 87.295 22.910 87.775 ;
        RECT 23.080 87.125 23.305 87.585 ;
        RECT 23.475 87.295 23.805 87.775 ;
        RECT 23.995 87.125 24.245 87.925 ;
        RECT 24.415 87.295 24.755 87.925 ;
        RECT 26.380 87.905 26.550 88.535 ;
        RECT 26.720 88.115 27.050 88.315 ;
        RECT 27.220 88.115 27.550 88.315 ;
        RECT 27.720 88.115 28.140 88.315 ;
        RECT 28.315 88.285 28.485 88.535 ;
        RECT 28.315 88.115 29.010 88.285 ;
        RECT 26.050 87.295 26.550 87.905 ;
        RECT 27.180 87.775 28.405 87.945 ;
        RECT 29.180 87.925 29.355 88.535 ;
        RECT 27.180 87.295 27.510 87.775 ;
        RECT 27.680 87.125 27.905 87.585 ;
        RECT 28.075 87.295 28.405 87.775 ;
        RECT 28.595 87.125 28.845 87.925 ;
        RECT 29.015 87.295 29.355 87.925 ;
        RECT 29.525 87.895 31.175 88.415 ;
        RECT 31.345 88.065 33.035 88.585 ;
        RECT 33.870 88.705 34.200 89.505 ;
        RECT 34.370 88.875 34.700 89.675 ;
        RECT 35.000 88.705 35.330 89.505 ;
        RECT 35.975 88.875 36.225 89.675 ;
        RECT 33.870 88.535 36.305 88.705 ;
        RECT 36.495 88.535 36.665 89.675 ;
        RECT 36.835 88.535 37.175 89.505 ;
        RECT 37.350 89.165 39.005 89.455 ;
        RECT 37.350 88.825 38.940 88.995 ;
        RECT 39.175 88.875 39.455 89.675 ;
        RECT 37.350 88.535 37.670 88.825 ;
        RECT 38.770 88.705 38.940 88.825 ;
        RECT 33.665 88.115 34.015 88.365 ;
        RECT 34.200 87.905 34.370 88.535 ;
        RECT 34.540 88.115 34.870 88.315 ;
        RECT 35.040 88.115 35.370 88.315 ;
        RECT 35.540 88.115 35.960 88.315 ;
        RECT 36.135 88.285 36.305 88.535 ;
        RECT 36.135 88.115 36.830 88.285 ;
        RECT 37.000 87.975 37.175 88.535 ;
        RECT 37.865 88.485 38.580 88.655 ;
        RECT 38.770 88.535 39.495 88.705 ;
        RECT 39.665 88.535 39.935 89.505 ;
        RECT 40.105 88.585 43.615 89.675 ;
        RECT 29.525 87.125 33.035 87.895 ;
        RECT 33.870 87.295 34.370 87.905 ;
        RECT 35.000 87.775 36.225 87.945 ;
        RECT 36.945 87.925 37.175 87.975 ;
        RECT 35.000 87.295 35.330 87.775 ;
        RECT 35.500 87.125 35.725 87.585 ;
        RECT 35.895 87.295 36.225 87.775 ;
        RECT 36.415 87.125 36.665 87.925 ;
        RECT 36.835 87.295 37.175 87.925 ;
        RECT 37.350 87.795 37.700 88.365 ;
        RECT 37.870 88.035 38.580 88.485 ;
        RECT 39.325 88.365 39.495 88.535 ;
        RECT 38.750 88.035 39.155 88.365 ;
        RECT 39.325 88.035 39.595 88.365 ;
        RECT 39.325 87.865 39.495 88.035 ;
        RECT 37.885 87.695 39.495 87.865 ;
        RECT 39.765 87.800 39.935 88.535 ;
        RECT 37.355 87.125 37.685 87.625 ;
        RECT 37.885 87.345 38.055 87.695 ;
        RECT 38.255 87.125 38.585 87.525 ;
        RECT 38.755 87.345 38.925 87.695 ;
        RECT 39.095 87.125 39.475 87.525 ;
        RECT 39.665 87.455 39.935 87.800 ;
        RECT 40.105 87.895 41.755 88.415 ;
        RECT 41.925 88.065 43.615 88.585 ;
        RECT 44.245 88.510 44.535 89.675 ;
        RECT 44.705 88.585 45.915 89.675 ;
        RECT 40.105 87.125 43.615 87.895 ;
        RECT 44.705 87.875 45.225 88.415 ;
        RECT 45.395 88.045 45.915 88.585 ;
        RECT 46.175 88.745 46.345 89.505 ;
        RECT 46.525 88.915 46.855 89.675 ;
        RECT 46.175 88.575 46.840 88.745 ;
        RECT 47.025 88.600 47.295 89.505 ;
        RECT 46.670 88.430 46.840 88.575 ;
        RECT 46.105 88.025 46.435 88.395 ;
        RECT 46.670 88.100 46.955 88.430 ;
        RECT 44.245 87.125 44.535 87.850 ;
        RECT 44.705 87.125 45.915 87.875 ;
        RECT 46.670 87.845 46.840 88.100 ;
        RECT 46.175 87.675 46.840 87.845 ;
        RECT 47.125 87.800 47.295 88.600 ;
        RECT 46.175 87.295 46.345 87.675 ;
        RECT 46.525 87.125 46.855 87.505 ;
        RECT 47.035 87.295 47.295 87.800 ;
        RECT 47.465 88.600 47.735 89.505 ;
        RECT 47.905 88.915 48.235 89.675 ;
        RECT 48.415 88.745 48.585 89.505 ;
        RECT 47.465 87.800 47.635 88.600 ;
        RECT 47.920 88.575 48.585 88.745 ;
        RECT 47.920 88.430 48.090 88.575 ;
        RECT 47.805 88.100 48.090 88.430 ;
        RECT 49.310 88.535 49.645 89.505 ;
        RECT 49.815 88.535 49.985 89.675 ;
        RECT 50.155 89.335 52.185 89.505 ;
        RECT 47.920 87.845 48.090 88.100 ;
        RECT 48.325 88.025 48.655 88.395 ;
        RECT 49.310 87.865 49.480 88.535 ;
        RECT 50.155 88.365 50.325 89.335 ;
        RECT 49.650 88.035 49.905 88.365 ;
        RECT 50.130 88.035 50.325 88.365 ;
        RECT 50.495 88.995 51.620 89.165 ;
        RECT 49.735 87.865 49.905 88.035 ;
        RECT 50.495 87.865 50.665 88.995 ;
        RECT 47.465 87.295 47.725 87.800 ;
        RECT 47.920 87.675 48.585 87.845 ;
        RECT 47.905 87.125 48.235 87.505 ;
        RECT 48.415 87.295 48.585 87.675 ;
        RECT 49.310 87.295 49.565 87.865 ;
        RECT 49.735 87.695 50.665 87.865 ;
        RECT 50.835 88.655 51.845 88.825 ;
        RECT 50.835 87.855 51.005 88.655 ;
        RECT 51.210 87.975 51.485 88.455 ;
        RECT 51.205 87.805 51.485 87.975 ;
        RECT 50.490 87.660 50.665 87.695 ;
        RECT 49.735 87.125 50.065 87.525 ;
        RECT 50.490 87.295 51.020 87.660 ;
        RECT 51.210 87.295 51.485 87.805 ;
        RECT 51.655 87.295 51.845 88.655 ;
        RECT 52.015 88.670 52.185 89.335 ;
        RECT 52.355 88.915 52.525 89.675 ;
        RECT 52.760 88.915 53.275 89.325 ;
        RECT 52.015 88.480 52.765 88.670 ;
        RECT 52.935 88.105 53.275 88.915 ;
        RECT 52.045 87.935 53.275 88.105 ;
        RECT 53.450 88.535 53.785 89.505 ;
        RECT 53.955 88.535 54.125 89.675 ;
        RECT 54.295 89.335 56.325 89.505 ;
        RECT 52.025 87.125 52.535 87.660 ;
        RECT 52.755 87.330 53.000 87.935 ;
        RECT 53.450 87.865 53.620 88.535 ;
        RECT 54.295 88.365 54.465 89.335 ;
        RECT 53.790 88.035 54.045 88.365 ;
        RECT 54.270 88.035 54.465 88.365 ;
        RECT 54.635 88.995 55.760 89.165 ;
        RECT 53.875 87.865 54.045 88.035 ;
        RECT 54.635 87.865 54.805 88.995 ;
        RECT 53.450 87.295 53.705 87.865 ;
        RECT 53.875 87.695 54.805 87.865 ;
        RECT 54.975 88.655 55.985 88.825 ;
        RECT 54.975 87.855 55.145 88.655 ;
        RECT 55.350 88.315 55.625 88.455 ;
        RECT 55.345 88.145 55.625 88.315 ;
        RECT 54.630 87.660 54.805 87.695 ;
        RECT 53.875 87.125 54.205 87.525 ;
        RECT 54.630 87.295 55.160 87.660 ;
        RECT 55.350 87.295 55.625 88.145 ;
        RECT 55.795 87.295 55.985 88.655 ;
        RECT 56.155 88.670 56.325 89.335 ;
        RECT 56.495 88.915 56.665 89.675 ;
        RECT 56.900 88.915 57.415 89.325 ;
        RECT 56.155 88.480 56.905 88.670 ;
        RECT 57.075 88.105 57.415 88.915 ;
        RECT 56.185 87.935 57.415 88.105 ;
        RECT 57.585 88.535 57.925 89.505 ;
        RECT 58.095 88.535 58.265 89.675 ;
        RECT 58.535 88.875 58.785 89.675 ;
        RECT 59.430 88.705 59.760 89.505 ;
        RECT 60.060 88.875 60.390 89.675 ;
        RECT 60.560 88.705 60.890 89.505 ;
        RECT 61.265 89.240 66.610 89.675 ;
        RECT 58.455 88.535 60.890 88.705 ;
        RECT 56.165 87.125 56.675 87.660 ;
        RECT 56.895 87.330 57.140 87.935 ;
        RECT 57.585 87.925 57.760 88.535 ;
        RECT 58.455 88.285 58.625 88.535 ;
        RECT 57.930 88.115 58.625 88.285 ;
        RECT 58.800 88.115 59.220 88.315 ;
        RECT 59.390 88.115 59.720 88.315 ;
        RECT 59.890 88.115 60.220 88.315 ;
        RECT 57.585 87.295 57.925 87.925 ;
        RECT 58.095 87.125 58.345 87.925 ;
        RECT 58.535 87.775 59.760 87.945 ;
        RECT 58.535 87.295 58.865 87.775 ;
        RECT 59.035 87.125 59.260 87.585 ;
        RECT 59.430 87.295 59.760 87.775 ;
        RECT 60.390 87.905 60.560 88.535 ;
        RECT 60.745 88.115 61.095 88.365 ;
        RECT 60.390 87.295 60.890 87.905 ;
        RECT 62.850 87.670 63.190 88.500 ;
        RECT 64.670 87.990 65.020 89.240 ;
        RECT 67.705 88.600 67.975 89.505 ;
        RECT 68.145 88.915 68.475 89.675 ;
        RECT 68.655 88.745 68.825 89.505 ;
        RECT 67.705 87.800 67.875 88.600 ;
        RECT 68.160 88.575 68.825 88.745 ;
        RECT 68.160 88.430 68.330 88.575 ;
        RECT 70.005 88.510 70.295 89.675 ;
        RECT 70.470 88.535 70.805 89.505 ;
        RECT 70.975 88.535 71.145 89.675 ;
        RECT 71.315 89.335 73.345 89.505 ;
        RECT 68.045 88.100 68.330 88.430 ;
        RECT 68.160 87.845 68.330 88.100 ;
        RECT 68.565 88.025 68.895 88.395 ;
        RECT 70.470 87.865 70.640 88.535 ;
        RECT 71.315 88.365 71.485 89.335 ;
        RECT 70.810 88.035 71.065 88.365 ;
        RECT 71.290 88.035 71.485 88.365 ;
        RECT 71.655 88.995 72.780 89.165 ;
        RECT 70.895 87.865 71.065 88.035 ;
        RECT 71.655 87.865 71.825 88.995 ;
        RECT 61.265 87.125 66.610 87.670 ;
        RECT 67.705 87.295 67.965 87.800 ;
        RECT 68.160 87.675 68.825 87.845 ;
        RECT 68.145 87.125 68.475 87.505 ;
        RECT 68.655 87.295 68.825 87.675 ;
        RECT 70.005 87.125 70.295 87.850 ;
        RECT 70.470 87.295 70.725 87.865 ;
        RECT 70.895 87.695 71.825 87.865 ;
        RECT 71.995 88.655 73.005 88.825 ;
        RECT 71.995 87.855 72.165 88.655 ;
        RECT 71.650 87.660 71.825 87.695 ;
        RECT 70.895 87.125 71.225 87.525 ;
        RECT 71.650 87.295 72.180 87.660 ;
        RECT 72.370 87.635 72.645 88.455 ;
        RECT 72.365 87.465 72.645 87.635 ;
        RECT 72.370 87.295 72.645 87.465 ;
        RECT 72.815 87.295 73.005 88.655 ;
        RECT 73.175 88.670 73.345 89.335 ;
        RECT 73.515 88.915 73.685 89.675 ;
        RECT 73.920 88.915 74.435 89.325 ;
        RECT 73.175 88.480 73.925 88.670 ;
        RECT 74.095 88.105 74.435 88.915 ;
        RECT 74.665 88.535 74.875 89.675 ;
        RECT 73.205 87.935 74.435 88.105 ;
        RECT 75.045 88.525 75.375 89.505 ;
        RECT 75.545 88.535 75.775 89.675 ;
        RECT 75.985 89.240 81.330 89.675 ;
        RECT 73.185 87.125 73.695 87.660 ;
        RECT 73.915 87.330 74.160 87.935 ;
        RECT 74.665 87.125 74.875 87.945 ;
        RECT 75.045 87.925 75.295 88.525 ;
        RECT 75.465 88.115 75.795 88.365 ;
        RECT 75.045 87.295 75.375 87.925 ;
        RECT 75.545 87.125 75.775 87.945 ;
        RECT 77.570 87.670 77.910 88.500 ;
        RECT 79.390 87.990 79.740 89.240 ;
        RECT 81.505 88.585 85.015 89.675 ;
        RECT 86.195 89.005 86.365 89.505 ;
        RECT 86.535 89.175 86.865 89.675 ;
        RECT 86.195 88.835 86.860 89.005 ;
        RECT 81.505 87.895 83.155 88.415 ;
        RECT 83.325 88.065 85.015 88.585 ;
        RECT 86.110 88.015 86.460 88.665 ;
        RECT 75.985 87.125 81.330 87.670 ;
        RECT 81.505 87.125 85.015 87.895 ;
        RECT 86.630 87.845 86.860 88.835 ;
        RECT 86.195 87.675 86.860 87.845 ;
        RECT 86.195 87.385 86.365 87.675 ;
        RECT 86.535 87.125 86.865 87.505 ;
        RECT 87.035 87.385 87.260 89.505 ;
        RECT 87.475 89.175 87.805 89.675 ;
        RECT 87.975 89.005 88.145 89.505 ;
        RECT 88.380 89.290 89.210 89.460 ;
        RECT 89.450 89.295 89.830 89.675 ;
        RECT 87.450 88.835 88.145 89.005 ;
        RECT 87.450 87.865 87.620 88.835 ;
        RECT 87.790 88.045 88.200 88.665 ;
        RECT 88.370 88.615 88.870 88.995 ;
        RECT 87.450 87.675 88.145 87.865 ;
        RECT 88.370 87.745 88.590 88.615 ;
        RECT 89.040 88.445 89.210 89.290 ;
        RECT 90.010 89.125 90.180 89.415 ;
        RECT 90.350 89.295 90.680 89.675 ;
        RECT 91.150 89.205 91.780 89.455 ;
        RECT 91.960 89.295 92.380 89.675 ;
        RECT 91.610 89.125 91.780 89.205 ;
        RECT 92.580 89.125 92.820 89.415 ;
        RECT 89.380 88.875 90.750 89.125 ;
        RECT 89.380 88.615 89.630 88.875 ;
        RECT 90.140 88.445 90.390 88.605 ;
        RECT 89.040 88.275 90.390 88.445 ;
        RECT 89.040 88.235 89.460 88.275 ;
        RECT 88.770 87.685 89.120 88.055 ;
        RECT 87.475 87.125 87.805 87.505 ;
        RECT 87.975 87.345 88.145 87.675 ;
        RECT 89.290 87.505 89.460 88.235 ;
        RECT 90.560 88.105 90.750 88.875 ;
        RECT 89.630 87.775 90.040 88.105 ;
        RECT 90.330 87.765 90.750 88.105 ;
        RECT 90.920 88.695 91.440 89.005 ;
        RECT 91.610 88.955 92.820 89.125 ;
        RECT 93.050 88.985 93.380 89.675 ;
        RECT 90.920 87.935 91.090 88.695 ;
        RECT 91.260 88.105 91.440 88.515 ;
        RECT 91.610 88.445 91.780 88.955 ;
        RECT 93.550 88.805 93.720 89.415 ;
        RECT 93.990 88.955 94.320 89.465 ;
        RECT 93.550 88.785 93.870 88.805 ;
        RECT 91.950 88.615 93.870 88.785 ;
        RECT 91.610 88.275 93.510 88.445 ;
        RECT 91.840 87.935 92.170 88.055 ;
        RECT 90.920 87.765 92.170 87.935 ;
        RECT 88.445 87.305 89.460 87.505 ;
        RECT 89.630 87.125 90.040 87.565 ;
        RECT 90.330 87.335 90.580 87.765 ;
        RECT 90.780 87.125 91.100 87.585 ;
        RECT 92.340 87.515 92.510 88.275 ;
        RECT 93.180 88.215 93.510 88.275 ;
        RECT 92.700 88.045 93.030 88.105 ;
        RECT 92.700 87.775 93.360 88.045 ;
        RECT 93.680 87.720 93.870 88.615 ;
        RECT 91.660 87.345 92.510 87.515 ;
        RECT 92.710 87.125 93.370 87.605 ;
        RECT 93.550 87.390 93.870 87.720 ;
        RECT 94.070 88.365 94.320 88.955 ;
        RECT 94.500 88.875 94.785 89.675 ;
        RECT 94.965 89.335 95.220 89.365 ;
        RECT 94.965 89.165 95.305 89.335 ;
        RECT 94.965 88.695 95.220 89.165 ;
        RECT 94.070 88.035 94.870 88.365 ;
        RECT 94.070 87.385 94.320 88.035 ;
        RECT 95.040 87.835 95.220 88.695 ;
        RECT 95.765 88.510 96.055 89.675 ;
        RECT 96.225 89.240 101.570 89.675 ;
        RECT 94.500 87.125 94.785 87.585 ;
        RECT 94.965 87.305 95.220 87.835 ;
        RECT 95.765 87.125 96.055 87.850 ;
        RECT 97.810 87.670 98.150 88.500 ;
        RECT 99.630 87.990 99.980 89.240 ;
        RECT 101.745 88.585 104.335 89.675 ;
        RECT 101.745 87.895 102.955 88.415 ;
        RECT 103.125 88.065 104.335 88.585 ;
        RECT 104.965 88.955 105.425 89.505 ;
        RECT 105.615 88.955 105.945 89.675 ;
        RECT 96.225 87.125 101.570 87.670 ;
        RECT 101.745 87.125 104.335 87.895 ;
        RECT 104.965 87.585 105.215 88.955 ;
        RECT 106.145 88.785 106.445 89.335 ;
        RECT 106.615 89.005 106.895 89.675 ;
        RECT 105.505 88.615 106.445 88.785 ;
        RECT 107.265 88.955 107.725 89.505 ;
        RECT 107.915 88.955 108.245 89.675 ;
        RECT 105.505 88.365 105.675 88.615 ;
        RECT 106.815 88.365 107.080 88.725 ;
        RECT 105.385 88.035 105.675 88.365 ;
        RECT 105.845 88.115 106.185 88.365 ;
        RECT 106.405 88.115 107.080 88.365 ;
        RECT 105.505 87.945 105.675 88.035 ;
        RECT 105.505 87.755 106.895 87.945 ;
        RECT 104.965 87.295 105.525 87.585 ;
        RECT 105.695 87.125 105.945 87.585 ;
        RECT 106.565 87.395 106.895 87.755 ;
        RECT 107.265 87.585 107.515 88.955 ;
        RECT 108.445 88.785 108.745 89.335 ;
        RECT 108.915 89.005 109.195 89.675 ;
        RECT 107.805 88.615 108.745 88.785 ;
        RECT 110.575 88.745 110.745 89.505 ;
        RECT 110.925 88.915 111.255 89.675 ;
        RECT 107.805 88.365 107.975 88.615 ;
        RECT 109.115 88.365 109.380 88.725 ;
        RECT 110.575 88.575 111.240 88.745 ;
        RECT 111.425 88.600 111.695 89.505 ;
        RECT 111.955 89.005 112.125 89.505 ;
        RECT 112.295 89.175 112.625 89.675 ;
        RECT 111.955 88.835 112.620 89.005 ;
        RECT 111.070 88.430 111.240 88.575 ;
        RECT 107.685 88.035 107.975 88.365 ;
        RECT 108.145 88.115 108.485 88.365 ;
        RECT 108.705 88.115 109.380 88.365 ;
        RECT 107.805 87.945 107.975 88.035 ;
        RECT 110.505 88.025 110.835 88.395 ;
        RECT 111.070 88.100 111.355 88.430 ;
        RECT 107.805 87.755 109.195 87.945 ;
        RECT 111.070 87.845 111.240 88.100 ;
        RECT 107.265 87.295 107.825 87.585 ;
        RECT 107.995 87.125 108.245 87.585 ;
        RECT 108.865 87.395 109.195 87.755 ;
        RECT 110.575 87.675 111.240 87.845 ;
        RECT 111.525 87.800 111.695 88.600 ;
        RECT 111.870 88.015 112.220 88.665 ;
        RECT 112.390 87.845 112.620 88.835 ;
        RECT 110.575 87.295 110.745 87.675 ;
        RECT 110.925 87.125 111.255 87.505 ;
        RECT 111.435 87.295 111.695 87.800 ;
        RECT 111.955 87.675 112.620 87.845 ;
        RECT 111.955 87.385 112.125 87.675 ;
        RECT 112.295 87.125 112.625 87.505 ;
        RECT 112.795 87.385 113.020 89.505 ;
        RECT 113.235 89.175 113.565 89.675 ;
        RECT 113.735 89.005 113.905 89.505 ;
        RECT 114.140 89.290 114.970 89.460 ;
        RECT 115.210 89.295 115.590 89.675 ;
        RECT 113.210 88.835 113.905 89.005 ;
        RECT 113.210 87.865 113.380 88.835 ;
        RECT 113.550 88.045 113.960 88.665 ;
        RECT 114.130 88.615 114.630 88.995 ;
        RECT 113.210 87.675 113.905 87.865 ;
        RECT 114.130 87.745 114.350 88.615 ;
        RECT 114.800 88.445 114.970 89.290 ;
        RECT 115.770 89.125 115.940 89.415 ;
        RECT 116.110 89.295 116.440 89.675 ;
        RECT 116.910 89.205 117.540 89.455 ;
        RECT 117.720 89.295 118.140 89.675 ;
        RECT 117.370 89.125 117.540 89.205 ;
        RECT 118.340 89.125 118.580 89.415 ;
        RECT 115.140 88.875 116.510 89.125 ;
        RECT 115.140 88.615 115.390 88.875 ;
        RECT 115.900 88.445 116.150 88.605 ;
        RECT 114.800 88.275 116.150 88.445 ;
        RECT 114.800 88.235 115.220 88.275 ;
        RECT 114.530 87.685 114.880 88.055 ;
        RECT 113.235 87.125 113.565 87.505 ;
        RECT 113.735 87.345 113.905 87.675 ;
        RECT 115.050 87.505 115.220 88.235 ;
        RECT 116.320 88.105 116.510 88.875 ;
        RECT 115.390 87.775 115.800 88.105 ;
        RECT 116.090 87.765 116.510 88.105 ;
        RECT 116.680 88.695 117.200 89.005 ;
        RECT 117.370 88.955 118.580 89.125 ;
        RECT 118.810 88.985 119.140 89.675 ;
        RECT 116.680 87.935 116.850 88.695 ;
        RECT 117.020 88.105 117.200 88.515 ;
        RECT 117.370 88.445 117.540 88.955 ;
        RECT 119.310 88.805 119.480 89.415 ;
        RECT 119.750 88.955 120.080 89.465 ;
        RECT 119.310 88.785 119.630 88.805 ;
        RECT 117.710 88.615 119.630 88.785 ;
        RECT 117.370 88.275 119.270 88.445 ;
        RECT 117.600 87.935 117.930 88.055 ;
        RECT 116.680 87.765 117.930 87.935 ;
        RECT 114.205 87.305 115.220 87.505 ;
        RECT 115.390 87.125 115.800 87.565 ;
        RECT 116.090 87.335 116.340 87.765 ;
        RECT 116.540 87.125 116.860 87.585 ;
        RECT 118.100 87.515 118.270 88.275 ;
        RECT 118.940 88.215 119.270 88.275 ;
        RECT 118.460 88.045 118.790 88.105 ;
        RECT 118.460 87.775 119.120 88.045 ;
        RECT 119.440 87.720 119.630 88.615 ;
        RECT 117.420 87.345 118.270 87.515 ;
        RECT 118.470 87.125 119.130 87.605 ;
        RECT 119.310 87.390 119.630 87.720 ;
        RECT 119.830 88.365 120.080 88.955 ;
        RECT 120.260 88.875 120.545 89.675 ;
        RECT 120.725 88.695 120.980 89.365 ;
        RECT 119.830 88.035 120.630 88.365 ;
        RECT 119.830 87.385 120.080 88.035 ;
        RECT 120.800 87.835 120.980 88.695 ;
        RECT 121.525 88.510 121.815 89.675 ;
        RECT 121.985 88.600 122.255 89.505 ;
        RECT 122.425 88.915 122.755 89.675 ;
        RECT 122.935 88.745 123.105 89.505 ;
        RECT 120.725 87.635 120.980 87.835 ;
        RECT 120.260 87.125 120.545 87.585 ;
        RECT 120.725 87.465 121.065 87.635 ;
        RECT 120.725 87.305 120.980 87.465 ;
        RECT 121.525 87.125 121.815 87.850 ;
        RECT 121.985 87.800 122.155 88.600 ;
        RECT 122.440 88.575 123.105 88.745 ;
        RECT 124.285 88.585 125.495 89.675 ;
        RECT 122.440 88.430 122.610 88.575 ;
        RECT 122.325 88.100 122.610 88.430 ;
        RECT 122.440 87.845 122.610 88.100 ;
        RECT 122.845 88.025 123.175 88.395 ;
        RECT 124.285 88.045 124.805 88.585 ;
        RECT 124.975 87.875 125.495 88.415 ;
        RECT 121.985 87.295 122.245 87.800 ;
        RECT 122.440 87.675 123.105 87.845 ;
        RECT 122.425 87.125 122.755 87.505 ;
        RECT 122.935 87.295 123.105 87.675 ;
        RECT 124.285 87.125 125.495 87.875 ;
        RECT 5.520 86.955 125.580 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 6.985 86.410 12.330 86.955 ;
        RECT 12.505 86.410 17.850 86.955 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 8.570 85.580 8.910 86.410 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 10.390 84.840 10.740 86.090 ;
        RECT 14.090 85.580 14.430 86.410 ;
        RECT 18.025 86.185 21.535 86.955 ;
        RECT 21.705 86.205 22.915 86.955 ;
        RECT 23.085 86.280 23.355 86.625 ;
        RECT 23.545 86.555 23.925 86.955 ;
        RECT 24.095 86.385 24.265 86.735 ;
        RECT 24.435 86.555 24.765 86.955 ;
        RECT 24.965 86.385 25.135 86.735 ;
        RECT 25.335 86.455 25.665 86.955 ;
        RECT 25.845 86.410 31.190 86.955 ;
        RECT 15.910 84.840 16.260 86.090 ;
        RECT 18.025 85.665 19.675 86.185 ;
        RECT 19.845 85.495 21.535 86.015 ;
        RECT 21.705 85.665 22.225 86.205 ;
        RECT 22.395 85.495 22.915 86.035 ;
        RECT 6.985 84.405 12.330 84.840 ;
        RECT 12.505 84.405 17.850 84.840 ;
        RECT 18.025 84.405 21.535 85.495 ;
        RECT 21.705 84.405 22.915 85.495 ;
        RECT 23.085 85.545 23.255 86.280 ;
        RECT 23.525 86.215 25.135 86.385 ;
        RECT 23.525 86.045 23.695 86.215 ;
        RECT 23.425 85.715 23.695 86.045 ;
        RECT 23.865 85.715 24.270 86.045 ;
        RECT 23.525 85.545 23.695 85.715 ;
        RECT 23.085 84.575 23.355 85.545 ;
        RECT 23.525 85.375 24.250 85.545 ;
        RECT 24.440 85.425 25.150 86.045 ;
        RECT 25.320 85.715 25.670 86.285 ;
        RECT 27.430 85.580 27.770 86.410 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 31.825 86.410 37.170 86.955 ;
        RECT 37.345 86.410 42.690 86.955 ;
        RECT 24.080 85.255 24.250 85.375 ;
        RECT 25.350 85.255 25.670 85.545 ;
        RECT 23.565 84.405 23.845 85.205 ;
        RECT 24.080 85.085 25.670 85.255 ;
        RECT 24.015 84.625 25.670 84.915 ;
        RECT 29.250 84.840 29.600 86.090 ;
        RECT 33.410 85.580 33.750 86.410 ;
        RECT 25.845 84.405 31.190 84.840 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 35.230 84.840 35.580 86.090 ;
        RECT 38.930 85.580 39.270 86.410 ;
        RECT 42.865 86.205 44.075 86.955 ;
        RECT 40.750 84.840 41.100 86.090 ;
        RECT 42.865 85.665 43.385 86.205 ;
        RECT 44.285 86.135 44.515 86.955 ;
        RECT 44.685 86.155 45.015 86.785 ;
        RECT 43.555 85.495 44.075 86.035 ;
        RECT 44.265 85.715 44.595 85.965 ;
        RECT 44.765 85.555 45.015 86.155 ;
        RECT 45.185 86.135 45.395 86.955 ;
        RECT 45.715 86.405 45.885 86.695 ;
        RECT 46.055 86.575 46.385 86.955 ;
        RECT 45.715 86.235 46.380 86.405 ;
        RECT 31.825 84.405 37.170 84.840 ;
        RECT 37.345 84.405 42.690 84.840 ;
        RECT 42.865 84.405 44.075 85.495 ;
        RECT 44.285 84.405 44.515 85.545 ;
        RECT 44.685 84.575 45.015 85.555 ;
        RECT 45.185 84.405 45.395 85.545 ;
        RECT 45.630 85.415 45.980 86.065 ;
        RECT 46.150 85.245 46.380 86.235 ;
        RECT 45.715 85.075 46.380 85.245 ;
        RECT 45.715 84.575 45.885 85.075 ;
        RECT 46.055 84.405 46.385 84.905 ;
        RECT 46.555 84.575 46.780 86.695 ;
        RECT 46.995 86.575 47.325 86.955 ;
        RECT 47.495 86.405 47.665 86.735 ;
        RECT 47.965 86.575 48.980 86.775 ;
        RECT 46.970 86.215 47.665 86.405 ;
        RECT 46.970 85.245 47.140 86.215 ;
        RECT 47.310 85.415 47.720 86.035 ;
        RECT 47.890 85.465 48.110 86.335 ;
        RECT 48.290 86.025 48.640 86.395 ;
        RECT 48.810 85.845 48.980 86.575 ;
        RECT 49.150 86.515 49.560 86.955 ;
        RECT 49.850 86.315 50.100 86.745 ;
        RECT 50.300 86.495 50.620 86.955 ;
        RECT 51.180 86.565 52.030 86.735 ;
        RECT 49.150 85.975 49.560 86.305 ;
        RECT 49.850 85.975 50.270 86.315 ;
        RECT 48.560 85.805 48.980 85.845 ;
        RECT 48.560 85.635 49.910 85.805 ;
        RECT 46.970 85.075 47.665 85.245 ;
        RECT 47.890 85.085 48.390 85.465 ;
        RECT 46.995 84.405 47.325 84.905 ;
        RECT 47.495 84.575 47.665 85.075 ;
        RECT 48.560 84.790 48.730 85.635 ;
        RECT 49.660 85.475 49.910 85.635 ;
        RECT 48.900 85.205 49.150 85.465 ;
        RECT 50.080 85.205 50.270 85.975 ;
        RECT 48.900 84.955 50.270 85.205 ;
        RECT 50.440 86.145 51.690 86.315 ;
        RECT 50.440 85.385 50.610 86.145 ;
        RECT 51.360 86.025 51.690 86.145 ;
        RECT 50.780 85.565 50.960 85.975 ;
        RECT 51.860 85.805 52.030 86.565 ;
        RECT 52.230 86.475 52.890 86.955 ;
        RECT 53.070 86.360 53.390 86.690 ;
        RECT 52.220 86.035 52.880 86.305 ;
        RECT 52.220 85.975 52.550 86.035 ;
        RECT 52.700 85.805 53.030 85.865 ;
        RECT 51.130 85.635 53.030 85.805 ;
        RECT 50.440 85.075 50.960 85.385 ;
        RECT 51.130 85.125 51.300 85.635 ;
        RECT 53.200 85.465 53.390 86.360 ;
        RECT 51.470 85.295 53.390 85.465 ;
        RECT 53.070 85.275 53.390 85.295 ;
        RECT 53.590 86.045 53.840 86.695 ;
        RECT 54.020 86.495 54.305 86.955 ;
        RECT 54.485 86.615 54.740 86.775 ;
        RECT 54.485 86.445 54.825 86.615 ;
        RECT 54.485 86.245 54.740 86.445 ;
        RECT 53.590 85.715 54.390 86.045 ;
        RECT 51.130 84.955 52.340 85.125 ;
        RECT 47.900 84.620 48.730 84.790 ;
        RECT 48.970 84.405 49.350 84.785 ;
        RECT 49.530 84.665 49.700 84.955 ;
        RECT 51.130 84.875 51.300 84.955 ;
        RECT 49.870 84.405 50.200 84.785 ;
        RECT 50.670 84.625 51.300 84.875 ;
        RECT 51.480 84.405 51.900 84.785 ;
        RECT 52.100 84.665 52.340 84.955 ;
        RECT 52.570 84.405 52.900 85.095 ;
        RECT 53.070 84.665 53.240 85.275 ;
        RECT 53.590 85.125 53.840 85.715 ;
        RECT 54.560 85.385 54.740 86.245 ;
        RECT 55.285 86.185 56.955 86.955 ;
        RECT 57.125 86.230 57.415 86.955 ;
        RECT 55.285 85.665 56.035 86.185 ;
        RECT 57.585 86.155 57.925 86.785 ;
        RECT 58.095 86.155 58.345 86.955 ;
        RECT 58.535 86.305 58.865 86.785 ;
        RECT 59.035 86.495 59.260 86.955 ;
        RECT 59.430 86.305 59.760 86.785 ;
        RECT 56.205 85.495 56.955 86.015 ;
        RECT 53.510 84.615 53.840 85.125 ;
        RECT 54.020 84.405 54.305 85.205 ;
        RECT 54.485 84.715 54.740 85.385 ;
        RECT 55.285 84.405 56.955 85.495 ;
        RECT 57.125 84.405 57.415 85.570 ;
        RECT 57.585 85.545 57.760 86.155 ;
        RECT 58.535 86.135 59.760 86.305 ;
        RECT 60.390 86.175 60.890 86.785 ;
        RECT 61.265 86.185 62.935 86.955 ;
        RECT 57.930 85.795 58.625 85.965 ;
        RECT 58.455 85.545 58.625 85.795 ;
        RECT 58.800 85.765 59.220 85.965 ;
        RECT 59.390 85.765 59.720 85.965 ;
        RECT 59.890 85.765 60.220 85.965 ;
        RECT 60.390 85.545 60.560 86.175 ;
        RECT 60.745 85.715 61.095 85.965 ;
        RECT 61.265 85.665 62.015 86.185 ;
        RECT 63.570 86.115 63.830 86.955 ;
        RECT 64.005 86.210 64.260 86.785 ;
        RECT 64.430 86.575 64.760 86.955 ;
        RECT 64.975 86.405 65.145 86.785 ;
        RECT 65.405 86.410 70.750 86.955 ;
        RECT 70.925 86.410 76.270 86.955 ;
        RECT 64.430 86.235 65.145 86.405 ;
        RECT 57.585 84.575 57.925 85.545 ;
        RECT 58.095 84.405 58.265 85.545 ;
        RECT 58.455 85.375 60.890 85.545 ;
        RECT 62.185 85.495 62.935 86.015 ;
        RECT 58.535 84.405 58.785 85.205 ;
        RECT 59.430 84.575 59.760 85.375 ;
        RECT 60.060 84.405 60.390 85.205 ;
        RECT 60.560 84.575 60.890 85.375 ;
        RECT 61.265 84.405 62.935 85.495 ;
        RECT 63.570 84.405 63.830 85.555 ;
        RECT 64.005 85.480 64.175 86.210 ;
        RECT 64.430 86.045 64.600 86.235 ;
        RECT 64.345 85.715 64.600 86.045 ;
        RECT 64.430 85.505 64.600 85.715 ;
        RECT 64.880 85.685 65.235 86.055 ;
        RECT 66.990 85.580 67.330 86.410 ;
        RECT 64.005 84.575 64.260 85.480 ;
        RECT 64.430 85.335 65.145 85.505 ;
        RECT 64.430 84.405 64.760 85.165 ;
        RECT 64.975 84.575 65.145 85.335 ;
        RECT 68.810 84.840 69.160 86.090 ;
        RECT 72.510 85.580 72.850 86.410 ;
        RECT 76.445 86.280 76.705 86.785 ;
        RECT 76.885 86.575 77.215 86.955 ;
        RECT 77.395 86.405 77.565 86.785 ;
        RECT 74.330 84.840 74.680 86.090 ;
        RECT 76.445 85.480 76.615 86.280 ;
        RECT 76.900 86.235 77.565 86.405 ;
        RECT 76.900 85.980 77.070 86.235 ;
        RECT 77.885 86.135 78.095 86.955 ;
        RECT 78.265 86.155 78.595 86.785 ;
        RECT 76.785 85.650 77.070 85.980 ;
        RECT 77.305 85.685 77.635 86.055 ;
        RECT 76.900 85.505 77.070 85.650 ;
        RECT 78.265 85.555 78.515 86.155 ;
        RECT 78.765 86.135 78.995 86.955 ;
        RECT 79.205 86.185 82.715 86.955 ;
        RECT 82.885 86.230 83.175 86.955 ;
        RECT 83.345 86.185 86.855 86.955 ;
        RECT 87.945 86.280 88.205 86.785 ;
        RECT 88.385 86.575 88.715 86.955 ;
        RECT 88.895 86.405 89.065 86.785 ;
        RECT 78.685 85.715 79.015 85.965 ;
        RECT 79.205 85.665 80.855 86.185 ;
        RECT 65.405 84.405 70.750 84.840 ;
        RECT 70.925 84.405 76.270 84.840 ;
        RECT 76.445 84.575 76.715 85.480 ;
        RECT 76.900 85.335 77.565 85.505 ;
        RECT 76.885 84.405 77.215 85.165 ;
        RECT 77.395 84.575 77.565 85.335 ;
        RECT 77.885 84.405 78.095 85.545 ;
        RECT 78.265 84.575 78.595 85.555 ;
        RECT 78.765 84.405 78.995 85.545 ;
        RECT 81.025 85.495 82.715 86.015 ;
        RECT 83.345 85.665 84.995 86.185 ;
        RECT 79.205 84.405 82.715 85.495 ;
        RECT 82.885 84.405 83.175 85.570 ;
        RECT 85.165 85.495 86.855 86.015 ;
        RECT 83.345 84.405 86.855 85.495 ;
        RECT 87.945 85.480 88.115 86.280 ;
        RECT 88.400 86.235 89.065 86.405 ;
        RECT 88.400 85.980 88.570 86.235 ;
        RECT 89.325 86.185 91.915 86.955 ;
        RECT 88.285 85.650 88.570 85.980 ;
        RECT 88.805 85.685 89.135 86.055 ;
        RECT 89.325 85.665 90.535 86.185 ;
        RECT 92.290 86.175 92.790 86.785 ;
        RECT 88.400 85.505 88.570 85.650 ;
        RECT 87.945 84.575 88.215 85.480 ;
        RECT 88.400 85.335 89.065 85.505 ;
        RECT 90.705 85.495 91.915 86.015 ;
        RECT 92.085 85.715 92.435 85.965 ;
        RECT 92.620 85.545 92.790 86.175 ;
        RECT 93.420 86.305 93.750 86.785 ;
        RECT 93.920 86.495 94.145 86.955 ;
        RECT 94.315 86.305 94.645 86.785 ;
        RECT 93.420 86.135 94.645 86.305 ;
        RECT 94.835 86.155 95.085 86.955 ;
        RECT 95.255 86.155 95.595 86.785 ;
        RECT 95.765 86.410 101.110 86.955 ;
        RECT 102.215 86.455 102.545 86.955 ;
        RECT 95.365 86.105 95.595 86.155 ;
        RECT 92.960 85.765 93.290 85.965 ;
        RECT 93.460 85.765 93.790 85.965 ;
        RECT 93.960 85.765 94.380 85.965 ;
        RECT 94.555 85.795 95.250 85.965 ;
        RECT 94.555 85.545 94.725 85.795 ;
        RECT 95.420 85.545 95.595 86.105 ;
        RECT 97.350 85.580 97.690 86.410 ;
        RECT 102.745 86.385 102.915 86.735 ;
        RECT 103.115 86.555 103.445 86.955 ;
        RECT 103.615 86.385 103.785 86.735 ;
        RECT 103.955 86.555 104.335 86.955 ;
        RECT 88.385 84.405 88.715 85.165 ;
        RECT 88.895 84.575 89.065 85.335 ;
        RECT 89.325 84.405 91.915 85.495 ;
        RECT 92.290 85.375 94.725 85.545 ;
        RECT 92.290 84.575 92.620 85.375 ;
        RECT 92.790 84.405 93.120 85.205 ;
        RECT 93.420 84.575 93.750 85.375 ;
        RECT 94.395 84.405 94.645 85.205 ;
        RECT 94.915 84.405 95.085 85.545 ;
        RECT 95.255 84.575 95.595 85.545 ;
        RECT 99.170 84.840 99.520 86.090 ;
        RECT 102.210 85.715 102.560 86.285 ;
        RECT 102.745 86.215 104.355 86.385 ;
        RECT 104.525 86.280 104.795 86.625 ;
        RECT 104.185 86.045 104.355 86.215 ;
        RECT 102.730 85.595 103.440 86.045 ;
        RECT 103.610 85.715 104.015 86.045 ;
        RECT 104.185 85.715 104.455 86.045 ;
        RECT 102.210 85.255 102.530 85.545 ;
        RECT 102.725 85.425 103.440 85.595 ;
        RECT 104.185 85.545 104.355 85.715 ;
        RECT 104.625 85.545 104.795 86.280 ;
        RECT 103.630 85.375 104.355 85.545 ;
        RECT 103.630 85.255 103.800 85.375 ;
        RECT 102.210 85.085 103.800 85.255 ;
        RECT 95.765 84.405 101.110 84.840 ;
        RECT 102.210 84.625 103.865 84.915 ;
        RECT 104.035 84.405 104.315 85.205 ;
        RECT 104.525 84.575 104.795 85.545 ;
        RECT 104.965 86.495 105.525 86.785 ;
        RECT 105.695 86.495 105.945 86.955 ;
        RECT 104.965 85.125 105.215 86.495 ;
        RECT 106.565 86.325 106.895 86.685 ;
        RECT 105.505 86.135 106.895 86.325 ;
        RECT 107.265 86.205 108.475 86.955 ;
        RECT 108.645 86.230 108.935 86.955 ;
        RECT 105.505 86.045 105.675 86.135 ;
        RECT 105.385 85.715 105.675 86.045 ;
        RECT 105.845 85.715 106.185 85.965 ;
        RECT 106.405 85.715 107.080 85.965 ;
        RECT 105.505 85.465 105.675 85.715 ;
        RECT 105.505 85.295 106.445 85.465 ;
        RECT 106.815 85.355 107.080 85.715 ;
        RECT 107.265 85.665 107.785 86.205 ;
        RECT 109.105 86.185 112.615 86.955 ;
        RECT 112.875 86.405 113.045 86.695 ;
        RECT 113.215 86.575 113.545 86.955 ;
        RECT 112.875 86.235 113.540 86.405 ;
        RECT 107.955 85.495 108.475 86.035 ;
        RECT 109.105 85.665 110.755 86.185 ;
        RECT 104.965 84.575 105.425 85.125 ;
        RECT 105.615 84.405 105.945 85.125 ;
        RECT 106.145 84.745 106.445 85.295 ;
        RECT 106.615 84.405 106.895 85.075 ;
        RECT 107.265 84.405 108.475 85.495 ;
        RECT 108.645 84.405 108.935 85.570 ;
        RECT 110.925 85.495 112.615 86.015 ;
        RECT 109.105 84.405 112.615 85.495 ;
        RECT 112.790 85.415 113.140 86.065 ;
        RECT 113.310 85.245 113.540 86.235 ;
        RECT 112.875 85.075 113.540 85.245 ;
        RECT 112.875 84.575 113.045 85.075 ;
        RECT 113.215 84.405 113.545 84.905 ;
        RECT 113.715 84.575 113.940 86.695 ;
        RECT 114.155 86.575 114.485 86.955 ;
        RECT 114.655 86.405 114.825 86.735 ;
        RECT 115.125 86.575 116.140 86.775 ;
        RECT 114.130 86.215 114.825 86.405 ;
        RECT 114.130 85.245 114.300 86.215 ;
        RECT 114.470 85.415 114.880 86.035 ;
        RECT 115.050 85.465 115.270 86.335 ;
        RECT 115.450 86.025 115.800 86.395 ;
        RECT 115.970 85.845 116.140 86.575 ;
        RECT 116.310 86.515 116.720 86.955 ;
        RECT 117.010 86.315 117.260 86.745 ;
        RECT 117.460 86.495 117.780 86.955 ;
        RECT 118.340 86.565 119.190 86.735 ;
        RECT 116.310 85.975 116.720 86.305 ;
        RECT 117.010 85.975 117.430 86.315 ;
        RECT 115.720 85.805 116.140 85.845 ;
        RECT 115.720 85.635 117.070 85.805 ;
        RECT 114.130 85.075 114.825 85.245 ;
        RECT 115.050 85.085 115.550 85.465 ;
        RECT 114.155 84.405 114.485 84.905 ;
        RECT 114.655 84.575 114.825 85.075 ;
        RECT 115.720 84.790 115.890 85.635 ;
        RECT 116.820 85.475 117.070 85.635 ;
        RECT 116.060 85.205 116.310 85.465 ;
        RECT 117.240 85.205 117.430 85.975 ;
        RECT 116.060 84.955 117.430 85.205 ;
        RECT 117.600 86.145 118.850 86.315 ;
        RECT 117.600 85.385 117.770 86.145 ;
        RECT 118.520 86.025 118.850 86.145 ;
        RECT 117.940 85.565 118.120 85.975 ;
        RECT 119.020 85.805 119.190 86.565 ;
        RECT 119.390 86.475 120.050 86.955 ;
        RECT 120.230 86.360 120.550 86.690 ;
        RECT 119.380 86.035 120.040 86.305 ;
        RECT 119.380 85.975 119.710 86.035 ;
        RECT 119.860 85.805 120.190 85.865 ;
        RECT 118.290 85.635 120.190 85.805 ;
        RECT 117.600 85.075 118.120 85.385 ;
        RECT 118.290 85.125 118.460 85.635 ;
        RECT 120.360 85.465 120.550 86.360 ;
        RECT 118.630 85.295 120.550 85.465 ;
        RECT 120.230 85.275 120.550 85.295 ;
        RECT 120.750 86.045 121.000 86.695 ;
        RECT 121.180 86.495 121.465 86.955 ;
        RECT 121.645 86.615 121.900 86.775 ;
        RECT 121.645 86.445 121.985 86.615 ;
        RECT 121.645 86.245 121.900 86.445 ;
        RECT 120.750 85.715 121.550 86.045 ;
        RECT 118.290 84.955 119.500 85.125 ;
        RECT 115.060 84.620 115.890 84.790 ;
        RECT 116.130 84.405 116.510 84.785 ;
        RECT 116.690 84.665 116.860 84.955 ;
        RECT 118.290 84.875 118.460 84.955 ;
        RECT 117.030 84.405 117.360 84.785 ;
        RECT 117.830 84.625 118.460 84.875 ;
        RECT 118.640 84.405 119.060 84.785 ;
        RECT 119.260 84.665 119.500 84.955 ;
        RECT 119.730 84.405 120.060 85.095 ;
        RECT 120.230 84.665 120.400 85.275 ;
        RECT 120.750 85.125 121.000 85.715 ;
        RECT 121.720 85.385 121.900 86.245 ;
        RECT 122.445 86.185 124.115 86.955 ;
        RECT 124.285 86.205 125.495 86.955 ;
        RECT 122.445 85.665 123.195 86.185 ;
        RECT 123.365 85.495 124.115 86.015 ;
        RECT 120.670 84.615 121.000 85.125 ;
        RECT 121.180 84.405 121.465 85.205 ;
        RECT 121.645 84.715 121.900 85.385 ;
        RECT 122.445 84.405 124.115 85.495 ;
        RECT 124.285 85.495 124.805 86.035 ;
        RECT 124.975 85.665 125.495 86.205 ;
        RECT 124.285 84.405 125.495 85.495 ;
        RECT 5.520 84.235 125.580 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 6.985 83.800 12.330 84.235 ;
        RECT 12.505 83.800 17.850 84.235 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 8.570 82.230 8.910 83.060 ;
        RECT 10.390 82.550 10.740 83.800 ;
        RECT 14.090 82.230 14.430 83.060 ;
        RECT 15.910 82.550 16.260 83.800 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 18.945 83.145 20.615 84.235 ;
        RECT 18.945 82.455 19.695 82.975 ;
        RECT 19.865 82.625 20.615 83.145 ;
        RECT 20.990 83.265 21.320 84.065 ;
        RECT 21.490 83.435 21.820 84.235 ;
        RECT 22.120 83.265 22.450 84.065 ;
        RECT 23.095 83.435 23.345 84.235 ;
        RECT 20.990 83.095 23.425 83.265 ;
        RECT 23.615 83.095 23.785 84.235 ;
        RECT 23.955 83.095 24.295 84.065 ;
        RECT 25.590 83.265 25.920 84.065 ;
        RECT 26.090 83.435 26.420 84.235 ;
        RECT 26.720 83.265 27.050 84.065 ;
        RECT 27.695 83.435 27.945 84.235 ;
        RECT 25.590 83.095 28.025 83.265 ;
        RECT 28.215 83.095 28.385 84.235 ;
        RECT 28.555 83.095 28.895 84.065 ;
        RECT 20.785 82.675 21.135 82.925 ;
        RECT 21.320 82.465 21.490 83.095 ;
        RECT 21.660 82.675 21.990 82.875 ;
        RECT 22.160 82.675 22.490 82.875 ;
        RECT 22.660 82.675 23.080 82.875 ;
        RECT 23.255 82.845 23.425 83.095 ;
        RECT 23.255 82.675 23.950 82.845 ;
        RECT 6.985 81.685 12.330 82.230 ;
        RECT 12.505 81.685 17.850 82.230 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 18.945 81.685 20.615 82.455 ;
        RECT 20.990 81.855 21.490 82.465 ;
        RECT 22.120 82.335 23.345 82.505 ;
        RECT 24.120 82.485 24.295 83.095 ;
        RECT 25.385 82.675 25.735 82.925 ;
        RECT 22.120 81.855 22.450 82.335 ;
        RECT 22.620 81.685 22.845 82.145 ;
        RECT 23.015 81.855 23.345 82.335 ;
        RECT 23.535 81.685 23.785 82.485 ;
        RECT 23.955 81.855 24.295 82.485 ;
        RECT 25.920 82.465 26.090 83.095 ;
        RECT 26.260 82.675 26.590 82.875 ;
        RECT 26.760 82.675 27.090 82.875 ;
        RECT 27.260 82.675 27.680 82.875 ;
        RECT 27.855 82.845 28.025 83.095 ;
        RECT 27.855 82.675 28.550 82.845 ;
        RECT 25.590 81.855 26.090 82.465 ;
        RECT 26.720 82.335 27.945 82.505 ;
        RECT 28.720 82.485 28.895 83.095 ;
        RECT 26.720 81.855 27.050 82.335 ;
        RECT 27.220 81.685 27.445 82.145 ;
        RECT 27.615 81.855 27.945 82.335 ;
        RECT 28.135 81.685 28.385 82.485 ;
        RECT 28.555 81.855 28.895 82.485 ;
        RECT 29.065 83.095 29.450 84.065 ;
        RECT 29.620 83.775 29.945 84.235 ;
        RECT 30.465 83.605 30.745 84.065 ;
        RECT 29.620 83.385 30.745 83.605 ;
        RECT 29.065 82.425 29.345 83.095 ;
        RECT 29.620 82.925 30.070 83.385 ;
        RECT 30.935 83.215 31.335 84.065 ;
        RECT 31.735 83.775 32.005 84.235 ;
        RECT 32.175 83.605 32.460 84.065 ;
        RECT 29.515 82.595 30.070 82.925 ;
        RECT 30.240 82.655 31.335 83.215 ;
        RECT 29.620 82.485 30.070 82.595 ;
        RECT 29.065 81.855 29.450 82.425 ;
        RECT 29.620 82.315 30.745 82.485 ;
        RECT 29.620 81.685 29.945 82.145 ;
        RECT 30.465 81.855 30.745 82.315 ;
        RECT 30.935 81.855 31.335 82.655 ;
        RECT 31.505 83.385 32.460 83.605 ;
        RECT 32.750 83.565 33.005 84.065 ;
        RECT 33.175 83.735 33.505 84.235 ;
        RECT 32.750 83.395 33.500 83.565 ;
        RECT 31.505 82.485 31.715 83.385 ;
        RECT 31.885 82.655 32.575 83.215 ;
        RECT 32.750 82.575 33.100 83.225 ;
        RECT 31.505 82.315 32.460 82.485 ;
        RECT 33.270 82.405 33.500 83.395 ;
        RECT 31.735 81.685 32.005 82.145 ;
        RECT 32.175 81.855 32.460 82.315 ;
        RECT 32.750 82.235 33.500 82.405 ;
        RECT 32.750 81.945 33.005 82.235 ;
        RECT 33.175 81.685 33.505 82.065 ;
        RECT 33.675 81.945 33.845 84.065 ;
        RECT 34.015 83.265 34.340 84.050 ;
        RECT 34.510 83.775 34.760 84.235 ;
        RECT 34.930 83.735 35.180 84.065 ;
        RECT 35.395 83.735 36.075 84.065 ;
        RECT 34.930 83.605 35.100 83.735 ;
        RECT 34.705 83.435 35.100 83.605 ;
        RECT 34.075 82.215 34.535 83.265 ;
        RECT 34.705 82.075 34.875 83.435 ;
        RECT 35.270 83.175 35.735 83.565 ;
        RECT 35.045 82.365 35.395 82.985 ;
        RECT 35.565 82.585 35.735 83.175 ;
        RECT 35.905 82.955 36.075 83.735 ;
        RECT 36.245 83.635 36.415 83.975 ;
        RECT 36.650 83.805 36.980 84.235 ;
        RECT 37.150 83.635 37.320 83.975 ;
        RECT 37.615 83.775 37.985 84.235 ;
        RECT 36.245 83.465 37.320 83.635 ;
        RECT 38.155 83.605 38.325 84.065 ;
        RECT 38.560 83.725 39.430 84.065 ;
        RECT 39.600 83.775 39.850 84.235 ;
        RECT 37.765 83.435 38.325 83.605 ;
        RECT 37.765 83.295 37.935 83.435 ;
        RECT 36.435 83.125 37.935 83.295 ;
        RECT 38.630 83.265 39.090 83.555 ;
        RECT 35.905 82.785 37.595 82.955 ;
        RECT 35.565 82.365 35.920 82.585 ;
        RECT 36.090 82.075 36.260 82.785 ;
        RECT 36.465 82.365 37.255 82.615 ;
        RECT 37.425 82.605 37.595 82.785 ;
        RECT 37.765 82.435 37.935 83.125 ;
        RECT 34.205 81.685 34.535 82.045 ;
        RECT 34.705 81.905 35.200 82.075 ;
        RECT 35.405 81.905 36.260 82.075 ;
        RECT 37.135 81.685 37.465 82.145 ;
        RECT 37.675 82.045 37.935 82.435 ;
        RECT 38.125 83.255 39.090 83.265 ;
        RECT 39.260 83.345 39.430 83.725 ;
        RECT 40.020 83.685 40.190 83.975 ;
        RECT 40.370 83.855 40.700 84.235 ;
        RECT 40.020 83.515 40.820 83.685 ;
        RECT 38.125 83.095 38.800 83.255 ;
        RECT 39.260 83.175 40.480 83.345 ;
        RECT 38.125 82.305 38.335 83.095 ;
        RECT 39.260 83.085 39.430 83.175 ;
        RECT 38.505 82.305 38.855 82.925 ;
        RECT 39.025 82.915 39.430 83.085 ;
        RECT 39.025 82.135 39.195 82.915 ;
        RECT 39.365 82.465 39.585 82.745 ;
        RECT 39.765 82.635 40.305 83.005 ;
        RECT 40.650 82.925 40.820 83.515 ;
        RECT 41.040 83.095 41.345 84.235 ;
        RECT 41.515 83.045 41.770 83.925 ;
        RECT 42.005 83.095 42.215 84.235 ;
        RECT 40.650 82.895 41.390 82.925 ;
        RECT 39.365 82.295 39.895 82.465 ;
        RECT 37.675 81.875 38.025 82.045 ;
        RECT 38.245 81.855 39.195 82.135 ;
        RECT 39.365 81.685 39.555 82.125 ;
        RECT 39.725 82.065 39.895 82.295 ;
        RECT 40.065 82.235 40.305 82.635 ;
        RECT 40.475 82.595 41.390 82.895 ;
        RECT 40.475 82.420 40.800 82.595 ;
        RECT 40.475 82.065 40.795 82.420 ;
        RECT 41.560 82.395 41.770 83.045 ;
        RECT 42.385 83.085 42.715 84.065 ;
        RECT 42.885 83.095 43.115 84.235 ;
        RECT 39.725 81.895 40.795 82.065 ;
        RECT 41.040 81.685 41.345 82.145 ;
        RECT 41.515 81.865 41.770 82.395 ;
        RECT 42.005 81.685 42.215 82.505 ;
        RECT 42.385 82.485 42.635 83.085 ;
        RECT 44.245 83.070 44.535 84.235 ;
        RECT 44.795 83.565 44.965 84.065 ;
        RECT 45.135 83.735 45.465 84.235 ;
        RECT 44.795 83.395 45.460 83.565 ;
        RECT 42.805 82.675 43.135 82.925 ;
        RECT 44.710 82.575 45.060 83.225 ;
        RECT 42.385 81.855 42.715 82.485 ;
        RECT 42.885 81.685 43.115 82.505 ;
        RECT 44.245 81.685 44.535 82.410 ;
        RECT 45.230 82.405 45.460 83.395 ;
        RECT 44.795 82.235 45.460 82.405 ;
        RECT 44.795 81.945 44.965 82.235 ;
        RECT 45.135 81.685 45.465 82.065 ;
        RECT 45.635 81.945 45.860 84.065 ;
        RECT 46.075 83.735 46.405 84.235 ;
        RECT 46.575 83.565 46.745 84.065 ;
        RECT 46.980 83.850 47.810 84.020 ;
        RECT 48.050 83.855 48.430 84.235 ;
        RECT 46.050 83.395 46.745 83.565 ;
        RECT 46.050 82.425 46.220 83.395 ;
        RECT 46.390 82.605 46.800 83.225 ;
        RECT 46.970 83.175 47.470 83.555 ;
        RECT 46.050 82.235 46.745 82.425 ;
        RECT 46.970 82.305 47.190 83.175 ;
        RECT 47.640 83.005 47.810 83.850 ;
        RECT 48.610 83.685 48.780 83.975 ;
        RECT 48.950 83.855 49.280 84.235 ;
        RECT 49.750 83.765 50.380 84.015 ;
        RECT 50.560 83.855 50.980 84.235 ;
        RECT 50.210 83.685 50.380 83.765 ;
        RECT 51.180 83.685 51.420 83.975 ;
        RECT 47.980 83.435 49.350 83.685 ;
        RECT 47.980 83.175 48.230 83.435 ;
        RECT 48.740 83.005 48.990 83.165 ;
        RECT 47.640 82.835 48.990 83.005 ;
        RECT 47.640 82.795 48.060 82.835 ;
        RECT 47.370 82.245 47.720 82.615 ;
        RECT 46.075 81.685 46.405 82.065 ;
        RECT 46.575 81.905 46.745 82.235 ;
        RECT 47.890 82.065 48.060 82.795 ;
        RECT 49.160 82.665 49.350 83.435 ;
        RECT 48.230 82.335 48.640 82.665 ;
        RECT 48.930 82.325 49.350 82.665 ;
        RECT 49.520 83.255 50.040 83.565 ;
        RECT 50.210 83.515 51.420 83.685 ;
        RECT 51.650 83.545 51.980 84.235 ;
        RECT 49.520 82.495 49.690 83.255 ;
        RECT 49.860 82.665 50.040 83.075 ;
        RECT 50.210 83.005 50.380 83.515 ;
        RECT 52.150 83.365 52.320 83.975 ;
        RECT 52.590 83.515 52.920 84.025 ;
        RECT 52.150 83.345 52.470 83.365 ;
        RECT 50.550 83.175 52.470 83.345 ;
        RECT 50.210 82.835 52.110 83.005 ;
        RECT 50.440 82.495 50.770 82.615 ;
        RECT 49.520 82.325 50.770 82.495 ;
        RECT 47.045 81.865 48.060 82.065 ;
        RECT 48.230 81.685 48.640 82.125 ;
        RECT 48.930 81.895 49.180 82.325 ;
        RECT 49.380 81.685 49.700 82.145 ;
        RECT 50.940 82.075 51.110 82.835 ;
        RECT 51.780 82.775 52.110 82.835 ;
        RECT 51.300 82.605 51.630 82.665 ;
        RECT 51.300 82.335 51.960 82.605 ;
        RECT 52.280 82.280 52.470 83.175 ;
        RECT 50.260 81.905 51.110 82.075 ;
        RECT 51.310 81.685 51.970 82.165 ;
        RECT 52.150 81.950 52.470 82.280 ;
        RECT 52.670 82.925 52.920 83.515 ;
        RECT 53.100 83.435 53.385 84.235 ;
        RECT 53.565 83.255 53.820 83.925 ;
        RECT 53.640 83.215 53.820 83.255 ;
        RECT 53.640 83.045 53.905 83.215 ;
        RECT 54.365 83.095 54.635 84.065 ;
        RECT 54.845 83.435 55.125 84.235 ;
        RECT 55.295 83.725 56.950 84.015 ;
        RECT 55.360 83.385 56.950 83.555 ;
        RECT 55.360 83.265 55.530 83.385 ;
        RECT 54.805 83.095 55.530 83.265 ;
        RECT 52.670 82.595 53.470 82.925 ;
        RECT 52.670 81.945 52.920 82.595 ;
        RECT 53.640 82.395 53.820 83.045 ;
        RECT 53.100 81.685 53.385 82.145 ;
        RECT 53.565 81.865 53.820 82.395 ;
        RECT 54.365 82.360 54.535 83.095 ;
        RECT 54.805 82.925 54.975 83.095 ;
        RECT 55.720 83.045 56.435 83.215 ;
        RECT 56.630 83.095 56.950 83.385 ;
        RECT 57.125 83.145 58.795 84.235 ;
        RECT 59.480 83.365 59.765 84.235 ;
        RECT 59.935 83.605 60.195 84.065 ;
        RECT 60.370 83.775 60.625 84.235 ;
        RECT 60.795 83.605 61.055 84.065 ;
        RECT 59.935 83.435 61.055 83.605 ;
        RECT 61.225 83.435 61.535 84.235 ;
        RECT 59.935 83.185 60.195 83.435 ;
        RECT 60.405 83.385 60.575 83.435 ;
        RECT 61.705 83.265 62.015 84.065 ;
        RECT 54.705 82.595 54.975 82.925 ;
        RECT 55.145 82.595 55.550 82.925 ;
        RECT 55.720 82.595 56.430 83.045 ;
        RECT 54.805 82.425 54.975 82.595 ;
        RECT 54.365 82.015 54.635 82.360 ;
        RECT 54.805 82.255 56.415 82.425 ;
        RECT 56.600 82.355 56.950 82.925 ;
        RECT 57.125 82.455 57.875 82.975 ;
        RECT 58.045 82.625 58.795 83.145 ;
        RECT 59.440 83.015 60.195 83.185 ;
        RECT 60.985 83.095 62.015 83.265 ;
        RECT 59.440 82.505 59.845 83.015 ;
        RECT 60.985 82.845 61.155 83.095 ;
        RECT 60.015 82.675 61.155 82.845 ;
        RECT 54.825 81.685 55.205 82.085 ;
        RECT 55.375 81.905 55.545 82.255 ;
        RECT 55.715 81.685 56.045 82.085 ;
        RECT 56.245 81.905 56.415 82.255 ;
        RECT 56.615 81.685 56.945 82.185 ;
        RECT 57.125 81.685 58.795 82.455 ;
        RECT 59.440 82.335 61.090 82.505 ;
        RECT 61.325 82.355 61.675 82.925 ;
        RECT 59.485 81.685 59.765 82.165 ;
        RECT 59.935 81.945 60.195 82.335 ;
        RECT 60.370 81.685 60.625 82.165 ;
        RECT 60.795 81.945 61.090 82.335 ;
        RECT 61.845 82.185 62.015 83.095 ;
        RECT 63.110 83.085 63.370 84.235 ;
        RECT 63.545 83.160 63.800 84.065 ;
        RECT 63.970 83.475 64.300 84.235 ;
        RECT 64.515 83.305 64.685 84.065 ;
        RECT 61.270 81.685 61.545 82.165 ;
        RECT 61.715 81.855 62.015 82.185 ;
        RECT 63.110 81.685 63.370 82.525 ;
        RECT 63.545 82.430 63.715 83.160 ;
        RECT 63.970 83.135 64.685 83.305 ;
        RECT 65.405 83.265 65.715 84.065 ;
        RECT 65.885 83.435 66.195 84.235 ;
        RECT 66.365 83.605 66.625 84.065 ;
        RECT 66.795 83.775 67.050 84.235 ;
        RECT 67.225 83.605 67.485 84.065 ;
        RECT 66.365 83.435 67.485 83.605 ;
        RECT 63.970 82.925 64.140 83.135 ;
        RECT 65.405 83.095 66.435 83.265 ;
        RECT 63.885 82.595 64.140 82.925 ;
        RECT 63.545 81.855 63.800 82.430 ;
        RECT 63.970 82.405 64.140 82.595 ;
        RECT 64.420 82.585 64.775 82.955 ;
        RECT 63.970 82.235 64.685 82.405 ;
        RECT 63.970 81.685 64.300 82.065 ;
        RECT 64.515 81.855 64.685 82.235 ;
        RECT 65.405 82.185 65.575 83.095 ;
        RECT 65.745 82.355 66.095 82.925 ;
        RECT 66.265 82.845 66.435 83.095 ;
        RECT 67.225 83.185 67.485 83.435 ;
        RECT 67.655 83.365 67.940 84.235 ;
        RECT 68.255 83.305 68.425 84.065 ;
        RECT 68.640 83.475 68.970 84.235 ;
        RECT 67.225 83.015 67.980 83.185 ;
        RECT 68.255 83.135 68.970 83.305 ;
        RECT 69.140 83.160 69.395 84.065 ;
        RECT 66.265 82.675 67.405 82.845 ;
        RECT 67.575 82.505 67.980 83.015 ;
        RECT 68.165 82.585 68.520 82.955 ;
        RECT 68.800 82.925 68.970 83.135 ;
        RECT 68.800 82.595 69.055 82.925 ;
        RECT 66.330 82.335 67.980 82.505 ;
        RECT 68.800 82.405 68.970 82.595 ;
        RECT 69.225 82.430 69.395 83.160 ;
        RECT 69.570 83.085 69.830 84.235 ;
        RECT 70.005 83.070 70.295 84.235 ;
        RECT 70.465 83.385 70.725 84.065 ;
        RECT 70.895 83.455 71.145 84.235 ;
        RECT 71.395 83.685 71.645 84.065 ;
        RECT 71.815 83.855 72.170 84.235 ;
        RECT 73.175 83.845 73.510 84.065 ;
        RECT 72.775 83.685 73.005 83.725 ;
        RECT 71.395 83.485 73.005 83.685 ;
        RECT 71.395 83.475 72.230 83.485 ;
        RECT 72.820 83.395 73.005 83.485 ;
        RECT 65.405 81.855 65.705 82.185 ;
        RECT 65.875 81.685 66.150 82.165 ;
        RECT 66.330 81.945 66.625 82.335 ;
        RECT 66.795 81.685 67.050 82.165 ;
        RECT 67.225 81.945 67.485 82.335 ;
        RECT 68.255 82.235 68.970 82.405 ;
        RECT 67.655 81.685 67.935 82.165 ;
        RECT 68.255 81.855 68.425 82.235 ;
        RECT 68.640 81.685 68.970 82.065 ;
        RECT 69.140 81.855 69.395 82.430 ;
        RECT 69.570 81.685 69.830 82.525 ;
        RECT 70.005 81.685 70.295 82.410 ;
        RECT 70.465 82.195 70.635 83.385 ;
        RECT 72.335 83.285 72.665 83.315 ;
        RECT 70.865 83.225 72.665 83.285 ;
        RECT 73.255 83.225 73.510 83.845 ;
        RECT 70.805 83.115 73.510 83.225 ;
        RECT 70.805 83.080 71.005 83.115 ;
        RECT 70.805 82.505 70.975 83.080 ;
        RECT 72.335 83.055 73.510 83.115 ;
        RECT 73.745 83.095 73.955 84.235 ;
        RECT 74.125 83.085 74.455 84.065 ;
        RECT 74.625 83.095 74.855 84.235 ;
        RECT 75.525 83.095 75.910 84.065 ;
        RECT 76.080 83.775 76.405 84.235 ;
        RECT 76.925 83.605 77.205 84.065 ;
        RECT 76.080 83.385 77.205 83.605 ;
        RECT 71.205 82.640 71.615 82.945 ;
        RECT 71.785 82.675 72.115 82.885 ;
        RECT 70.805 82.385 71.075 82.505 ;
        RECT 70.805 82.340 71.650 82.385 ;
        RECT 70.895 82.215 71.650 82.340 ;
        RECT 71.905 82.275 72.115 82.675 ;
        RECT 72.360 82.675 72.835 82.885 ;
        RECT 73.025 82.675 73.515 82.875 ;
        RECT 72.360 82.275 72.580 82.675 ;
        RECT 70.465 82.185 70.695 82.195 ;
        RECT 70.465 81.855 70.725 82.185 ;
        RECT 71.480 82.065 71.650 82.215 ;
        RECT 70.895 81.685 71.225 82.045 ;
        RECT 71.480 81.855 72.780 82.065 ;
        RECT 73.055 81.685 73.510 82.450 ;
        RECT 73.745 81.685 73.955 82.505 ;
        RECT 74.125 82.485 74.375 83.085 ;
        RECT 74.545 82.675 74.875 82.925 ;
        RECT 74.125 81.855 74.455 82.485 ;
        RECT 74.625 81.685 74.855 82.505 ;
        RECT 75.525 82.425 75.805 83.095 ;
        RECT 76.080 82.925 76.530 83.385 ;
        RECT 77.395 83.215 77.795 84.065 ;
        RECT 78.195 83.775 78.465 84.235 ;
        RECT 78.635 83.605 78.920 84.065 ;
        RECT 75.975 82.595 76.530 82.925 ;
        RECT 76.700 82.655 77.795 83.215 ;
        RECT 76.080 82.485 76.530 82.595 ;
        RECT 75.525 81.855 75.910 82.425 ;
        RECT 76.080 82.315 77.205 82.485 ;
        RECT 76.080 81.685 76.405 82.145 ;
        RECT 76.925 81.855 77.205 82.315 ;
        RECT 77.395 81.855 77.795 82.655 ;
        RECT 77.965 83.385 78.920 83.605 ;
        RECT 77.965 82.485 78.175 83.385 ;
        RECT 80.330 83.265 80.660 84.065 ;
        RECT 80.830 83.435 81.160 84.235 ;
        RECT 81.460 83.265 81.790 84.065 ;
        RECT 82.435 83.435 82.685 84.235 ;
        RECT 78.345 82.655 79.035 83.215 ;
        RECT 80.330 83.095 82.765 83.265 ;
        RECT 82.955 83.095 83.125 84.235 ;
        RECT 83.295 83.095 83.635 84.065 ;
        RECT 83.805 83.145 85.475 84.235 ;
        RECT 86.195 83.565 86.365 84.065 ;
        RECT 86.535 83.735 86.865 84.235 ;
        RECT 86.195 83.395 86.860 83.565 ;
        RECT 80.125 82.675 80.475 82.925 ;
        RECT 77.965 82.315 78.920 82.485 ;
        RECT 80.660 82.465 80.830 83.095 ;
        RECT 81.000 82.675 81.330 82.875 ;
        RECT 81.500 82.675 81.830 82.875 ;
        RECT 82.000 82.675 82.420 82.875 ;
        RECT 82.595 82.845 82.765 83.095 ;
        RECT 82.595 82.675 83.290 82.845 ;
        RECT 78.195 81.685 78.465 82.145 ;
        RECT 78.635 81.855 78.920 82.315 ;
        RECT 80.330 81.855 80.830 82.465 ;
        RECT 81.460 82.335 82.685 82.505 ;
        RECT 83.460 82.485 83.635 83.095 ;
        RECT 81.460 81.855 81.790 82.335 ;
        RECT 81.960 81.685 82.185 82.145 ;
        RECT 82.355 81.855 82.685 82.335 ;
        RECT 82.875 81.685 83.125 82.485 ;
        RECT 83.295 81.855 83.635 82.485 ;
        RECT 83.805 82.455 84.555 82.975 ;
        RECT 84.725 82.625 85.475 83.145 ;
        RECT 86.110 82.575 86.460 83.225 ;
        RECT 83.805 81.685 85.475 82.455 ;
        RECT 86.630 82.405 86.860 83.395 ;
        RECT 86.195 82.235 86.860 82.405 ;
        RECT 86.195 81.945 86.365 82.235 ;
        RECT 86.535 81.685 86.865 82.065 ;
        RECT 87.035 81.945 87.260 84.065 ;
        RECT 87.475 83.735 87.805 84.235 ;
        RECT 87.975 83.565 88.145 84.065 ;
        RECT 88.380 83.850 89.210 84.020 ;
        RECT 89.450 83.855 89.830 84.235 ;
        RECT 87.450 83.395 88.145 83.565 ;
        RECT 87.450 82.425 87.620 83.395 ;
        RECT 87.790 82.605 88.200 83.225 ;
        RECT 88.370 83.175 88.870 83.555 ;
        RECT 87.450 82.235 88.145 82.425 ;
        RECT 88.370 82.305 88.590 83.175 ;
        RECT 89.040 83.005 89.210 83.850 ;
        RECT 90.010 83.685 90.180 83.975 ;
        RECT 90.350 83.855 90.680 84.235 ;
        RECT 91.150 83.765 91.780 84.015 ;
        RECT 91.960 83.855 92.380 84.235 ;
        RECT 91.610 83.685 91.780 83.765 ;
        RECT 92.580 83.685 92.820 83.975 ;
        RECT 89.380 83.435 90.750 83.685 ;
        RECT 89.380 83.175 89.630 83.435 ;
        RECT 90.140 83.005 90.390 83.165 ;
        RECT 89.040 82.835 90.390 83.005 ;
        RECT 89.040 82.795 89.460 82.835 ;
        RECT 88.770 82.245 89.120 82.615 ;
        RECT 87.475 81.685 87.805 82.065 ;
        RECT 87.975 81.905 88.145 82.235 ;
        RECT 89.290 82.065 89.460 82.795 ;
        RECT 90.560 82.665 90.750 83.435 ;
        RECT 89.630 82.335 90.040 82.665 ;
        RECT 90.330 82.325 90.750 82.665 ;
        RECT 90.920 83.255 91.440 83.565 ;
        RECT 91.610 83.515 92.820 83.685 ;
        RECT 93.050 83.545 93.380 84.235 ;
        RECT 90.920 82.495 91.090 83.255 ;
        RECT 91.260 82.665 91.440 83.075 ;
        RECT 91.610 83.005 91.780 83.515 ;
        RECT 93.550 83.365 93.720 83.975 ;
        RECT 93.990 83.515 94.320 84.025 ;
        RECT 93.550 83.345 93.870 83.365 ;
        RECT 91.950 83.175 93.870 83.345 ;
        RECT 91.610 82.835 93.510 83.005 ;
        RECT 91.840 82.495 92.170 82.615 ;
        RECT 90.920 82.325 92.170 82.495 ;
        RECT 88.445 81.865 89.460 82.065 ;
        RECT 89.630 81.685 90.040 82.125 ;
        RECT 90.330 81.895 90.580 82.325 ;
        RECT 90.780 81.685 91.100 82.145 ;
        RECT 92.340 82.075 92.510 82.835 ;
        RECT 93.180 82.775 93.510 82.835 ;
        RECT 92.700 82.605 93.030 82.665 ;
        RECT 92.700 82.335 93.360 82.605 ;
        RECT 93.680 82.280 93.870 83.175 ;
        RECT 91.660 81.905 92.510 82.075 ;
        RECT 92.710 81.685 93.370 82.165 ;
        RECT 93.550 81.950 93.870 82.280 ;
        RECT 94.070 82.925 94.320 83.515 ;
        RECT 94.500 83.435 94.785 84.235 ;
        RECT 94.965 83.255 95.220 83.925 ;
        RECT 94.070 82.595 94.870 82.925 ;
        RECT 94.070 81.945 94.320 82.595 ;
        RECT 95.040 82.395 95.220 83.255 ;
        RECT 95.765 83.070 96.055 84.235 ;
        RECT 96.430 83.265 96.760 84.065 ;
        RECT 96.930 83.435 97.260 84.235 ;
        RECT 97.560 83.265 97.890 84.065 ;
        RECT 98.535 83.435 98.785 84.235 ;
        RECT 96.430 83.095 98.865 83.265 ;
        RECT 99.055 83.095 99.225 84.235 ;
        RECT 99.395 83.095 99.735 84.065 ;
        RECT 99.905 83.145 101.575 84.235 ;
        RECT 102.210 83.725 103.865 84.015 ;
        RECT 96.225 82.675 96.575 82.925 ;
        RECT 96.760 82.465 96.930 83.095 ;
        RECT 97.100 82.675 97.430 82.875 ;
        RECT 97.600 82.675 97.930 82.875 ;
        RECT 98.100 82.675 98.520 82.875 ;
        RECT 98.695 82.845 98.865 83.095 ;
        RECT 98.695 82.675 99.390 82.845 ;
        RECT 99.560 82.535 99.735 83.095 ;
        RECT 94.965 82.195 95.220 82.395 ;
        RECT 94.500 81.685 94.785 82.145 ;
        RECT 94.965 82.025 95.305 82.195 ;
        RECT 94.965 81.865 95.220 82.025 ;
        RECT 95.765 81.685 96.055 82.410 ;
        RECT 96.430 81.855 96.930 82.465 ;
        RECT 97.560 82.335 98.785 82.505 ;
        RECT 99.505 82.485 99.735 82.535 ;
        RECT 97.560 81.855 97.890 82.335 ;
        RECT 98.060 81.685 98.285 82.145 ;
        RECT 98.455 81.855 98.785 82.335 ;
        RECT 98.975 81.685 99.225 82.485 ;
        RECT 99.395 81.855 99.735 82.485 ;
        RECT 99.905 82.455 100.655 82.975 ;
        RECT 100.825 82.625 101.575 83.145 ;
        RECT 102.210 83.385 103.800 83.555 ;
        RECT 104.035 83.435 104.315 84.235 ;
        RECT 102.210 83.095 102.530 83.385 ;
        RECT 103.630 83.265 103.800 83.385 ;
        RECT 99.905 81.685 101.575 82.455 ;
        RECT 102.210 82.355 102.560 82.925 ;
        RECT 102.730 82.595 103.440 83.215 ;
        RECT 103.630 83.095 104.355 83.265 ;
        RECT 104.525 83.095 104.795 84.065 ;
        RECT 104.970 83.725 106.625 84.015 ;
        RECT 104.970 83.385 106.560 83.555 ;
        RECT 106.795 83.435 107.075 84.235 ;
        RECT 104.970 83.095 105.290 83.385 ;
        RECT 106.390 83.265 106.560 83.385 ;
        RECT 104.185 82.925 104.355 83.095 ;
        RECT 103.610 82.595 104.015 82.925 ;
        RECT 104.185 82.595 104.455 82.925 ;
        RECT 104.185 82.425 104.355 82.595 ;
        RECT 102.745 82.255 104.355 82.425 ;
        RECT 104.625 82.360 104.795 83.095 ;
        RECT 102.215 81.685 102.545 82.185 ;
        RECT 102.745 81.905 102.915 82.255 ;
        RECT 103.115 81.685 103.445 82.085 ;
        RECT 103.615 81.905 103.785 82.255 ;
        RECT 103.955 81.685 104.335 82.085 ;
        RECT 104.525 82.015 104.795 82.360 ;
        RECT 104.970 82.355 105.320 82.925 ;
        RECT 105.490 82.595 106.200 83.215 ;
        RECT 106.390 83.095 107.115 83.265 ;
        RECT 107.285 83.095 107.555 84.065 ;
        RECT 107.725 83.800 113.070 84.235 ;
        RECT 106.945 82.925 107.115 83.095 ;
        RECT 106.370 82.595 106.775 82.925 ;
        RECT 106.945 82.595 107.215 82.925 ;
        RECT 106.945 82.425 107.115 82.595 ;
        RECT 105.505 82.255 107.115 82.425 ;
        RECT 107.385 82.360 107.555 83.095 ;
        RECT 104.975 81.685 105.305 82.185 ;
        RECT 105.505 81.905 105.675 82.255 ;
        RECT 105.875 81.685 106.205 82.085 ;
        RECT 106.375 81.905 106.545 82.255 ;
        RECT 106.715 81.685 107.095 82.085 ;
        RECT 107.285 82.015 107.555 82.360 ;
        RECT 109.310 82.230 109.650 83.060 ;
        RECT 111.130 82.550 111.480 83.800 ;
        RECT 113.245 83.145 116.755 84.235 ;
        RECT 113.245 82.455 114.895 82.975 ;
        RECT 115.065 82.625 116.755 83.145 ;
        RECT 117.445 83.095 117.655 84.235 ;
        RECT 117.825 83.085 118.155 84.065 ;
        RECT 118.325 83.095 118.555 84.235 ;
        RECT 118.765 83.145 121.355 84.235 ;
        RECT 107.725 81.685 113.070 82.230 ;
        RECT 113.245 81.685 116.755 82.455 ;
        RECT 117.445 81.685 117.655 82.505 ;
        RECT 117.825 82.485 118.075 83.085 ;
        RECT 118.245 82.675 118.575 82.925 ;
        RECT 117.825 81.855 118.155 82.485 ;
        RECT 118.325 81.685 118.555 82.505 ;
        RECT 118.765 82.455 119.975 82.975 ;
        RECT 120.145 82.625 121.355 83.145 ;
        RECT 121.525 83.070 121.815 84.235 ;
        RECT 121.985 83.145 123.655 84.235 ;
        RECT 121.985 82.455 122.735 82.975 ;
        RECT 122.905 82.625 123.655 83.145 ;
        RECT 124.285 83.145 125.495 84.235 ;
        RECT 124.285 82.605 124.805 83.145 ;
        RECT 118.765 81.685 121.355 82.455 ;
        RECT 121.525 81.685 121.815 82.410 ;
        RECT 121.985 81.685 123.655 82.455 ;
        RECT 124.975 82.435 125.495 82.975 ;
        RECT 124.285 81.685 125.495 82.435 ;
        RECT 5.520 81.515 125.580 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.985 80.745 8.655 81.515 ;
        RECT 8.825 80.840 9.085 81.345 ;
        RECT 9.265 81.135 9.595 81.515 ;
        RECT 9.775 80.965 9.945 81.345 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 6.985 80.225 7.735 80.745 ;
        RECT 7.905 80.055 8.655 80.575 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 6.985 78.965 8.655 80.055 ;
        RECT 8.825 80.040 8.995 80.840 ;
        RECT 9.280 80.795 9.945 80.965 ;
        RECT 10.205 80.840 10.465 81.345 ;
        RECT 10.645 81.135 10.975 81.515 ;
        RECT 11.155 80.965 11.325 81.345 ;
        RECT 9.280 80.540 9.450 80.795 ;
        RECT 9.165 80.210 9.450 80.540 ;
        RECT 9.685 80.245 10.015 80.615 ;
        RECT 9.280 80.065 9.450 80.210 ;
        RECT 8.825 79.135 9.095 80.040 ;
        RECT 9.280 79.895 9.945 80.065 ;
        RECT 9.265 78.965 9.595 79.725 ;
        RECT 9.775 79.135 9.945 79.895 ;
        RECT 10.205 80.040 10.375 80.840 ;
        RECT 10.660 80.795 11.325 80.965 ;
        RECT 10.660 80.540 10.830 80.795 ;
        RECT 11.590 80.775 11.845 81.345 ;
        RECT 12.015 81.115 12.345 81.515 ;
        RECT 12.770 80.980 13.300 81.345 ;
        RECT 12.770 80.945 12.945 80.980 ;
        RECT 12.015 80.775 12.945 80.945 ;
        RECT 13.490 80.835 13.765 81.345 ;
        RECT 10.545 80.210 10.830 80.540 ;
        RECT 11.065 80.245 11.395 80.615 ;
        RECT 10.660 80.065 10.830 80.210 ;
        RECT 11.590 80.105 11.760 80.775 ;
        RECT 12.015 80.605 12.185 80.775 ;
        RECT 11.930 80.275 12.185 80.605 ;
        RECT 12.410 80.275 12.605 80.605 ;
        RECT 10.205 79.135 10.475 80.040 ;
        RECT 10.660 79.895 11.325 80.065 ;
        RECT 10.645 78.965 10.975 79.725 ;
        RECT 11.155 79.135 11.325 79.895 ;
        RECT 11.590 79.135 11.925 80.105 ;
        RECT 12.095 78.965 12.265 80.105 ;
        RECT 12.435 79.305 12.605 80.275 ;
        RECT 12.775 79.645 12.945 80.775 ;
        RECT 13.115 79.985 13.285 80.785 ;
        RECT 13.485 80.665 13.765 80.835 ;
        RECT 13.490 80.185 13.765 80.665 ;
        RECT 13.935 79.985 14.125 81.345 ;
        RECT 14.305 80.980 14.815 81.515 ;
        RECT 15.035 80.705 15.280 81.310 ;
        RECT 15.730 80.775 15.985 81.345 ;
        RECT 16.155 81.115 16.485 81.515 ;
        RECT 16.910 80.980 17.440 81.345 ;
        RECT 17.630 81.175 17.905 81.345 ;
        RECT 17.625 81.005 17.905 81.175 ;
        RECT 16.910 80.945 17.085 80.980 ;
        RECT 16.155 80.775 17.085 80.945 ;
        RECT 14.325 80.535 15.555 80.705 ;
        RECT 13.115 79.815 14.125 79.985 ;
        RECT 14.295 79.970 15.045 80.160 ;
        RECT 12.775 79.475 13.900 79.645 ;
        RECT 14.295 79.305 14.465 79.970 ;
        RECT 15.215 79.725 15.555 80.535 ;
        RECT 12.435 79.135 14.465 79.305 ;
        RECT 14.635 78.965 14.805 79.725 ;
        RECT 15.040 79.315 15.555 79.725 ;
        RECT 15.730 80.105 15.900 80.775 ;
        RECT 16.155 80.605 16.325 80.775 ;
        RECT 16.070 80.275 16.325 80.605 ;
        RECT 16.550 80.275 16.745 80.605 ;
        RECT 15.730 79.135 16.065 80.105 ;
        RECT 16.235 78.965 16.405 80.105 ;
        RECT 16.575 79.305 16.745 80.275 ;
        RECT 16.915 79.645 17.085 80.775 ;
        RECT 17.255 79.985 17.425 80.785 ;
        RECT 17.630 80.185 17.905 81.005 ;
        RECT 18.075 79.985 18.265 81.345 ;
        RECT 18.445 80.980 18.955 81.515 ;
        RECT 19.175 80.705 19.420 81.310 ;
        RECT 19.865 80.765 21.075 81.515 ;
        RECT 18.465 80.535 19.695 80.705 ;
        RECT 17.255 79.815 18.265 79.985 ;
        RECT 18.435 79.970 19.185 80.160 ;
        RECT 16.915 79.475 18.040 79.645 ;
        RECT 18.435 79.305 18.605 79.970 ;
        RECT 19.355 79.725 19.695 80.535 ;
        RECT 19.865 80.225 20.385 80.765 ;
        RECT 21.450 80.735 21.950 81.345 ;
        RECT 20.555 80.055 21.075 80.595 ;
        RECT 21.245 80.275 21.595 80.525 ;
        RECT 21.780 80.105 21.950 80.735 ;
        RECT 22.580 80.865 22.910 81.345 ;
        RECT 23.080 81.055 23.305 81.515 ;
        RECT 23.475 80.865 23.805 81.345 ;
        RECT 22.580 80.695 23.805 80.865 ;
        RECT 23.995 80.715 24.245 81.515 ;
        RECT 24.415 80.715 24.755 81.345 ;
        RECT 24.935 81.015 25.265 81.515 ;
        RECT 25.465 80.945 25.635 81.295 ;
        RECT 25.835 81.115 26.165 81.515 ;
        RECT 26.335 80.945 26.505 81.295 ;
        RECT 26.675 81.115 27.055 81.515 ;
        RECT 24.525 80.665 24.755 80.715 ;
        RECT 22.120 80.325 22.450 80.525 ;
        RECT 22.620 80.325 22.950 80.525 ;
        RECT 23.120 80.325 23.540 80.525 ;
        RECT 23.715 80.355 24.410 80.525 ;
        RECT 23.715 80.105 23.885 80.355 ;
        RECT 24.580 80.105 24.755 80.665 ;
        RECT 24.930 80.275 25.280 80.845 ;
        RECT 25.465 80.775 27.075 80.945 ;
        RECT 27.245 80.840 27.515 81.185 ;
        RECT 26.905 80.605 27.075 80.775 ;
        RECT 16.575 79.135 18.605 79.305 ;
        RECT 18.775 78.965 18.945 79.725 ;
        RECT 19.180 79.315 19.695 79.725 ;
        RECT 19.865 78.965 21.075 80.055 ;
        RECT 21.450 79.935 23.885 80.105 ;
        RECT 21.450 79.135 21.780 79.935 ;
        RECT 21.950 78.965 22.280 79.765 ;
        RECT 22.580 79.135 22.910 79.935 ;
        RECT 23.555 78.965 23.805 79.765 ;
        RECT 24.075 78.965 24.245 80.105 ;
        RECT 24.415 79.135 24.755 80.105 ;
        RECT 24.930 79.815 25.250 80.105 ;
        RECT 25.450 79.985 26.160 80.605 ;
        RECT 26.330 80.275 26.735 80.605 ;
        RECT 26.905 80.275 27.175 80.605 ;
        RECT 26.905 80.105 27.075 80.275 ;
        RECT 27.345 80.105 27.515 80.840 ;
        RECT 26.350 79.935 27.075 80.105 ;
        RECT 26.350 79.815 26.520 79.935 ;
        RECT 24.930 79.645 26.520 79.815 ;
        RECT 24.930 79.185 26.585 79.475 ;
        RECT 26.755 78.965 27.035 79.765 ;
        RECT 27.245 79.135 27.515 80.105 ;
        RECT 27.685 80.840 27.955 81.185 ;
        RECT 28.145 81.115 28.525 81.515 ;
        RECT 28.695 80.945 28.865 81.295 ;
        RECT 29.035 81.115 29.365 81.515 ;
        RECT 29.565 80.945 29.735 81.295 ;
        RECT 29.935 81.015 30.265 81.515 ;
        RECT 27.685 80.105 27.855 80.840 ;
        RECT 28.125 80.775 29.735 80.945 ;
        RECT 28.125 80.605 28.295 80.775 ;
        RECT 28.025 80.275 28.295 80.605 ;
        RECT 28.465 80.275 28.870 80.605 ;
        RECT 28.125 80.105 28.295 80.275 ;
        RECT 27.685 79.135 27.955 80.105 ;
        RECT 28.125 79.935 28.850 80.105 ;
        RECT 29.040 79.985 29.750 80.605 ;
        RECT 29.920 80.275 30.270 80.845 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 31.825 80.745 35.335 81.515 ;
        RECT 35.505 80.840 35.765 81.345 ;
        RECT 35.945 81.135 36.275 81.515 ;
        RECT 36.455 80.965 36.625 81.345 ;
        RECT 31.825 80.225 33.475 80.745 ;
        RECT 28.680 79.815 28.850 79.935 ;
        RECT 29.950 79.815 30.270 80.105 ;
        RECT 28.165 78.965 28.445 79.765 ;
        RECT 28.680 79.645 30.270 79.815 ;
        RECT 28.615 79.185 30.270 79.475 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 33.645 80.055 35.335 80.575 ;
        RECT 31.825 78.965 35.335 80.055 ;
        RECT 35.505 80.040 35.675 80.840 ;
        RECT 35.960 80.795 36.625 80.965 ;
        RECT 35.960 80.540 36.130 80.795 ;
        RECT 37.350 80.775 37.605 81.345 ;
        RECT 37.775 81.115 38.105 81.515 ;
        RECT 38.530 80.980 39.060 81.345 ;
        RECT 39.250 81.175 39.525 81.345 ;
        RECT 39.245 81.005 39.525 81.175 ;
        RECT 38.530 80.945 38.705 80.980 ;
        RECT 37.775 80.775 38.705 80.945 ;
        RECT 35.845 80.210 36.130 80.540 ;
        RECT 36.365 80.245 36.695 80.615 ;
        RECT 35.960 80.065 36.130 80.210 ;
        RECT 37.350 80.105 37.520 80.775 ;
        RECT 37.775 80.605 37.945 80.775 ;
        RECT 37.690 80.275 37.945 80.605 ;
        RECT 38.170 80.275 38.365 80.605 ;
        RECT 35.505 79.135 35.775 80.040 ;
        RECT 35.960 79.895 36.625 80.065 ;
        RECT 35.945 78.965 36.275 79.725 ;
        RECT 36.455 79.135 36.625 79.895 ;
        RECT 37.350 79.135 37.685 80.105 ;
        RECT 37.855 78.965 38.025 80.105 ;
        RECT 38.195 79.305 38.365 80.275 ;
        RECT 38.535 79.645 38.705 80.775 ;
        RECT 38.875 79.985 39.045 80.785 ;
        RECT 39.250 80.185 39.525 81.005 ;
        RECT 39.695 79.985 39.885 81.345 ;
        RECT 40.065 80.980 40.575 81.515 ;
        RECT 40.795 80.705 41.040 81.310 ;
        RECT 41.485 80.970 46.830 81.515 ;
        RECT 40.085 80.535 41.315 80.705 ;
        RECT 38.875 79.815 39.885 79.985 ;
        RECT 40.055 79.970 40.805 80.160 ;
        RECT 38.535 79.475 39.660 79.645 ;
        RECT 40.055 79.305 40.225 79.970 ;
        RECT 40.975 79.725 41.315 80.535 ;
        RECT 43.070 80.140 43.410 80.970 ;
        RECT 47.965 80.695 48.195 81.515 ;
        RECT 48.365 80.715 48.695 81.345 ;
        RECT 38.195 79.135 40.225 79.305 ;
        RECT 40.395 78.965 40.565 79.725 ;
        RECT 40.800 79.315 41.315 79.725 ;
        RECT 44.890 79.400 45.240 80.650 ;
        RECT 47.945 80.275 48.275 80.525 ;
        RECT 48.445 80.115 48.695 80.715 ;
        RECT 48.865 80.695 49.075 81.515 ;
        RECT 49.305 80.970 54.650 81.515 ;
        RECT 50.890 80.140 51.230 80.970 ;
        RECT 54.825 80.745 56.495 81.515 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 57.585 80.745 61.095 81.515 ;
        RECT 61.265 80.755 61.975 81.345 ;
        RECT 62.485 80.985 62.815 81.345 ;
        RECT 63.015 81.155 63.345 81.515 ;
        RECT 63.515 80.985 63.845 81.345 ;
        RECT 62.485 80.775 63.845 80.985 ;
        RECT 41.485 78.965 46.830 79.400 ;
        RECT 47.965 78.965 48.195 80.105 ;
        RECT 48.365 79.135 48.695 80.115 ;
        RECT 48.865 78.965 49.075 80.105 ;
        RECT 52.710 79.400 53.060 80.650 ;
        RECT 54.825 80.225 55.575 80.745 ;
        RECT 55.745 80.055 56.495 80.575 ;
        RECT 57.585 80.225 59.235 80.745 ;
        RECT 49.305 78.965 54.650 79.400 ;
        RECT 54.825 78.965 56.495 80.055 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 59.405 80.055 61.095 80.575 ;
        RECT 57.585 78.965 61.095 80.055 ;
        RECT 61.265 79.785 61.470 80.755 ;
        RECT 64.030 80.675 64.290 81.515 ;
        RECT 64.465 80.770 64.720 81.345 ;
        RECT 64.890 81.135 65.220 81.515 ;
        RECT 65.435 80.965 65.605 81.345 ;
        RECT 64.890 80.795 65.605 80.965 ;
        RECT 65.955 80.965 66.125 81.345 ;
        RECT 66.340 81.135 66.670 81.515 ;
        RECT 65.955 80.795 66.670 80.965 ;
        RECT 61.640 79.985 61.970 80.525 ;
        RECT 62.145 80.275 62.640 80.605 ;
        RECT 62.960 80.275 63.335 80.605 ;
        RECT 63.545 80.275 63.855 80.605 ;
        RECT 62.145 79.985 62.470 80.275 ;
        RECT 62.665 79.785 62.995 80.005 ;
        RECT 61.265 79.555 62.995 79.785 ;
        RECT 61.265 79.135 61.965 79.555 ;
        RECT 62.165 78.965 62.495 79.325 ;
        RECT 62.665 79.155 62.995 79.555 ;
        RECT 63.165 79.350 63.335 80.275 ;
        RECT 63.515 78.965 63.845 80.025 ;
        RECT 64.030 78.965 64.290 80.115 ;
        RECT 64.465 80.040 64.635 80.770 ;
        RECT 64.890 80.605 65.060 80.795 ;
        RECT 64.805 80.275 65.060 80.605 ;
        RECT 64.890 80.065 65.060 80.275 ;
        RECT 65.340 80.245 65.695 80.615 ;
        RECT 65.865 80.245 66.220 80.615 ;
        RECT 66.500 80.605 66.670 80.795 ;
        RECT 66.840 80.770 67.095 81.345 ;
        RECT 66.500 80.275 66.755 80.605 ;
        RECT 66.500 80.065 66.670 80.275 ;
        RECT 64.465 79.135 64.720 80.040 ;
        RECT 64.890 79.895 65.605 80.065 ;
        RECT 64.890 78.965 65.220 79.725 ;
        RECT 65.435 79.135 65.605 79.895 ;
        RECT 65.955 79.895 66.670 80.065 ;
        RECT 66.925 80.040 67.095 80.770 ;
        RECT 67.270 80.675 67.530 81.515 ;
        RECT 68.715 80.965 68.885 81.255 ;
        RECT 69.055 81.135 69.385 81.515 ;
        RECT 68.715 80.795 69.380 80.965 ;
        RECT 65.955 79.135 66.125 79.895 ;
        RECT 66.340 78.965 66.670 79.725 ;
        RECT 66.840 79.135 67.095 80.040 ;
        RECT 67.270 78.965 67.530 80.115 ;
        RECT 68.630 79.975 68.980 80.625 ;
        RECT 69.150 79.805 69.380 80.795 ;
        RECT 68.715 79.635 69.380 79.805 ;
        RECT 68.715 79.135 68.885 79.635 ;
        RECT 69.055 78.965 69.385 79.465 ;
        RECT 69.555 79.135 69.780 81.255 ;
        RECT 69.995 81.135 70.325 81.515 ;
        RECT 70.495 80.965 70.665 81.295 ;
        RECT 70.965 81.135 71.980 81.335 ;
        RECT 69.970 80.775 70.665 80.965 ;
        RECT 69.970 79.805 70.140 80.775 ;
        RECT 70.310 79.975 70.720 80.595 ;
        RECT 70.890 80.025 71.110 80.895 ;
        RECT 71.290 80.585 71.640 80.955 ;
        RECT 71.810 80.405 71.980 81.135 ;
        RECT 72.150 81.075 72.560 81.515 ;
        RECT 72.850 80.875 73.100 81.305 ;
        RECT 73.300 81.055 73.620 81.515 ;
        RECT 74.180 81.125 75.030 81.295 ;
        RECT 72.150 80.535 72.560 80.865 ;
        RECT 72.850 80.535 73.270 80.875 ;
        RECT 71.560 80.365 71.980 80.405 ;
        RECT 71.560 80.195 72.910 80.365 ;
        RECT 69.970 79.635 70.665 79.805 ;
        RECT 70.890 79.645 71.390 80.025 ;
        RECT 69.995 78.965 70.325 79.465 ;
        RECT 70.495 79.135 70.665 79.635 ;
        RECT 71.560 79.350 71.730 80.195 ;
        RECT 72.660 80.035 72.910 80.195 ;
        RECT 71.900 79.765 72.150 80.025 ;
        RECT 73.080 79.765 73.270 80.535 ;
        RECT 71.900 79.515 73.270 79.765 ;
        RECT 73.440 80.705 74.690 80.875 ;
        RECT 73.440 79.945 73.610 80.705 ;
        RECT 74.360 80.585 74.690 80.705 ;
        RECT 73.780 80.125 73.960 80.535 ;
        RECT 74.860 80.365 75.030 81.125 ;
        RECT 75.230 81.035 75.890 81.515 ;
        RECT 76.070 80.920 76.390 81.250 ;
        RECT 75.220 80.595 75.880 80.865 ;
        RECT 75.220 80.535 75.550 80.595 ;
        RECT 75.700 80.365 76.030 80.425 ;
        RECT 74.130 80.195 76.030 80.365 ;
        RECT 73.440 79.635 73.960 79.945 ;
        RECT 74.130 79.685 74.300 80.195 ;
        RECT 76.200 80.025 76.390 80.920 ;
        RECT 74.470 79.855 76.390 80.025 ;
        RECT 76.070 79.835 76.390 79.855 ;
        RECT 76.590 80.605 76.840 81.255 ;
        RECT 77.020 81.055 77.305 81.515 ;
        RECT 77.485 81.175 77.740 81.335 ;
        RECT 77.485 81.005 77.825 81.175 ;
        RECT 77.485 80.805 77.740 81.005 ;
        RECT 76.590 80.275 77.390 80.605 ;
        RECT 74.130 79.515 75.340 79.685 ;
        RECT 70.900 79.180 71.730 79.350 ;
        RECT 71.970 78.965 72.350 79.345 ;
        RECT 72.530 79.225 72.700 79.515 ;
        RECT 74.130 79.435 74.300 79.515 ;
        RECT 72.870 78.965 73.200 79.345 ;
        RECT 73.670 79.185 74.300 79.435 ;
        RECT 74.480 78.965 74.900 79.345 ;
        RECT 75.100 79.225 75.340 79.515 ;
        RECT 75.570 78.965 75.900 79.655 ;
        RECT 76.070 79.225 76.240 79.835 ;
        RECT 76.590 79.685 76.840 80.275 ;
        RECT 77.560 79.945 77.740 80.805 ;
        RECT 76.510 79.175 76.840 79.685 ;
        RECT 77.020 78.965 77.305 79.765 ;
        RECT 77.485 79.275 77.740 79.945 ;
        RECT 79.205 80.715 79.545 81.345 ;
        RECT 79.715 80.715 79.965 81.515 ;
        RECT 80.155 80.865 80.485 81.345 ;
        RECT 80.655 81.055 80.880 81.515 ;
        RECT 81.050 80.865 81.380 81.345 ;
        RECT 79.205 80.155 79.380 80.715 ;
        RECT 80.155 80.695 81.380 80.865 ;
        RECT 82.010 80.735 82.510 81.345 ;
        RECT 82.885 80.790 83.175 81.515 ;
        RECT 83.350 80.775 83.605 81.345 ;
        RECT 83.775 81.115 84.105 81.515 ;
        RECT 84.530 80.980 85.060 81.345 ;
        RECT 84.530 80.945 84.705 80.980 ;
        RECT 83.775 80.775 84.705 80.945 ;
        RECT 85.250 80.835 85.525 81.345 ;
        RECT 79.550 80.355 80.245 80.525 ;
        RECT 79.205 80.105 79.435 80.155 ;
        RECT 80.075 80.105 80.245 80.355 ;
        RECT 80.420 80.325 80.840 80.525 ;
        RECT 81.010 80.325 81.340 80.525 ;
        RECT 81.510 80.325 81.840 80.525 ;
        RECT 82.010 80.105 82.180 80.735 ;
        RECT 82.365 80.275 82.715 80.525 ;
        RECT 79.205 79.135 79.545 80.105 ;
        RECT 79.715 78.965 79.885 80.105 ;
        RECT 80.075 79.935 82.510 80.105 ;
        RECT 80.155 78.965 80.405 79.765 ;
        RECT 81.050 79.135 81.380 79.935 ;
        RECT 81.680 78.965 82.010 79.765 ;
        RECT 82.180 79.135 82.510 79.935 ;
        RECT 82.885 78.965 83.175 80.130 ;
        RECT 83.350 80.105 83.520 80.775 ;
        RECT 83.775 80.605 83.945 80.775 ;
        RECT 83.690 80.275 83.945 80.605 ;
        RECT 84.170 80.275 84.365 80.605 ;
        RECT 83.350 79.135 83.685 80.105 ;
        RECT 83.855 78.965 84.025 80.105 ;
        RECT 84.195 79.305 84.365 80.275 ;
        RECT 84.535 79.645 84.705 80.775 ;
        RECT 84.875 79.985 85.045 80.785 ;
        RECT 85.245 80.665 85.525 80.835 ;
        RECT 85.250 80.185 85.525 80.665 ;
        RECT 85.695 79.985 85.885 81.345 ;
        RECT 86.065 80.980 86.575 81.515 ;
        RECT 86.795 80.705 87.040 81.310 ;
        RECT 87.950 80.775 88.205 81.345 ;
        RECT 88.375 81.115 88.705 81.515 ;
        RECT 89.130 80.980 89.660 81.345 ;
        RECT 89.850 81.175 90.125 81.345 ;
        RECT 89.845 81.005 90.125 81.175 ;
        RECT 89.130 80.945 89.305 80.980 ;
        RECT 88.375 80.775 89.305 80.945 ;
        RECT 86.085 80.535 87.315 80.705 ;
        RECT 84.875 79.815 85.885 79.985 ;
        RECT 86.055 79.970 86.805 80.160 ;
        RECT 84.535 79.475 85.660 79.645 ;
        RECT 86.055 79.305 86.225 79.970 ;
        RECT 86.975 79.725 87.315 80.535 ;
        RECT 84.195 79.135 86.225 79.305 ;
        RECT 86.395 78.965 86.565 79.725 ;
        RECT 86.800 79.315 87.315 79.725 ;
        RECT 87.950 80.105 88.120 80.775 ;
        RECT 88.375 80.605 88.545 80.775 ;
        RECT 88.290 80.275 88.545 80.605 ;
        RECT 88.770 80.275 88.965 80.605 ;
        RECT 87.950 79.135 88.285 80.105 ;
        RECT 88.455 78.965 88.625 80.105 ;
        RECT 88.795 79.305 88.965 80.275 ;
        RECT 89.135 79.645 89.305 80.775 ;
        RECT 89.475 79.985 89.645 80.785 ;
        RECT 89.850 80.185 90.125 81.005 ;
        RECT 90.295 79.985 90.485 81.345 ;
        RECT 90.665 80.980 91.175 81.515 ;
        RECT 91.395 80.705 91.640 81.310 ;
        RECT 90.685 80.535 91.915 80.705 ;
        RECT 92.145 80.695 92.355 81.515 ;
        RECT 92.525 80.715 92.855 81.345 ;
        RECT 89.475 79.815 90.485 79.985 ;
        RECT 90.655 79.970 91.405 80.160 ;
        RECT 89.135 79.475 90.260 79.645 ;
        RECT 90.655 79.305 90.825 79.970 ;
        RECT 91.575 79.725 91.915 80.535 ;
        RECT 92.525 80.115 92.775 80.715 ;
        RECT 93.025 80.695 93.255 81.515 ;
        RECT 93.465 80.745 96.055 81.515 ;
        RECT 96.695 81.015 97.025 81.515 ;
        RECT 97.225 80.945 97.395 81.295 ;
        RECT 97.595 81.115 97.925 81.515 ;
        RECT 98.095 80.945 98.265 81.295 ;
        RECT 98.435 81.115 98.815 81.515 ;
        RECT 92.945 80.275 93.275 80.525 ;
        RECT 93.465 80.225 94.675 80.745 ;
        RECT 88.795 79.135 90.825 79.305 ;
        RECT 90.995 78.965 91.165 79.725 ;
        RECT 91.400 79.315 91.915 79.725 ;
        RECT 92.145 78.965 92.355 80.105 ;
        RECT 92.525 79.135 92.855 80.115 ;
        RECT 93.025 78.965 93.255 80.105 ;
        RECT 94.845 80.055 96.055 80.575 ;
        RECT 96.690 80.275 97.040 80.845 ;
        RECT 97.225 80.775 98.835 80.945 ;
        RECT 99.005 80.840 99.275 81.185 ;
        RECT 99.445 80.970 104.790 81.515 ;
        RECT 98.665 80.605 98.835 80.775 ;
        RECT 97.210 80.155 97.920 80.605 ;
        RECT 98.090 80.275 98.495 80.605 ;
        RECT 98.665 80.275 98.935 80.605 ;
        RECT 93.465 78.965 96.055 80.055 ;
        RECT 96.690 79.815 97.010 80.105 ;
        RECT 97.205 79.985 97.920 80.155 ;
        RECT 98.665 80.105 98.835 80.275 ;
        RECT 99.105 80.105 99.275 80.840 ;
        RECT 101.030 80.140 101.370 80.970 ;
        RECT 104.965 80.745 108.475 81.515 ;
        RECT 108.645 80.790 108.935 81.515 ;
        RECT 109.105 80.970 114.450 81.515 ;
        RECT 114.625 80.970 119.970 81.515 ;
        RECT 98.110 79.935 98.835 80.105 ;
        RECT 98.110 79.815 98.280 79.935 ;
        RECT 96.690 79.645 98.280 79.815 ;
        RECT 96.690 79.185 98.345 79.475 ;
        RECT 98.515 78.965 98.795 79.765 ;
        RECT 99.005 79.135 99.275 80.105 ;
        RECT 102.850 79.400 103.200 80.650 ;
        RECT 104.965 80.225 106.615 80.745 ;
        RECT 106.785 80.055 108.475 80.575 ;
        RECT 110.690 80.140 111.030 80.970 ;
        RECT 99.445 78.965 104.790 79.400 ;
        RECT 104.965 78.965 108.475 80.055 ;
        RECT 108.645 78.965 108.935 80.130 ;
        RECT 112.510 79.400 112.860 80.650 ;
        RECT 116.210 80.140 116.550 80.970 ;
        RECT 120.145 80.745 123.655 81.515 ;
        RECT 124.285 80.765 125.495 81.515 ;
        RECT 118.030 79.400 118.380 80.650 ;
        RECT 120.145 80.225 121.795 80.745 ;
        RECT 121.965 80.055 123.655 80.575 ;
        RECT 109.105 78.965 114.450 79.400 ;
        RECT 114.625 78.965 119.970 79.400 ;
        RECT 120.145 78.965 123.655 80.055 ;
        RECT 124.285 80.055 124.805 80.595 ;
        RECT 124.975 80.225 125.495 80.765 ;
        RECT 124.285 78.965 125.495 80.055 ;
        RECT 5.520 78.795 125.580 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 7.535 78.125 7.705 78.625 ;
        RECT 7.875 78.295 8.205 78.795 ;
        RECT 7.535 77.955 8.200 78.125 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 7.450 77.135 7.800 77.785 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 7.970 76.965 8.200 77.955 ;
        RECT 7.535 76.795 8.200 76.965 ;
        RECT 7.535 76.505 7.705 76.795 ;
        RECT 7.875 76.245 8.205 76.625 ;
        RECT 8.375 76.505 8.600 78.625 ;
        RECT 8.815 78.295 9.145 78.795 ;
        RECT 9.315 78.125 9.485 78.625 ;
        RECT 9.720 78.410 10.550 78.580 ;
        RECT 10.790 78.415 11.170 78.795 ;
        RECT 8.790 77.955 9.485 78.125 ;
        RECT 8.790 76.985 8.960 77.955 ;
        RECT 9.130 77.165 9.540 77.785 ;
        RECT 9.710 77.735 10.210 78.115 ;
        RECT 8.790 76.795 9.485 76.985 ;
        RECT 9.710 76.865 9.930 77.735 ;
        RECT 10.380 77.565 10.550 78.410 ;
        RECT 11.350 78.245 11.520 78.535 ;
        RECT 11.690 78.415 12.020 78.795 ;
        RECT 12.490 78.325 13.120 78.575 ;
        RECT 13.300 78.415 13.720 78.795 ;
        RECT 12.950 78.245 13.120 78.325 ;
        RECT 13.920 78.245 14.160 78.535 ;
        RECT 10.720 77.995 12.090 78.245 ;
        RECT 10.720 77.735 10.970 77.995 ;
        RECT 11.480 77.565 11.730 77.725 ;
        RECT 10.380 77.395 11.730 77.565 ;
        RECT 10.380 77.355 10.800 77.395 ;
        RECT 10.110 76.805 10.460 77.175 ;
        RECT 8.815 76.245 9.145 76.625 ;
        RECT 9.315 76.465 9.485 76.795 ;
        RECT 10.630 76.625 10.800 77.355 ;
        RECT 11.900 77.225 12.090 77.995 ;
        RECT 10.970 76.895 11.380 77.225 ;
        RECT 11.670 76.885 12.090 77.225 ;
        RECT 12.260 77.815 12.780 78.125 ;
        RECT 12.950 78.075 14.160 78.245 ;
        RECT 14.390 78.105 14.720 78.795 ;
        RECT 12.260 77.055 12.430 77.815 ;
        RECT 12.600 77.225 12.780 77.635 ;
        RECT 12.950 77.565 13.120 78.075 ;
        RECT 14.890 77.925 15.060 78.535 ;
        RECT 15.330 78.075 15.660 78.585 ;
        RECT 14.890 77.905 15.210 77.925 ;
        RECT 13.290 77.735 15.210 77.905 ;
        RECT 12.950 77.395 14.850 77.565 ;
        RECT 13.180 77.055 13.510 77.175 ;
        RECT 12.260 76.885 13.510 77.055 ;
        RECT 9.785 76.425 10.800 76.625 ;
        RECT 10.970 76.245 11.380 76.685 ;
        RECT 11.670 76.455 11.920 76.885 ;
        RECT 12.120 76.245 12.440 76.705 ;
        RECT 13.680 76.635 13.850 77.395 ;
        RECT 14.520 77.335 14.850 77.395 ;
        RECT 14.040 77.165 14.370 77.225 ;
        RECT 14.040 76.895 14.700 77.165 ;
        RECT 15.020 76.840 15.210 77.735 ;
        RECT 13.000 76.465 13.850 76.635 ;
        RECT 14.050 76.245 14.710 76.725 ;
        RECT 14.890 76.510 15.210 76.840 ;
        RECT 15.410 77.485 15.660 78.075 ;
        RECT 15.840 77.995 16.125 78.795 ;
        RECT 16.305 78.455 16.560 78.485 ;
        RECT 16.305 78.285 16.645 78.455 ;
        RECT 16.305 77.815 16.560 78.285 ;
        RECT 15.410 77.155 16.210 77.485 ;
        RECT 15.410 76.505 15.660 77.155 ;
        RECT 16.380 76.955 16.560 77.815 ;
        RECT 17.165 77.655 17.375 78.795 ;
        RECT 17.545 77.645 17.875 78.625 ;
        RECT 18.045 77.655 18.275 78.795 ;
        RECT 15.840 76.245 16.125 76.705 ;
        RECT 16.305 76.425 16.560 76.955 ;
        RECT 17.165 76.245 17.375 77.065 ;
        RECT 17.545 77.045 17.795 77.645 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 18.945 77.655 19.330 78.625 ;
        RECT 19.500 78.335 19.825 78.795 ;
        RECT 20.345 78.165 20.625 78.625 ;
        RECT 19.500 77.945 20.625 78.165 ;
        RECT 17.965 77.235 18.295 77.485 ;
        RECT 17.545 76.415 17.875 77.045 ;
        RECT 18.045 76.245 18.275 77.065 ;
        RECT 18.945 76.985 19.225 77.655 ;
        RECT 19.500 77.485 19.950 77.945 ;
        RECT 20.815 77.775 21.215 78.625 ;
        RECT 21.615 78.335 21.885 78.795 ;
        RECT 22.055 78.165 22.340 78.625 ;
        RECT 19.395 77.155 19.950 77.485 ;
        RECT 20.120 77.215 21.215 77.775 ;
        RECT 19.500 77.045 19.950 77.155 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 18.945 76.415 19.330 76.985 ;
        RECT 19.500 76.875 20.625 77.045 ;
        RECT 19.500 76.245 19.825 76.705 ;
        RECT 20.345 76.415 20.625 76.875 ;
        RECT 20.815 76.415 21.215 77.215 ;
        RECT 21.385 77.945 22.340 78.165 ;
        RECT 21.385 77.045 21.595 77.945 ;
        RECT 21.765 77.215 22.455 77.775 ;
        RECT 22.685 77.655 22.895 78.795 ;
        RECT 23.065 77.645 23.395 78.625 ;
        RECT 23.565 77.655 23.795 78.795 ;
        RECT 24.005 78.360 29.350 78.795 ;
        RECT 29.525 78.360 34.870 78.795 ;
        RECT 35.045 78.360 40.390 78.795 ;
        RECT 21.385 76.875 22.340 77.045 ;
        RECT 21.615 76.245 21.885 76.705 ;
        RECT 22.055 76.415 22.340 76.875 ;
        RECT 22.685 76.245 22.895 77.065 ;
        RECT 23.065 77.045 23.315 77.645 ;
        RECT 23.485 77.235 23.815 77.485 ;
        RECT 23.065 76.415 23.395 77.045 ;
        RECT 23.565 76.245 23.795 77.065 ;
        RECT 25.590 76.790 25.930 77.620 ;
        RECT 27.410 77.110 27.760 78.360 ;
        RECT 31.110 76.790 31.450 77.620 ;
        RECT 32.930 77.110 33.280 78.360 ;
        RECT 36.630 76.790 36.970 77.620 ;
        RECT 38.450 77.110 38.800 78.360 ;
        RECT 40.565 77.705 44.075 78.795 ;
        RECT 40.565 77.015 42.215 77.535 ;
        RECT 42.385 77.185 44.075 77.705 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.705 78.360 50.050 78.795 ;
        RECT 50.225 78.360 55.570 78.795 ;
        RECT 55.745 78.360 61.090 78.795 ;
        RECT 24.005 76.245 29.350 76.790 ;
        RECT 29.525 76.245 34.870 76.790 ;
        RECT 35.045 76.245 40.390 76.790 ;
        RECT 40.565 76.245 44.075 77.015 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 46.290 76.790 46.630 77.620 ;
        RECT 48.110 77.110 48.460 78.360 ;
        RECT 51.810 76.790 52.150 77.620 ;
        RECT 53.630 77.110 53.980 78.360 ;
        RECT 57.330 76.790 57.670 77.620 ;
        RECT 59.150 77.110 59.500 78.360 ;
        RECT 61.265 77.705 62.935 78.795 ;
        RECT 61.265 77.015 62.015 77.535 ;
        RECT 62.185 77.185 62.935 77.705 ;
        RECT 63.195 77.865 63.365 78.625 ;
        RECT 63.580 78.035 63.910 78.795 ;
        RECT 63.195 77.695 63.910 77.865 ;
        RECT 64.080 77.720 64.335 78.625 ;
        RECT 63.105 77.145 63.460 77.515 ;
        RECT 63.740 77.485 63.910 77.695 ;
        RECT 63.740 77.155 63.995 77.485 ;
        RECT 44.705 76.245 50.050 76.790 ;
        RECT 50.225 76.245 55.570 76.790 ;
        RECT 55.745 76.245 61.090 76.790 ;
        RECT 61.265 76.245 62.935 77.015 ;
        RECT 63.740 76.965 63.910 77.155 ;
        RECT 64.165 76.990 64.335 77.720 ;
        RECT 64.510 77.645 64.770 78.795 ;
        RECT 64.945 77.705 68.455 78.795 ;
        RECT 68.625 77.705 69.835 78.795 ;
        RECT 63.195 76.795 63.910 76.965 ;
        RECT 63.195 76.415 63.365 76.795 ;
        RECT 63.580 76.245 63.910 76.625 ;
        RECT 64.080 76.415 64.335 76.990 ;
        RECT 64.510 76.245 64.770 77.085 ;
        RECT 64.945 77.015 66.595 77.535 ;
        RECT 66.765 77.185 68.455 77.705 ;
        RECT 64.945 76.245 68.455 77.015 ;
        RECT 68.625 76.995 69.145 77.535 ;
        RECT 69.315 77.165 69.835 77.705 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.465 77.705 72.135 78.795 ;
        RECT 72.855 78.125 73.025 78.625 ;
        RECT 73.195 78.295 73.525 78.795 ;
        RECT 72.855 77.955 73.520 78.125 ;
        RECT 70.465 77.015 71.215 77.535 ;
        RECT 71.385 77.185 72.135 77.705 ;
        RECT 72.770 77.135 73.120 77.785 ;
        RECT 68.625 76.245 69.835 76.995 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 70.465 76.245 72.135 77.015 ;
        RECT 73.290 76.965 73.520 77.955 ;
        RECT 72.855 76.795 73.520 76.965 ;
        RECT 72.855 76.505 73.025 76.795 ;
        RECT 73.195 76.245 73.525 76.625 ;
        RECT 73.695 76.505 73.920 78.625 ;
        RECT 74.135 78.295 74.465 78.795 ;
        RECT 74.635 78.125 74.805 78.625 ;
        RECT 75.040 78.410 75.870 78.580 ;
        RECT 76.110 78.415 76.490 78.795 ;
        RECT 74.110 77.955 74.805 78.125 ;
        RECT 74.110 76.985 74.280 77.955 ;
        RECT 74.450 77.165 74.860 77.785 ;
        RECT 75.030 77.735 75.530 78.115 ;
        RECT 74.110 76.795 74.805 76.985 ;
        RECT 75.030 76.865 75.250 77.735 ;
        RECT 75.700 77.565 75.870 78.410 ;
        RECT 76.670 78.245 76.840 78.535 ;
        RECT 77.010 78.415 77.340 78.795 ;
        RECT 77.810 78.325 78.440 78.575 ;
        RECT 78.620 78.415 79.040 78.795 ;
        RECT 78.270 78.245 78.440 78.325 ;
        RECT 79.240 78.245 79.480 78.535 ;
        RECT 76.040 77.995 77.410 78.245 ;
        RECT 76.040 77.735 76.290 77.995 ;
        RECT 76.800 77.565 77.050 77.725 ;
        RECT 75.700 77.395 77.050 77.565 ;
        RECT 75.700 77.355 76.120 77.395 ;
        RECT 75.430 76.805 75.780 77.175 ;
        RECT 74.135 76.245 74.465 76.625 ;
        RECT 74.635 76.465 74.805 76.795 ;
        RECT 75.950 76.625 76.120 77.355 ;
        RECT 77.220 77.225 77.410 77.995 ;
        RECT 76.290 76.895 76.700 77.225 ;
        RECT 76.990 76.885 77.410 77.225 ;
        RECT 77.580 77.815 78.100 78.125 ;
        RECT 78.270 78.075 79.480 78.245 ;
        RECT 79.710 78.105 80.040 78.795 ;
        RECT 77.580 77.055 77.750 77.815 ;
        RECT 77.920 77.225 78.100 77.635 ;
        RECT 78.270 77.565 78.440 78.075 ;
        RECT 80.210 77.925 80.380 78.535 ;
        RECT 80.650 78.075 80.980 78.585 ;
        RECT 80.210 77.905 80.530 77.925 ;
        RECT 78.610 77.735 80.530 77.905 ;
        RECT 78.270 77.395 80.170 77.565 ;
        RECT 78.500 77.055 78.830 77.175 ;
        RECT 77.580 76.885 78.830 77.055 ;
        RECT 75.105 76.425 76.120 76.625 ;
        RECT 76.290 76.245 76.700 76.685 ;
        RECT 76.990 76.455 77.240 76.885 ;
        RECT 77.440 76.245 77.760 76.705 ;
        RECT 79.000 76.635 79.170 77.395 ;
        RECT 79.840 77.335 80.170 77.395 ;
        RECT 79.360 77.165 79.690 77.225 ;
        RECT 79.360 76.895 80.020 77.165 ;
        RECT 80.340 76.840 80.530 77.735 ;
        RECT 78.320 76.465 79.170 76.635 ;
        RECT 79.370 76.245 80.030 76.725 ;
        RECT 80.210 76.510 80.530 76.840 ;
        RECT 80.730 77.485 80.980 78.075 ;
        RECT 81.160 77.995 81.445 78.795 ;
        RECT 81.625 78.455 81.880 78.485 ;
        RECT 81.625 78.285 81.965 78.455 ;
        RECT 82.425 78.360 87.770 78.795 ;
        RECT 87.945 78.360 93.290 78.795 ;
        RECT 81.625 77.815 81.880 78.285 ;
        RECT 80.730 77.155 81.530 77.485 ;
        RECT 80.730 76.505 80.980 77.155 ;
        RECT 81.700 76.955 81.880 77.815 ;
        RECT 81.160 76.245 81.445 76.705 ;
        RECT 81.625 76.425 81.880 76.955 ;
        RECT 84.010 76.790 84.350 77.620 ;
        RECT 85.830 77.110 86.180 78.360 ;
        RECT 89.530 76.790 89.870 77.620 ;
        RECT 91.350 77.110 91.700 78.360 ;
        RECT 93.465 77.705 95.135 78.795 ;
        RECT 93.465 77.015 94.215 77.535 ;
        RECT 94.385 77.185 95.135 77.705 ;
        RECT 95.765 77.630 96.055 78.795 ;
        RECT 96.225 77.705 99.735 78.795 ;
        RECT 99.905 77.705 101.115 78.795 ;
        RECT 96.225 77.015 97.875 77.535 ;
        RECT 98.045 77.185 99.735 77.705 ;
        RECT 82.425 76.245 87.770 76.790 ;
        RECT 87.945 76.245 93.290 76.790 ;
        RECT 93.465 76.245 95.135 77.015 ;
        RECT 95.765 76.245 96.055 76.970 ;
        RECT 96.225 76.245 99.735 77.015 ;
        RECT 99.905 76.995 100.425 77.535 ;
        RECT 100.595 77.165 101.115 77.705 ;
        RECT 101.490 77.825 101.820 78.625 ;
        RECT 101.990 77.995 102.320 78.795 ;
        RECT 102.620 77.825 102.950 78.625 ;
        RECT 103.595 77.995 103.845 78.795 ;
        RECT 101.490 77.655 103.925 77.825 ;
        RECT 104.115 77.655 104.285 78.795 ;
        RECT 104.455 77.655 104.795 78.625 ;
        RECT 101.285 77.235 101.635 77.485 ;
        RECT 101.820 77.025 101.990 77.655 ;
        RECT 102.160 77.235 102.490 77.435 ;
        RECT 102.660 77.235 102.990 77.435 ;
        RECT 103.160 77.235 103.580 77.435 ;
        RECT 103.755 77.405 103.925 77.655 ;
        RECT 103.755 77.235 104.450 77.405 ;
        RECT 99.905 76.245 101.115 76.995 ;
        RECT 101.490 76.415 101.990 77.025 ;
        RECT 102.620 76.895 103.845 77.065 ;
        RECT 104.620 77.045 104.795 77.655 ;
        RECT 102.620 76.415 102.950 76.895 ;
        RECT 103.120 76.245 103.345 76.705 ;
        RECT 103.515 76.415 103.845 76.895 ;
        RECT 104.035 76.245 104.285 77.045 ;
        RECT 104.455 76.415 104.795 77.045 ;
        RECT 104.965 77.655 105.305 78.625 ;
        RECT 105.475 77.655 105.645 78.795 ;
        RECT 105.915 77.995 106.165 78.795 ;
        RECT 106.810 77.825 107.140 78.625 ;
        RECT 107.440 77.995 107.770 78.795 ;
        RECT 107.940 77.825 108.270 78.625 ;
        RECT 105.835 77.655 108.270 77.825 ;
        RECT 108.645 77.705 110.315 78.795 ;
        RECT 104.965 77.045 105.140 77.655 ;
        RECT 105.835 77.405 106.005 77.655 ;
        RECT 105.310 77.235 106.005 77.405 ;
        RECT 106.180 77.235 106.600 77.435 ;
        RECT 106.770 77.235 107.100 77.435 ;
        RECT 107.270 77.235 107.600 77.435 ;
        RECT 104.965 76.415 105.305 77.045 ;
        RECT 105.475 76.245 105.725 77.045 ;
        RECT 105.915 76.895 107.140 77.065 ;
        RECT 105.915 76.415 106.245 76.895 ;
        RECT 106.415 76.245 106.640 76.705 ;
        RECT 106.810 76.415 107.140 76.895 ;
        RECT 107.770 77.025 107.940 77.655 ;
        RECT 108.125 77.235 108.475 77.485 ;
        RECT 107.770 76.415 108.270 77.025 ;
        RECT 108.645 77.015 109.395 77.535 ;
        RECT 109.565 77.185 110.315 77.705 ;
        RECT 110.575 77.865 110.745 78.625 ;
        RECT 110.925 78.035 111.255 78.795 ;
        RECT 110.575 77.695 111.240 77.865 ;
        RECT 111.425 77.720 111.695 78.625 ;
        RECT 111.955 78.125 112.125 78.625 ;
        RECT 112.295 78.295 112.625 78.795 ;
        RECT 111.955 77.955 112.620 78.125 ;
        RECT 111.070 77.550 111.240 77.695 ;
        RECT 110.505 77.145 110.835 77.515 ;
        RECT 111.070 77.220 111.355 77.550 ;
        RECT 108.645 76.245 110.315 77.015 ;
        RECT 111.070 76.965 111.240 77.220 ;
        RECT 110.575 76.795 111.240 76.965 ;
        RECT 111.525 76.920 111.695 77.720 ;
        RECT 111.870 77.135 112.220 77.785 ;
        RECT 112.390 76.965 112.620 77.955 ;
        RECT 110.575 76.415 110.745 76.795 ;
        RECT 110.925 76.245 111.255 76.625 ;
        RECT 111.435 76.415 111.695 76.920 ;
        RECT 111.955 76.795 112.620 76.965 ;
        RECT 111.955 76.505 112.125 76.795 ;
        RECT 112.295 76.245 112.625 76.625 ;
        RECT 112.795 76.505 113.020 78.625 ;
        RECT 113.235 78.295 113.565 78.795 ;
        RECT 113.735 78.125 113.905 78.625 ;
        RECT 114.140 78.410 114.970 78.580 ;
        RECT 115.210 78.415 115.590 78.795 ;
        RECT 113.210 77.955 113.905 78.125 ;
        RECT 113.210 76.985 113.380 77.955 ;
        RECT 113.550 77.165 113.960 77.785 ;
        RECT 114.130 77.735 114.630 78.115 ;
        RECT 113.210 76.795 113.905 76.985 ;
        RECT 114.130 76.865 114.350 77.735 ;
        RECT 114.800 77.565 114.970 78.410 ;
        RECT 115.770 78.245 115.940 78.535 ;
        RECT 116.110 78.415 116.440 78.795 ;
        RECT 116.910 78.325 117.540 78.575 ;
        RECT 117.720 78.415 118.140 78.795 ;
        RECT 117.370 78.245 117.540 78.325 ;
        RECT 118.340 78.245 118.580 78.535 ;
        RECT 115.140 77.995 116.510 78.245 ;
        RECT 115.140 77.735 115.390 77.995 ;
        RECT 115.900 77.565 116.150 77.725 ;
        RECT 114.800 77.395 116.150 77.565 ;
        RECT 114.800 77.355 115.220 77.395 ;
        RECT 114.530 76.805 114.880 77.175 ;
        RECT 113.235 76.245 113.565 76.625 ;
        RECT 113.735 76.465 113.905 76.795 ;
        RECT 115.050 76.625 115.220 77.355 ;
        RECT 116.320 77.225 116.510 77.995 ;
        RECT 115.390 76.895 115.800 77.225 ;
        RECT 116.090 76.885 116.510 77.225 ;
        RECT 116.680 77.815 117.200 78.125 ;
        RECT 117.370 78.075 118.580 78.245 ;
        RECT 118.810 78.105 119.140 78.795 ;
        RECT 116.680 77.055 116.850 77.815 ;
        RECT 117.020 77.225 117.200 77.635 ;
        RECT 117.370 77.565 117.540 78.075 ;
        RECT 119.310 77.925 119.480 78.535 ;
        RECT 119.750 78.075 120.080 78.585 ;
        RECT 119.310 77.905 119.630 77.925 ;
        RECT 117.710 77.735 119.630 77.905 ;
        RECT 117.370 77.395 119.270 77.565 ;
        RECT 117.600 77.055 117.930 77.175 ;
        RECT 116.680 76.885 117.930 77.055 ;
        RECT 114.205 76.425 115.220 76.625 ;
        RECT 115.390 76.245 115.800 76.685 ;
        RECT 116.090 76.455 116.340 76.885 ;
        RECT 116.540 76.245 116.860 76.705 ;
        RECT 118.100 76.635 118.270 77.395 ;
        RECT 118.940 77.335 119.270 77.395 ;
        RECT 118.460 77.165 118.790 77.225 ;
        RECT 118.460 76.895 119.120 77.165 ;
        RECT 119.440 76.840 119.630 77.735 ;
        RECT 117.420 76.465 118.270 76.635 ;
        RECT 118.470 76.245 119.130 76.725 ;
        RECT 119.310 76.510 119.630 76.840 ;
        RECT 119.830 77.485 120.080 78.075 ;
        RECT 120.260 77.995 120.545 78.795 ;
        RECT 120.725 77.815 120.980 78.485 ;
        RECT 119.830 77.155 120.630 77.485 ;
        RECT 119.830 76.505 120.080 77.155 ;
        RECT 120.800 76.955 120.980 77.815 ;
        RECT 121.525 77.630 121.815 78.795 ;
        RECT 121.985 77.705 123.655 78.795 ;
        RECT 121.985 77.015 122.735 77.535 ;
        RECT 122.905 77.185 123.655 77.705 ;
        RECT 124.285 77.705 125.495 78.795 ;
        RECT 124.285 77.165 124.805 77.705 ;
        RECT 120.725 76.755 120.980 76.955 ;
        RECT 120.260 76.245 120.545 76.705 ;
        RECT 120.725 76.585 121.065 76.755 ;
        RECT 120.725 76.425 120.980 76.585 ;
        RECT 121.525 76.245 121.815 76.970 ;
        RECT 121.985 76.245 123.655 77.015 ;
        RECT 124.975 76.995 125.495 77.535 ;
        RECT 124.285 76.245 125.495 76.995 ;
        RECT 5.520 76.075 125.580 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 6.985 75.325 8.195 76.075 ;
        RECT 8.370 75.525 8.625 75.815 ;
        RECT 8.795 75.695 9.125 76.075 ;
        RECT 8.370 75.355 9.120 75.525 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 6.985 74.785 7.505 75.325 ;
        RECT 7.675 74.615 8.195 75.155 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 6.985 73.525 8.195 74.615 ;
        RECT 8.370 74.535 8.720 75.185 ;
        RECT 8.890 74.365 9.120 75.355 ;
        RECT 8.370 74.195 9.120 74.365 ;
        RECT 8.370 73.695 8.625 74.195 ;
        RECT 8.795 73.525 9.125 74.025 ;
        RECT 9.295 73.695 9.465 75.815 ;
        RECT 9.825 75.715 10.155 76.075 ;
        RECT 10.325 75.685 10.820 75.855 ;
        RECT 11.025 75.685 11.880 75.855 ;
        RECT 9.695 74.495 10.155 75.545 ;
        RECT 9.635 73.710 9.960 74.495 ;
        RECT 10.325 74.325 10.495 75.685 ;
        RECT 10.665 74.775 11.015 75.395 ;
        RECT 11.185 75.175 11.540 75.395 ;
        RECT 11.185 74.585 11.355 75.175 ;
        RECT 11.710 74.975 11.880 75.685 ;
        RECT 12.755 75.615 13.085 76.075 ;
        RECT 13.295 75.715 13.645 75.885 ;
        RECT 12.085 75.145 12.875 75.395 ;
        RECT 13.295 75.325 13.555 75.715 ;
        RECT 13.865 75.625 14.815 75.905 ;
        RECT 14.985 75.635 15.175 76.075 ;
        RECT 15.345 75.695 16.415 75.865 ;
        RECT 13.045 74.975 13.215 75.155 ;
        RECT 10.325 74.155 10.720 74.325 ;
        RECT 10.890 74.195 11.355 74.585 ;
        RECT 11.525 74.805 13.215 74.975 ;
        RECT 10.550 74.025 10.720 74.155 ;
        RECT 11.525 74.025 11.695 74.805 ;
        RECT 13.385 74.635 13.555 75.325 ;
        RECT 12.055 74.465 13.555 74.635 ;
        RECT 13.745 74.665 13.955 75.455 ;
        RECT 14.125 74.835 14.475 75.455 ;
        RECT 14.645 74.845 14.815 75.625 ;
        RECT 15.345 75.465 15.515 75.695 ;
        RECT 14.985 75.295 15.515 75.465 ;
        RECT 14.985 75.015 15.205 75.295 ;
        RECT 15.685 75.125 15.925 75.525 ;
        RECT 14.645 74.675 15.050 74.845 ;
        RECT 15.385 74.755 15.925 75.125 ;
        RECT 16.095 75.340 16.415 75.695 ;
        RECT 16.660 75.615 16.965 76.075 ;
        RECT 17.135 75.365 17.390 75.895 ;
        RECT 16.095 75.165 16.420 75.340 ;
        RECT 16.095 74.865 17.010 75.165 ;
        RECT 16.270 74.835 17.010 74.865 ;
        RECT 13.745 74.505 14.420 74.665 ;
        RECT 14.880 74.585 15.050 74.675 ;
        RECT 13.745 74.495 14.710 74.505 ;
        RECT 13.385 74.325 13.555 74.465 ;
        RECT 10.130 73.525 10.380 73.985 ;
        RECT 10.550 73.695 10.800 74.025 ;
        RECT 11.015 73.695 11.695 74.025 ;
        RECT 11.865 74.125 12.940 74.295 ;
        RECT 13.385 74.155 13.945 74.325 ;
        RECT 14.250 74.205 14.710 74.495 ;
        RECT 14.880 74.415 16.100 74.585 ;
        RECT 11.865 73.785 12.035 74.125 ;
        RECT 12.270 73.525 12.600 73.955 ;
        RECT 12.770 73.785 12.940 74.125 ;
        RECT 13.235 73.525 13.605 73.985 ;
        RECT 13.775 73.695 13.945 74.155 ;
        RECT 14.880 74.035 15.050 74.415 ;
        RECT 16.270 74.245 16.440 74.835 ;
        RECT 17.180 74.715 17.390 75.365 ;
        RECT 17.715 75.275 18.045 76.075 ;
        RECT 18.215 75.425 18.385 75.905 ;
        RECT 18.555 75.595 18.885 76.075 ;
        RECT 19.055 75.425 19.225 75.905 ;
        RECT 19.475 75.595 19.715 76.075 ;
        RECT 19.895 75.425 20.065 75.905 ;
        RECT 14.180 73.695 15.050 74.035 ;
        RECT 15.640 74.075 16.440 74.245 ;
        RECT 15.220 73.525 15.470 73.985 ;
        RECT 15.640 73.785 15.810 74.075 ;
        RECT 15.990 73.525 16.320 73.905 ;
        RECT 16.660 73.525 16.965 74.665 ;
        RECT 17.135 73.835 17.390 74.715 ;
        RECT 18.215 75.255 19.225 75.425 ;
        RECT 19.430 75.255 20.065 75.425 ;
        RECT 20.530 75.295 21.030 75.905 ;
        RECT 18.215 75.055 18.710 75.255 ;
        RECT 19.430 75.085 19.600 75.255 ;
        RECT 18.215 74.885 18.715 75.055 ;
        RECT 19.100 74.915 19.600 75.085 ;
        RECT 18.215 74.715 18.710 74.885 ;
        RECT 17.715 73.525 18.045 74.675 ;
        RECT 18.215 74.545 19.225 74.715 ;
        RECT 18.215 73.695 18.385 74.545 ;
        RECT 18.555 73.525 18.885 74.325 ;
        RECT 19.055 73.695 19.225 74.545 ;
        RECT 19.430 74.675 19.600 74.915 ;
        RECT 19.770 74.845 20.150 75.085 ;
        RECT 20.325 74.835 20.675 75.085 ;
        RECT 19.430 74.505 20.145 74.675 ;
        RECT 20.860 74.665 21.030 75.295 ;
        RECT 21.660 75.425 21.990 75.905 ;
        RECT 22.160 75.615 22.385 76.075 ;
        RECT 22.555 75.425 22.885 75.905 ;
        RECT 21.660 75.255 22.885 75.425 ;
        RECT 23.075 75.275 23.325 76.075 ;
        RECT 23.495 75.275 23.835 75.905 ;
        RECT 24.210 75.295 24.710 75.905 ;
        RECT 21.200 74.885 21.530 75.085 ;
        RECT 21.700 74.885 22.030 75.085 ;
        RECT 22.200 74.885 22.620 75.085 ;
        RECT 22.795 74.915 23.490 75.085 ;
        RECT 22.795 74.665 22.965 74.915 ;
        RECT 23.660 74.665 23.835 75.275 ;
        RECT 24.005 74.835 24.355 75.085 ;
        RECT 24.540 74.665 24.710 75.295 ;
        RECT 25.340 75.425 25.670 75.905 ;
        RECT 25.840 75.615 26.065 76.075 ;
        RECT 26.235 75.425 26.565 75.905 ;
        RECT 25.340 75.255 26.565 75.425 ;
        RECT 26.755 75.275 27.005 76.075 ;
        RECT 27.175 75.275 27.515 75.905 ;
        RECT 27.890 75.295 28.390 75.905 ;
        RECT 24.880 74.885 25.210 75.085 ;
        RECT 25.380 74.885 25.710 75.085 ;
        RECT 25.880 74.885 26.300 75.085 ;
        RECT 26.475 74.915 27.170 75.085 ;
        RECT 26.475 74.665 26.645 74.915 ;
        RECT 27.340 74.665 27.515 75.275 ;
        RECT 27.685 74.835 28.035 75.085 ;
        RECT 28.220 74.665 28.390 75.295 ;
        RECT 29.020 75.425 29.350 75.905 ;
        RECT 29.520 75.615 29.745 76.075 ;
        RECT 29.915 75.425 30.245 75.905 ;
        RECT 29.020 75.255 30.245 75.425 ;
        RECT 30.435 75.275 30.685 76.075 ;
        RECT 30.855 75.275 31.195 75.905 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 28.560 74.885 28.890 75.085 ;
        RECT 29.060 74.885 29.390 75.085 ;
        RECT 29.560 74.885 29.980 75.085 ;
        RECT 30.155 74.915 30.850 75.085 ;
        RECT 30.155 74.665 30.325 74.915 ;
        RECT 31.020 74.665 31.195 75.275 ;
        RECT 31.825 75.305 34.415 76.075 ;
        RECT 31.825 74.785 33.035 75.305 ;
        RECT 34.790 75.295 35.290 75.905 ;
        RECT 19.405 73.525 19.645 74.325 ;
        RECT 19.815 73.695 20.145 74.505 ;
        RECT 20.530 74.495 22.965 74.665 ;
        RECT 20.530 73.695 20.860 74.495 ;
        RECT 21.030 73.525 21.360 74.325 ;
        RECT 21.660 73.695 21.990 74.495 ;
        RECT 22.635 73.525 22.885 74.325 ;
        RECT 23.155 73.525 23.325 74.665 ;
        RECT 23.495 73.695 23.835 74.665 ;
        RECT 24.210 74.495 26.645 74.665 ;
        RECT 24.210 73.695 24.540 74.495 ;
        RECT 24.710 73.525 25.040 74.325 ;
        RECT 25.340 73.695 25.670 74.495 ;
        RECT 26.315 73.525 26.565 74.325 ;
        RECT 26.835 73.525 27.005 74.665 ;
        RECT 27.175 73.695 27.515 74.665 ;
        RECT 27.890 74.495 30.325 74.665 ;
        RECT 27.890 73.695 28.220 74.495 ;
        RECT 28.390 73.525 28.720 74.325 ;
        RECT 29.020 73.695 29.350 74.495 ;
        RECT 29.995 73.525 30.245 74.325 ;
        RECT 30.515 73.525 30.685 74.665 ;
        RECT 30.855 73.695 31.195 74.665 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 33.205 74.615 34.415 75.135 ;
        RECT 34.585 74.835 34.935 75.085 ;
        RECT 35.120 74.665 35.290 75.295 ;
        RECT 35.920 75.425 36.250 75.905 ;
        RECT 36.420 75.615 36.645 76.075 ;
        RECT 36.815 75.425 37.145 75.905 ;
        RECT 35.920 75.255 37.145 75.425 ;
        RECT 37.335 75.275 37.585 76.075 ;
        RECT 37.755 75.275 38.095 75.905 ;
        RECT 35.460 74.885 35.790 75.085 ;
        RECT 35.960 74.885 36.290 75.085 ;
        RECT 36.460 74.885 36.880 75.085 ;
        RECT 37.055 74.915 37.750 75.085 ;
        RECT 37.055 74.665 37.225 74.915 ;
        RECT 37.920 74.665 38.095 75.275 ;
        RECT 31.825 73.525 34.415 74.615 ;
        RECT 34.790 74.495 37.225 74.665 ;
        RECT 34.790 73.695 35.120 74.495 ;
        RECT 35.290 73.525 35.620 74.325 ;
        RECT 35.920 73.695 36.250 74.495 ;
        RECT 36.895 73.525 37.145 74.325 ;
        RECT 37.415 73.525 37.585 74.665 ;
        RECT 37.755 73.695 38.095 74.665 ;
        RECT 38.270 75.335 38.525 75.905 ;
        RECT 38.695 75.675 39.025 76.075 ;
        RECT 39.450 75.540 39.980 75.905 ;
        RECT 39.450 75.505 39.625 75.540 ;
        RECT 38.695 75.335 39.625 75.505 ;
        RECT 40.170 75.395 40.445 75.905 ;
        RECT 38.270 74.665 38.440 75.335 ;
        RECT 38.695 75.165 38.865 75.335 ;
        RECT 38.610 74.835 38.865 75.165 ;
        RECT 39.090 74.835 39.285 75.165 ;
        RECT 38.270 73.695 38.605 74.665 ;
        RECT 38.775 73.525 38.945 74.665 ;
        RECT 39.115 73.865 39.285 74.835 ;
        RECT 39.455 74.205 39.625 75.335 ;
        RECT 39.795 74.545 39.965 75.345 ;
        RECT 40.165 75.225 40.445 75.395 ;
        RECT 40.170 74.745 40.445 75.225 ;
        RECT 40.615 74.545 40.805 75.905 ;
        RECT 40.985 75.540 41.495 76.075 ;
        RECT 41.715 75.265 41.960 75.870 ;
        RECT 42.405 75.530 47.750 76.075 ;
        RECT 41.005 75.095 42.235 75.265 ;
        RECT 39.795 74.375 40.805 74.545 ;
        RECT 40.975 74.530 41.725 74.720 ;
        RECT 39.455 74.035 40.580 74.205 ;
        RECT 40.975 73.865 41.145 74.530 ;
        RECT 41.895 74.285 42.235 75.095 ;
        RECT 43.990 74.700 44.330 75.530 ;
        RECT 47.925 75.325 49.135 76.075 ;
        RECT 39.115 73.695 41.145 73.865 ;
        RECT 41.315 73.525 41.485 74.285 ;
        RECT 41.720 73.875 42.235 74.285 ;
        RECT 45.810 73.960 46.160 75.210 ;
        RECT 47.925 74.785 48.445 75.325 ;
        RECT 49.345 75.255 49.575 76.075 ;
        RECT 49.745 75.275 50.075 75.905 ;
        RECT 48.615 74.615 49.135 75.155 ;
        RECT 49.325 74.835 49.655 75.085 ;
        RECT 49.825 74.675 50.075 75.275 ;
        RECT 50.245 75.255 50.455 76.075 ;
        RECT 50.685 75.305 53.275 76.075 ;
        RECT 50.685 74.785 51.895 75.305 ;
        RECT 53.650 75.295 54.150 75.905 ;
        RECT 42.405 73.525 47.750 73.960 ;
        RECT 47.925 73.525 49.135 74.615 ;
        RECT 49.345 73.525 49.575 74.665 ;
        RECT 49.745 73.695 50.075 74.675 ;
        RECT 50.245 73.525 50.455 74.665 ;
        RECT 52.065 74.615 53.275 75.135 ;
        RECT 53.445 74.835 53.795 75.085 ;
        RECT 53.980 74.665 54.150 75.295 ;
        RECT 54.780 75.425 55.110 75.905 ;
        RECT 55.280 75.615 55.505 76.075 ;
        RECT 55.675 75.425 56.005 75.905 ;
        RECT 54.780 75.255 56.005 75.425 ;
        RECT 56.195 75.275 56.445 76.075 ;
        RECT 56.615 75.275 56.955 75.905 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 54.320 74.885 54.650 75.085 ;
        RECT 54.820 74.885 55.150 75.085 ;
        RECT 55.320 74.885 55.740 75.085 ;
        RECT 55.915 74.915 56.610 75.085 ;
        RECT 55.915 74.665 56.085 74.915 ;
        RECT 56.780 74.665 56.955 75.275 ;
        RECT 57.585 75.275 57.925 75.905 ;
        RECT 58.095 75.275 58.345 76.075 ;
        RECT 58.535 75.425 58.865 75.905 ;
        RECT 59.035 75.615 59.260 76.075 ;
        RECT 59.430 75.425 59.760 75.905 ;
        RECT 50.685 73.525 53.275 74.615 ;
        RECT 53.650 74.495 56.085 74.665 ;
        RECT 53.650 73.695 53.980 74.495 ;
        RECT 54.150 73.525 54.480 74.325 ;
        RECT 54.780 73.695 55.110 74.495 ;
        RECT 55.755 73.525 56.005 74.325 ;
        RECT 56.275 73.525 56.445 74.665 ;
        RECT 56.615 73.695 56.955 74.665 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 57.585 74.665 57.760 75.275 ;
        RECT 58.535 75.255 59.760 75.425 ;
        RECT 60.390 75.295 60.890 75.905 ;
        RECT 61.265 75.305 64.775 76.075 ;
        RECT 64.945 75.565 65.250 76.075 ;
        RECT 57.930 74.915 58.625 75.085 ;
        RECT 58.455 74.665 58.625 74.915 ;
        RECT 58.800 74.885 59.220 75.085 ;
        RECT 59.390 74.885 59.720 75.085 ;
        RECT 59.890 74.885 60.220 75.085 ;
        RECT 60.390 74.665 60.560 75.295 ;
        RECT 60.745 74.835 61.095 75.085 ;
        RECT 61.265 74.785 62.915 75.305 ;
        RECT 57.585 73.695 57.925 74.665 ;
        RECT 58.095 73.525 58.265 74.665 ;
        RECT 58.455 74.495 60.890 74.665 ;
        RECT 63.085 74.615 64.775 75.135 ;
        RECT 64.945 74.835 65.260 75.395 ;
        RECT 65.430 75.085 65.680 75.895 ;
        RECT 65.850 75.550 66.110 76.075 ;
        RECT 66.290 75.085 66.540 75.895 ;
        RECT 66.710 75.515 66.970 76.075 ;
        RECT 67.140 75.425 67.400 75.880 ;
        RECT 67.570 75.595 67.830 76.075 ;
        RECT 68.000 75.425 68.260 75.880 ;
        RECT 68.430 75.595 68.690 76.075 ;
        RECT 68.860 75.425 69.120 75.880 ;
        RECT 69.290 75.595 69.535 76.075 ;
        RECT 69.705 75.425 69.980 75.880 ;
        RECT 70.150 75.595 70.395 76.075 ;
        RECT 70.565 75.425 70.825 75.880 ;
        RECT 71.005 75.595 71.255 76.075 ;
        RECT 71.425 75.425 71.685 75.880 ;
        RECT 71.865 75.595 72.115 76.075 ;
        RECT 72.285 75.425 72.545 75.880 ;
        RECT 72.725 75.595 72.985 76.075 ;
        RECT 73.155 75.425 73.415 75.880 ;
        RECT 73.585 75.595 73.885 76.075 ;
        RECT 74.145 75.530 79.490 76.075 ;
        RECT 67.140 75.395 73.885 75.425 ;
        RECT 67.140 75.255 73.915 75.395 ;
        RECT 72.720 75.225 73.915 75.255 ;
        RECT 65.430 74.835 72.550 75.085 ;
        RECT 58.535 73.525 58.785 74.325 ;
        RECT 59.430 73.695 59.760 74.495 ;
        RECT 60.060 73.525 60.390 74.325 ;
        RECT 60.560 73.695 60.890 74.495 ;
        RECT 61.265 73.525 64.775 74.615 ;
        RECT 64.955 73.525 65.250 74.335 ;
        RECT 65.430 73.695 65.675 74.835 ;
        RECT 65.850 73.525 66.110 74.335 ;
        RECT 66.290 73.700 66.540 74.835 ;
        RECT 72.720 74.665 73.885 75.225 ;
        RECT 75.730 74.700 76.070 75.530 ;
        RECT 79.665 75.305 82.255 76.075 ;
        RECT 82.885 75.350 83.175 76.075 ;
        RECT 83.345 75.530 88.690 76.075 ;
        RECT 67.140 74.440 73.885 74.665 ;
        RECT 67.140 74.425 72.545 74.440 ;
        RECT 66.710 73.530 66.970 74.325 ;
        RECT 67.140 73.700 67.400 74.425 ;
        RECT 67.570 73.530 67.830 74.255 ;
        RECT 68.000 73.700 68.260 74.425 ;
        RECT 68.430 73.530 68.690 74.255 ;
        RECT 68.860 73.700 69.120 74.425 ;
        RECT 69.290 73.530 69.550 74.255 ;
        RECT 69.720 73.700 69.980 74.425 ;
        RECT 70.150 73.530 70.395 74.255 ;
        RECT 70.565 73.700 70.825 74.425 ;
        RECT 71.010 73.530 71.255 74.255 ;
        RECT 71.425 73.700 71.685 74.425 ;
        RECT 71.870 73.530 72.115 74.255 ;
        RECT 72.285 73.700 72.545 74.425 ;
        RECT 72.730 73.530 72.985 74.255 ;
        RECT 73.155 73.700 73.445 74.440 ;
        RECT 66.710 73.525 72.985 73.530 ;
        RECT 73.615 73.525 73.885 74.270 ;
        RECT 77.550 73.960 77.900 75.210 ;
        RECT 79.665 74.785 80.875 75.305 ;
        RECT 81.045 74.615 82.255 75.135 ;
        RECT 84.930 74.700 85.270 75.530 ;
        RECT 88.865 75.305 90.535 76.075 ;
        RECT 74.145 73.525 79.490 73.960 ;
        RECT 79.665 73.525 82.255 74.615 ;
        RECT 82.885 73.525 83.175 74.690 ;
        RECT 86.750 73.960 87.100 75.210 ;
        RECT 88.865 74.785 89.615 75.305 ;
        RECT 91.370 75.295 91.870 75.905 ;
        RECT 89.785 74.615 90.535 75.135 ;
        RECT 91.165 74.835 91.515 75.085 ;
        RECT 91.700 74.665 91.870 75.295 ;
        RECT 92.500 75.425 92.830 75.905 ;
        RECT 93.000 75.615 93.225 76.075 ;
        RECT 93.395 75.425 93.725 75.905 ;
        RECT 92.500 75.255 93.725 75.425 ;
        RECT 93.915 75.275 94.165 76.075 ;
        RECT 94.335 75.275 94.675 75.905 ;
        RECT 92.040 74.885 92.370 75.085 ;
        RECT 92.540 74.885 92.870 75.085 ;
        RECT 93.040 74.885 93.460 75.085 ;
        RECT 93.635 74.915 94.330 75.085 ;
        RECT 93.635 74.665 93.805 74.915 ;
        RECT 94.500 74.665 94.675 75.275 ;
        RECT 94.845 75.305 96.515 76.075 ;
        RECT 96.685 75.335 97.070 75.905 ;
        RECT 97.240 75.615 97.565 76.075 ;
        RECT 98.085 75.445 98.365 75.905 ;
        RECT 94.845 74.785 95.595 75.305 ;
        RECT 83.345 73.525 88.690 73.960 ;
        RECT 88.865 73.525 90.535 74.615 ;
        RECT 91.370 74.495 93.805 74.665 ;
        RECT 91.370 73.695 91.700 74.495 ;
        RECT 91.870 73.525 92.200 74.325 ;
        RECT 92.500 73.695 92.830 74.495 ;
        RECT 93.475 73.525 93.725 74.325 ;
        RECT 93.995 73.525 94.165 74.665 ;
        RECT 94.335 73.695 94.675 74.665 ;
        RECT 95.765 74.615 96.515 75.135 ;
        RECT 94.845 73.525 96.515 74.615 ;
        RECT 96.685 74.665 96.965 75.335 ;
        RECT 97.240 75.275 98.365 75.445 ;
        RECT 97.240 75.165 97.690 75.275 ;
        RECT 97.135 74.835 97.690 75.165 ;
        RECT 98.555 75.105 98.955 75.905 ;
        RECT 99.355 75.615 99.625 76.075 ;
        RECT 99.795 75.445 100.080 75.905 ;
        RECT 96.685 73.695 97.070 74.665 ;
        RECT 97.240 74.375 97.690 74.835 ;
        RECT 97.860 74.545 98.955 75.105 ;
        RECT 97.240 74.155 98.365 74.375 ;
        RECT 97.240 73.525 97.565 73.985 ;
        RECT 98.085 73.695 98.365 74.155 ;
        RECT 98.555 73.695 98.955 74.545 ;
        RECT 99.125 75.275 100.080 75.445 ;
        RECT 100.365 75.305 102.035 76.075 ;
        RECT 99.125 74.375 99.335 75.275 ;
        RECT 99.505 74.545 100.195 75.105 ;
        RECT 100.365 74.785 101.115 75.305 ;
        RECT 102.870 75.295 103.370 75.905 ;
        RECT 101.285 74.615 102.035 75.135 ;
        RECT 102.665 74.835 103.015 75.085 ;
        RECT 103.200 74.665 103.370 75.295 ;
        RECT 104.000 75.425 104.330 75.905 ;
        RECT 104.500 75.615 104.725 76.075 ;
        RECT 104.895 75.425 105.225 75.905 ;
        RECT 104.000 75.255 105.225 75.425 ;
        RECT 105.415 75.275 105.665 76.075 ;
        RECT 105.835 75.275 106.175 75.905 ;
        RECT 103.540 74.885 103.870 75.085 ;
        RECT 104.040 74.885 104.370 75.085 ;
        RECT 104.540 74.885 104.960 75.085 ;
        RECT 105.135 74.915 105.830 75.085 ;
        RECT 105.135 74.665 105.305 74.915 ;
        RECT 106.000 74.665 106.175 75.275 ;
        RECT 106.345 75.305 108.015 76.075 ;
        RECT 108.645 75.350 108.935 76.075 ;
        RECT 106.345 74.785 107.095 75.305 ;
        RECT 109.840 75.265 110.085 75.870 ;
        RECT 110.305 75.540 110.815 76.075 ;
        RECT 99.125 74.155 100.080 74.375 ;
        RECT 99.355 73.525 99.625 73.985 ;
        RECT 99.795 73.695 100.080 74.155 ;
        RECT 100.365 73.525 102.035 74.615 ;
        RECT 102.870 74.495 105.305 74.665 ;
        RECT 102.870 73.695 103.200 74.495 ;
        RECT 103.370 73.525 103.700 74.325 ;
        RECT 104.000 73.695 104.330 74.495 ;
        RECT 104.975 73.525 105.225 74.325 ;
        RECT 105.495 73.525 105.665 74.665 ;
        RECT 105.835 73.695 106.175 74.665 ;
        RECT 107.265 74.615 108.015 75.135 ;
        RECT 109.565 75.095 110.795 75.265 ;
        RECT 106.345 73.525 108.015 74.615 ;
        RECT 108.645 73.525 108.935 74.690 ;
        RECT 109.565 74.285 109.905 75.095 ;
        RECT 110.075 74.530 110.825 74.720 ;
        RECT 109.565 73.875 110.080 74.285 ;
        RECT 110.315 73.525 110.485 74.285 ;
        RECT 110.655 73.865 110.825 74.530 ;
        RECT 110.995 74.545 111.185 75.905 ;
        RECT 111.355 75.055 111.630 75.905 ;
        RECT 111.820 75.540 112.350 75.905 ;
        RECT 112.775 75.675 113.105 76.075 ;
        RECT 112.175 75.505 112.350 75.540 ;
        RECT 111.355 74.885 111.635 75.055 ;
        RECT 111.355 74.745 111.630 74.885 ;
        RECT 111.835 74.545 112.005 75.345 ;
        RECT 110.995 74.375 112.005 74.545 ;
        RECT 112.175 75.335 113.105 75.505 ;
        RECT 113.275 75.335 113.530 75.905 ;
        RECT 112.175 74.205 112.345 75.335 ;
        RECT 112.935 75.165 113.105 75.335 ;
        RECT 111.220 74.035 112.345 74.205 ;
        RECT 112.515 74.835 112.710 75.165 ;
        RECT 112.935 74.835 113.190 75.165 ;
        RECT 112.515 73.865 112.685 74.835 ;
        RECT 113.360 74.665 113.530 75.335 ;
        RECT 113.705 75.305 116.295 76.075 ;
        RECT 113.705 74.785 114.915 75.305 ;
        RECT 116.505 75.255 116.735 76.075 ;
        RECT 116.905 75.275 117.235 75.905 ;
        RECT 110.655 73.695 112.685 73.865 ;
        RECT 112.855 73.525 113.025 74.665 ;
        RECT 113.195 73.695 113.530 74.665 ;
        RECT 115.085 74.615 116.295 75.135 ;
        RECT 116.485 74.835 116.815 75.085 ;
        RECT 116.985 74.675 117.235 75.275 ;
        RECT 117.405 75.255 117.615 76.075 ;
        RECT 117.845 75.400 118.105 75.905 ;
        RECT 118.285 75.695 118.615 76.075 ;
        RECT 118.795 75.525 118.965 75.905 ;
        RECT 113.705 73.525 116.295 74.615 ;
        RECT 116.505 73.525 116.735 74.665 ;
        RECT 116.905 73.695 117.235 74.675 ;
        RECT 117.405 73.525 117.615 74.665 ;
        RECT 117.845 74.600 118.015 75.400 ;
        RECT 118.300 75.355 118.965 75.525 ;
        RECT 118.300 75.100 118.470 75.355 ;
        RECT 119.225 75.305 122.735 76.075 ;
        RECT 122.905 75.325 124.115 76.075 ;
        RECT 124.285 75.325 125.495 76.075 ;
        RECT 118.185 74.770 118.470 75.100 ;
        RECT 118.705 74.805 119.035 75.175 ;
        RECT 119.225 74.785 120.875 75.305 ;
        RECT 118.300 74.625 118.470 74.770 ;
        RECT 117.845 73.695 118.115 74.600 ;
        RECT 118.300 74.455 118.965 74.625 ;
        RECT 121.045 74.615 122.735 75.135 ;
        RECT 122.905 74.785 123.425 75.325 ;
        RECT 123.595 74.615 124.115 75.155 ;
        RECT 118.285 73.525 118.615 74.285 ;
        RECT 118.795 73.695 118.965 74.455 ;
        RECT 119.225 73.525 122.735 74.615 ;
        RECT 122.905 73.525 124.115 74.615 ;
        RECT 124.285 74.615 124.805 75.155 ;
        RECT 124.975 74.785 125.495 75.325 ;
        RECT 124.285 73.525 125.495 74.615 ;
        RECT 5.520 73.355 125.580 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 6.985 72.920 12.330 73.355 ;
        RECT 12.505 72.920 17.850 73.355 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 8.570 71.350 8.910 72.180 ;
        RECT 10.390 71.670 10.740 72.920 ;
        RECT 14.090 71.350 14.430 72.180 ;
        RECT 15.910 71.670 16.260 72.920 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.265 20.155 73.355 ;
        RECT 18.945 71.555 19.465 72.095 ;
        RECT 19.635 71.725 20.155 72.265 ;
        RECT 20.530 72.385 20.860 73.185 ;
        RECT 21.030 72.555 21.360 73.355 ;
        RECT 21.660 72.385 21.990 73.185 ;
        RECT 22.635 72.555 22.885 73.355 ;
        RECT 20.530 72.215 22.965 72.385 ;
        RECT 23.155 72.215 23.325 73.355 ;
        RECT 23.495 72.215 23.835 73.185 ;
        RECT 24.210 72.385 24.540 73.185 ;
        RECT 24.710 72.555 25.040 73.355 ;
        RECT 25.340 72.385 25.670 73.185 ;
        RECT 26.315 72.555 26.565 73.355 ;
        RECT 24.210 72.215 26.645 72.385 ;
        RECT 26.835 72.215 27.005 73.355 ;
        RECT 27.175 72.215 27.515 73.185 ;
        RECT 27.685 72.920 33.030 73.355 ;
        RECT 20.325 71.795 20.675 72.045 ;
        RECT 20.860 71.585 21.030 72.215 ;
        RECT 21.200 71.795 21.530 71.995 ;
        RECT 21.700 71.795 22.030 71.995 ;
        RECT 22.200 71.795 22.620 71.995 ;
        RECT 22.795 71.965 22.965 72.215 ;
        RECT 22.795 71.795 23.490 71.965 ;
        RECT 6.985 70.805 12.330 71.350 ;
        RECT 12.505 70.805 17.850 71.350 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 18.945 70.805 20.155 71.555 ;
        RECT 20.530 70.975 21.030 71.585 ;
        RECT 21.660 71.455 22.885 71.625 ;
        RECT 23.660 71.605 23.835 72.215 ;
        RECT 24.005 71.795 24.355 72.045 ;
        RECT 21.660 70.975 21.990 71.455 ;
        RECT 22.160 70.805 22.385 71.265 ;
        RECT 22.555 70.975 22.885 71.455 ;
        RECT 23.075 70.805 23.325 71.605 ;
        RECT 23.495 70.975 23.835 71.605 ;
        RECT 24.540 71.585 24.710 72.215 ;
        RECT 24.880 71.795 25.210 71.995 ;
        RECT 25.380 71.795 25.710 71.995 ;
        RECT 25.880 71.795 26.300 71.995 ;
        RECT 26.475 71.965 26.645 72.215 ;
        RECT 26.475 71.795 27.170 71.965 ;
        RECT 24.210 70.975 24.710 71.585 ;
        RECT 25.340 71.455 26.565 71.625 ;
        RECT 27.340 71.605 27.515 72.215 ;
        RECT 25.340 70.975 25.670 71.455 ;
        RECT 25.840 70.805 26.065 71.265 ;
        RECT 26.235 70.975 26.565 71.455 ;
        RECT 26.755 70.805 27.005 71.605 ;
        RECT 27.175 70.975 27.515 71.605 ;
        RECT 29.270 71.350 29.610 72.180 ;
        RECT 31.090 71.670 31.440 72.920 ;
        RECT 33.295 72.425 33.465 73.185 ;
        RECT 33.645 72.595 33.975 73.355 ;
        RECT 33.295 72.255 33.960 72.425 ;
        RECT 34.145 72.280 34.415 73.185 ;
        RECT 34.675 72.685 34.845 73.185 ;
        RECT 35.015 72.855 35.345 73.355 ;
        RECT 34.675 72.515 35.340 72.685 ;
        RECT 33.790 72.110 33.960 72.255 ;
        RECT 33.225 71.705 33.555 72.075 ;
        RECT 33.790 71.780 34.075 72.110 ;
        RECT 33.790 71.525 33.960 71.780 ;
        RECT 33.295 71.355 33.960 71.525 ;
        RECT 34.245 71.480 34.415 72.280 ;
        RECT 34.590 71.695 34.940 72.345 ;
        RECT 35.110 71.525 35.340 72.515 ;
        RECT 27.685 70.805 33.030 71.350 ;
        RECT 33.295 70.975 33.465 71.355 ;
        RECT 33.645 70.805 33.975 71.185 ;
        RECT 34.155 70.975 34.415 71.480 ;
        RECT 34.675 71.355 35.340 71.525 ;
        RECT 34.675 71.065 34.845 71.355 ;
        RECT 35.015 70.805 35.345 71.185 ;
        RECT 35.515 71.065 35.740 73.185 ;
        RECT 35.955 72.855 36.285 73.355 ;
        RECT 36.455 72.685 36.625 73.185 ;
        RECT 36.860 72.970 37.690 73.140 ;
        RECT 37.930 72.975 38.310 73.355 ;
        RECT 35.930 72.515 36.625 72.685 ;
        RECT 35.930 71.545 36.100 72.515 ;
        RECT 36.270 71.725 36.680 72.345 ;
        RECT 36.850 72.295 37.350 72.675 ;
        RECT 35.930 71.355 36.625 71.545 ;
        RECT 36.850 71.425 37.070 72.295 ;
        RECT 37.520 72.125 37.690 72.970 ;
        RECT 38.490 72.805 38.660 73.095 ;
        RECT 38.830 72.975 39.160 73.355 ;
        RECT 39.630 72.885 40.260 73.135 ;
        RECT 40.440 72.975 40.860 73.355 ;
        RECT 40.090 72.805 40.260 72.885 ;
        RECT 41.060 72.805 41.300 73.095 ;
        RECT 37.860 72.555 39.230 72.805 ;
        RECT 37.860 72.295 38.110 72.555 ;
        RECT 38.620 72.125 38.870 72.285 ;
        RECT 37.520 71.955 38.870 72.125 ;
        RECT 37.520 71.915 37.940 71.955 ;
        RECT 37.250 71.365 37.600 71.735 ;
        RECT 35.955 70.805 36.285 71.185 ;
        RECT 36.455 71.025 36.625 71.355 ;
        RECT 37.770 71.185 37.940 71.915 ;
        RECT 39.040 71.785 39.230 72.555 ;
        RECT 38.110 71.455 38.520 71.785 ;
        RECT 38.810 71.445 39.230 71.785 ;
        RECT 39.400 72.375 39.920 72.685 ;
        RECT 40.090 72.635 41.300 72.805 ;
        RECT 41.530 72.665 41.860 73.355 ;
        RECT 39.400 71.615 39.570 72.375 ;
        RECT 39.740 71.785 39.920 72.195 ;
        RECT 40.090 72.125 40.260 72.635 ;
        RECT 42.030 72.485 42.200 73.095 ;
        RECT 42.470 72.635 42.800 73.145 ;
        RECT 42.030 72.465 42.350 72.485 ;
        RECT 40.430 72.295 42.350 72.465 ;
        RECT 40.090 71.955 41.990 72.125 ;
        RECT 40.320 71.615 40.650 71.735 ;
        RECT 39.400 71.445 40.650 71.615 ;
        RECT 36.925 70.985 37.940 71.185 ;
        RECT 38.110 70.805 38.520 71.245 ;
        RECT 38.810 71.015 39.060 71.445 ;
        RECT 39.260 70.805 39.580 71.265 ;
        RECT 40.820 71.195 40.990 71.955 ;
        RECT 41.660 71.895 41.990 71.955 ;
        RECT 41.180 71.725 41.510 71.785 ;
        RECT 41.180 71.455 41.840 71.725 ;
        RECT 42.160 71.400 42.350 72.295 ;
        RECT 40.140 71.025 40.990 71.195 ;
        RECT 41.190 70.805 41.850 71.285 ;
        RECT 42.030 71.070 42.350 71.400 ;
        RECT 42.550 72.045 42.800 72.635 ;
        RECT 42.980 72.555 43.265 73.355 ;
        RECT 43.445 73.015 43.700 73.045 ;
        RECT 43.445 72.845 43.785 73.015 ;
        RECT 43.445 72.375 43.700 72.845 ;
        RECT 42.550 71.715 43.350 72.045 ;
        RECT 42.550 71.065 42.800 71.715 ;
        RECT 43.520 71.515 43.700 72.375 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.765 72.215 44.975 73.355 ;
        RECT 45.145 72.205 45.475 73.185 ;
        RECT 45.645 72.215 45.875 73.355 ;
        RECT 46.175 72.685 46.345 73.185 ;
        RECT 46.515 72.855 46.845 73.355 ;
        RECT 46.175 72.515 46.840 72.685 ;
        RECT 42.980 70.805 43.265 71.265 ;
        RECT 43.445 70.985 43.700 71.515 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.765 70.805 44.975 71.625 ;
        RECT 45.145 71.605 45.395 72.205 ;
        RECT 45.565 71.795 45.895 72.045 ;
        RECT 46.090 71.695 46.440 72.345 ;
        RECT 45.145 70.975 45.475 71.605 ;
        RECT 45.645 70.805 45.875 71.625 ;
        RECT 46.610 71.525 46.840 72.515 ;
        RECT 46.175 71.355 46.840 71.525 ;
        RECT 46.175 71.065 46.345 71.355 ;
        RECT 46.515 70.805 46.845 71.185 ;
        RECT 47.015 71.065 47.240 73.185 ;
        RECT 47.455 72.855 47.785 73.355 ;
        RECT 47.955 72.685 48.125 73.185 ;
        RECT 48.360 72.970 49.190 73.140 ;
        RECT 49.430 72.975 49.810 73.355 ;
        RECT 47.430 72.515 48.125 72.685 ;
        RECT 47.430 71.545 47.600 72.515 ;
        RECT 47.770 71.725 48.180 72.345 ;
        RECT 48.350 72.295 48.850 72.675 ;
        RECT 47.430 71.355 48.125 71.545 ;
        RECT 48.350 71.425 48.570 72.295 ;
        RECT 49.020 72.125 49.190 72.970 ;
        RECT 49.990 72.805 50.160 73.095 ;
        RECT 50.330 72.975 50.660 73.355 ;
        RECT 51.130 72.885 51.760 73.135 ;
        RECT 51.940 72.975 52.360 73.355 ;
        RECT 51.590 72.805 51.760 72.885 ;
        RECT 52.560 72.805 52.800 73.095 ;
        RECT 49.360 72.555 50.730 72.805 ;
        RECT 49.360 72.295 49.610 72.555 ;
        RECT 50.120 72.125 50.370 72.285 ;
        RECT 49.020 71.955 50.370 72.125 ;
        RECT 49.020 71.915 49.440 71.955 ;
        RECT 48.750 71.365 49.100 71.735 ;
        RECT 47.455 70.805 47.785 71.185 ;
        RECT 47.955 71.025 48.125 71.355 ;
        RECT 49.270 71.185 49.440 71.915 ;
        RECT 50.540 71.785 50.730 72.555 ;
        RECT 49.610 71.455 50.020 71.785 ;
        RECT 50.310 71.445 50.730 71.785 ;
        RECT 50.900 72.375 51.420 72.685 ;
        RECT 51.590 72.635 52.800 72.805 ;
        RECT 53.030 72.665 53.360 73.355 ;
        RECT 50.900 71.615 51.070 72.375 ;
        RECT 51.240 71.785 51.420 72.195 ;
        RECT 51.590 72.125 51.760 72.635 ;
        RECT 53.530 72.485 53.700 73.095 ;
        RECT 53.970 72.635 54.300 73.145 ;
        RECT 53.530 72.465 53.850 72.485 ;
        RECT 51.930 72.295 53.850 72.465 ;
        RECT 51.590 71.955 53.490 72.125 ;
        RECT 51.820 71.615 52.150 71.735 ;
        RECT 50.900 71.445 52.150 71.615 ;
        RECT 48.425 70.985 49.440 71.185 ;
        RECT 49.610 70.805 50.020 71.245 ;
        RECT 50.310 71.015 50.560 71.445 ;
        RECT 50.760 70.805 51.080 71.265 ;
        RECT 52.320 71.195 52.490 71.955 ;
        RECT 53.160 71.895 53.490 71.955 ;
        RECT 52.680 71.725 53.010 71.785 ;
        RECT 52.680 71.455 53.340 71.725 ;
        RECT 53.660 71.400 53.850 72.295 ;
        RECT 51.640 71.025 52.490 71.195 ;
        RECT 52.690 70.805 53.350 71.285 ;
        RECT 53.530 71.070 53.850 71.400 ;
        RECT 54.050 72.045 54.300 72.635 ;
        RECT 54.480 72.555 54.765 73.355 ;
        RECT 54.945 72.675 55.200 73.045 ;
        RECT 54.945 72.505 55.285 72.675 ;
        RECT 54.945 72.375 55.200 72.505 ;
        RECT 54.050 71.715 54.850 72.045 ;
        RECT 54.050 71.065 54.300 71.715 ;
        RECT 55.020 71.515 55.200 72.375 ;
        RECT 55.950 72.385 56.280 73.185 ;
        RECT 56.450 72.555 56.780 73.355 ;
        RECT 57.080 72.385 57.410 73.185 ;
        RECT 58.055 72.555 58.305 73.355 ;
        RECT 55.950 72.215 58.385 72.385 ;
        RECT 58.575 72.215 58.745 73.355 ;
        RECT 58.915 72.215 59.255 73.185 ;
        RECT 55.745 71.795 56.095 72.045 ;
        RECT 56.280 71.585 56.450 72.215 ;
        RECT 56.620 71.795 56.950 71.995 ;
        RECT 57.120 71.795 57.450 71.995 ;
        RECT 57.620 71.795 58.040 71.995 ;
        RECT 58.215 71.965 58.385 72.215 ;
        RECT 58.215 71.795 58.910 71.965 ;
        RECT 54.480 70.805 54.765 71.265 ;
        RECT 54.945 70.985 55.200 71.515 ;
        RECT 55.950 70.975 56.450 71.585 ;
        RECT 57.080 71.455 58.305 71.625 ;
        RECT 59.080 71.605 59.255 72.215 ;
        RECT 57.080 70.975 57.410 71.455 ;
        RECT 57.580 70.805 57.805 71.265 ;
        RECT 57.975 70.975 58.305 71.455 ;
        RECT 58.495 70.805 58.745 71.605 ;
        RECT 58.915 70.975 59.255 71.605 ;
        RECT 59.425 72.215 59.765 73.185 ;
        RECT 59.935 72.215 60.105 73.355 ;
        RECT 60.375 72.555 60.625 73.355 ;
        RECT 61.270 72.385 61.600 73.185 ;
        RECT 61.900 72.555 62.230 73.355 ;
        RECT 62.400 72.385 62.730 73.185 ;
        RECT 60.295 72.215 62.730 72.385 ;
        RECT 63.195 72.425 63.365 73.185 ;
        RECT 63.580 72.595 63.910 73.355 ;
        RECT 63.195 72.255 63.910 72.425 ;
        RECT 64.080 72.280 64.335 73.185 ;
        RECT 59.425 71.605 59.600 72.215 ;
        RECT 60.295 71.965 60.465 72.215 ;
        RECT 59.770 71.795 60.465 71.965 ;
        RECT 60.640 71.795 61.060 71.995 ;
        RECT 61.230 71.795 61.560 71.995 ;
        RECT 61.730 71.795 62.060 71.995 ;
        RECT 59.425 70.975 59.765 71.605 ;
        RECT 59.935 70.805 60.185 71.605 ;
        RECT 60.375 71.455 61.600 71.625 ;
        RECT 60.375 70.975 60.705 71.455 ;
        RECT 60.875 70.805 61.100 71.265 ;
        RECT 61.270 70.975 61.600 71.455 ;
        RECT 62.230 71.585 62.400 72.215 ;
        RECT 62.585 71.795 62.935 72.045 ;
        RECT 63.105 71.705 63.460 72.075 ;
        RECT 63.740 72.045 63.910 72.255 ;
        RECT 63.740 71.715 63.995 72.045 ;
        RECT 62.230 70.975 62.730 71.585 ;
        RECT 63.740 71.525 63.910 71.715 ;
        RECT 64.165 71.550 64.335 72.280 ;
        RECT 64.510 72.205 64.770 73.355 ;
        RECT 64.945 72.265 68.455 73.355 ;
        RECT 68.625 72.265 69.835 73.355 ;
        RECT 63.195 71.355 63.910 71.525 ;
        RECT 63.195 70.975 63.365 71.355 ;
        RECT 63.580 70.805 63.910 71.185 ;
        RECT 64.080 70.975 64.335 71.550 ;
        RECT 64.510 70.805 64.770 71.645 ;
        RECT 64.945 71.575 66.595 72.095 ;
        RECT 66.765 71.745 68.455 72.265 ;
        RECT 64.945 70.805 68.455 71.575 ;
        RECT 68.625 71.555 69.145 72.095 ;
        RECT 69.315 71.725 69.835 72.265 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 70.475 72.375 70.805 73.185 ;
        RECT 70.975 72.555 71.215 73.355 ;
        RECT 70.475 72.205 71.190 72.375 ;
        RECT 70.470 71.795 70.850 72.035 ;
        RECT 71.020 71.965 71.190 72.205 ;
        RECT 71.395 72.335 71.565 73.185 ;
        RECT 71.735 72.555 72.065 73.355 ;
        RECT 72.235 72.335 72.405 73.185 ;
        RECT 71.395 72.165 72.405 72.335 ;
        RECT 72.575 72.205 72.905 73.355 ;
        RECT 73.225 72.265 75.815 73.355 ;
        RECT 71.910 71.995 72.405 72.165 ;
        RECT 71.020 71.795 71.520 71.965 ;
        RECT 71.905 71.825 72.405 71.995 ;
        RECT 71.020 71.625 71.190 71.795 ;
        RECT 71.910 71.625 72.405 71.825 ;
        RECT 68.625 70.805 69.835 71.555 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 70.555 71.455 71.190 71.625 ;
        RECT 71.395 71.455 72.405 71.625 ;
        RECT 70.555 70.975 70.725 71.455 ;
        RECT 70.905 70.805 71.145 71.285 ;
        RECT 71.395 70.975 71.565 71.455 ;
        RECT 71.735 70.805 72.065 71.285 ;
        RECT 72.235 70.975 72.405 71.455 ;
        RECT 72.575 70.805 72.905 71.605 ;
        RECT 73.225 71.575 74.435 72.095 ;
        RECT 74.605 71.745 75.815 72.265 ;
        RECT 76.650 72.385 76.980 73.185 ;
        RECT 77.150 72.555 77.480 73.355 ;
        RECT 77.780 72.385 78.110 73.185 ;
        RECT 78.755 72.555 79.005 73.355 ;
        RECT 76.650 72.215 79.085 72.385 ;
        RECT 79.275 72.215 79.445 73.355 ;
        RECT 79.615 72.215 79.955 73.185 ;
        RECT 80.330 72.385 80.660 73.185 ;
        RECT 80.830 72.555 81.160 73.355 ;
        RECT 81.460 72.385 81.790 73.185 ;
        RECT 82.435 72.555 82.685 73.355 ;
        RECT 80.330 72.215 82.765 72.385 ;
        RECT 82.955 72.215 83.125 73.355 ;
        RECT 83.295 72.215 83.635 73.185 ;
        RECT 76.445 71.795 76.795 72.045 ;
        RECT 76.980 71.585 77.150 72.215 ;
        RECT 77.320 71.795 77.650 71.995 ;
        RECT 77.820 71.795 78.150 71.995 ;
        RECT 78.320 71.795 78.740 71.995 ;
        RECT 78.915 71.965 79.085 72.215 ;
        RECT 78.915 71.795 79.610 71.965 ;
        RECT 73.225 70.805 75.815 71.575 ;
        RECT 76.650 70.975 77.150 71.585 ;
        RECT 77.780 71.455 79.005 71.625 ;
        RECT 79.780 71.605 79.955 72.215 ;
        RECT 80.125 71.795 80.475 72.045 ;
        RECT 77.780 70.975 78.110 71.455 ;
        RECT 78.280 70.805 78.505 71.265 ;
        RECT 78.675 70.975 79.005 71.455 ;
        RECT 79.195 70.805 79.445 71.605 ;
        RECT 79.615 70.975 79.955 71.605 ;
        RECT 80.660 71.585 80.830 72.215 ;
        RECT 81.000 71.795 81.330 71.995 ;
        RECT 81.500 71.795 81.830 71.995 ;
        RECT 82.000 71.795 82.420 71.995 ;
        RECT 82.595 71.965 82.765 72.215 ;
        RECT 82.595 71.795 83.290 71.965 ;
        RECT 80.330 70.975 80.830 71.585 ;
        RECT 81.460 71.455 82.685 71.625 ;
        RECT 83.460 71.605 83.635 72.215 ;
        RECT 81.460 70.975 81.790 71.455 ;
        RECT 81.960 70.805 82.185 71.265 ;
        RECT 82.355 70.975 82.685 71.455 ;
        RECT 82.875 70.805 83.125 71.605 ;
        RECT 83.295 70.975 83.635 71.605 ;
        RECT 83.805 72.215 84.145 73.185 ;
        RECT 84.315 72.215 84.485 73.355 ;
        RECT 84.755 72.555 85.005 73.355 ;
        RECT 85.650 72.385 85.980 73.185 ;
        RECT 86.280 72.555 86.610 73.355 ;
        RECT 86.780 72.385 87.110 73.185 ;
        RECT 84.675 72.215 87.110 72.385 ;
        RECT 87.485 72.215 87.825 73.185 ;
        RECT 87.995 72.215 88.165 73.355 ;
        RECT 88.435 72.555 88.685 73.355 ;
        RECT 89.330 72.385 89.660 73.185 ;
        RECT 89.960 72.555 90.290 73.355 ;
        RECT 90.460 72.385 90.790 73.185 ;
        RECT 88.355 72.215 90.790 72.385 ;
        RECT 91.165 72.215 91.505 73.185 ;
        RECT 91.675 72.215 91.845 73.355 ;
        RECT 92.115 72.555 92.365 73.355 ;
        RECT 93.010 72.385 93.340 73.185 ;
        RECT 93.640 72.555 93.970 73.355 ;
        RECT 94.140 72.385 94.470 73.185 ;
        RECT 92.035 72.215 94.470 72.385 ;
        RECT 83.805 71.605 83.980 72.215 ;
        RECT 84.675 71.965 84.845 72.215 ;
        RECT 84.150 71.795 84.845 71.965 ;
        RECT 85.020 71.795 85.440 71.995 ;
        RECT 85.610 71.795 85.940 71.995 ;
        RECT 86.110 71.795 86.440 71.995 ;
        RECT 83.805 70.975 84.145 71.605 ;
        RECT 84.315 70.805 84.565 71.605 ;
        RECT 84.755 71.455 85.980 71.625 ;
        RECT 84.755 70.975 85.085 71.455 ;
        RECT 85.255 70.805 85.480 71.265 ;
        RECT 85.650 70.975 85.980 71.455 ;
        RECT 86.610 71.585 86.780 72.215 ;
        RECT 86.965 71.795 87.315 72.045 ;
        RECT 87.485 71.605 87.660 72.215 ;
        RECT 88.355 71.965 88.525 72.215 ;
        RECT 87.830 71.795 88.525 71.965 ;
        RECT 88.700 71.795 89.120 71.995 ;
        RECT 89.290 71.795 89.620 71.995 ;
        RECT 89.790 71.795 90.120 71.995 ;
        RECT 86.610 70.975 87.110 71.585 ;
        RECT 87.485 70.975 87.825 71.605 ;
        RECT 87.995 70.805 88.245 71.605 ;
        RECT 88.435 71.455 89.660 71.625 ;
        RECT 88.435 70.975 88.765 71.455 ;
        RECT 88.935 70.805 89.160 71.265 ;
        RECT 89.330 70.975 89.660 71.455 ;
        RECT 90.290 71.585 90.460 72.215 ;
        RECT 90.645 71.795 90.995 72.045 ;
        RECT 91.165 71.605 91.340 72.215 ;
        RECT 92.035 71.965 92.205 72.215 ;
        RECT 91.510 71.795 92.205 71.965 ;
        RECT 92.380 71.795 92.800 71.995 ;
        RECT 92.970 71.795 93.300 71.995 ;
        RECT 93.470 71.795 93.800 71.995 ;
        RECT 90.290 70.975 90.790 71.585 ;
        RECT 91.165 70.975 91.505 71.605 ;
        RECT 91.675 70.805 91.925 71.605 ;
        RECT 92.115 71.455 93.340 71.625 ;
        RECT 92.115 70.975 92.445 71.455 ;
        RECT 92.615 70.805 92.840 71.265 ;
        RECT 93.010 70.975 93.340 71.455 ;
        RECT 93.970 71.585 94.140 72.215 ;
        RECT 95.765 72.190 96.055 73.355 ;
        RECT 96.225 72.215 96.565 73.185 ;
        RECT 96.735 72.215 96.905 73.355 ;
        RECT 97.175 72.555 97.425 73.355 ;
        RECT 98.070 72.385 98.400 73.185 ;
        RECT 98.700 72.555 99.030 73.355 ;
        RECT 99.200 72.385 99.530 73.185 ;
        RECT 97.095 72.215 99.530 72.385 ;
        RECT 99.995 72.425 100.165 73.185 ;
        RECT 100.345 72.595 100.675 73.355 ;
        RECT 99.995 72.255 100.660 72.425 ;
        RECT 100.845 72.280 101.115 73.185 ;
        RECT 101.375 72.685 101.545 73.185 ;
        RECT 101.715 72.855 102.045 73.355 ;
        RECT 101.375 72.515 102.040 72.685 ;
        RECT 94.325 71.795 94.675 72.045 ;
        RECT 96.225 71.605 96.400 72.215 ;
        RECT 97.095 71.965 97.265 72.215 ;
        RECT 96.570 71.795 97.265 71.965 ;
        RECT 97.440 71.795 97.860 71.995 ;
        RECT 98.030 71.795 98.360 71.995 ;
        RECT 98.530 71.795 98.860 71.995 ;
        RECT 93.970 70.975 94.470 71.585 ;
        RECT 95.765 70.805 96.055 71.530 ;
        RECT 96.225 70.975 96.565 71.605 ;
        RECT 96.735 70.805 96.985 71.605 ;
        RECT 97.175 71.455 98.400 71.625 ;
        RECT 97.175 70.975 97.505 71.455 ;
        RECT 97.675 70.805 97.900 71.265 ;
        RECT 98.070 70.975 98.400 71.455 ;
        RECT 99.030 71.585 99.200 72.215 ;
        RECT 100.490 72.110 100.660 72.255 ;
        RECT 99.385 71.795 99.735 72.045 ;
        RECT 99.925 71.705 100.255 72.075 ;
        RECT 100.490 71.780 100.775 72.110 ;
        RECT 99.030 70.975 99.530 71.585 ;
        RECT 100.490 71.525 100.660 71.780 ;
        RECT 99.995 71.355 100.660 71.525 ;
        RECT 100.945 71.480 101.115 72.280 ;
        RECT 101.290 71.695 101.640 72.345 ;
        RECT 101.810 71.525 102.040 72.515 ;
        RECT 99.995 70.975 100.165 71.355 ;
        RECT 100.345 70.805 100.675 71.185 ;
        RECT 100.855 70.975 101.115 71.480 ;
        RECT 101.375 71.355 102.040 71.525 ;
        RECT 101.375 71.065 101.545 71.355 ;
        RECT 101.715 70.805 102.045 71.185 ;
        RECT 102.215 71.065 102.440 73.185 ;
        RECT 102.655 72.855 102.985 73.355 ;
        RECT 103.155 72.685 103.325 73.185 ;
        RECT 103.560 72.970 104.390 73.140 ;
        RECT 104.630 72.975 105.010 73.355 ;
        RECT 102.630 72.515 103.325 72.685 ;
        RECT 102.630 71.545 102.800 72.515 ;
        RECT 102.970 71.725 103.380 72.345 ;
        RECT 103.550 72.295 104.050 72.675 ;
        RECT 102.630 71.355 103.325 71.545 ;
        RECT 103.550 71.425 103.770 72.295 ;
        RECT 104.220 72.125 104.390 72.970 ;
        RECT 105.190 72.805 105.360 73.095 ;
        RECT 105.530 72.975 105.860 73.355 ;
        RECT 106.330 72.885 106.960 73.135 ;
        RECT 107.140 72.975 107.560 73.355 ;
        RECT 106.790 72.805 106.960 72.885 ;
        RECT 107.760 72.805 108.000 73.095 ;
        RECT 104.560 72.555 105.930 72.805 ;
        RECT 104.560 72.295 104.810 72.555 ;
        RECT 105.320 72.125 105.570 72.285 ;
        RECT 104.220 71.955 105.570 72.125 ;
        RECT 104.220 71.915 104.640 71.955 ;
        RECT 103.950 71.365 104.300 71.735 ;
        RECT 102.655 70.805 102.985 71.185 ;
        RECT 103.155 71.025 103.325 71.355 ;
        RECT 104.470 71.185 104.640 71.915 ;
        RECT 105.740 71.785 105.930 72.555 ;
        RECT 104.810 71.455 105.220 71.785 ;
        RECT 105.510 71.445 105.930 71.785 ;
        RECT 106.100 72.375 106.620 72.685 ;
        RECT 106.790 72.635 108.000 72.805 ;
        RECT 108.230 72.665 108.560 73.355 ;
        RECT 106.100 71.615 106.270 72.375 ;
        RECT 106.440 71.785 106.620 72.195 ;
        RECT 106.790 72.125 106.960 72.635 ;
        RECT 108.730 72.485 108.900 73.095 ;
        RECT 109.170 72.635 109.500 73.145 ;
        RECT 108.730 72.465 109.050 72.485 ;
        RECT 107.130 72.295 109.050 72.465 ;
        RECT 106.790 71.955 108.690 72.125 ;
        RECT 107.020 71.615 107.350 71.735 ;
        RECT 106.100 71.445 107.350 71.615 ;
        RECT 103.625 70.985 104.640 71.185 ;
        RECT 104.810 70.805 105.220 71.245 ;
        RECT 105.510 71.015 105.760 71.445 ;
        RECT 105.960 70.805 106.280 71.265 ;
        RECT 107.520 71.195 107.690 71.955 ;
        RECT 108.360 71.895 108.690 71.955 ;
        RECT 107.880 71.725 108.210 71.785 ;
        RECT 107.880 71.455 108.540 71.725 ;
        RECT 108.860 71.400 109.050 72.295 ;
        RECT 106.840 71.025 107.690 71.195 ;
        RECT 107.890 70.805 108.550 71.285 ;
        RECT 108.730 71.070 109.050 71.400 ;
        RECT 109.250 72.045 109.500 72.635 ;
        RECT 109.680 72.555 109.965 73.355 ;
        RECT 110.145 72.375 110.400 73.045 ;
        RECT 111.955 72.685 112.125 73.185 ;
        RECT 112.295 72.855 112.625 73.355 ;
        RECT 111.955 72.515 112.620 72.685 ;
        RECT 109.250 71.715 110.050 72.045 ;
        RECT 109.250 71.065 109.500 71.715 ;
        RECT 110.220 71.515 110.400 72.375 ;
        RECT 111.870 71.695 112.220 72.345 ;
        RECT 112.390 71.525 112.620 72.515 ;
        RECT 110.145 71.315 110.400 71.515 ;
        RECT 111.955 71.355 112.620 71.525 ;
        RECT 109.680 70.805 109.965 71.265 ;
        RECT 110.145 71.145 110.485 71.315 ;
        RECT 110.145 70.985 110.400 71.145 ;
        RECT 111.955 71.065 112.125 71.355 ;
        RECT 112.295 70.805 112.625 71.185 ;
        RECT 112.795 71.065 113.020 73.185 ;
        RECT 113.235 72.855 113.565 73.355 ;
        RECT 113.735 72.685 113.905 73.185 ;
        RECT 114.140 72.970 114.970 73.140 ;
        RECT 115.210 72.975 115.590 73.355 ;
        RECT 113.210 72.515 113.905 72.685 ;
        RECT 113.210 71.545 113.380 72.515 ;
        RECT 113.550 71.725 113.960 72.345 ;
        RECT 114.130 72.295 114.630 72.675 ;
        RECT 113.210 71.355 113.905 71.545 ;
        RECT 114.130 71.425 114.350 72.295 ;
        RECT 114.800 72.125 114.970 72.970 ;
        RECT 115.770 72.805 115.940 73.095 ;
        RECT 116.110 72.975 116.440 73.355 ;
        RECT 116.910 72.885 117.540 73.135 ;
        RECT 117.720 72.975 118.140 73.355 ;
        RECT 117.370 72.805 117.540 72.885 ;
        RECT 118.340 72.805 118.580 73.095 ;
        RECT 115.140 72.555 116.510 72.805 ;
        RECT 115.140 72.295 115.390 72.555 ;
        RECT 115.900 72.125 116.150 72.285 ;
        RECT 114.800 71.955 116.150 72.125 ;
        RECT 114.800 71.915 115.220 71.955 ;
        RECT 114.530 71.365 114.880 71.735 ;
        RECT 113.235 70.805 113.565 71.185 ;
        RECT 113.735 71.025 113.905 71.355 ;
        RECT 115.050 71.185 115.220 71.915 ;
        RECT 116.320 71.785 116.510 72.555 ;
        RECT 115.390 71.455 115.800 71.785 ;
        RECT 116.090 71.445 116.510 71.785 ;
        RECT 116.680 72.375 117.200 72.685 ;
        RECT 117.370 72.635 118.580 72.805 ;
        RECT 118.810 72.665 119.140 73.355 ;
        RECT 116.680 71.615 116.850 72.375 ;
        RECT 117.020 71.785 117.200 72.195 ;
        RECT 117.370 72.125 117.540 72.635 ;
        RECT 119.310 72.485 119.480 73.095 ;
        RECT 119.750 72.635 120.080 73.145 ;
        RECT 119.310 72.465 119.630 72.485 ;
        RECT 117.710 72.295 119.630 72.465 ;
        RECT 117.370 71.955 119.270 72.125 ;
        RECT 117.600 71.615 117.930 71.735 ;
        RECT 116.680 71.445 117.930 71.615 ;
        RECT 114.205 70.985 115.220 71.185 ;
        RECT 115.390 70.805 115.800 71.245 ;
        RECT 116.090 71.015 116.340 71.445 ;
        RECT 116.540 70.805 116.860 71.265 ;
        RECT 118.100 71.195 118.270 71.955 ;
        RECT 118.940 71.895 119.270 71.955 ;
        RECT 118.460 71.725 118.790 71.785 ;
        RECT 118.460 71.455 119.120 71.725 ;
        RECT 119.440 71.400 119.630 72.295 ;
        RECT 117.420 71.025 118.270 71.195 ;
        RECT 118.470 70.805 119.130 71.285 ;
        RECT 119.310 71.070 119.630 71.400 ;
        RECT 119.830 72.045 120.080 72.635 ;
        RECT 120.260 72.555 120.545 73.355 ;
        RECT 120.725 72.375 120.980 73.045 ;
        RECT 119.830 71.715 120.630 72.045 ;
        RECT 119.830 71.065 120.080 71.715 ;
        RECT 120.800 71.515 120.980 72.375 ;
        RECT 121.525 72.190 121.815 73.355 ;
        RECT 122.025 72.215 122.255 73.355 ;
        RECT 122.425 72.205 122.755 73.185 ;
        RECT 122.925 72.215 123.135 73.355 ;
        RECT 124.285 72.265 125.495 73.355 ;
        RECT 122.005 71.795 122.335 72.045 ;
        RECT 120.725 71.315 120.980 71.515 ;
        RECT 120.260 70.805 120.545 71.265 ;
        RECT 120.725 71.145 121.065 71.315 ;
        RECT 120.725 70.985 120.980 71.145 ;
        RECT 121.525 70.805 121.815 71.530 ;
        RECT 122.025 70.805 122.255 71.625 ;
        RECT 122.505 71.605 122.755 72.205 ;
        RECT 124.285 71.725 124.805 72.265 ;
        RECT 122.425 70.975 122.755 71.605 ;
        RECT 122.925 70.805 123.135 71.625 ;
        RECT 124.975 71.555 125.495 72.095 ;
        RECT 124.285 70.805 125.495 71.555 ;
        RECT 5.520 70.635 125.580 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 6.985 70.090 12.330 70.635 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 8.570 69.260 8.910 70.090 ;
        RECT 12.505 69.885 13.715 70.635 ;
        RECT 13.975 69.985 14.145 70.465 ;
        RECT 14.325 70.155 14.565 70.635 ;
        RECT 14.815 69.985 14.985 70.465 ;
        RECT 15.155 70.155 15.485 70.635 ;
        RECT 15.655 69.985 15.825 70.465 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 10.390 68.520 10.740 69.770 ;
        RECT 12.505 69.345 13.025 69.885 ;
        RECT 13.975 69.815 14.610 69.985 ;
        RECT 14.815 69.815 15.825 69.985 ;
        RECT 15.995 69.835 16.325 70.635 ;
        RECT 16.645 70.090 21.990 70.635 ;
        RECT 22.165 70.090 27.510 70.635 ;
        RECT 13.195 69.175 13.715 69.715 ;
        RECT 14.440 69.645 14.610 69.815 ;
        RECT 15.325 69.785 15.825 69.815 ;
        RECT 13.890 69.405 14.270 69.645 ;
        RECT 14.440 69.475 14.940 69.645 ;
        RECT 14.440 69.235 14.610 69.475 ;
        RECT 15.330 69.275 15.825 69.785 ;
        RECT 6.985 68.085 12.330 68.520 ;
        RECT 12.505 68.085 13.715 69.175 ;
        RECT 13.895 69.065 14.610 69.235 ;
        RECT 14.815 69.105 15.825 69.275 ;
        RECT 18.230 69.260 18.570 70.090 ;
        RECT 13.895 68.255 14.225 69.065 ;
        RECT 14.395 68.085 14.635 68.885 ;
        RECT 14.815 68.255 14.985 69.105 ;
        RECT 15.155 68.085 15.485 68.885 ;
        RECT 15.655 68.255 15.825 69.105 ;
        RECT 15.995 68.085 16.325 69.235 ;
        RECT 20.050 68.520 20.400 69.770 ;
        RECT 23.750 69.260 24.090 70.090 ;
        RECT 27.685 69.865 29.355 70.635 ;
        RECT 30.075 70.085 30.245 70.465 ;
        RECT 30.425 70.255 30.755 70.635 ;
        RECT 30.075 69.915 30.740 70.085 ;
        RECT 30.935 69.960 31.195 70.465 ;
        RECT 25.570 68.520 25.920 69.770 ;
        RECT 27.685 69.345 28.435 69.865 ;
        RECT 28.605 69.175 29.355 69.695 ;
        RECT 30.005 69.365 30.335 69.735 ;
        RECT 30.570 69.660 30.740 69.915 ;
        RECT 30.570 69.330 30.855 69.660 ;
        RECT 30.570 69.185 30.740 69.330 ;
        RECT 16.645 68.085 21.990 68.520 ;
        RECT 22.165 68.085 27.510 68.520 ;
        RECT 27.685 68.085 29.355 69.175 ;
        RECT 30.075 69.015 30.740 69.185 ;
        RECT 31.025 69.160 31.195 69.960 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 31.915 70.085 32.085 70.375 ;
        RECT 32.255 70.255 32.585 70.635 ;
        RECT 31.915 69.915 32.580 70.085 ;
        RECT 30.075 68.255 30.245 69.015 ;
        RECT 30.425 68.085 30.755 68.845 ;
        RECT 30.925 68.255 31.195 69.160 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 31.830 69.095 32.180 69.745 ;
        RECT 32.350 68.925 32.580 69.915 ;
        RECT 31.915 68.755 32.580 68.925 ;
        RECT 31.915 68.255 32.085 68.755 ;
        RECT 32.255 68.085 32.585 68.585 ;
        RECT 32.755 68.255 32.980 70.375 ;
        RECT 33.195 70.255 33.525 70.635 ;
        RECT 33.695 70.085 33.865 70.415 ;
        RECT 34.165 70.255 35.180 70.455 ;
        RECT 33.170 69.895 33.865 70.085 ;
        RECT 33.170 68.925 33.340 69.895 ;
        RECT 33.510 69.095 33.920 69.715 ;
        RECT 34.090 69.145 34.310 70.015 ;
        RECT 34.490 69.705 34.840 70.075 ;
        RECT 35.010 69.525 35.180 70.255 ;
        RECT 35.350 70.195 35.760 70.635 ;
        RECT 36.050 69.995 36.300 70.425 ;
        RECT 36.500 70.175 36.820 70.635 ;
        RECT 37.380 70.245 38.230 70.415 ;
        RECT 35.350 69.655 35.760 69.985 ;
        RECT 36.050 69.655 36.470 69.995 ;
        RECT 34.760 69.485 35.180 69.525 ;
        RECT 34.760 69.315 36.110 69.485 ;
        RECT 33.170 68.755 33.865 68.925 ;
        RECT 34.090 68.765 34.590 69.145 ;
        RECT 33.195 68.085 33.525 68.585 ;
        RECT 33.695 68.255 33.865 68.755 ;
        RECT 34.760 68.470 34.930 69.315 ;
        RECT 35.860 69.155 36.110 69.315 ;
        RECT 35.100 68.885 35.350 69.145 ;
        RECT 36.280 68.885 36.470 69.655 ;
        RECT 35.100 68.635 36.470 68.885 ;
        RECT 36.640 69.825 37.890 69.995 ;
        RECT 36.640 69.065 36.810 69.825 ;
        RECT 37.560 69.705 37.890 69.825 ;
        RECT 36.980 69.245 37.160 69.655 ;
        RECT 38.060 69.485 38.230 70.245 ;
        RECT 38.430 70.155 39.090 70.635 ;
        RECT 39.270 70.040 39.590 70.370 ;
        RECT 38.420 69.715 39.080 69.985 ;
        RECT 38.420 69.655 38.750 69.715 ;
        RECT 38.900 69.485 39.230 69.545 ;
        RECT 37.330 69.315 39.230 69.485 ;
        RECT 36.640 68.755 37.160 69.065 ;
        RECT 37.330 68.805 37.500 69.315 ;
        RECT 39.400 69.145 39.590 70.040 ;
        RECT 37.670 68.975 39.590 69.145 ;
        RECT 39.270 68.955 39.590 68.975 ;
        RECT 39.790 69.725 40.040 70.375 ;
        RECT 40.220 70.175 40.505 70.635 ;
        RECT 40.685 69.925 40.940 70.455 ;
        RECT 41.485 70.090 46.830 70.635 ;
        RECT 39.790 69.395 40.590 69.725 ;
        RECT 37.330 68.635 38.540 68.805 ;
        RECT 34.100 68.300 34.930 68.470 ;
        RECT 35.170 68.085 35.550 68.465 ;
        RECT 35.730 68.345 35.900 68.635 ;
        RECT 37.330 68.555 37.500 68.635 ;
        RECT 36.070 68.085 36.400 68.465 ;
        RECT 36.870 68.305 37.500 68.555 ;
        RECT 37.680 68.085 38.100 68.465 ;
        RECT 38.300 68.345 38.540 68.635 ;
        RECT 38.770 68.085 39.100 68.775 ;
        RECT 39.270 68.345 39.440 68.955 ;
        RECT 39.790 68.805 40.040 69.395 ;
        RECT 40.760 69.275 40.940 69.925 ;
        RECT 40.760 69.105 41.025 69.275 ;
        RECT 43.070 69.260 43.410 70.090 ;
        RECT 47.005 69.865 48.675 70.635 ;
        RECT 48.845 69.960 49.105 70.465 ;
        RECT 49.285 70.255 49.615 70.635 ;
        RECT 49.795 70.085 49.965 70.465 ;
        RECT 40.760 69.065 40.940 69.105 ;
        RECT 39.710 68.295 40.040 68.805 ;
        RECT 40.220 68.085 40.505 68.885 ;
        RECT 40.685 68.395 40.940 69.065 ;
        RECT 44.890 68.520 45.240 69.770 ;
        RECT 47.005 69.345 47.755 69.865 ;
        RECT 47.925 69.175 48.675 69.695 ;
        RECT 41.485 68.085 46.830 68.520 ;
        RECT 47.005 68.085 48.675 69.175 ;
        RECT 48.845 69.160 49.015 69.960 ;
        RECT 49.300 69.915 49.965 70.085 ;
        RECT 49.300 69.660 49.470 69.915 ;
        RECT 50.230 69.895 50.485 70.465 ;
        RECT 50.655 70.235 50.985 70.635 ;
        RECT 51.410 70.100 51.940 70.465 ;
        RECT 52.130 70.295 52.405 70.465 ;
        RECT 52.125 70.125 52.405 70.295 ;
        RECT 51.410 70.065 51.585 70.100 ;
        RECT 50.655 69.895 51.585 70.065 ;
        RECT 49.185 69.330 49.470 69.660 ;
        RECT 49.705 69.365 50.035 69.735 ;
        RECT 49.300 69.185 49.470 69.330 ;
        RECT 50.230 69.225 50.400 69.895 ;
        RECT 50.655 69.725 50.825 69.895 ;
        RECT 50.570 69.395 50.825 69.725 ;
        RECT 51.050 69.395 51.245 69.725 ;
        RECT 48.845 68.255 49.115 69.160 ;
        RECT 49.300 69.015 49.965 69.185 ;
        RECT 49.285 68.085 49.615 68.845 ;
        RECT 49.795 68.255 49.965 69.015 ;
        RECT 50.230 68.255 50.565 69.225 ;
        RECT 50.735 68.085 50.905 69.225 ;
        RECT 51.075 68.425 51.245 69.395 ;
        RECT 51.415 68.765 51.585 69.895 ;
        RECT 51.755 69.105 51.925 69.905 ;
        RECT 52.130 69.305 52.405 70.125 ;
        RECT 52.575 69.105 52.765 70.465 ;
        RECT 52.945 70.100 53.455 70.635 ;
        RECT 53.675 69.825 53.920 70.430 ;
        RECT 54.365 69.865 56.955 70.635 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 57.585 69.865 61.095 70.635 ;
        RECT 52.965 69.655 54.195 69.825 ;
        RECT 51.755 68.935 52.765 69.105 ;
        RECT 52.935 69.090 53.685 69.280 ;
        RECT 51.415 68.595 52.540 68.765 ;
        RECT 52.935 68.425 53.105 69.090 ;
        RECT 53.855 68.845 54.195 69.655 ;
        RECT 54.365 69.345 55.575 69.865 ;
        RECT 55.745 69.175 56.955 69.695 ;
        RECT 57.585 69.345 59.235 69.865 ;
        RECT 62.190 69.795 62.450 70.635 ;
        RECT 62.625 69.890 62.880 70.465 ;
        RECT 63.050 70.255 63.380 70.635 ;
        RECT 63.595 70.085 63.765 70.465 ;
        RECT 63.050 69.915 63.765 70.085 ;
        RECT 51.075 68.255 53.105 68.425 ;
        RECT 53.275 68.085 53.445 68.845 ;
        RECT 53.680 68.435 54.195 68.845 ;
        RECT 54.365 68.085 56.955 69.175 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 59.405 69.175 61.095 69.695 ;
        RECT 57.585 68.085 61.095 69.175 ;
        RECT 62.190 68.085 62.450 69.235 ;
        RECT 62.625 69.160 62.795 69.890 ;
        RECT 63.050 69.725 63.220 69.915 ;
        RECT 64.030 69.795 64.290 70.635 ;
        RECT 64.465 69.890 64.720 70.465 ;
        RECT 64.890 70.255 65.220 70.635 ;
        RECT 65.435 70.085 65.605 70.465 ;
        RECT 64.890 69.915 65.605 70.085 ;
        RECT 65.955 70.085 66.125 70.465 ;
        RECT 66.340 70.255 66.670 70.635 ;
        RECT 65.955 69.915 66.670 70.085 ;
        RECT 62.965 69.395 63.220 69.725 ;
        RECT 63.050 69.185 63.220 69.395 ;
        RECT 63.500 69.365 63.855 69.735 ;
        RECT 62.625 68.255 62.880 69.160 ;
        RECT 63.050 69.015 63.765 69.185 ;
        RECT 63.050 68.085 63.380 68.845 ;
        RECT 63.595 68.255 63.765 69.015 ;
        RECT 64.030 68.085 64.290 69.235 ;
        RECT 64.465 69.160 64.635 69.890 ;
        RECT 64.890 69.725 65.060 69.915 ;
        RECT 64.805 69.395 65.060 69.725 ;
        RECT 64.890 69.185 65.060 69.395 ;
        RECT 65.340 69.365 65.695 69.735 ;
        RECT 65.865 69.365 66.220 69.735 ;
        RECT 66.500 69.725 66.670 69.915 ;
        RECT 66.840 69.890 67.095 70.465 ;
        RECT 66.500 69.395 66.755 69.725 ;
        RECT 66.500 69.185 66.670 69.395 ;
        RECT 64.465 68.255 64.720 69.160 ;
        RECT 64.890 69.015 65.605 69.185 ;
        RECT 64.890 68.085 65.220 68.845 ;
        RECT 65.435 68.255 65.605 69.015 ;
        RECT 65.955 69.015 66.670 69.185 ;
        RECT 66.925 69.160 67.095 69.890 ;
        RECT 67.270 69.795 67.530 70.635 ;
        RECT 67.795 70.085 67.965 70.465 ;
        RECT 68.180 70.255 68.510 70.635 ;
        RECT 67.795 69.915 68.510 70.085 ;
        RECT 67.705 69.365 68.060 69.735 ;
        RECT 68.340 69.725 68.510 69.915 ;
        RECT 68.680 69.890 68.935 70.465 ;
        RECT 68.340 69.395 68.595 69.725 ;
        RECT 65.955 68.255 66.125 69.015 ;
        RECT 66.340 68.085 66.670 68.845 ;
        RECT 66.840 68.255 67.095 69.160 ;
        RECT 67.270 68.085 67.530 69.235 ;
        RECT 68.340 69.185 68.510 69.395 ;
        RECT 67.795 69.015 68.510 69.185 ;
        RECT 68.765 69.160 68.935 69.890 ;
        RECT 69.110 69.795 69.370 70.635 ;
        RECT 69.545 69.865 73.055 70.635 ;
        RECT 73.690 69.895 73.945 70.465 ;
        RECT 74.115 70.235 74.445 70.635 ;
        RECT 74.870 70.100 75.400 70.465 ;
        RECT 74.870 70.065 75.045 70.100 ;
        RECT 74.115 69.895 75.045 70.065 ;
        RECT 75.590 69.955 75.865 70.465 ;
        RECT 69.545 69.345 71.195 69.865 ;
        RECT 67.795 68.255 67.965 69.015 ;
        RECT 68.180 68.085 68.510 68.845 ;
        RECT 68.680 68.255 68.935 69.160 ;
        RECT 69.110 68.085 69.370 69.235 ;
        RECT 71.365 69.175 73.055 69.695 ;
        RECT 69.545 68.085 73.055 69.175 ;
        RECT 73.690 69.225 73.860 69.895 ;
        RECT 74.115 69.725 74.285 69.895 ;
        RECT 74.030 69.395 74.285 69.725 ;
        RECT 74.510 69.395 74.705 69.725 ;
        RECT 73.690 68.255 74.025 69.225 ;
        RECT 74.195 68.085 74.365 69.225 ;
        RECT 74.535 68.425 74.705 69.395 ;
        RECT 74.875 68.765 75.045 69.895 ;
        RECT 75.215 69.105 75.385 69.905 ;
        RECT 75.585 69.785 75.865 69.955 ;
        RECT 75.590 69.305 75.865 69.785 ;
        RECT 76.035 69.105 76.225 70.465 ;
        RECT 76.405 70.100 76.915 70.635 ;
        RECT 77.135 69.825 77.380 70.430 ;
        RECT 77.825 69.865 81.335 70.635 ;
        RECT 81.505 69.885 82.715 70.635 ;
        RECT 82.885 69.910 83.175 70.635 ;
        RECT 83.345 69.895 83.730 70.465 ;
        RECT 83.900 70.175 84.225 70.635 ;
        RECT 84.745 70.005 85.025 70.465 ;
        RECT 76.425 69.655 77.655 69.825 ;
        RECT 75.215 68.935 76.225 69.105 ;
        RECT 76.395 69.090 77.145 69.280 ;
        RECT 74.875 68.595 76.000 68.765 ;
        RECT 76.395 68.425 76.565 69.090 ;
        RECT 77.315 68.845 77.655 69.655 ;
        RECT 77.825 69.345 79.475 69.865 ;
        RECT 79.645 69.175 81.335 69.695 ;
        RECT 81.505 69.345 82.025 69.885 ;
        RECT 82.195 69.175 82.715 69.715 ;
        RECT 74.535 68.255 76.565 68.425 ;
        RECT 76.735 68.085 76.905 68.845 ;
        RECT 77.140 68.435 77.655 68.845 ;
        RECT 77.825 68.085 81.335 69.175 ;
        RECT 81.505 68.085 82.715 69.175 ;
        RECT 82.885 68.085 83.175 69.250 ;
        RECT 83.345 69.225 83.625 69.895 ;
        RECT 83.900 69.835 85.025 70.005 ;
        RECT 83.900 69.725 84.350 69.835 ;
        RECT 83.795 69.395 84.350 69.725 ;
        RECT 85.215 69.665 85.615 70.465 ;
        RECT 86.015 70.175 86.285 70.635 ;
        RECT 86.455 70.005 86.740 70.465 ;
        RECT 83.345 68.255 83.730 69.225 ;
        RECT 83.900 68.935 84.350 69.395 ;
        RECT 84.520 69.105 85.615 69.665 ;
        RECT 83.900 68.715 85.025 68.935 ;
        RECT 83.900 68.085 84.225 68.545 ;
        RECT 84.745 68.255 85.025 68.715 ;
        RECT 85.215 68.255 85.615 69.105 ;
        RECT 85.785 69.835 86.740 70.005 ;
        RECT 87.025 69.895 87.410 70.465 ;
        RECT 87.580 70.175 87.905 70.635 ;
        RECT 88.425 70.005 88.705 70.465 ;
        RECT 85.785 68.935 85.995 69.835 ;
        RECT 86.165 69.105 86.855 69.665 ;
        RECT 87.025 69.225 87.305 69.895 ;
        RECT 87.580 69.835 88.705 70.005 ;
        RECT 87.580 69.725 88.030 69.835 ;
        RECT 87.475 69.395 88.030 69.725 ;
        RECT 88.895 69.665 89.295 70.465 ;
        RECT 89.695 70.175 89.965 70.635 ;
        RECT 90.135 70.005 90.420 70.465 ;
        RECT 85.785 68.715 86.740 68.935 ;
        RECT 86.015 68.085 86.285 68.545 ;
        RECT 86.455 68.255 86.740 68.715 ;
        RECT 87.025 68.255 87.410 69.225 ;
        RECT 87.580 68.935 88.030 69.395 ;
        RECT 88.200 69.105 89.295 69.665 ;
        RECT 87.580 68.715 88.705 68.935 ;
        RECT 87.580 68.085 87.905 68.545 ;
        RECT 88.425 68.255 88.705 68.715 ;
        RECT 88.895 68.255 89.295 69.105 ;
        RECT 89.465 69.835 90.420 70.005 ;
        RECT 90.705 69.865 94.215 70.635 ;
        RECT 89.465 68.935 89.675 69.835 ;
        RECT 89.845 69.105 90.535 69.665 ;
        RECT 90.705 69.345 92.355 69.865 ;
        RECT 94.660 69.825 94.905 70.430 ;
        RECT 95.125 70.100 95.635 70.635 ;
        RECT 92.525 69.175 94.215 69.695 ;
        RECT 89.465 68.715 90.420 68.935 ;
        RECT 89.695 68.085 89.965 68.545 ;
        RECT 90.135 68.255 90.420 68.715 ;
        RECT 90.705 68.085 94.215 69.175 ;
        RECT 94.385 69.655 95.615 69.825 ;
        RECT 94.385 68.845 94.725 69.655 ;
        RECT 94.895 69.090 95.645 69.280 ;
        RECT 94.385 68.435 94.900 68.845 ;
        RECT 95.135 68.085 95.305 68.845 ;
        RECT 95.475 68.425 95.645 69.090 ;
        RECT 95.815 69.105 96.005 70.465 ;
        RECT 96.175 70.295 96.450 70.465 ;
        RECT 96.175 70.125 96.455 70.295 ;
        RECT 96.175 69.305 96.450 70.125 ;
        RECT 96.640 70.100 97.170 70.465 ;
        RECT 97.595 70.235 97.925 70.635 ;
        RECT 96.995 70.065 97.170 70.100 ;
        RECT 96.655 69.105 96.825 69.905 ;
        RECT 95.815 68.935 96.825 69.105 ;
        RECT 96.995 69.895 97.925 70.065 ;
        RECT 98.095 69.895 98.350 70.465 ;
        RECT 96.995 68.765 97.165 69.895 ;
        RECT 97.755 69.725 97.925 69.895 ;
        RECT 96.040 68.595 97.165 68.765 ;
        RECT 97.335 69.395 97.530 69.725 ;
        RECT 97.755 69.395 98.010 69.725 ;
        RECT 97.335 68.425 97.505 69.395 ;
        RECT 98.180 69.225 98.350 69.895 ;
        RECT 95.475 68.255 97.505 68.425 ;
        RECT 97.675 68.085 97.845 69.225 ;
        RECT 98.015 68.255 98.350 69.225 ;
        RECT 98.525 69.960 98.785 70.465 ;
        RECT 98.965 70.255 99.295 70.635 ;
        RECT 99.475 70.085 99.645 70.465 ;
        RECT 98.525 69.160 98.695 69.960 ;
        RECT 98.980 69.915 99.645 70.085 ;
        RECT 98.980 69.660 99.150 69.915 ;
        RECT 99.905 69.885 101.115 70.635 ;
        RECT 101.290 69.895 101.545 70.465 ;
        RECT 101.715 70.235 102.045 70.635 ;
        RECT 102.470 70.100 103.000 70.465 ;
        RECT 103.190 70.295 103.465 70.465 ;
        RECT 103.185 70.125 103.465 70.295 ;
        RECT 102.470 70.065 102.645 70.100 ;
        RECT 101.715 69.895 102.645 70.065 ;
        RECT 98.865 69.330 99.150 69.660 ;
        RECT 99.385 69.365 99.715 69.735 ;
        RECT 99.905 69.345 100.425 69.885 ;
        RECT 98.980 69.185 99.150 69.330 ;
        RECT 98.525 68.255 98.795 69.160 ;
        RECT 98.980 69.015 99.645 69.185 ;
        RECT 100.595 69.175 101.115 69.715 ;
        RECT 98.965 68.085 99.295 68.845 ;
        RECT 99.475 68.255 99.645 69.015 ;
        RECT 99.905 68.085 101.115 69.175 ;
        RECT 101.290 69.225 101.460 69.895 ;
        RECT 101.715 69.725 101.885 69.895 ;
        RECT 101.630 69.395 101.885 69.725 ;
        RECT 102.110 69.395 102.305 69.725 ;
        RECT 101.290 68.255 101.625 69.225 ;
        RECT 101.795 68.085 101.965 69.225 ;
        RECT 102.135 68.425 102.305 69.395 ;
        RECT 102.475 68.765 102.645 69.895 ;
        RECT 102.815 69.105 102.985 69.905 ;
        RECT 103.190 69.305 103.465 70.125 ;
        RECT 103.635 69.105 103.825 70.465 ;
        RECT 104.005 70.100 104.515 70.635 ;
        RECT 104.735 69.825 104.980 70.430 ;
        RECT 104.025 69.655 105.255 69.825 ;
        RECT 106.405 69.815 106.615 70.635 ;
        RECT 106.785 69.835 107.115 70.465 ;
        RECT 102.815 68.935 103.825 69.105 ;
        RECT 103.995 69.090 104.745 69.280 ;
        RECT 102.475 68.595 103.600 68.765 ;
        RECT 103.995 68.425 104.165 69.090 ;
        RECT 104.915 68.845 105.255 69.655 ;
        RECT 106.785 69.235 107.035 69.835 ;
        RECT 107.285 69.815 107.515 70.635 ;
        RECT 108.645 69.910 108.935 70.635 ;
        RECT 109.105 70.090 114.450 70.635 ;
        RECT 107.205 69.395 107.535 69.645 ;
        RECT 110.690 69.260 111.030 70.090 ;
        RECT 115.360 69.825 115.605 70.430 ;
        RECT 115.825 70.100 116.335 70.635 ;
        RECT 102.135 68.255 104.165 68.425 ;
        RECT 104.335 68.085 104.505 68.845 ;
        RECT 104.740 68.435 105.255 68.845 ;
        RECT 106.405 68.085 106.615 69.225 ;
        RECT 106.785 68.255 107.115 69.235 ;
        RECT 107.285 68.085 107.515 69.225 ;
        RECT 108.645 68.085 108.935 69.250 ;
        RECT 112.510 68.520 112.860 69.770 ;
        RECT 115.085 69.655 116.315 69.825 ;
        RECT 115.085 68.845 115.425 69.655 ;
        RECT 115.595 69.090 116.345 69.280 ;
        RECT 109.105 68.085 114.450 68.520 ;
        RECT 115.085 68.435 115.600 68.845 ;
        RECT 115.835 68.085 116.005 68.845 ;
        RECT 116.175 68.425 116.345 69.090 ;
        RECT 116.515 69.105 116.705 70.465 ;
        RECT 116.875 69.615 117.150 70.465 ;
        RECT 117.340 70.100 117.870 70.465 ;
        RECT 118.295 70.235 118.625 70.635 ;
        RECT 117.695 70.065 117.870 70.100 ;
        RECT 116.875 69.445 117.155 69.615 ;
        RECT 116.875 69.305 117.150 69.445 ;
        RECT 117.355 69.105 117.525 69.905 ;
        RECT 116.515 68.935 117.525 69.105 ;
        RECT 117.695 69.895 118.625 70.065 ;
        RECT 118.795 69.895 119.050 70.465 ;
        RECT 117.695 68.765 117.865 69.895 ;
        RECT 118.455 69.725 118.625 69.895 ;
        RECT 116.740 68.595 117.865 68.765 ;
        RECT 118.035 69.395 118.230 69.725 ;
        RECT 118.455 69.395 118.710 69.725 ;
        RECT 118.035 68.425 118.205 69.395 ;
        RECT 118.880 69.225 119.050 69.895 ;
        RECT 119.225 69.865 122.735 70.635 ;
        RECT 122.905 69.885 124.115 70.635 ;
        RECT 124.285 69.885 125.495 70.635 ;
        RECT 119.225 69.345 120.875 69.865 ;
        RECT 116.175 68.255 118.205 68.425 ;
        RECT 118.375 68.085 118.545 69.225 ;
        RECT 118.715 68.255 119.050 69.225 ;
        RECT 121.045 69.175 122.735 69.695 ;
        RECT 122.905 69.345 123.425 69.885 ;
        RECT 123.595 69.175 124.115 69.715 ;
        RECT 119.225 68.085 122.735 69.175 ;
        RECT 122.905 68.085 124.115 69.175 ;
        RECT 124.285 69.175 124.805 69.715 ;
        RECT 124.975 69.345 125.495 69.885 ;
        RECT 124.285 68.085 125.495 69.175 ;
        RECT 5.520 67.915 125.580 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 6.985 66.825 10.495 67.915 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 6.985 66.135 8.635 66.655 ;
        RECT 8.805 66.305 10.495 66.825 ;
        RECT 10.665 66.775 11.050 67.745 ;
        RECT 11.220 67.455 11.545 67.915 ;
        RECT 12.065 67.285 12.345 67.745 ;
        RECT 11.220 67.065 12.345 67.285 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 6.985 65.365 10.495 66.135 ;
        RECT 10.665 66.105 10.945 66.775 ;
        RECT 11.220 66.605 11.670 67.065 ;
        RECT 12.535 66.895 12.935 67.745 ;
        RECT 13.335 67.455 13.605 67.915 ;
        RECT 13.775 67.285 14.060 67.745 ;
        RECT 11.115 66.275 11.670 66.605 ;
        RECT 11.840 66.335 12.935 66.895 ;
        RECT 11.220 66.165 11.670 66.275 ;
        RECT 10.665 65.535 11.050 66.105 ;
        RECT 11.220 65.995 12.345 66.165 ;
        RECT 11.220 65.365 11.545 65.825 ;
        RECT 12.065 65.535 12.345 65.995 ;
        RECT 12.535 65.535 12.935 66.335 ;
        RECT 13.105 67.065 14.060 67.285 ;
        RECT 13.105 66.165 13.315 67.065 ;
        RECT 13.485 66.335 14.175 66.895 ;
        RECT 14.350 66.775 14.685 67.745 ;
        RECT 14.855 66.775 15.025 67.915 ;
        RECT 15.195 67.575 17.225 67.745 ;
        RECT 13.105 65.995 14.060 66.165 ;
        RECT 13.335 65.365 13.605 65.825 ;
        RECT 13.775 65.535 14.060 65.995 ;
        RECT 14.350 66.105 14.520 66.775 ;
        RECT 15.195 66.605 15.365 67.575 ;
        RECT 14.690 66.275 14.945 66.605 ;
        RECT 15.170 66.275 15.365 66.605 ;
        RECT 15.535 67.235 16.660 67.405 ;
        RECT 14.775 66.105 14.945 66.275 ;
        RECT 15.535 66.105 15.705 67.235 ;
        RECT 14.350 65.535 14.605 66.105 ;
        RECT 14.775 65.935 15.705 66.105 ;
        RECT 15.875 66.895 16.885 67.065 ;
        RECT 15.875 66.095 16.045 66.895 ;
        RECT 16.250 66.555 16.525 66.695 ;
        RECT 16.245 66.385 16.525 66.555 ;
        RECT 15.530 65.900 15.705 65.935 ;
        RECT 14.775 65.365 15.105 65.765 ;
        RECT 15.530 65.535 16.060 65.900 ;
        RECT 16.250 65.535 16.525 66.385 ;
        RECT 16.695 65.535 16.885 66.895 ;
        RECT 17.055 66.910 17.225 67.575 ;
        RECT 17.395 67.155 17.565 67.915 ;
        RECT 17.800 67.155 18.315 67.565 ;
        RECT 17.055 66.720 17.805 66.910 ;
        RECT 17.975 66.345 18.315 67.155 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.950 66.775 19.285 67.745 ;
        RECT 19.455 66.775 19.625 67.915 ;
        RECT 19.795 67.575 21.825 67.745 ;
        RECT 17.085 66.175 18.315 66.345 ;
        RECT 17.065 65.365 17.575 65.900 ;
        RECT 17.795 65.570 18.040 66.175 ;
        RECT 18.950 66.105 19.120 66.775 ;
        RECT 19.795 66.605 19.965 67.575 ;
        RECT 19.290 66.275 19.545 66.605 ;
        RECT 19.770 66.275 19.965 66.605 ;
        RECT 20.135 67.235 21.260 67.405 ;
        RECT 19.375 66.105 19.545 66.275 ;
        RECT 20.135 66.105 20.305 67.235 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 18.950 65.535 19.205 66.105 ;
        RECT 19.375 65.935 20.305 66.105 ;
        RECT 20.475 66.895 21.485 67.065 ;
        RECT 20.475 66.095 20.645 66.895 ;
        RECT 20.850 66.555 21.125 66.695 ;
        RECT 20.845 66.385 21.125 66.555 ;
        RECT 20.130 65.900 20.305 65.935 ;
        RECT 19.375 65.365 19.705 65.765 ;
        RECT 20.130 65.535 20.660 65.900 ;
        RECT 20.850 65.535 21.125 66.385 ;
        RECT 21.295 65.535 21.485 66.895 ;
        RECT 21.655 66.910 21.825 67.575 ;
        RECT 21.995 67.155 22.165 67.915 ;
        RECT 22.400 67.155 22.915 67.565 ;
        RECT 21.655 66.720 22.405 66.910 ;
        RECT 22.575 66.345 22.915 67.155 ;
        RECT 24.120 67.285 24.405 67.745 ;
        RECT 24.575 67.455 24.845 67.915 ;
        RECT 24.120 67.065 25.075 67.285 ;
        RECT 21.685 66.175 22.915 66.345 ;
        RECT 24.005 66.335 24.695 66.895 ;
        RECT 21.665 65.365 22.175 65.900 ;
        RECT 22.395 65.570 22.640 66.175 ;
        RECT 24.865 66.165 25.075 67.065 ;
        RECT 24.120 65.995 25.075 66.165 ;
        RECT 25.245 66.895 25.645 67.745 ;
        RECT 25.835 67.285 26.115 67.745 ;
        RECT 26.635 67.455 26.960 67.915 ;
        RECT 25.835 67.065 26.960 67.285 ;
        RECT 25.245 66.335 26.340 66.895 ;
        RECT 26.510 66.605 26.960 67.065 ;
        RECT 27.130 66.775 27.515 67.745 ;
        RECT 27.800 67.285 28.085 67.745 ;
        RECT 28.255 67.455 28.525 67.915 ;
        RECT 27.800 67.065 28.755 67.285 ;
        RECT 24.120 65.535 24.405 65.995 ;
        RECT 24.575 65.365 24.845 65.825 ;
        RECT 25.245 65.535 25.645 66.335 ;
        RECT 26.510 66.275 27.065 66.605 ;
        RECT 26.510 66.165 26.960 66.275 ;
        RECT 25.835 65.995 26.960 66.165 ;
        RECT 27.235 66.105 27.515 66.775 ;
        RECT 27.685 66.335 28.375 66.895 ;
        RECT 28.545 66.165 28.755 67.065 ;
        RECT 25.835 65.535 26.115 65.995 ;
        RECT 26.635 65.365 26.960 65.825 ;
        RECT 27.130 65.535 27.515 66.105 ;
        RECT 27.800 65.995 28.755 66.165 ;
        RECT 28.925 66.895 29.325 67.745 ;
        RECT 29.515 67.285 29.795 67.745 ;
        RECT 30.315 67.455 30.640 67.915 ;
        RECT 29.515 67.065 30.640 67.285 ;
        RECT 28.925 66.335 30.020 66.895 ;
        RECT 30.190 66.605 30.640 67.065 ;
        RECT 30.810 66.775 31.195 67.745 ;
        RECT 27.800 65.535 28.085 65.995 ;
        RECT 28.255 65.365 28.525 65.825 ;
        RECT 28.925 65.535 29.325 66.335 ;
        RECT 30.190 66.275 30.745 66.605 ;
        RECT 30.190 66.165 30.640 66.275 ;
        RECT 29.515 65.995 30.640 66.165 ;
        RECT 30.915 66.105 31.195 66.775 ;
        RECT 29.515 65.535 29.795 65.995 ;
        RECT 30.315 65.365 30.640 65.825 ;
        RECT 30.810 65.535 31.195 66.105 ;
        RECT 31.370 66.775 31.705 67.745 ;
        RECT 31.875 66.775 32.045 67.915 ;
        RECT 32.215 67.575 34.245 67.745 ;
        RECT 31.370 66.105 31.540 66.775 ;
        RECT 32.215 66.605 32.385 67.575 ;
        RECT 31.710 66.275 31.965 66.605 ;
        RECT 32.190 66.275 32.385 66.605 ;
        RECT 32.555 67.235 33.680 67.405 ;
        RECT 31.795 66.105 31.965 66.275 ;
        RECT 32.555 66.105 32.725 67.235 ;
        RECT 31.370 65.535 31.625 66.105 ;
        RECT 31.795 65.935 32.725 66.105 ;
        RECT 32.895 66.895 33.905 67.065 ;
        RECT 32.895 66.095 33.065 66.895 ;
        RECT 32.550 65.900 32.725 65.935 ;
        RECT 31.795 65.365 32.125 65.765 ;
        RECT 32.550 65.535 33.080 65.900 ;
        RECT 33.270 65.875 33.545 66.695 ;
        RECT 33.265 65.705 33.545 65.875 ;
        RECT 33.270 65.535 33.545 65.705 ;
        RECT 33.715 65.535 33.905 66.895 ;
        RECT 34.075 66.910 34.245 67.575 ;
        RECT 34.415 67.155 34.585 67.915 ;
        RECT 34.820 67.155 35.335 67.565 ;
        RECT 34.075 66.720 34.825 66.910 ;
        RECT 34.995 66.345 35.335 67.155 ;
        RECT 35.545 66.775 35.775 67.915 ;
        RECT 35.945 66.765 36.275 67.745 ;
        RECT 36.445 66.775 36.655 67.915 ;
        RECT 36.885 67.480 42.230 67.915 ;
        RECT 35.525 66.355 35.855 66.605 ;
        RECT 34.105 66.175 35.335 66.345 ;
        RECT 34.085 65.365 34.595 65.900 ;
        RECT 34.815 65.570 35.060 66.175 ;
        RECT 35.545 65.365 35.775 66.185 ;
        RECT 36.025 66.165 36.275 66.765 ;
        RECT 35.945 65.535 36.275 66.165 ;
        RECT 36.445 65.365 36.655 66.185 ;
        RECT 38.470 65.910 38.810 66.740 ;
        RECT 40.290 66.230 40.640 67.480 ;
        RECT 42.405 66.825 44.075 67.915 ;
        RECT 42.405 66.135 43.155 66.655 ;
        RECT 43.325 66.305 44.075 66.825 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.745 66.775 44.975 67.915 ;
        RECT 45.145 66.765 45.475 67.745 ;
        RECT 45.645 66.775 45.855 67.915 ;
        RECT 46.085 66.825 47.295 67.915 ;
        RECT 44.725 66.355 45.055 66.605 ;
        RECT 36.885 65.365 42.230 65.910 ;
        RECT 42.405 65.365 44.075 66.135 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 44.745 65.365 44.975 66.185 ;
        RECT 45.225 66.165 45.475 66.765 ;
        RECT 45.145 65.535 45.475 66.165 ;
        RECT 45.645 65.365 45.855 66.185 ;
        RECT 46.085 66.115 46.605 66.655 ;
        RECT 46.775 66.285 47.295 66.825 ;
        RECT 47.505 66.775 47.735 67.915 ;
        RECT 47.905 66.765 48.235 67.745 ;
        RECT 48.405 66.775 48.615 67.915 ;
        RECT 48.845 66.840 49.115 67.745 ;
        RECT 49.285 67.155 49.615 67.915 ;
        RECT 49.795 66.985 49.965 67.745 ;
        RECT 47.485 66.355 47.815 66.605 ;
        RECT 46.085 65.365 47.295 66.115 ;
        RECT 47.505 65.365 47.735 66.185 ;
        RECT 47.985 66.165 48.235 66.765 ;
        RECT 47.905 65.535 48.235 66.165 ;
        RECT 48.405 65.365 48.615 66.185 ;
        RECT 48.845 66.040 49.015 66.840 ;
        RECT 49.300 66.815 49.965 66.985 ;
        RECT 49.300 66.670 49.470 66.815 ;
        RECT 49.185 66.340 49.470 66.670 ;
        RECT 51.150 66.775 51.485 67.745 ;
        RECT 51.655 66.775 51.825 67.915 ;
        RECT 51.995 67.575 54.025 67.745 ;
        RECT 49.300 66.085 49.470 66.340 ;
        RECT 49.705 66.265 50.035 66.635 ;
        RECT 51.150 66.105 51.320 66.775 ;
        RECT 51.995 66.605 52.165 67.575 ;
        RECT 51.490 66.275 51.745 66.605 ;
        RECT 51.970 66.275 52.165 66.605 ;
        RECT 52.335 67.235 53.460 67.405 ;
        RECT 51.575 66.105 51.745 66.275 ;
        RECT 52.335 66.105 52.505 67.235 ;
        RECT 48.845 65.535 49.105 66.040 ;
        RECT 49.300 65.915 49.965 66.085 ;
        RECT 49.285 65.365 49.615 65.745 ;
        RECT 49.795 65.535 49.965 65.915 ;
        RECT 51.150 65.535 51.405 66.105 ;
        RECT 51.575 65.935 52.505 66.105 ;
        RECT 52.675 66.895 53.685 67.065 ;
        RECT 52.675 66.095 52.845 66.895 ;
        RECT 53.050 66.555 53.325 66.695 ;
        RECT 53.045 66.385 53.325 66.555 ;
        RECT 52.330 65.900 52.505 65.935 ;
        RECT 51.575 65.365 51.905 65.765 ;
        RECT 52.330 65.535 52.860 65.900 ;
        RECT 53.050 65.535 53.325 66.385 ;
        RECT 53.495 65.535 53.685 66.895 ;
        RECT 53.855 66.910 54.025 67.575 ;
        RECT 54.195 67.155 54.365 67.915 ;
        RECT 54.600 67.155 55.115 67.565 ;
        RECT 55.285 67.480 60.630 67.915 ;
        RECT 53.855 66.720 54.605 66.910 ;
        RECT 54.775 66.345 55.115 67.155 ;
        RECT 53.885 66.175 55.115 66.345 ;
        RECT 53.865 65.365 54.375 65.900 ;
        RECT 54.595 65.570 54.840 66.175 ;
        RECT 56.870 65.910 57.210 66.740 ;
        RECT 58.690 66.230 59.040 67.480 ;
        RECT 61.355 66.985 61.525 67.745 ;
        RECT 61.740 67.155 62.070 67.915 ;
        RECT 61.355 66.815 62.070 66.985 ;
        RECT 62.240 66.840 62.495 67.745 ;
        RECT 61.265 66.265 61.620 66.635 ;
        RECT 61.900 66.605 62.070 66.815 ;
        RECT 61.900 66.275 62.155 66.605 ;
        RECT 61.900 66.085 62.070 66.275 ;
        RECT 62.325 66.110 62.495 66.840 ;
        RECT 62.670 66.765 62.930 67.915 ;
        RECT 63.115 66.935 63.445 67.745 ;
        RECT 63.615 67.115 63.855 67.915 ;
        RECT 63.115 66.765 63.830 66.935 ;
        RECT 63.110 66.355 63.490 66.595 ;
        RECT 63.660 66.525 63.830 66.765 ;
        RECT 64.035 66.895 64.205 67.745 ;
        RECT 64.375 67.115 64.705 67.915 ;
        RECT 64.875 66.895 65.045 67.745 ;
        RECT 64.035 66.725 65.045 66.895 ;
        RECT 65.215 66.765 65.545 67.915 ;
        RECT 65.865 66.945 66.175 67.745 ;
        RECT 66.345 67.115 66.655 67.915 ;
        RECT 66.825 67.285 67.085 67.745 ;
        RECT 67.255 67.455 67.510 67.915 ;
        RECT 67.685 67.285 67.945 67.745 ;
        RECT 66.825 67.115 67.945 67.285 ;
        RECT 65.865 66.775 66.895 66.945 ;
        RECT 64.550 66.555 65.045 66.725 ;
        RECT 63.660 66.355 64.160 66.525 ;
        RECT 64.545 66.385 65.045 66.555 ;
        RECT 61.355 65.915 62.070 66.085 ;
        RECT 55.285 65.365 60.630 65.910 ;
        RECT 61.355 65.535 61.525 65.915 ;
        RECT 61.740 65.365 62.070 65.745 ;
        RECT 62.240 65.535 62.495 66.110 ;
        RECT 62.670 65.365 62.930 66.205 ;
        RECT 63.660 66.185 63.830 66.355 ;
        RECT 64.550 66.185 65.045 66.385 ;
        RECT 63.195 66.015 63.830 66.185 ;
        RECT 64.035 66.015 65.045 66.185 ;
        RECT 63.195 65.535 63.365 66.015 ;
        RECT 63.545 65.365 63.785 65.845 ;
        RECT 64.035 65.535 64.205 66.015 ;
        RECT 64.375 65.365 64.705 65.845 ;
        RECT 64.875 65.535 65.045 66.015 ;
        RECT 65.215 65.365 65.545 66.165 ;
        RECT 65.865 65.865 66.035 66.775 ;
        RECT 66.205 66.035 66.555 66.605 ;
        RECT 66.725 66.525 66.895 66.775 ;
        RECT 67.685 66.865 67.945 67.115 ;
        RECT 68.115 67.045 68.400 67.915 ;
        RECT 68.715 66.985 68.885 67.745 ;
        RECT 69.065 67.155 69.395 67.915 ;
        RECT 67.685 66.695 68.440 66.865 ;
        RECT 68.715 66.815 69.380 66.985 ;
        RECT 69.565 66.840 69.835 67.745 ;
        RECT 66.725 66.355 67.865 66.525 ;
        RECT 68.035 66.185 68.440 66.695 ;
        RECT 69.210 66.670 69.380 66.815 ;
        RECT 68.645 66.265 68.975 66.635 ;
        RECT 69.210 66.340 69.495 66.670 ;
        RECT 66.790 66.015 68.440 66.185 ;
        RECT 69.210 66.085 69.380 66.340 ;
        RECT 65.865 65.535 66.165 65.865 ;
        RECT 66.335 65.365 66.610 65.845 ;
        RECT 66.790 65.625 67.085 66.015 ;
        RECT 67.255 65.365 67.510 65.845 ;
        RECT 67.685 65.625 67.945 66.015 ;
        RECT 68.715 65.915 69.380 66.085 ;
        RECT 69.665 66.040 69.835 66.840 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 70.470 67.245 70.725 67.745 ;
        RECT 70.895 67.415 71.225 67.915 ;
        RECT 70.470 67.075 71.220 67.245 ;
        RECT 70.470 66.255 70.820 66.905 ;
        RECT 68.115 65.365 68.395 65.845 ;
        RECT 68.715 65.535 68.885 65.915 ;
        RECT 69.065 65.365 69.395 65.745 ;
        RECT 69.575 65.535 69.835 66.040 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 70.990 66.085 71.220 67.075 ;
        RECT 70.470 65.915 71.220 66.085 ;
        RECT 70.470 65.625 70.725 65.915 ;
        RECT 70.895 65.365 71.225 65.745 ;
        RECT 71.395 65.625 71.565 67.745 ;
        RECT 71.735 66.945 72.060 67.730 ;
        RECT 72.230 67.455 72.480 67.915 ;
        RECT 72.650 67.415 72.900 67.745 ;
        RECT 73.115 67.415 73.795 67.745 ;
        RECT 72.650 67.285 72.820 67.415 ;
        RECT 72.425 67.115 72.820 67.285 ;
        RECT 71.795 65.895 72.255 66.945 ;
        RECT 72.425 65.755 72.595 67.115 ;
        RECT 72.990 66.855 73.455 67.245 ;
        RECT 72.765 66.045 73.115 66.665 ;
        RECT 73.285 66.265 73.455 66.855 ;
        RECT 73.625 66.635 73.795 67.415 ;
        RECT 73.965 67.315 74.135 67.655 ;
        RECT 74.370 67.485 74.700 67.915 ;
        RECT 74.870 67.315 75.040 67.655 ;
        RECT 75.335 67.455 75.705 67.915 ;
        RECT 73.965 67.145 75.040 67.315 ;
        RECT 75.875 67.285 76.045 67.745 ;
        RECT 76.280 67.405 77.150 67.745 ;
        RECT 77.320 67.455 77.570 67.915 ;
        RECT 75.485 67.115 76.045 67.285 ;
        RECT 75.485 66.975 75.655 67.115 ;
        RECT 74.155 66.805 75.655 66.975 ;
        RECT 76.350 66.945 76.810 67.235 ;
        RECT 73.625 66.465 75.315 66.635 ;
        RECT 73.285 66.045 73.640 66.265 ;
        RECT 73.810 65.755 73.980 66.465 ;
        RECT 74.185 66.045 74.975 66.295 ;
        RECT 75.145 66.285 75.315 66.465 ;
        RECT 75.485 66.115 75.655 66.805 ;
        RECT 71.925 65.365 72.255 65.725 ;
        RECT 72.425 65.585 72.920 65.755 ;
        RECT 73.125 65.585 73.980 65.755 ;
        RECT 74.855 65.365 75.185 65.825 ;
        RECT 75.395 65.725 75.655 66.115 ;
        RECT 75.845 66.935 76.810 66.945 ;
        RECT 76.980 67.025 77.150 67.405 ;
        RECT 77.740 67.365 77.910 67.655 ;
        RECT 78.090 67.535 78.420 67.915 ;
        RECT 77.740 67.195 78.540 67.365 ;
        RECT 75.845 66.775 76.520 66.935 ;
        RECT 76.980 66.855 78.200 67.025 ;
        RECT 75.845 65.985 76.055 66.775 ;
        RECT 76.980 66.765 77.150 66.855 ;
        RECT 76.225 65.985 76.575 66.605 ;
        RECT 76.745 66.595 77.150 66.765 ;
        RECT 76.745 65.815 76.915 66.595 ;
        RECT 77.085 66.145 77.305 66.425 ;
        RECT 77.485 66.315 78.025 66.685 ;
        RECT 78.370 66.605 78.540 67.195 ;
        RECT 78.760 66.775 79.065 67.915 ;
        RECT 79.235 66.725 79.490 67.605 ;
        RECT 78.370 66.575 79.110 66.605 ;
        RECT 77.085 65.975 77.615 66.145 ;
        RECT 75.395 65.555 75.745 65.725 ;
        RECT 75.965 65.535 76.915 65.815 ;
        RECT 77.085 65.365 77.275 65.805 ;
        RECT 77.445 65.745 77.615 65.975 ;
        RECT 77.785 65.915 78.025 66.315 ;
        RECT 78.195 66.275 79.110 66.575 ;
        RECT 78.195 66.100 78.520 66.275 ;
        RECT 78.195 65.745 78.515 66.100 ;
        RECT 79.280 66.075 79.490 66.725 ;
        RECT 77.445 65.575 78.515 65.745 ;
        RECT 78.760 65.365 79.065 65.825 ;
        RECT 79.235 65.545 79.490 66.075 ;
        RECT 79.670 66.775 80.005 67.745 ;
        RECT 80.175 66.775 80.345 67.915 ;
        RECT 80.515 67.575 82.545 67.745 ;
        RECT 79.670 66.105 79.840 66.775 ;
        RECT 80.515 66.605 80.685 67.575 ;
        RECT 80.010 66.275 80.265 66.605 ;
        RECT 80.490 66.275 80.685 66.605 ;
        RECT 80.855 67.235 81.980 67.405 ;
        RECT 80.095 66.105 80.265 66.275 ;
        RECT 80.855 66.105 81.025 67.235 ;
        RECT 79.670 65.535 79.925 66.105 ;
        RECT 80.095 65.935 81.025 66.105 ;
        RECT 81.195 66.895 82.205 67.065 ;
        RECT 81.195 66.095 81.365 66.895 ;
        RECT 81.570 66.555 81.845 66.695 ;
        RECT 81.565 66.385 81.845 66.555 ;
        RECT 80.850 65.900 81.025 65.935 ;
        RECT 80.095 65.365 80.425 65.765 ;
        RECT 80.850 65.535 81.380 65.900 ;
        RECT 81.570 65.535 81.845 66.385 ;
        RECT 82.015 65.535 82.205 66.895 ;
        RECT 82.375 66.910 82.545 67.575 ;
        RECT 82.715 67.155 82.885 67.915 ;
        RECT 83.120 67.155 83.635 67.565 ;
        RECT 82.375 66.720 83.125 66.910 ;
        RECT 83.295 66.345 83.635 67.155 ;
        RECT 82.405 66.175 83.635 66.345 ;
        RECT 83.805 66.775 84.190 67.745 ;
        RECT 84.360 67.455 84.685 67.915 ;
        RECT 85.205 67.285 85.485 67.745 ;
        RECT 84.360 67.065 85.485 67.285 ;
        RECT 82.385 65.365 82.895 65.900 ;
        RECT 83.115 65.570 83.360 66.175 ;
        RECT 83.805 66.105 84.085 66.775 ;
        RECT 84.360 66.605 84.810 67.065 ;
        RECT 85.675 66.895 86.075 67.745 ;
        RECT 86.475 67.455 86.745 67.915 ;
        RECT 86.915 67.285 87.200 67.745 ;
        RECT 84.255 66.275 84.810 66.605 ;
        RECT 84.980 66.335 86.075 66.895 ;
        RECT 84.360 66.165 84.810 66.275 ;
        RECT 83.805 65.535 84.190 66.105 ;
        RECT 84.360 65.995 85.485 66.165 ;
        RECT 84.360 65.365 84.685 65.825 ;
        RECT 85.205 65.535 85.485 65.995 ;
        RECT 85.675 65.535 86.075 66.335 ;
        RECT 86.245 67.065 87.200 67.285 ;
        RECT 87.485 67.155 88.000 67.565 ;
        RECT 88.235 67.155 88.405 67.915 ;
        RECT 88.575 67.575 90.605 67.745 ;
        RECT 86.245 66.165 86.455 67.065 ;
        RECT 86.625 66.335 87.315 66.895 ;
        RECT 87.485 66.345 87.825 67.155 ;
        RECT 88.575 66.910 88.745 67.575 ;
        RECT 89.140 67.235 90.265 67.405 ;
        RECT 87.995 66.720 88.745 66.910 ;
        RECT 88.915 66.895 89.925 67.065 ;
        RECT 87.485 66.175 88.715 66.345 ;
        RECT 86.245 65.995 87.200 66.165 ;
        RECT 86.475 65.365 86.745 65.825 ;
        RECT 86.915 65.535 87.200 65.995 ;
        RECT 87.760 65.570 88.005 66.175 ;
        RECT 88.225 65.365 88.735 65.900 ;
        RECT 88.915 65.535 89.105 66.895 ;
        RECT 89.275 65.875 89.550 66.695 ;
        RECT 89.755 66.095 89.925 66.895 ;
        RECT 90.095 66.105 90.265 67.235 ;
        RECT 90.435 66.605 90.605 67.575 ;
        RECT 90.775 66.775 90.945 67.915 ;
        RECT 91.115 66.775 91.450 67.745 ;
        RECT 91.740 67.285 92.025 67.745 ;
        RECT 92.195 67.455 92.465 67.915 ;
        RECT 91.740 67.065 92.695 67.285 ;
        RECT 90.435 66.275 90.630 66.605 ;
        RECT 90.855 66.275 91.110 66.605 ;
        RECT 90.855 66.105 91.025 66.275 ;
        RECT 91.280 66.105 91.450 66.775 ;
        RECT 91.625 66.335 92.315 66.895 ;
        RECT 92.485 66.165 92.695 67.065 ;
        RECT 90.095 65.935 91.025 66.105 ;
        RECT 90.095 65.900 90.270 65.935 ;
        RECT 89.275 65.705 89.555 65.875 ;
        RECT 89.275 65.535 89.550 65.705 ;
        RECT 89.740 65.535 90.270 65.900 ;
        RECT 90.695 65.365 91.025 65.765 ;
        RECT 91.195 65.535 91.450 66.105 ;
        RECT 91.740 65.995 92.695 66.165 ;
        RECT 92.865 66.895 93.265 67.745 ;
        RECT 93.455 67.285 93.735 67.745 ;
        RECT 94.255 67.455 94.580 67.915 ;
        RECT 93.455 67.065 94.580 67.285 ;
        RECT 92.865 66.335 93.960 66.895 ;
        RECT 94.130 66.605 94.580 67.065 ;
        RECT 94.750 66.775 95.135 67.745 ;
        RECT 91.740 65.535 92.025 65.995 ;
        RECT 92.195 65.365 92.465 65.825 ;
        RECT 92.865 65.535 93.265 66.335 ;
        RECT 94.130 66.275 94.685 66.605 ;
        RECT 94.130 66.165 94.580 66.275 ;
        RECT 93.455 65.995 94.580 66.165 ;
        RECT 94.855 66.105 95.135 66.775 ;
        RECT 95.765 66.750 96.055 67.915 ;
        RECT 96.315 67.245 96.485 67.745 ;
        RECT 96.655 67.415 96.985 67.915 ;
        RECT 96.315 67.075 96.980 67.245 ;
        RECT 96.230 66.255 96.580 66.905 ;
        RECT 93.455 65.535 93.735 65.995 ;
        RECT 94.255 65.365 94.580 65.825 ;
        RECT 94.750 65.535 95.135 66.105 ;
        RECT 95.765 65.365 96.055 66.090 ;
        RECT 96.750 66.085 96.980 67.075 ;
        RECT 96.315 65.915 96.980 66.085 ;
        RECT 96.315 65.625 96.485 65.915 ;
        RECT 96.655 65.365 96.985 65.745 ;
        RECT 97.155 65.625 97.380 67.745 ;
        RECT 97.595 67.415 97.925 67.915 ;
        RECT 98.095 67.245 98.265 67.745 ;
        RECT 98.500 67.530 99.330 67.700 ;
        RECT 99.570 67.535 99.950 67.915 ;
        RECT 97.570 67.075 98.265 67.245 ;
        RECT 97.570 66.105 97.740 67.075 ;
        RECT 97.910 66.285 98.320 66.905 ;
        RECT 98.490 66.855 98.990 67.235 ;
        RECT 97.570 65.915 98.265 66.105 ;
        RECT 98.490 65.985 98.710 66.855 ;
        RECT 99.160 66.685 99.330 67.530 ;
        RECT 100.130 67.365 100.300 67.655 ;
        RECT 100.470 67.535 100.800 67.915 ;
        RECT 101.270 67.445 101.900 67.695 ;
        RECT 102.080 67.535 102.500 67.915 ;
        RECT 101.730 67.365 101.900 67.445 ;
        RECT 102.700 67.365 102.940 67.655 ;
        RECT 99.500 67.115 100.870 67.365 ;
        RECT 99.500 66.855 99.750 67.115 ;
        RECT 100.260 66.685 100.510 66.845 ;
        RECT 99.160 66.515 100.510 66.685 ;
        RECT 99.160 66.475 99.580 66.515 ;
        RECT 98.890 65.925 99.240 66.295 ;
        RECT 97.595 65.365 97.925 65.745 ;
        RECT 98.095 65.585 98.265 65.915 ;
        RECT 99.410 65.745 99.580 66.475 ;
        RECT 100.680 66.345 100.870 67.115 ;
        RECT 99.750 66.015 100.160 66.345 ;
        RECT 100.450 66.005 100.870 66.345 ;
        RECT 101.040 66.935 101.560 67.245 ;
        RECT 101.730 67.195 102.940 67.365 ;
        RECT 103.170 67.225 103.500 67.915 ;
        RECT 101.040 66.175 101.210 66.935 ;
        RECT 101.380 66.345 101.560 66.755 ;
        RECT 101.730 66.685 101.900 67.195 ;
        RECT 103.670 67.045 103.840 67.655 ;
        RECT 104.110 67.195 104.440 67.705 ;
        RECT 103.670 67.025 103.990 67.045 ;
        RECT 102.070 66.855 103.990 67.025 ;
        RECT 101.730 66.515 103.630 66.685 ;
        RECT 101.960 66.175 102.290 66.295 ;
        RECT 101.040 66.005 102.290 66.175 ;
        RECT 98.565 65.545 99.580 65.745 ;
        RECT 99.750 65.365 100.160 65.805 ;
        RECT 100.450 65.575 100.700 66.005 ;
        RECT 100.900 65.365 101.220 65.825 ;
        RECT 102.460 65.755 102.630 66.515 ;
        RECT 103.300 66.455 103.630 66.515 ;
        RECT 102.820 66.285 103.150 66.345 ;
        RECT 102.820 66.015 103.480 66.285 ;
        RECT 103.800 65.960 103.990 66.855 ;
        RECT 101.780 65.585 102.630 65.755 ;
        RECT 102.830 65.365 103.490 65.845 ;
        RECT 103.670 65.630 103.990 65.960 ;
        RECT 104.190 66.605 104.440 67.195 ;
        RECT 104.620 67.115 104.905 67.915 ;
        RECT 105.085 67.575 105.340 67.605 ;
        RECT 105.085 67.405 105.425 67.575 ;
        RECT 105.885 67.480 111.230 67.915 ;
        RECT 105.085 66.935 105.340 67.405 ;
        RECT 104.190 66.275 104.990 66.605 ;
        RECT 104.190 65.625 104.440 66.275 ;
        RECT 105.160 66.075 105.340 66.935 ;
        RECT 104.620 65.365 104.905 65.825 ;
        RECT 105.085 65.545 105.340 66.075 ;
        RECT 107.470 65.910 107.810 66.740 ;
        RECT 109.290 66.230 109.640 67.480 ;
        RECT 111.405 66.825 113.995 67.915 ;
        RECT 111.405 66.135 112.615 66.655 ;
        RECT 112.785 66.305 113.995 66.825 ;
        RECT 114.625 67.155 115.140 67.565 ;
        RECT 115.375 67.155 115.545 67.915 ;
        RECT 115.715 67.575 117.745 67.745 ;
        RECT 114.625 66.345 114.965 67.155 ;
        RECT 115.715 66.910 115.885 67.575 ;
        RECT 116.280 67.235 117.405 67.405 ;
        RECT 115.135 66.720 115.885 66.910 ;
        RECT 116.055 66.895 117.065 67.065 ;
        RECT 114.625 66.175 115.855 66.345 ;
        RECT 105.885 65.365 111.230 65.910 ;
        RECT 111.405 65.365 113.995 66.135 ;
        RECT 114.900 65.570 115.145 66.175 ;
        RECT 115.365 65.365 115.875 65.900 ;
        RECT 116.055 65.535 116.245 66.895 ;
        RECT 116.415 66.555 116.690 66.695 ;
        RECT 116.415 66.385 116.695 66.555 ;
        RECT 116.415 65.535 116.690 66.385 ;
        RECT 116.895 66.095 117.065 66.895 ;
        RECT 117.235 66.105 117.405 67.235 ;
        RECT 117.575 66.605 117.745 67.575 ;
        RECT 117.915 66.775 118.085 67.915 ;
        RECT 118.255 66.775 118.590 67.745 ;
        RECT 117.575 66.275 117.770 66.605 ;
        RECT 117.995 66.275 118.250 66.605 ;
        RECT 117.995 66.105 118.165 66.275 ;
        RECT 118.420 66.105 118.590 66.775 ;
        RECT 117.235 65.935 118.165 66.105 ;
        RECT 117.235 65.900 117.410 65.935 ;
        RECT 116.880 65.535 117.410 65.900 ;
        RECT 117.835 65.365 118.165 65.765 ;
        RECT 118.335 65.535 118.590 66.105 ;
        RECT 118.765 66.840 119.035 67.745 ;
        RECT 119.205 67.155 119.535 67.915 ;
        RECT 119.715 66.985 119.885 67.745 ;
        RECT 118.765 66.040 118.935 66.840 ;
        RECT 119.220 66.815 119.885 66.985 ;
        RECT 119.220 66.670 119.390 66.815 ;
        RECT 120.205 66.775 120.415 67.915 ;
        RECT 119.105 66.340 119.390 66.670 ;
        RECT 120.585 66.765 120.915 67.745 ;
        RECT 121.085 66.775 121.315 67.915 ;
        RECT 119.220 66.085 119.390 66.340 ;
        RECT 119.625 66.265 119.955 66.635 ;
        RECT 118.765 65.535 119.025 66.040 ;
        RECT 119.220 65.915 119.885 66.085 ;
        RECT 119.205 65.365 119.535 65.745 ;
        RECT 119.715 65.535 119.885 65.915 ;
        RECT 120.205 65.365 120.415 66.185 ;
        RECT 120.585 66.165 120.835 66.765 ;
        RECT 121.525 66.750 121.815 67.915 ;
        RECT 121.985 66.825 123.655 67.915 ;
        RECT 121.005 66.355 121.335 66.605 ;
        RECT 120.585 65.535 120.915 66.165 ;
        RECT 121.085 65.365 121.315 66.185 ;
        RECT 121.985 66.135 122.735 66.655 ;
        RECT 122.905 66.305 123.655 66.825 ;
        RECT 124.285 66.825 125.495 67.915 ;
        RECT 124.285 66.285 124.805 66.825 ;
        RECT 121.525 65.365 121.815 66.090 ;
        RECT 121.985 65.365 123.655 66.135 ;
        RECT 124.975 66.115 125.495 66.655 ;
        RECT 124.285 65.365 125.495 66.115 ;
        RECT 5.520 65.195 125.580 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.985 64.425 9.575 65.195 ;
        RECT 9.745 64.520 10.005 65.025 ;
        RECT 10.185 64.815 10.515 65.195 ;
        RECT 10.695 64.645 10.865 65.025 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 6.985 63.905 8.195 64.425 ;
        RECT 8.365 63.735 9.575 64.255 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 6.985 62.645 9.575 63.735 ;
        RECT 9.745 63.720 9.915 64.520 ;
        RECT 10.200 64.475 10.865 64.645 ;
        RECT 11.215 64.645 11.385 65.025 ;
        RECT 11.565 64.815 11.895 65.195 ;
        RECT 11.215 64.475 11.880 64.645 ;
        RECT 12.075 64.520 12.335 65.025 ;
        RECT 10.200 64.220 10.370 64.475 ;
        RECT 10.085 63.890 10.370 64.220 ;
        RECT 10.605 63.925 10.935 64.295 ;
        RECT 11.145 63.925 11.475 64.295 ;
        RECT 11.710 64.220 11.880 64.475 ;
        RECT 10.200 63.745 10.370 63.890 ;
        RECT 11.710 63.890 11.995 64.220 ;
        RECT 11.710 63.745 11.880 63.890 ;
        RECT 9.745 62.815 10.015 63.720 ;
        RECT 10.200 63.575 10.865 63.745 ;
        RECT 10.185 62.645 10.515 63.405 ;
        RECT 10.695 62.815 10.865 63.575 ;
        RECT 11.215 63.575 11.880 63.745 ;
        RECT 12.165 63.720 12.335 64.520 ;
        RECT 12.510 64.645 12.765 64.935 ;
        RECT 12.935 64.815 13.265 65.195 ;
        RECT 12.510 64.475 13.260 64.645 ;
        RECT 11.215 62.815 11.385 63.575 ;
        RECT 11.565 62.645 11.895 63.405 ;
        RECT 12.065 62.815 12.335 63.720 ;
        RECT 12.510 63.655 12.860 64.305 ;
        RECT 13.030 63.485 13.260 64.475 ;
        RECT 12.510 63.315 13.260 63.485 ;
        RECT 12.510 62.815 12.765 63.315 ;
        RECT 12.935 62.645 13.265 63.145 ;
        RECT 13.435 62.815 13.605 64.935 ;
        RECT 13.965 64.835 14.295 65.195 ;
        RECT 14.465 64.805 14.960 64.975 ;
        RECT 15.165 64.805 16.020 64.975 ;
        RECT 13.835 63.615 14.295 64.665 ;
        RECT 13.775 62.830 14.100 63.615 ;
        RECT 14.465 63.445 14.635 64.805 ;
        RECT 14.805 63.895 15.155 64.515 ;
        RECT 15.325 64.295 15.680 64.515 ;
        RECT 15.325 63.705 15.495 64.295 ;
        RECT 15.850 64.095 16.020 64.805 ;
        RECT 16.895 64.735 17.225 65.195 ;
        RECT 17.435 64.835 17.785 65.005 ;
        RECT 16.225 64.265 17.015 64.515 ;
        RECT 17.435 64.445 17.695 64.835 ;
        RECT 18.005 64.745 18.955 65.025 ;
        RECT 19.125 64.755 19.315 65.195 ;
        RECT 19.485 64.815 20.555 64.985 ;
        RECT 17.185 64.095 17.355 64.275 ;
        RECT 14.465 63.275 14.860 63.445 ;
        RECT 15.030 63.315 15.495 63.705 ;
        RECT 15.665 63.925 17.355 64.095 ;
        RECT 14.690 63.145 14.860 63.275 ;
        RECT 15.665 63.145 15.835 63.925 ;
        RECT 17.525 63.755 17.695 64.445 ;
        RECT 16.195 63.585 17.695 63.755 ;
        RECT 17.885 63.785 18.095 64.575 ;
        RECT 18.265 63.955 18.615 64.575 ;
        RECT 18.785 63.965 18.955 64.745 ;
        RECT 19.485 64.585 19.655 64.815 ;
        RECT 19.125 64.415 19.655 64.585 ;
        RECT 19.125 64.135 19.345 64.415 ;
        RECT 19.825 64.245 20.065 64.645 ;
        RECT 18.785 63.795 19.190 63.965 ;
        RECT 19.525 63.875 20.065 64.245 ;
        RECT 20.235 64.460 20.555 64.815 ;
        RECT 20.800 64.735 21.105 65.195 ;
        RECT 21.275 64.485 21.530 65.015 ;
        RECT 22.180 64.670 22.475 65.195 ;
        RECT 20.235 64.285 20.560 64.460 ;
        RECT 20.235 63.985 21.150 64.285 ;
        RECT 20.410 63.955 21.150 63.985 ;
        RECT 17.885 63.625 18.560 63.785 ;
        RECT 19.020 63.705 19.190 63.795 ;
        RECT 17.885 63.615 18.850 63.625 ;
        RECT 17.525 63.445 17.695 63.585 ;
        RECT 14.270 62.645 14.520 63.105 ;
        RECT 14.690 62.815 14.940 63.145 ;
        RECT 15.155 62.815 15.835 63.145 ;
        RECT 16.005 63.245 17.080 63.415 ;
        RECT 17.525 63.275 18.085 63.445 ;
        RECT 18.390 63.325 18.850 63.615 ;
        RECT 19.020 63.535 20.240 63.705 ;
        RECT 16.005 62.905 16.175 63.245 ;
        RECT 16.410 62.645 16.740 63.075 ;
        RECT 16.910 62.905 17.080 63.245 ;
        RECT 17.375 62.645 17.745 63.105 ;
        RECT 17.915 62.815 18.085 63.275 ;
        RECT 19.020 63.155 19.190 63.535 ;
        RECT 20.410 63.365 20.580 63.955 ;
        RECT 21.320 63.835 21.530 64.485 ;
        RECT 22.645 64.555 22.870 65.000 ;
        RECT 23.040 64.725 23.370 65.195 ;
        RECT 22.645 64.385 23.375 64.555 ;
        RECT 24.740 64.385 24.985 64.990 ;
        RECT 25.205 64.660 25.715 65.195 ;
        RECT 21.705 63.990 22.925 64.215 ;
        RECT 18.320 62.815 19.190 63.155 ;
        RECT 19.780 63.195 20.580 63.365 ;
        RECT 19.360 62.645 19.610 63.105 ;
        RECT 19.780 62.905 19.950 63.195 ;
        RECT 20.130 62.645 20.460 63.025 ;
        RECT 20.800 62.645 21.105 63.785 ;
        RECT 21.275 62.955 21.530 63.835 ;
        RECT 23.095 63.820 23.375 64.385 ;
        RECT 21.775 63.650 23.375 63.820 ;
        RECT 24.465 64.215 25.695 64.385 ;
        RECT 21.775 62.845 22.030 63.650 ;
        RECT 22.200 62.645 22.460 63.480 ;
        RECT 22.630 62.845 22.890 63.650 ;
        RECT 23.060 62.645 23.315 63.480 ;
        RECT 24.465 63.405 24.805 64.215 ;
        RECT 24.975 63.650 25.725 63.840 ;
        RECT 24.465 62.995 24.980 63.405 ;
        RECT 25.215 62.645 25.385 63.405 ;
        RECT 25.555 62.985 25.725 63.650 ;
        RECT 25.895 63.665 26.085 65.025 ;
        RECT 26.255 64.855 26.530 65.025 ;
        RECT 26.255 64.685 26.535 64.855 ;
        RECT 26.255 63.865 26.530 64.685 ;
        RECT 26.720 64.660 27.250 65.025 ;
        RECT 27.675 64.795 28.005 65.195 ;
        RECT 27.075 64.625 27.250 64.660 ;
        RECT 26.735 63.665 26.905 64.465 ;
        RECT 25.895 63.495 26.905 63.665 ;
        RECT 27.075 64.455 28.005 64.625 ;
        RECT 28.175 64.455 28.430 65.025 ;
        RECT 27.075 63.325 27.245 64.455 ;
        RECT 27.835 64.285 28.005 64.455 ;
        RECT 26.120 63.155 27.245 63.325 ;
        RECT 27.415 63.955 27.610 64.285 ;
        RECT 27.835 63.955 28.090 64.285 ;
        RECT 27.415 62.985 27.585 63.955 ;
        RECT 28.260 63.785 28.430 64.455 ;
        RECT 25.555 62.815 27.585 62.985 ;
        RECT 27.755 62.645 27.925 63.785 ;
        RECT 28.095 62.815 28.430 63.785 ;
        RECT 28.605 64.520 28.865 65.025 ;
        RECT 29.045 64.815 29.375 65.195 ;
        RECT 29.555 64.645 29.725 65.025 ;
        RECT 28.605 63.720 28.775 64.520 ;
        RECT 29.060 64.475 29.725 64.645 ;
        RECT 29.060 64.220 29.230 64.475 ;
        RECT 29.985 64.445 31.195 65.195 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 31.825 64.445 33.035 65.195 ;
        RECT 33.205 64.455 33.590 65.025 ;
        RECT 33.760 64.735 34.085 65.195 ;
        RECT 34.605 64.565 34.885 65.025 ;
        RECT 28.945 63.890 29.230 64.220 ;
        RECT 29.465 63.925 29.795 64.295 ;
        RECT 29.985 63.905 30.505 64.445 ;
        RECT 29.060 63.745 29.230 63.890 ;
        RECT 28.605 62.815 28.875 63.720 ;
        RECT 29.060 63.575 29.725 63.745 ;
        RECT 30.675 63.735 31.195 64.275 ;
        RECT 31.825 63.905 32.345 64.445 ;
        RECT 29.045 62.645 29.375 63.405 ;
        RECT 29.555 62.815 29.725 63.575 ;
        RECT 29.985 62.645 31.195 63.735 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 32.515 63.735 33.035 64.275 ;
        RECT 31.825 62.645 33.035 63.735 ;
        RECT 33.205 63.785 33.485 64.455 ;
        RECT 33.760 64.395 34.885 64.565 ;
        RECT 33.760 64.285 34.210 64.395 ;
        RECT 33.655 63.955 34.210 64.285 ;
        RECT 35.075 64.225 35.475 65.025 ;
        RECT 35.875 64.735 36.145 65.195 ;
        RECT 36.315 64.565 36.600 65.025 ;
        RECT 33.205 62.815 33.590 63.785 ;
        RECT 33.760 63.495 34.210 63.955 ;
        RECT 34.380 63.665 35.475 64.225 ;
        RECT 33.760 63.275 34.885 63.495 ;
        RECT 33.760 62.645 34.085 63.105 ;
        RECT 34.605 62.815 34.885 63.275 ;
        RECT 35.075 62.815 35.475 63.665 ;
        RECT 35.645 64.395 36.600 64.565 ;
        RECT 36.885 64.425 40.395 65.195 ;
        RECT 41.485 64.455 41.870 65.025 ;
        RECT 42.040 64.735 42.365 65.195 ;
        RECT 42.885 64.565 43.165 65.025 ;
        RECT 35.645 63.495 35.855 64.395 ;
        RECT 36.025 63.665 36.715 64.225 ;
        RECT 36.885 63.905 38.535 64.425 ;
        RECT 38.705 63.735 40.395 64.255 ;
        RECT 35.645 63.275 36.600 63.495 ;
        RECT 35.875 62.645 36.145 63.105 ;
        RECT 36.315 62.815 36.600 63.275 ;
        RECT 36.885 62.645 40.395 63.735 ;
        RECT 41.485 63.785 41.765 64.455 ;
        RECT 42.040 64.395 43.165 64.565 ;
        RECT 42.040 64.285 42.490 64.395 ;
        RECT 41.935 63.955 42.490 64.285 ;
        RECT 43.355 64.225 43.755 65.025 ;
        RECT 44.155 64.735 44.425 65.195 ;
        RECT 44.595 64.565 44.880 65.025 ;
        RECT 41.485 62.815 41.870 63.785 ;
        RECT 42.040 63.495 42.490 63.955 ;
        RECT 42.660 63.665 43.755 64.225 ;
        RECT 42.040 63.275 43.165 63.495 ;
        RECT 42.040 62.645 42.365 63.105 ;
        RECT 42.885 62.815 43.165 63.275 ;
        RECT 43.355 62.815 43.755 63.665 ;
        RECT 43.925 64.395 44.880 64.565 ;
        RECT 46.175 64.645 46.345 64.935 ;
        RECT 46.515 64.815 46.845 65.195 ;
        RECT 46.175 64.475 46.840 64.645 ;
        RECT 43.925 63.495 44.135 64.395 ;
        RECT 44.305 63.665 44.995 64.225 ;
        RECT 46.090 63.655 46.440 64.305 ;
        RECT 43.925 63.275 44.880 63.495 ;
        RECT 46.610 63.485 46.840 64.475 ;
        RECT 44.155 62.645 44.425 63.105 ;
        RECT 44.595 62.815 44.880 63.275 ;
        RECT 46.175 63.315 46.840 63.485 ;
        RECT 46.175 62.815 46.345 63.315 ;
        RECT 46.515 62.645 46.845 63.145 ;
        RECT 47.015 62.815 47.240 64.935 ;
        RECT 47.455 64.815 47.785 65.195 ;
        RECT 47.955 64.645 48.125 64.975 ;
        RECT 48.425 64.815 49.440 65.015 ;
        RECT 47.430 64.455 48.125 64.645 ;
        RECT 47.430 63.485 47.600 64.455 ;
        RECT 47.770 63.655 48.180 64.275 ;
        RECT 48.350 63.705 48.570 64.575 ;
        RECT 48.750 64.265 49.100 64.635 ;
        RECT 49.270 64.085 49.440 64.815 ;
        RECT 49.610 64.755 50.020 65.195 ;
        RECT 50.310 64.555 50.560 64.985 ;
        RECT 50.760 64.735 51.080 65.195 ;
        RECT 51.640 64.805 52.490 64.975 ;
        RECT 49.610 64.215 50.020 64.545 ;
        RECT 50.310 64.215 50.730 64.555 ;
        RECT 49.020 64.045 49.440 64.085 ;
        RECT 49.020 63.875 50.370 64.045 ;
        RECT 47.430 63.315 48.125 63.485 ;
        RECT 48.350 63.325 48.850 63.705 ;
        RECT 47.455 62.645 47.785 63.145 ;
        RECT 47.955 62.815 48.125 63.315 ;
        RECT 49.020 63.030 49.190 63.875 ;
        RECT 50.120 63.715 50.370 63.875 ;
        RECT 49.360 63.445 49.610 63.705 ;
        RECT 50.540 63.445 50.730 64.215 ;
        RECT 49.360 63.195 50.730 63.445 ;
        RECT 50.900 64.385 52.150 64.555 ;
        RECT 50.900 63.625 51.070 64.385 ;
        RECT 51.820 64.265 52.150 64.385 ;
        RECT 51.240 63.805 51.420 64.215 ;
        RECT 52.320 64.045 52.490 64.805 ;
        RECT 52.690 64.715 53.350 65.195 ;
        RECT 53.530 64.600 53.850 64.930 ;
        RECT 52.680 64.275 53.340 64.545 ;
        RECT 52.680 64.215 53.010 64.275 ;
        RECT 53.160 64.045 53.490 64.105 ;
        RECT 51.590 63.875 53.490 64.045 ;
        RECT 50.900 63.315 51.420 63.625 ;
        RECT 51.590 63.365 51.760 63.875 ;
        RECT 53.660 63.705 53.850 64.600 ;
        RECT 51.930 63.535 53.850 63.705 ;
        RECT 53.530 63.515 53.850 63.535 ;
        RECT 54.050 64.285 54.300 64.935 ;
        RECT 54.480 64.735 54.765 65.195 ;
        RECT 54.945 64.855 55.200 65.015 ;
        RECT 54.945 64.685 55.285 64.855 ;
        RECT 54.945 64.485 55.200 64.685 ;
        RECT 54.050 63.955 54.850 64.285 ;
        RECT 51.590 63.195 52.800 63.365 ;
        RECT 48.360 62.860 49.190 63.030 ;
        RECT 49.430 62.645 49.810 63.025 ;
        RECT 49.990 62.905 50.160 63.195 ;
        RECT 51.590 63.115 51.760 63.195 ;
        RECT 50.330 62.645 50.660 63.025 ;
        RECT 51.130 62.865 51.760 63.115 ;
        RECT 51.940 62.645 52.360 63.025 ;
        RECT 52.560 62.905 52.800 63.195 ;
        RECT 53.030 62.645 53.360 63.335 ;
        RECT 53.530 62.905 53.700 63.515 ;
        RECT 54.050 63.365 54.300 63.955 ;
        RECT 55.020 63.625 55.200 64.485 ;
        RECT 55.745 64.445 56.955 65.195 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 57.590 64.455 57.845 65.025 ;
        RECT 58.015 64.795 58.345 65.195 ;
        RECT 58.770 64.660 59.300 65.025 ;
        RECT 58.770 64.625 58.945 64.660 ;
        RECT 58.015 64.455 58.945 64.625 ;
        RECT 55.745 63.905 56.265 64.445 ;
        RECT 56.435 63.735 56.955 64.275 ;
        RECT 53.970 62.855 54.300 63.365 ;
        RECT 54.480 62.645 54.765 63.445 ;
        RECT 54.945 62.955 55.200 63.625 ;
        RECT 55.745 62.645 56.955 63.735 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 57.590 63.785 57.760 64.455 ;
        RECT 58.015 64.285 58.185 64.455 ;
        RECT 57.930 63.955 58.185 64.285 ;
        RECT 58.410 63.955 58.605 64.285 ;
        RECT 57.590 62.815 57.925 63.785 ;
        RECT 58.095 62.645 58.265 63.785 ;
        RECT 58.435 62.985 58.605 63.955 ;
        RECT 58.775 63.325 58.945 64.455 ;
        RECT 59.115 63.665 59.285 64.465 ;
        RECT 59.490 64.175 59.765 65.025 ;
        RECT 59.485 64.005 59.765 64.175 ;
        RECT 59.490 63.865 59.765 64.005 ;
        RECT 59.935 63.665 60.125 65.025 ;
        RECT 60.305 64.660 60.815 65.195 ;
        RECT 61.035 64.385 61.280 64.990 ;
        RECT 61.725 64.435 62.435 65.025 ;
        RECT 62.945 64.665 63.275 65.025 ;
        RECT 63.475 64.835 63.805 65.195 ;
        RECT 63.975 64.665 64.305 65.025 ;
        RECT 62.945 64.455 64.305 64.665 ;
        RECT 64.485 64.650 69.830 65.195 ;
        RECT 60.325 64.215 61.555 64.385 ;
        RECT 59.115 63.495 60.125 63.665 ;
        RECT 60.295 63.650 61.045 63.840 ;
        RECT 58.775 63.155 59.900 63.325 ;
        RECT 60.295 62.985 60.465 63.650 ;
        RECT 61.215 63.405 61.555 64.215 ;
        RECT 58.435 62.815 60.465 62.985 ;
        RECT 60.635 62.645 60.805 63.405 ;
        RECT 61.040 62.995 61.555 63.405 ;
        RECT 61.725 63.465 61.930 64.435 ;
        RECT 62.100 63.665 62.430 64.205 ;
        RECT 62.605 63.955 63.100 64.285 ;
        RECT 63.420 63.955 63.795 64.285 ;
        RECT 64.005 63.955 64.315 64.285 ;
        RECT 62.605 63.665 62.930 63.955 ;
        RECT 63.125 63.465 63.455 63.685 ;
        RECT 61.725 63.235 63.455 63.465 ;
        RECT 61.725 62.815 62.425 63.235 ;
        RECT 62.625 62.645 62.955 63.005 ;
        RECT 63.125 62.835 63.455 63.235 ;
        RECT 63.625 62.985 63.795 63.955 ;
        RECT 66.070 63.820 66.410 64.650 ;
        RECT 70.985 64.375 71.195 65.195 ;
        RECT 71.365 64.395 71.695 65.025 ;
        RECT 63.975 62.645 64.305 63.705 ;
        RECT 67.890 63.080 68.240 64.330 ;
        RECT 71.365 63.795 71.615 64.395 ;
        RECT 71.865 64.375 72.095 65.195 ;
        RECT 72.310 64.645 72.565 64.935 ;
        RECT 72.735 64.815 73.065 65.195 ;
        RECT 72.310 64.475 73.060 64.645 ;
        RECT 71.785 63.955 72.115 64.205 ;
        RECT 64.485 62.645 69.830 63.080 ;
        RECT 70.985 62.645 71.195 63.785 ;
        RECT 71.365 62.815 71.695 63.795 ;
        RECT 71.865 62.645 72.095 63.785 ;
        RECT 72.310 63.655 72.660 64.305 ;
        RECT 72.830 63.485 73.060 64.475 ;
        RECT 72.310 63.315 73.060 63.485 ;
        RECT 72.310 62.815 72.565 63.315 ;
        RECT 72.735 62.645 73.065 63.145 ;
        RECT 73.235 62.815 73.405 64.935 ;
        RECT 73.765 64.835 74.095 65.195 ;
        RECT 74.265 64.805 74.760 64.975 ;
        RECT 74.965 64.805 75.820 64.975 ;
        RECT 73.635 63.615 74.095 64.665 ;
        RECT 73.575 62.830 73.900 63.615 ;
        RECT 74.265 63.445 74.435 64.805 ;
        RECT 74.605 63.895 74.955 64.515 ;
        RECT 75.125 64.295 75.480 64.515 ;
        RECT 75.125 63.705 75.295 64.295 ;
        RECT 75.650 64.095 75.820 64.805 ;
        RECT 76.695 64.735 77.025 65.195 ;
        RECT 77.235 64.835 77.585 65.005 ;
        RECT 76.025 64.265 76.815 64.515 ;
        RECT 77.235 64.445 77.495 64.835 ;
        RECT 77.805 64.745 78.755 65.025 ;
        RECT 78.925 64.755 79.115 65.195 ;
        RECT 79.285 64.815 80.355 64.985 ;
        RECT 76.985 64.095 77.155 64.275 ;
        RECT 74.265 63.275 74.660 63.445 ;
        RECT 74.830 63.315 75.295 63.705 ;
        RECT 75.465 63.925 77.155 64.095 ;
        RECT 74.490 63.145 74.660 63.275 ;
        RECT 75.465 63.145 75.635 63.925 ;
        RECT 77.325 63.755 77.495 64.445 ;
        RECT 75.995 63.585 77.495 63.755 ;
        RECT 77.685 63.785 77.895 64.575 ;
        RECT 78.065 63.955 78.415 64.575 ;
        RECT 78.585 63.965 78.755 64.745 ;
        RECT 79.285 64.585 79.455 64.815 ;
        RECT 78.925 64.415 79.455 64.585 ;
        RECT 78.925 64.135 79.145 64.415 ;
        RECT 79.625 64.245 79.865 64.645 ;
        RECT 78.585 63.795 78.990 63.965 ;
        RECT 79.325 63.875 79.865 64.245 ;
        RECT 80.035 64.460 80.355 64.815 ;
        RECT 80.600 64.735 80.905 65.195 ;
        RECT 81.075 64.485 81.330 65.015 ;
        RECT 80.035 64.285 80.360 64.460 ;
        RECT 80.035 63.985 80.950 64.285 ;
        RECT 80.210 63.955 80.950 63.985 ;
        RECT 77.685 63.625 78.360 63.785 ;
        RECT 78.820 63.705 78.990 63.795 ;
        RECT 77.685 63.615 78.650 63.625 ;
        RECT 77.325 63.445 77.495 63.585 ;
        RECT 74.070 62.645 74.320 63.105 ;
        RECT 74.490 62.815 74.740 63.145 ;
        RECT 74.955 62.815 75.635 63.145 ;
        RECT 75.805 63.245 76.880 63.415 ;
        RECT 77.325 63.275 77.885 63.445 ;
        RECT 78.190 63.325 78.650 63.615 ;
        RECT 78.820 63.535 80.040 63.705 ;
        RECT 75.805 62.905 75.975 63.245 ;
        RECT 76.210 62.645 76.540 63.075 ;
        RECT 76.710 62.905 76.880 63.245 ;
        RECT 77.175 62.645 77.545 63.105 ;
        RECT 77.715 62.815 77.885 63.275 ;
        RECT 78.820 63.155 78.990 63.535 ;
        RECT 80.210 63.365 80.380 63.955 ;
        RECT 81.120 63.835 81.330 64.485 ;
        RECT 78.120 62.815 78.990 63.155 ;
        RECT 79.580 63.195 80.380 63.365 ;
        RECT 79.160 62.645 79.410 63.105 ;
        RECT 79.580 62.905 79.750 63.195 ;
        RECT 79.930 62.645 80.260 63.025 ;
        RECT 80.600 62.645 80.905 63.785 ;
        RECT 81.075 62.955 81.330 63.835 ;
        RECT 81.505 64.520 81.765 65.025 ;
        RECT 81.945 64.815 82.275 65.195 ;
        RECT 82.455 64.645 82.625 65.025 ;
        RECT 81.505 63.720 81.675 64.520 ;
        RECT 81.960 64.475 82.625 64.645 ;
        RECT 81.960 64.220 82.130 64.475 ;
        RECT 82.885 64.470 83.175 65.195 ;
        RECT 83.350 64.455 83.605 65.025 ;
        RECT 83.775 64.795 84.105 65.195 ;
        RECT 84.530 64.660 85.060 65.025 ;
        RECT 85.250 64.855 85.525 65.025 ;
        RECT 85.245 64.685 85.525 64.855 ;
        RECT 84.530 64.625 84.705 64.660 ;
        RECT 83.775 64.455 84.705 64.625 ;
        RECT 81.845 63.890 82.130 64.220 ;
        RECT 82.365 63.925 82.695 64.295 ;
        RECT 81.960 63.745 82.130 63.890 ;
        RECT 81.505 62.815 81.775 63.720 ;
        RECT 81.960 63.575 82.625 63.745 ;
        RECT 81.945 62.645 82.275 63.405 ;
        RECT 82.455 62.815 82.625 63.575 ;
        RECT 82.885 62.645 83.175 63.810 ;
        RECT 83.350 63.785 83.520 64.455 ;
        RECT 83.775 64.285 83.945 64.455 ;
        RECT 83.690 63.955 83.945 64.285 ;
        RECT 84.170 63.955 84.365 64.285 ;
        RECT 83.350 62.815 83.685 63.785 ;
        RECT 83.855 62.645 84.025 63.785 ;
        RECT 84.195 62.985 84.365 63.955 ;
        RECT 84.535 63.325 84.705 64.455 ;
        RECT 84.875 63.665 85.045 64.465 ;
        RECT 85.250 63.865 85.525 64.685 ;
        RECT 85.695 63.665 85.885 65.025 ;
        RECT 86.065 64.660 86.575 65.195 ;
        RECT 86.795 64.385 87.040 64.990 ;
        RECT 87.950 64.645 88.205 64.935 ;
        RECT 88.375 64.815 88.705 65.195 ;
        RECT 87.950 64.475 88.700 64.645 ;
        RECT 86.085 64.215 87.315 64.385 ;
        RECT 84.875 63.495 85.885 63.665 ;
        RECT 86.055 63.650 86.805 63.840 ;
        RECT 84.535 63.155 85.660 63.325 ;
        RECT 86.055 62.985 86.225 63.650 ;
        RECT 86.975 63.405 87.315 64.215 ;
        RECT 87.950 63.655 88.300 64.305 ;
        RECT 88.470 63.485 88.700 64.475 ;
        RECT 84.195 62.815 86.225 62.985 ;
        RECT 86.395 62.645 86.565 63.405 ;
        RECT 86.800 62.995 87.315 63.405 ;
        RECT 87.950 63.315 88.700 63.485 ;
        RECT 87.950 62.815 88.205 63.315 ;
        RECT 88.375 62.645 88.705 63.145 ;
        RECT 88.875 62.815 89.045 64.935 ;
        RECT 89.405 64.835 89.735 65.195 ;
        RECT 89.905 64.805 90.400 64.975 ;
        RECT 90.605 64.805 91.460 64.975 ;
        RECT 89.275 63.615 89.735 64.665 ;
        RECT 89.215 62.830 89.540 63.615 ;
        RECT 89.905 63.445 90.075 64.805 ;
        RECT 90.245 63.895 90.595 64.515 ;
        RECT 90.765 64.295 91.120 64.515 ;
        RECT 90.765 63.705 90.935 64.295 ;
        RECT 91.290 64.095 91.460 64.805 ;
        RECT 92.335 64.735 92.665 65.195 ;
        RECT 92.875 64.835 93.225 65.005 ;
        RECT 91.665 64.265 92.455 64.515 ;
        RECT 92.875 64.445 93.135 64.835 ;
        RECT 93.445 64.745 94.395 65.025 ;
        RECT 94.565 64.755 94.755 65.195 ;
        RECT 94.925 64.815 95.995 64.985 ;
        RECT 92.625 64.095 92.795 64.275 ;
        RECT 89.905 63.275 90.300 63.445 ;
        RECT 90.470 63.315 90.935 63.705 ;
        RECT 91.105 63.925 92.795 64.095 ;
        RECT 90.130 63.145 90.300 63.275 ;
        RECT 91.105 63.145 91.275 63.925 ;
        RECT 92.965 63.755 93.135 64.445 ;
        RECT 91.635 63.585 93.135 63.755 ;
        RECT 93.325 63.785 93.535 64.575 ;
        RECT 93.705 63.955 94.055 64.575 ;
        RECT 94.225 63.965 94.395 64.745 ;
        RECT 94.925 64.585 95.095 64.815 ;
        RECT 94.565 64.415 95.095 64.585 ;
        RECT 94.565 64.135 94.785 64.415 ;
        RECT 95.265 64.245 95.505 64.645 ;
        RECT 94.225 63.795 94.630 63.965 ;
        RECT 94.965 63.875 95.505 64.245 ;
        RECT 95.675 64.460 95.995 64.815 ;
        RECT 96.240 64.735 96.545 65.195 ;
        RECT 96.715 64.485 96.970 65.015 ;
        RECT 95.675 64.285 96.000 64.460 ;
        RECT 95.675 63.985 96.590 64.285 ;
        RECT 95.850 63.955 96.590 63.985 ;
        RECT 93.325 63.625 94.000 63.785 ;
        RECT 94.460 63.705 94.630 63.795 ;
        RECT 93.325 63.615 94.290 63.625 ;
        RECT 92.965 63.445 93.135 63.585 ;
        RECT 89.710 62.645 89.960 63.105 ;
        RECT 90.130 62.815 90.380 63.145 ;
        RECT 90.595 62.815 91.275 63.145 ;
        RECT 91.445 63.245 92.520 63.415 ;
        RECT 92.965 63.275 93.525 63.445 ;
        RECT 93.830 63.325 94.290 63.615 ;
        RECT 94.460 63.535 95.680 63.705 ;
        RECT 91.445 62.905 91.615 63.245 ;
        RECT 91.850 62.645 92.180 63.075 ;
        RECT 92.350 62.905 92.520 63.245 ;
        RECT 92.815 62.645 93.185 63.105 ;
        RECT 93.355 62.815 93.525 63.275 ;
        RECT 94.460 63.155 94.630 63.535 ;
        RECT 95.850 63.365 96.020 63.955 ;
        RECT 96.760 63.835 96.970 64.485 ;
        RECT 97.260 64.565 97.545 65.025 ;
        RECT 97.715 64.735 97.985 65.195 ;
        RECT 97.260 64.395 98.215 64.565 ;
        RECT 93.760 62.815 94.630 63.155 ;
        RECT 95.220 63.195 96.020 63.365 ;
        RECT 94.800 62.645 95.050 63.105 ;
        RECT 95.220 62.905 95.390 63.195 ;
        RECT 95.570 62.645 95.900 63.025 ;
        RECT 96.240 62.645 96.545 63.785 ;
        RECT 96.715 62.955 96.970 63.835 ;
        RECT 97.145 63.665 97.835 64.225 ;
        RECT 98.005 63.495 98.215 64.395 ;
        RECT 97.260 63.275 98.215 63.495 ;
        RECT 98.385 64.225 98.785 65.025 ;
        RECT 98.975 64.565 99.255 65.025 ;
        RECT 99.775 64.735 100.100 65.195 ;
        RECT 98.975 64.395 100.100 64.565 ;
        RECT 100.270 64.455 100.655 65.025 ;
        RECT 99.650 64.285 100.100 64.395 ;
        RECT 98.385 63.665 99.480 64.225 ;
        RECT 99.650 63.955 100.205 64.285 ;
        RECT 97.260 62.815 97.545 63.275 ;
        RECT 97.715 62.645 97.985 63.105 ;
        RECT 98.385 62.815 98.785 63.665 ;
        RECT 99.650 63.495 100.100 63.955 ;
        RECT 100.375 63.785 100.655 64.455 ;
        RECT 100.865 64.375 101.095 65.195 ;
        RECT 101.265 64.395 101.595 65.025 ;
        RECT 100.845 63.955 101.175 64.205 ;
        RECT 101.345 63.795 101.595 64.395 ;
        RECT 101.765 64.375 101.975 65.195 ;
        RECT 102.205 64.425 105.715 65.195 ;
        RECT 105.885 64.445 107.095 65.195 ;
        RECT 107.355 64.645 107.525 65.025 ;
        RECT 107.705 64.815 108.035 65.195 ;
        RECT 107.355 64.475 108.020 64.645 ;
        RECT 108.215 64.520 108.475 65.025 ;
        RECT 102.205 63.905 103.855 64.425 ;
        RECT 98.975 63.275 100.100 63.495 ;
        RECT 98.975 62.815 99.255 63.275 ;
        RECT 99.775 62.645 100.100 63.105 ;
        RECT 100.270 62.815 100.655 63.785 ;
        RECT 100.865 62.645 101.095 63.785 ;
        RECT 101.265 62.815 101.595 63.795 ;
        RECT 101.765 62.645 101.975 63.785 ;
        RECT 104.025 63.735 105.715 64.255 ;
        RECT 105.885 63.905 106.405 64.445 ;
        RECT 106.575 63.735 107.095 64.275 ;
        RECT 107.285 63.925 107.615 64.295 ;
        RECT 107.850 64.220 108.020 64.475 ;
        RECT 107.850 63.890 108.135 64.220 ;
        RECT 107.850 63.745 108.020 63.890 ;
        RECT 102.205 62.645 105.715 63.735 ;
        RECT 105.885 62.645 107.095 63.735 ;
        RECT 107.355 63.575 108.020 63.745 ;
        RECT 108.305 63.720 108.475 64.520 ;
        RECT 108.645 64.470 108.935 65.195 ;
        RECT 109.110 64.455 109.365 65.025 ;
        RECT 109.535 64.795 109.865 65.195 ;
        RECT 110.290 64.660 110.820 65.025 ;
        RECT 111.010 64.855 111.285 65.025 ;
        RECT 111.005 64.685 111.285 64.855 ;
        RECT 110.290 64.625 110.465 64.660 ;
        RECT 109.535 64.455 110.465 64.625 ;
        RECT 107.355 62.815 107.525 63.575 ;
        RECT 107.705 62.645 108.035 63.405 ;
        RECT 108.205 62.815 108.475 63.720 ;
        RECT 108.645 62.645 108.935 63.810 ;
        RECT 109.110 63.785 109.280 64.455 ;
        RECT 109.535 64.285 109.705 64.455 ;
        RECT 109.450 63.955 109.705 64.285 ;
        RECT 109.930 63.955 110.125 64.285 ;
        RECT 109.110 62.815 109.445 63.785 ;
        RECT 109.615 62.645 109.785 63.785 ;
        RECT 109.955 62.985 110.125 63.955 ;
        RECT 110.295 63.325 110.465 64.455 ;
        RECT 110.635 63.665 110.805 64.465 ;
        RECT 111.010 63.865 111.285 64.685 ;
        RECT 111.455 63.665 111.645 65.025 ;
        RECT 111.825 64.660 112.335 65.195 ;
        RECT 112.555 64.385 112.800 64.990 ;
        RECT 113.335 64.645 113.505 64.935 ;
        RECT 113.675 64.815 114.005 65.195 ;
        RECT 113.335 64.475 114.000 64.645 ;
        RECT 111.845 64.215 113.075 64.385 ;
        RECT 110.635 63.495 111.645 63.665 ;
        RECT 111.815 63.650 112.565 63.840 ;
        RECT 110.295 63.155 111.420 63.325 ;
        RECT 111.815 62.985 111.985 63.650 ;
        RECT 112.735 63.405 113.075 64.215 ;
        RECT 113.250 63.655 113.600 64.305 ;
        RECT 113.770 63.485 114.000 64.475 ;
        RECT 109.955 62.815 111.985 62.985 ;
        RECT 112.155 62.645 112.325 63.405 ;
        RECT 112.560 62.995 113.075 63.405 ;
        RECT 113.335 63.315 114.000 63.485 ;
        RECT 113.335 62.815 113.505 63.315 ;
        RECT 113.675 62.645 114.005 63.145 ;
        RECT 114.175 62.815 114.400 64.935 ;
        RECT 114.615 64.815 114.945 65.195 ;
        RECT 115.115 64.645 115.285 64.975 ;
        RECT 115.585 64.815 116.600 65.015 ;
        RECT 114.590 64.455 115.285 64.645 ;
        RECT 114.590 63.485 114.760 64.455 ;
        RECT 114.930 63.655 115.340 64.275 ;
        RECT 115.510 63.705 115.730 64.575 ;
        RECT 115.910 64.265 116.260 64.635 ;
        RECT 116.430 64.085 116.600 64.815 ;
        RECT 116.770 64.755 117.180 65.195 ;
        RECT 117.470 64.555 117.720 64.985 ;
        RECT 117.920 64.735 118.240 65.195 ;
        RECT 118.800 64.805 119.650 64.975 ;
        RECT 116.770 64.215 117.180 64.545 ;
        RECT 117.470 64.215 117.890 64.555 ;
        RECT 116.180 64.045 116.600 64.085 ;
        RECT 116.180 63.875 117.530 64.045 ;
        RECT 114.590 63.315 115.285 63.485 ;
        RECT 115.510 63.325 116.010 63.705 ;
        RECT 114.615 62.645 114.945 63.145 ;
        RECT 115.115 62.815 115.285 63.315 ;
        RECT 116.180 63.030 116.350 63.875 ;
        RECT 117.280 63.715 117.530 63.875 ;
        RECT 116.520 63.445 116.770 63.705 ;
        RECT 117.700 63.445 117.890 64.215 ;
        RECT 116.520 63.195 117.890 63.445 ;
        RECT 118.060 64.385 119.310 64.555 ;
        RECT 118.060 63.625 118.230 64.385 ;
        RECT 118.980 64.265 119.310 64.385 ;
        RECT 118.400 63.805 118.580 64.215 ;
        RECT 119.480 64.045 119.650 64.805 ;
        RECT 119.850 64.715 120.510 65.195 ;
        RECT 120.690 64.600 121.010 64.930 ;
        RECT 119.840 64.275 120.500 64.545 ;
        RECT 119.840 64.215 120.170 64.275 ;
        RECT 120.320 64.045 120.650 64.105 ;
        RECT 118.750 63.875 120.650 64.045 ;
        RECT 118.060 63.315 118.580 63.625 ;
        RECT 118.750 63.365 118.920 63.875 ;
        RECT 120.820 63.705 121.010 64.600 ;
        RECT 119.090 63.535 121.010 63.705 ;
        RECT 120.690 63.515 121.010 63.535 ;
        RECT 121.210 64.285 121.460 64.935 ;
        RECT 121.640 64.735 121.925 65.195 ;
        RECT 122.105 64.855 122.360 65.015 ;
        RECT 122.105 64.685 122.445 64.855 ;
        RECT 122.105 64.485 122.360 64.685 ;
        RECT 121.210 63.955 122.010 64.285 ;
        RECT 118.750 63.195 119.960 63.365 ;
        RECT 115.520 62.860 116.350 63.030 ;
        RECT 116.590 62.645 116.970 63.025 ;
        RECT 117.150 62.905 117.320 63.195 ;
        RECT 118.750 63.115 118.920 63.195 ;
        RECT 117.490 62.645 117.820 63.025 ;
        RECT 118.290 62.865 118.920 63.115 ;
        RECT 119.100 62.645 119.520 63.025 ;
        RECT 119.720 62.905 119.960 63.195 ;
        RECT 120.190 62.645 120.520 63.335 ;
        RECT 120.690 62.905 120.860 63.515 ;
        RECT 121.210 63.365 121.460 63.955 ;
        RECT 122.180 63.625 122.360 64.485 ;
        RECT 122.905 64.445 124.115 65.195 ;
        RECT 124.285 64.445 125.495 65.195 ;
        RECT 122.905 63.905 123.425 64.445 ;
        RECT 123.595 63.735 124.115 64.275 ;
        RECT 121.130 62.855 121.460 63.365 ;
        RECT 121.640 62.645 121.925 63.445 ;
        RECT 122.105 62.955 122.360 63.625 ;
        RECT 122.905 62.645 124.115 63.735 ;
        RECT 124.285 63.735 124.805 64.275 ;
        RECT 124.975 63.905 125.495 64.445 ;
        RECT 124.285 62.645 125.495 63.735 ;
        RECT 5.520 62.475 125.580 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 6.985 61.385 8.195 62.475 ;
        RECT 8.370 61.805 8.625 62.305 ;
        RECT 8.795 61.975 9.125 62.475 ;
        RECT 8.370 61.635 9.120 61.805 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 6.985 60.675 7.505 61.215 ;
        RECT 7.675 60.845 8.195 61.385 ;
        RECT 8.370 60.815 8.720 61.465 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 6.985 59.925 8.195 60.675 ;
        RECT 8.890 60.645 9.120 61.635 ;
        RECT 8.370 60.475 9.120 60.645 ;
        RECT 8.370 60.185 8.625 60.475 ;
        RECT 8.795 59.925 9.125 60.305 ;
        RECT 9.295 60.185 9.465 62.305 ;
        RECT 9.635 61.505 9.960 62.290 ;
        RECT 10.130 62.015 10.380 62.475 ;
        RECT 10.550 61.975 10.800 62.305 ;
        RECT 11.015 61.975 11.695 62.305 ;
        RECT 10.550 61.845 10.720 61.975 ;
        RECT 10.325 61.675 10.720 61.845 ;
        RECT 9.695 60.455 10.155 61.505 ;
        RECT 10.325 60.315 10.495 61.675 ;
        RECT 10.890 61.415 11.355 61.805 ;
        RECT 10.665 60.605 11.015 61.225 ;
        RECT 11.185 60.825 11.355 61.415 ;
        RECT 11.525 61.195 11.695 61.975 ;
        RECT 11.865 61.875 12.035 62.215 ;
        RECT 12.270 62.045 12.600 62.475 ;
        RECT 12.770 61.875 12.940 62.215 ;
        RECT 13.235 62.015 13.605 62.475 ;
        RECT 11.865 61.705 12.940 61.875 ;
        RECT 13.775 61.845 13.945 62.305 ;
        RECT 14.180 61.965 15.050 62.305 ;
        RECT 15.220 62.015 15.470 62.475 ;
        RECT 13.385 61.675 13.945 61.845 ;
        RECT 13.385 61.535 13.555 61.675 ;
        RECT 12.055 61.365 13.555 61.535 ;
        RECT 14.250 61.505 14.710 61.795 ;
        RECT 11.525 61.025 13.215 61.195 ;
        RECT 11.185 60.605 11.540 60.825 ;
        RECT 11.710 60.315 11.880 61.025 ;
        RECT 12.085 60.605 12.875 60.855 ;
        RECT 13.045 60.845 13.215 61.025 ;
        RECT 13.385 60.675 13.555 61.365 ;
        RECT 9.825 59.925 10.155 60.285 ;
        RECT 10.325 60.145 10.820 60.315 ;
        RECT 11.025 60.145 11.880 60.315 ;
        RECT 12.755 59.925 13.085 60.385 ;
        RECT 13.295 60.285 13.555 60.675 ;
        RECT 13.745 61.495 14.710 61.505 ;
        RECT 14.880 61.585 15.050 61.965 ;
        RECT 15.640 61.925 15.810 62.215 ;
        RECT 15.990 62.095 16.320 62.475 ;
        RECT 15.640 61.755 16.440 61.925 ;
        RECT 13.745 61.335 14.420 61.495 ;
        RECT 14.880 61.415 16.100 61.585 ;
        RECT 13.745 60.545 13.955 61.335 ;
        RECT 14.880 61.325 15.050 61.415 ;
        RECT 14.125 60.545 14.475 61.165 ;
        RECT 14.645 61.155 15.050 61.325 ;
        RECT 14.645 60.375 14.815 61.155 ;
        RECT 14.985 60.705 15.205 60.985 ;
        RECT 15.385 60.875 15.925 61.245 ;
        RECT 16.270 61.165 16.440 61.755 ;
        RECT 16.660 61.335 16.965 62.475 ;
        RECT 17.135 61.285 17.390 62.165 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 18.950 61.335 19.285 62.305 ;
        RECT 19.455 61.335 19.625 62.475 ;
        RECT 19.795 62.135 21.825 62.305 ;
        RECT 16.270 61.135 17.010 61.165 ;
        RECT 14.985 60.535 15.515 60.705 ;
        RECT 13.295 60.115 13.645 60.285 ;
        RECT 13.865 60.095 14.815 60.375 ;
        RECT 14.985 59.925 15.175 60.365 ;
        RECT 15.345 60.305 15.515 60.535 ;
        RECT 15.685 60.475 15.925 60.875 ;
        RECT 16.095 60.835 17.010 61.135 ;
        RECT 16.095 60.660 16.420 60.835 ;
        RECT 16.095 60.305 16.415 60.660 ;
        RECT 17.180 60.635 17.390 61.285 ;
        RECT 18.950 60.665 19.120 61.335 ;
        RECT 19.795 61.165 19.965 62.135 ;
        RECT 19.290 60.835 19.545 61.165 ;
        RECT 19.770 60.835 19.965 61.165 ;
        RECT 20.135 61.795 21.260 61.965 ;
        RECT 19.375 60.665 19.545 60.835 ;
        RECT 20.135 60.665 20.305 61.795 ;
        RECT 15.345 60.135 16.415 60.305 ;
        RECT 16.660 59.925 16.965 60.385 ;
        RECT 17.135 60.105 17.390 60.635 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 18.950 60.095 19.205 60.665 ;
        RECT 19.375 60.495 20.305 60.665 ;
        RECT 20.475 61.455 21.485 61.625 ;
        RECT 20.475 60.655 20.645 61.455 ;
        RECT 20.850 60.775 21.125 61.255 ;
        RECT 20.845 60.605 21.125 60.775 ;
        RECT 20.130 60.460 20.305 60.495 ;
        RECT 19.375 59.925 19.705 60.325 ;
        RECT 20.130 60.095 20.660 60.460 ;
        RECT 20.850 60.095 21.125 60.605 ;
        RECT 21.295 60.095 21.485 61.455 ;
        RECT 21.655 61.470 21.825 62.135 ;
        RECT 21.995 61.715 22.165 62.475 ;
        RECT 22.400 61.715 22.915 62.125 ;
        RECT 21.655 61.280 22.405 61.470 ;
        RECT 22.575 60.905 22.915 61.715 ;
        RECT 24.010 61.805 24.265 62.305 ;
        RECT 24.435 61.975 24.765 62.475 ;
        RECT 24.010 61.635 24.760 61.805 ;
        RECT 21.685 60.735 22.915 60.905 ;
        RECT 24.010 60.815 24.360 61.465 ;
        RECT 21.665 59.925 22.175 60.460 ;
        RECT 22.395 60.130 22.640 60.735 ;
        RECT 24.530 60.645 24.760 61.635 ;
        RECT 24.010 60.475 24.760 60.645 ;
        RECT 24.010 60.185 24.265 60.475 ;
        RECT 24.435 59.925 24.765 60.305 ;
        RECT 24.935 60.185 25.105 62.305 ;
        RECT 25.275 61.505 25.600 62.290 ;
        RECT 25.770 62.015 26.020 62.475 ;
        RECT 26.190 61.975 26.440 62.305 ;
        RECT 26.655 61.975 27.335 62.305 ;
        RECT 26.190 61.845 26.360 61.975 ;
        RECT 25.965 61.675 26.360 61.845 ;
        RECT 25.335 60.455 25.795 61.505 ;
        RECT 25.965 60.315 26.135 61.675 ;
        RECT 26.530 61.415 26.995 61.805 ;
        RECT 26.305 60.605 26.655 61.225 ;
        RECT 26.825 60.825 26.995 61.415 ;
        RECT 27.165 61.195 27.335 61.975 ;
        RECT 27.505 61.875 27.675 62.215 ;
        RECT 27.910 62.045 28.240 62.475 ;
        RECT 28.410 61.875 28.580 62.215 ;
        RECT 28.875 62.015 29.245 62.475 ;
        RECT 27.505 61.705 28.580 61.875 ;
        RECT 29.415 61.845 29.585 62.305 ;
        RECT 29.820 61.965 30.690 62.305 ;
        RECT 30.860 62.015 31.110 62.475 ;
        RECT 29.025 61.675 29.585 61.845 ;
        RECT 29.025 61.535 29.195 61.675 ;
        RECT 27.695 61.365 29.195 61.535 ;
        RECT 29.890 61.505 30.350 61.795 ;
        RECT 27.165 61.025 28.855 61.195 ;
        RECT 26.825 60.605 27.180 60.825 ;
        RECT 27.350 60.315 27.520 61.025 ;
        RECT 27.725 60.605 28.515 60.855 ;
        RECT 28.685 60.845 28.855 61.025 ;
        RECT 29.025 60.675 29.195 61.365 ;
        RECT 25.465 59.925 25.795 60.285 ;
        RECT 25.965 60.145 26.460 60.315 ;
        RECT 26.665 60.145 27.520 60.315 ;
        RECT 28.395 59.925 28.725 60.385 ;
        RECT 28.935 60.285 29.195 60.675 ;
        RECT 29.385 61.495 30.350 61.505 ;
        RECT 30.520 61.585 30.690 61.965 ;
        RECT 31.280 61.925 31.450 62.215 ;
        RECT 31.630 62.095 31.960 62.475 ;
        RECT 31.280 61.755 32.080 61.925 ;
        RECT 29.385 61.335 30.060 61.495 ;
        RECT 30.520 61.415 31.740 61.585 ;
        RECT 29.385 60.545 29.595 61.335 ;
        RECT 30.520 61.325 30.690 61.415 ;
        RECT 29.765 60.545 30.115 61.165 ;
        RECT 30.285 61.155 30.690 61.325 ;
        RECT 30.285 60.375 30.455 61.155 ;
        RECT 30.625 60.705 30.845 60.985 ;
        RECT 31.025 60.875 31.565 61.245 ;
        RECT 31.910 61.165 32.080 61.755 ;
        RECT 32.300 61.335 32.605 62.475 ;
        RECT 32.775 61.285 33.030 62.165 ;
        RECT 33.265 61.335 33.475 62.475 ;
        RECT 31.910 61.135 32.650 61.165 ;
        RECT 30.625 60.535 31.155 60.705 ;
        RECT 28.935 60.115 29.285 60.285 ;
        RECT 29.505 60.095 30.455 60.375 ;
        RECT 30.625 59.925 30.815 60.365 ;
        RECT 30.985 60.305 31.155 60.535 ;
        RECT 31.325 60.475 31.565 60.875 ;
        RECT 31.735 60.835 32.650 61.135 ;
        RECT 31.735 60.660 32.060 60.835 ;
        RECT 31.735 60.305 32.055 60.660 ;
        RECT 32.820 60.635 33.030 61.285 ;
        RECT 33.645 61.325 33.975 62.305 ;
        RECT 34.145 61.335 34.375 62.475 ;
        RECT 34.585 61.385 38.095 62.475 ;
        RECT 30.985 60.135 32.055 60.305 ;
        RECT 32.300 59.925 32.605 60.385 ;
        RECT 32.775 60.105 33.030 60.635 ;
        RECT 33.265 59.925 33.475 60.745 ;
        RECT 33.645 60.725 33.895 61.325 ;
        RECT 34.065 60.915 34.395 61.165 ;
        RECT 33.645 60.095 33.975 60.725 ;
        RECT 34.145 59.925 34.375 60.745 ;
        RECT 34.585 60.695 36.235 61.215 ;
        RECT 36.405 60.865 38.095 61.385 ;
        RECT 38.270 61.335 38.605 62.305 ;
        RECT 38.775 61.335 38.945 62.475 ;
        RECT 39.115 62.135 41.145 62.305 ;
        RECT 34.585 59.925 38.095 60.695 ;
        RECT 38.270 60.665 38.440 61.335 ;
        RECT 39.115 61.165 39.285 62.135 ;
        RECT 38.610 60.835 38.865 61.165 ;
        RECT 39.090 60.835 39.285 61.165 ;
        RECT 39.455 61.795 40.580 61.965 ;
        RECT 38.695 60.665 38.865 60.835 ;
        RECT 39.455 60.665 39.625 61.795 ;
        RECT 38.270 60.095 38.525 60.665 ;
        RECT 38.695 60.495 39.625 60.665 ;
        RECT 39.795 61.455 40.805 61.625 ;
        RECT 39.795 60.655 39.965 61.455 ;
        RECT 39.450 60.460 39.625 60.495 ;
        RECT 38.695 59.925 39.025 60.325 ;
        RECT 39.450 60.095 39.980 60.460 ;
        RECT 40.170 60.435 40.445 61.255 ;
        RECT 40.165 60.265 40.445 60.435 ;
        RECT 40.170 60.095 40.445 60.265 ;
        RECT 40.615 60.095 40.805 61.455 ;
        RECT 40.975 61.470 41.145 62.135 ;
        RECT 41.315 61.715 41.485 62.475 ;
        RECT 41.720 61.715 42.235 62.125 ;
        RECT 40.975 61.280 41.725 61.470 ;
        RECT 41.895 60.905 42.235 61.715 ;
        RECT 42.405 61.385 44.075 62.475 ;
        RECT 41.005 60.735 42.235 60.905 ;
        RECT 40.985 59.925 41.495 60.460 ;
        RECT 41.715 60.130 41.960 60.735 ;
        RECT 42.405 60.695 43.155 61.215 ;
        RECT 43.325 60.865 44.075 61.385 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 44.795 61.805 44.965 62.305 ;
        RECT 45.135 61.975 45.465 62.475 ;
        RECT 44.795 61.635 45.460 61.805 ;
        RECT 44.710 60.815 45.060 61.465 ;
        RECT 42.405 59.925 44.075 60.695 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 45.230 60.645 45.460 61.635 ;
        RECT 44.795 60.475 45.460 60.645 ;
        RECT 44.795 60.185 44.965 60.475 ;
        RECT 45.135 59.925 45.465 60.305 ;
        RECT 45.635 60.185 45.860 62.305 ;
        RECT 46.075 61.975 46.405 62.475 ;
        RECT 46.575 61.805 46.745 62.305 ;
        RECT 46.980 62.090 47.810 62.260 ;
        RECT 48.050 62.095 48.430 62.475 ;
        RECT 46.050 61.635 46.745 61.805 ;
        RECT 46.050 60.665 46.220 61.635 ;
        RECT 46.390 60.845 46.800 61.465 ;
        RECT 46.970 61.415 47.470 61.795 ;
        RECT 46.050 60.475 46.745 60.665 ;
        RECT 46.970 60.545 47.190 61.415 ;
        RECT 47.640 61.245 47.810 62.090 ;
        RECT 48.610 61.925 48.780 62.215 ;
        RECT 48.950 62.095 49.280 62.475 ;
        RECT 49.750 62.005 50.380 62.255 ;
        RECT 50.560 62.095 50.980 62.475 ;
        RECT 50.210 61.925 50.380 62.005 ;
        RECT 51.180 61.925 51.420 62.215 ;
        RECT 47.980 61.675 49.350 61.925 ;
        RECT 47.980 61.415 48.230 61.675 ;
        RECT 48.740 61.245 48.990 61.405 ;
        RECT 47.640 61.075 48.990 61.245 ;
        RECT 47.640 61.035 48.060 61.075 ;
        RECT 47.370 60.485 47.720 60.855 ;
        RECT 46.075 59.925 46.405 60.305 ;
        RECT 46.575 60.145 46.745 60.475 ;
        RECT 47.890 60.305 48.060 61.035 ;
        RECT 49.160 60.905 49.350 61.675 ;
        RECT 48.230 60.575 48.640 60.905 ;
        RECT 48.930 60.565 49.350 60.905 ;
        RECT 49.520 61.495 50.040 61.805 ;
        RECT 50.210 61.755 51.420 61.925 ;
        RECT 51.650 61.785 51.980 62.475 ;
        RECT 49.520 60.735 49.690 61.495 ;
        RECT 49.860 60.905 50.040 61.315 ;
        RECT 50.210 61.245 50.380 61.755 ;
        RECT 52.150 61.605 52.320 62.215 ;
        RECT 52.590 61.755 52.920 62.265 ;
        RECT 52.150 61.585 52.470 61.605 ;
        RECT 50.550 61.415 52.470 61.585 ;
        RECT 50.210 61.075 52.110 61.245 ;
        RECT 50.440 60.735 50.770 60.855 ;
        RECT 49.520 60.565 50.770 60.735 ;
        RECT 47.045 60.105 48.060 60.305 ;
        RECT 48.230 59.925 48.640 60.365 ;
        RECT 48.930 60.135 49.180 60.565 ;
        RECT 49.380 59.925 49.700 60.385 ;
        RECT 50.940 60.315 51.110 61.075 ;
        RECT 51.780 61.015 52.110 61.075 ;
        RECT 51.300 60.845 51.630 60.905 ;
        RECT 51.300 60.575 51.960 60.845 ;
        RECT 52.280 60.520 52.470 61.415 ;
        RECT 50.260 60.145 51.110 60.315 ;
        RECT 51.310 59.925 51.970 60.405 ;
        RECT 52.150 60.190 52.470 60.520 ;
        RECT 52.670 61.165 52.920 61.755 ;
        RECT 53.100 61.675 53.385 62.475 ;
        RECT 53.565 61.495 53.820 62.165 ;
        RECT 52.670 60.835 53.470 61.165 ;
        RECT 52.670 60.185 52.920 60.835 ;
        RECT 53.640 60.635 53.820 61.495 ;
        RECT 54.365 61.385 57.875 62.475 ;
        RECT 58.045 61.385 59.255 62.475 ;
        RECT 59.480 61.605 59.765 62.475 ;
        RECT 59.935 61.845 60.195 62.305 ;
        RECT 60.370 62.015 60.625 62.475 ;
        RECT 60.795 61.845 61.055 62.305 ;
        RECT 59.935 61.675 61.055 61.845 ;
        RECT 61.225 61.675 61.535 62.475 ;
        RECT 59.935 61.425 60.195 61.675 ;
        RECT 61.705 61.505 62.015 62.305 ;
        RECT 53.565 60.435 53.820 60.635 ;
        RECT 54.365 60.695 56.015 61.215 ;
        RECT 56.185 60.865 57.875 61.385 ;
        RECT 53.100 59.925 53.385 60.385 ;
        RECT 53.565 60.265 53.905 60.435 ;
        RECT 53.565 60.105 53.820 60.265 ;
        RECT 54.365 59.925 57.875 60.695 ;
        RECT 58.045 60.675 58.565 61.215 ;
        RECT 58.735 60.845 59.255 61.385 ;
        RECT 59.440 61.255 60.195 61.425 ;
        RECT 60.985 61.335 62.015 61.505 ;
        RECT 62.185 61.385 65.695 62.475 ;
        RECT 59.440 60.745 59.845 61.255 ;
        RECT 60.985 61.085 61.155 61.335 ;
        RECT 60.015 60.915 61.155 61.085 ;
        RECT 58.045 59.925 59.255 60.675 ;
        RECT 59.440 60.575 61.090 60.745 ;
        RECT 61.325 60.595 61.675 61.165 ;
        RECT 59.485 59.925 59.765 60.405 ;
        RECT 59.935 60.185 60.195 60.575 ;
        RECT 60.370 59.925 60.625 60.405 ;
        RECT 60.795 60.185 61.090 60.575 ;
        RECT 61.845 60.425 62.015 61.335 ;
        RECT 61.270 59.925 61.545 60.405 ;
        RECT 61.715 60.095 62.015 60.425 ;
        RECT 62.185 60.695 63.835 61.215 ;
        RECT 64.005 60.865 65.695 61.385 ;
        RECT 65.875 61.495 66.205 62.305 ;
        RECT 66.375 61.675 66.615 62.475 ;
        RECT 65.875 61.325 66.590 61.495 ;
        RECT 65.870 60.915 66.250 61.155 ;
        RECT 66.420 61.085 66.590 61.325 ;
        RECT 66.795 61.455 66.965 62.305 ;
        RECT 67.135 61.675 67.465 62.475 ;
        RECT 67.635 61.455 67.805 62.305 ;
        RECT 66.795 61.285 67.805 61.455 ;
        RECT 67.975 61.325 68.305 62.475 ;
        RECT 68.625 61.385 69.835 62.475 ;
        RECT 66.420 60.915 66.920 61.085 ;
        RECT 66.420 60.745 66.590 60.915 ;
        RECT 67.310 60.745 67.805 61.285 ;
        RECT 62.185 59.925 65.695 60.695 ;
        RECT 65.955 60.575 66.590 60.745 ;
        RECT 66.795 60.575 67.805 60.745 ;
        RECT 65.955 60.095 66.125 60.575 ;
        RECT 66.305 59.925 66.545 60.405 ;
        RECT 66.795 60.095 66.965 60.575 ;
        RECT 67.135 59.925 67.465 60.405 ;
        RECT 67.635 60.095 67.805 60.575 ;
        RECT 67.975 59.925 68.305 60.725 ;
        RECT 68.625 60.675 69.145 61.215 ;
        RECT 69.315 60.845 69.835 61.385 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.465 61.385 73.975 62.475 ;
        RECT 70.465 60.695 72.115 61.215 ;
        RECT 72.285 60.865 73.975 61.385 ;
        RECT 74.145 61.400 74.415 62.305 ;
        RECT 74.585 61.715 74.915 62.475 ;
        RECT 75.095 61.545 75.265 62.305 ;
        RECT 68.625 59.925 69.835 60.675 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 70.465 59.925 73.975 60.695 ;
        RECT 74.145 60.600 74.315 61.400 ;
        RECT 74.600 61.375 75.265 61.545 ;
        RECT 75.525 61.385 77.195 62.475 ;
        RECT 74.600 61.230 74.770 61.375 ;
        RECT 74.485 60.900 74.770 61.230 ;
        RECT 74.600 60.645 74.770 60.900 ;
        RECT 75.005 60.825 75.335 61.195 ;
        RECT 75.525 60.695 76.275 61.215 ;
        RECT 76.445 60.865 77.195 61.385 ;
        RECT 77.405 61.335 77.635 62.475 ;
        RECT 77.805 61.325 78.135 62.305 ;
        RECT 78.305 61.335 78.515 62.475 ;
        RECT 79.210 61.805 79.465 62.305 ;
        RECT 79.635 61.975 79.965 62.475 ;
        RECT 79.210 61.635 79.960 61.805 ;
        RECT 77.385 60.915 77.715 61.165 ;
        RECT 74.145 60.095 74.405 60.600 ;
        RECT 74.600 60.475 75.265 60.645 ;
        RECT 74.585 59.925 74.915 60.305 ;
        RECT 75.095 60.095 75.265 60.475 ;
        RECT 75.525 59.925 77.195 60.695 ;
        RECT 77.405 59.925 77.635 60.745 ;
        RECT 77.885 60.725 78.135 61.325 ;
        RECT 79.210 60.815 79.560 61.465 ;
        RECT 77.805 60.095 78.135 60.725 ;
        RECT 78.305 59.925 78.515 60.745 ;
        RECT 79.730 60.645 79.960 61.635 ;
        RECT 79.210 60.475 79.960 60.645 ;
        RECT 79.210 60.185 79.465 60.475 ;
        RECT 79.635 59.925 79.965 60.305 ;
        RECT 80.135 60.185 80.305 62.305 ;
        RECT 80.475 61.505 80.800 62.290 ;
        RECT 80.970 62.015 81.220 62.475 ;
        RECT 81.390 61.975 81.640 62.305 ;
        RECT 81.855 61.975 82.535 62.305 ;
        RECT 81.390 61.845 81.560 61.975 ;
        RECT 81.165 61.675 81.560 61.845 ;
        RECT 80.535 60.455 80.995 61.505 ;
        RECT 81.165 60.315 81.335 61.675 ;
        RECT 81.730 61.415 82.195 61.805 ;
        RECT 81.505 60.605 81.855 61.225 ;
        RECT 82.025 60.825 82.195 61.415 ;
        RECT 82.365 61.195 82.535 61.975 ;
        RECT 82.705 61.875 82.875 62.215 ;
        RECT 83.110 62.045 83.440 62.475 ;
        RECT 83.610 61.875 83.780 62.215 ;
        RECT 84.075 62.015 84.445 62.475 ;
        RECT 82.705 61.705 83.780 61.875 ;
        RECT 84.615 61.845 84.785 62.305 ;
        RECT 85.020 61.965 85.890 62.305 ;
        RECT 86.060 62.015 86.310 62.475 ;
        RECT 84.225 61.675 84.785 61.845 ;
        RECT 84.225 61.535 84.395 61.675 ;
        RECT 82.895 61.365 84.395 61.535 ;
        RECT 85.090 61.505 85.550 61.795 ;
        RECT 82.365 61.025 84.055 61.195 ;
        RECT 82.025 60.605 82.380 60.825 ;
        RECT 82.550 60.315 82.720 61.025 ;
        RECT 82.925 60.605 83.715 60.855 ;
        RECT 83.885 60.845 84.055 61.025 ;
        RECT 84.225 60.675 84.395 61.365 ;
        RECT 80.665 59.925 80.995 60.285 ;
        RECT 81.165 60.145 81.660 60.315 ;
        RECT 81.865 60.145 82.720 60.315 ;
        RECT 83.595 59.925 83.925 60.385 ;
        RECT 84.135 60.285 84.395 60.675 ;
        RECT 84.585 61.495 85.550 61.505 ;
        RECT 85.720 61.585 85.890 61.965 ;
        RECT 86.480 61.925 86.650 62.215 ;
        RECT 86.830 62.095 87.160 62.475 ;
        RECT 86.480 61.755 87.280 61.925 ;
        RECT 84.585 61.335 85.260 61.495 ;
        RECT 85.720 61.415 86.940 61.585 ;
        RECT 84.585 60.545 84.795 61.335 ;
        RECT 85.720 61.325 85.890 61.415 ;
        RECT 84.965 60.545 85.315 61.165 ;
        RECT 85.485 61.155 85.890 61.325 ;
        RECT 85.485 60.375 85.655 61.155 ;
        RECT 85.825 60.705 86.045 60.985 ;
        RECT 86.225 60.875 86.765 61.245 ;
        RECT 87.110 61.165 87.280 61.755 ;
        RECT 87.500 61.335 87.805 62.475 ;
        RECT 87.975 61.285 88.230 62.165 ;
        RECT 87.110 61.135 87.850 61.165 ;
        RECT 85.825 60.535 86.355 60.705 ;
        RECT 84.135 60.115 84.485 60.285 ;
        RECT 84.705 60.095 85.655 60.375 ;
        RECT 85.825 59.925 86.015 60.365 ;
        RECT 86.185 60.305 86.355 60.535 ;
        RECT 86.525 60.475 86.765 60.875 ;
        RECT 86.935 60.835 87.850 61.135 ;
        RECT 86.935 60.660 87.260 60.835 ;
        RECT 86.935 60.305 87.255 60.660 ;
        RECT 88.020 60.635 88.230 61.285 ;
        RECT 86.185 60.135 87.255 60.305 ;
        RECT 87.500 59.925 87.805 60.385 ;
        RECT 87.975 60.105 88.230 60.635 ;
        RECT 88.865 61.335 89.250 62.305 ;
        RECT 89.420 62.015 89.745 62.475 ;
        RECT 90.265 61.845 90.545 62.305 ;
        RECT 89.420 61.625 90.545 61.845 ;
        RECT 88.865 60.665 89.145 61.335 ;
        RECT 89.420 61.165 89.870 61.625 ;
        RECT 90.735 61.455 91.135 62.305 ;
        RECT 91.535 62.015 91.805 62.475 ;
        RECT 91.975 61.845 92.260 62.305 ;
        RECT 89.315 60.835 89.870 61.165 ;
        RECT 90.040 60.895 91.135 61.455 ;
        RECT 89.420 60.725 89.870 60.835 ;
        RECT 88.865 60.095 89.250 60.665 ;
        RECT 89.420 60.555 90.545 60.725 ;
        RECT 89.420 59.925 89.745 60.385 ;
        RECT 90.265 60.095 90.545 60.555 ;
        RECT 90.735 60.095 91.135 60.895 ;
        RECT 91.305 61.625 92.260 61.845 ;
        RECT 91.305 60.725 91.515 61.625 ;
        RECT 91.685 60.895 92.375 61.455 ;
        RECT 92.605 61.335 92.815 62.475 ;
        RECT 92.985 61.325 93.315 62.305 ;
        RECT 93.485 61.335 93.715 62.475 ;
        RECT 93.925 61.400 94.195 62.305 ;
        RECT 94.365 61.715 94.695 62.475 ;
        RECT 94.875 61.545 95.045 62.305 ;
        RECT 91.305 60.555 92.260 60.725 ;
        RECT 91.535 59.925 91.805 60.385 ;
        RECT 91.975 60.095 92.260 60.555 ;
        RECT 92.605 59.925 92.815 60.745 ;
        RECT 92.985 60.725 93.235 61.325 ;
        RECT 93.405 60.915 93.735 61.165 ;
        RECT 92.985 60.095 93.315 60.725 ;
        RECT 93.485 59.925 93.715 60.745 ;
        RECT 93.925 60.600 94.095 61.400 ;
        RECT 94.380 61.375 95.045 61.545 ;
        RECT 94.380 61.230 94.550 61.375 ;
        RECT 95.765 61.310 96.055 62.475 ;
        RECT 96.285 61.335 96.495 62.475 ;
        RECT 96.665 61.325 96.995 62.305 ;
        RECT 97.165 61.335 97.395 62.475 ;
        RECT 97.605 62.040 102.950 62.475 ;
        RECT 94.265 60.900 94.550 61.230 ;
        RECT 94.380 60.645 94.550 60.900 ;
        RECT 94.785 60.825 95.115 61.195 ;
        RECT 93.925 60.095 94.185 60.600 ;
        RECT 94.380 60.475 95.045 60.645 ;
        RECT 94.365 59.925 94.695 60.305 ;
        RECT 94.875 60.095 95.045 60.475 ;
        RECT 95.765 59.925 96.055 60.650 ;
        RECT 96.285 59.925 96.495 60.745 ;
        RECT 96.665 60.725 96.915 61.325 ;
        RECT 97.085 60.915 97.415 61.165 ;
        RECT 96.665 60.095 96.995 60.725 ;
        RECT 97.165 59.925 97.395 60.745 ;
        RECT 99.190 60.470 99.530 61.300 ;
        RECT 101.010 60.790 101.360 62.040 ;
        RECT 103.125 61.385 105.715 62.475 ;
        RECT 103.125 60.695 104.335 61.215 ;
        RECT 104.505 60.865 105.715 61.385 ;
        RECT 106.350 61.285 106.605 62.165 ;
        RECT 106.775 61.335 107.080 62.475 ;
        RECT 107.420 62.095 107.750 62.475 ;
        RECT 107.930 61.925 108.100 62.215 ;
        RECT 108.270 62.015 108.520 62.475 ;
        RECT 107.300 61.755 108.100 61.925 ;
        RECT 108.690 61.965 109.560 62.305 ;
        RECT 97.605 59.925 102.950 60.470 ;
        RECT 103.125 59.925 105.715 60.695 ;
        RECT 106.350 60.635 106.560 61.285 ;
        RECT 107.300 61.165 107.470 61.755 ;
        RECT 108.690 61.585 108.860 61.965 ;
        RECT 109.795 61.845 109.965 62.305 ;
        RECT 110.135 62.015 110.505 62.475 ;
        RECT 110.800 61.875 110.970 62.215 ;
        RECT 111.140 62.045 111.470 62.475 ;
        RECT 111.705 61.875 111.875 62.215 ;
        RECT 107.640 61.415 108.860 61.585 ;
        RECT 109.030 61.505 109.490 61.795 ;
        RECT 109.795 61.675 110.355 61.845 ;
        RECT 110.800 61.705 111.875 61.875 ;
        RECT 112.045 61.975 112.725 62.305 ;
        RECT 112.940 61.975 113.190 62.305 ;
        RECT 113.360 62.015 113.610 62.475 ;
        RECT 110.185 61.535 110.355 61.675 ;
        RECT 109.030 61.495 109.995 61.505 ;
        RECT 108.690 61.325 108.860 61.415 ;
        RECT 109.320 61.335 109.995 61.495 ;
        RECT 106.730 61.135 107.470 61.165 ;
        RECT 106.730 60.835 107.645 61.135 ;
        RECT 107.320 60.660 107.645 60.835 ;
        RECT 106.350 60.105 106.605 60.635 ;
        RECT 106.775 59.925 107.080 60.385 ;
        RECT 107.325 60.305 107.645 60.660 ;
        RECT 107.815 60.875 108.355 61.245 ;
        RECT 108.690 61.155 109.095 61.325 ;
        RECT 107.815 60.475 108.055 60.875 ;
        RECT 108.535 60.705 108.755 60.985 ;
        RECT 108.225 60.535 108.755 60.705 ;
        RECT 108.225 60.305 108.395 60.535 ;
        RECT 108.925 60.375 109.095 61.155 ;
        RECT 109.265 60.545 109.615 61.165 ;
        RECT 109.785 60.545 109.995 61.335 ;
        RECT 110.185 61.365 111.685 61.535 ;
        RECT 110.185 60.675 110.355 61.365 ;
        RECT 112.045 61.195 112.215 61.975 ;
        RECT 113.020 61.845 113.190 61.975 ;
        RECT 110.525 61.025 112.215 61.195 ;
        RECT 112.385 61.415 112.850 61.805 ;
        RECT 113.020 61.675 113.415 61.845 ;
        RECT 110.525 60.845 110.695 61.025 ;
        RECT 107.325 60.135 108.395 60.305 ;
        RECT 108.565 59.925 108.755 60.365 ;
        RECT 108.925 60.095 109.875 60.375 ;
        RECT 110.185 60.285 110.445 60.675 ;
        RECT 110.865 60.605 111.655 60.855 ;
        RECT 110.095 60.115 110.445 60.285 ;
        RECT 110.655 59.925 110.985 60.385 ;
        RECT 111.860 60.315 112.030 61.025 ;
        RECT 112.385 60.825 112.555 61.415 ;
        RECT 112.200 60.605 112.555 60.825 ;
        RECT 112.725 60.605 113.075 61.225 ;
        RECT 113.245 60.315 113.415 61.675 ;
        RECT 113.780 61.505 114.105 62.290 ;
        RECT 113.585 60.455 114.045 61.505 ;
        RECT 111.860 60.145 112.715 60.315 ;
        RECT 112.920 60.145 113.415 60.315 ;
        RECT 113.585 59.925 113.915 60.285 ;
        RECT 114.275 60.185 114.445 62.305 ;
        RECT 114.615 61.975 114.945 62.475 ;
        RECT 115.115 61.805 115.370 62.305 ;
        RECT 115.545 62.040 120.890 62.475 ;
        RECT 114.620 61.635 115.370 61.805 ;
        RECT 114.620 60.645 114.850 61.635 ;
        RECT 115.020 60.815 115.370 61.465 ;
        RECT 114.620 60.475 115.370 60.645 ;
        RECT 114.615 59.925 114.945 60.305 ;
        RECT 115.115 60.185 115.370 60.475 ;
        RECT 117.130 60.470 117.470 61.300 ;
        RECT 118.950 60.790 119.300 62.040 ;
        RECT 121.525 61.310 121.815 62.475 ;
        RECT 121.985 61.385 123.655 62.475 ;
        RECT 121.985 60.695 122.735 61.215 ;
        RECT 122.905 60.865 123.655 61.385 ;
        RECT 124.285 61.385 125.495 62.475 ;
        RECT 124.285 60.845 124.805 61.385 ;
        RECT 115.545 59.925 120.890 60.470 ;
        RECT 121.525 59.925 121.815 60.650 ;
        RECT 121.985 59.925 123.655 60.695 ;
        RECT 124.975 60.675 125.495 61.215 ;
        RECT 124.285 59.925 125.495 60.675 ;
        RECT 5.520 59.755 125.580 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.985 58.985 10.495 59.755 ;
        RECT 10.665 59.080 10.925 59.585 ;
        RECT 11.105 59.375 11.435 59.755 ;
        RECT 11.615 59.205 11.785 59.585 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 6.985 58.465 8.635 58.985 ;
        RECT 8.805 58.295 10.495 58.815 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 6.985 57.205 10.495 58.295 ;
        RECT 10.665 58.280 10.835 59.080 ;
        RECT 11.120 59.035 11.785 59.205 ;
        RECT 11.120 58.780 11.290 59.035 ;
        RECT 12.105 58.935 12.315 59.755 ;
        RECT 12.485 58.955 12.815 59.585 ;
        RECT 11.005 58.450 11.290 58.780 ;
        RECT 11.525 58.485 11.855 58.855 ;
        RECT 11.120 58.305 11.290 58.450 ;
        RECT 12.485 58.355 12.735 58.955 ;
        RECT 12.985 58.935 13.215 59.755 ;
        RECT 13.425 59.015 13.810 59.585 ;
        RECT 13.980 59.295 14.305 59.755 ;
        RECT 14.825 59.125 15.105 59.585 ;
        RECT 12.905 58.515 13.235 58.765 ;
        RECT 10.665 57.375 10.935 58.280 ;
        RECT 11.120 58.135 11.785 58.305 ;
        RECT 11.105 57.205 11.435 57.965 ;
        RECT 11.615 57.375 11.785 58.135 ;
        RECT 12.105 57.205 12.315 58.345 ;
        RECT 12.485 57.375 12.815 58.355 ;
        RECT 13.425 58.345 13.705 59.015 ;
        RECT 13.980 58.955 15.105 59.125 ;
        RECT 13.980 58.845 14.430 58.955 ;
        RECT 13.875 58.515 14.430 58.845 ;
        RECT 15.295 58.785 15.695 59.585 ;
        RECT 16.095 59.295 16.365 59.755 ;
        RECT 16.535 59.125 16.820 59.585 ;
        RECT 12.985 57.205 13.215 58.345 ;
        RECT 13.425 57.375 13.810 58.345 ;
        RECT 13.980 58.055 14.430 58.515 ;
        RECT 14.600 58.225 15.695 58.785 ;
        RECT 13.980 57.835 15.105 58.055 ;
        RECT 13.980 57.205 14.305 57.665 ;
        RECT 14.825 57.375 15.105 57.835 ;
        RECT 15.295 57.375 15.695 58.225 ;
        RECT 15.865 58.955 16.820 59.125 ;
        RECT 17.105 59.015 17.490 59.585 ;
        RECT 17.660 59.295 17.985 59.755 ;
        RECT 18.505 59.125 18.785 59.585 ;
        RECT 15.865 58.055 16.075 58.955 ;
        RECT 16.245 58.225 16.935 58.785 ;
        RECT 17.105 58.345 17.385 59.015 ;
        RECT 17.660 58.955 18.785 59.125 ;
        RECT 17.660 58.845 18.110 58.955 ;
        RECT 17.555 58.515 18.110 58.845 ;
        RECT 18.975 58.785 19.375 59.585 ;
        RECT 19.775 59.295 20.045 59.755 ;
        RECT 20.215 59.125 20.500 59.585 ;
        RECT 15.865 57.835 16.820 58.055 ;
        RECT 16.095 57.205 16.365 57.665 ;
        RECT 16.535 57.375 16.820 57.835 ;
        RECT 17.105 57.375 17.490 58.345 ;
        RECT 17.660 58.055 18.110 58.515 ;
        RECT 18.280 58.225 19.375 58.785 ;
        RECT 17.660 57.835 18.785 58.055 ;
        RECT 17.660 57.205 17.985 57.665 ;
        RECT 18.505 57.375 18.785 57.835 ;
        RECT 18.975 57.375 19.375 58.225 ;
        RECT 19.545 58.955 20.500 59.125 ;
        RECT 19.545 58.055 19.755 58.955 ;
        RECT 20.845 58.935 21.055 59.755 ;
        RECT 21.225 58.955 21.555 59.585 ;
        RECT 19.925 58.225 20.615 58.785 ;
        RECT 21.225 58.355 21.475 58.955 ;
        RECT 21.725 58.935 21.955 59.755 ;
        RECT 22.255 59.275 22.555 59.755 ;
        RECT 22.725 59.105 22.985 59.560 ;
        RECT 23.155 59.275 23.415 59.755 ;
        RECT 23.595 59.105 23.855 59.560 ;
        RECT 24.025 59.275 24.275 59.755 ;
        RECT 24.455 59.105 24.715 59.560 ;
        RECT 24.885 59.275 25.135 59.755 ;
        RECT 25.315 59.105 25.575 59.560 ;
        RECT 25.745 59.275 25.990 59.755 ;
        RECT 26.160 59.105 26.435 59.560 ;
        RECT 26.605 59.275 26.850 59.755 ;
        RECT 27.020 59.105 27.280 59.560 ;
        RECT 27.450 59.275 27.710 59.755 ;
        RECT 27.880 59.105 28.140 59.560 ;
        RECT 28.310 59.275 28.570 59.755 ;
        RECT 28.740 59.105 29.000 59.560 ;
        RECT 29.170 59.195 29.430 59.755 ;
        RECT 22.255 58.935 29.000 59.105 ;
        RECT 21.645 58.515 21.975 58.765 ;
        RECT 19.545 57.835 20.500 58.055 ;
        RECT 19.775 57.205 20.045 57.665 ;
        RECT 20.215 57.375 20.500 57.835 ;
        RECT 20.845 57.205 21.055 58.345 ;
        RECT 21.225 57.375 21.555 58.355 ;
        RECT 22.255 58.345 23.420 58.935 ;
        RECT 29.600 58.765 29.850 59.575 ;
        RECT 30.030 59.230 30.290 59.755 ;
        RECT 30.460 58.765 30.710 59.575 ;
        RECT 30.890 59.245 31.195 59.755 ;
        RECT 23.590 58.515 30.710 58.765 ;
        RECT 30.880 58.515 31.195 59.075 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.825 59.005 33.035 59.755 ;
        RECT 33.210 59.205 33.465 59.495 ;
        RECT 33.635 59.375 33.965 59.755 ;
        RECT 33.210 59.035 33.960 59.205 ;
        RECT 21.725 57.205 21.955 58.345 ;
        RECT 22.255 58.120 29.000 58.345 ;
        RECT 22.255 57.205 22.525 57.950 ;
        RECT 22.695 57.380 22.985 58.120 ;
        RECT 23.595 58.105 29.000 58.120 ;
        RECT 23.155 57.210 23.410 57.935 ;
        RECT 23.595 57.380 23.855 58.105 ;
        RECT 24.025 57.210 24.270 57.935 ;
        RECT 24.455 57.380 24.715 58.105 ;
        RECT 24.885 57.210 25.130 57.935 ;
        RECT 25.315 57.380 25.575 58.105 ;
        RECT 25.745 57.210 25.990 57.935 ;
        RECT 26.160 57.380 26.420 58.105 ;
        RECT 26.590 57.210 26.850 57.935 ;
        RECT 27.020 57.380 27.280 58.105 ;
        RECT 27.450 57.210 27.710 57.935 ;
        RECT 27.880 57.380 28.140 58.105 ;
        RECT 28.310 57.210 28.570 57.935 ;
        RECT 28.740 57.380 29.000 58.105 ;
        RECT 29.170 57.210 29.430 58.005 ;
        RECT 29.600 57.380 29.850 58.515 ;
        RECT 23.155 57.205 29.430 57.210 ;
        RECT 30.030 57.205 30.290 58.015 ;
        RECT 30.465 57.375 30.710 58.515 ;
        RECT 31.825 58.465 32.345 59.005 ;
        RECT 30.890 57.205 31.185 58.015 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 32.515 58.295 33.035 58.835 ;
        RECT 31.825 57.205 33.035 58.295 ;
        RECT 33.210 58.215 33.560 58.865 ;
        RECT 33.730 58.045 33.960 59.035 ;
        RECT 33.210 57.875 33.960 58.045 ;
        RECT 33.210 57.375 33.465 57.875 ;
        RECT 33.635 57.205 33.965 57.705 ;
        RECT 34.135 57.375 34.305 59.495 ;
        RECT 34.665 59.395 34.995 59.755 ;
        RECT 35.165 59.365 35.660 59.535 ;
        RECT 35.865 59.365 36.720 59.535 ;
        RECT 34.535 58.175 34.995 59.225 ;
        RECT 34.475 57.390 34.800 58.175 ;
        RECT 35.165 58.005 35.335 59.365 ;
        RECT 35.505 58.455 35.855 59.075 ;
        RECT 36.025 58.855 36.380 59.075 ;
        RECT 36.025 58.265 36.195 58.855 ;
        RECT 36.550 58.655 36.720 59.365 ;
        RECT 37.595 59.295 37.925 59.755 ;
        RECT 38.135 59.395 38.485 59.565 ;
        RECT 36.925 58.825 37.715 59.075 ;
        RECT 38.135 59.005 38.395 59.395 ;
        RECT 38.705 59.305 39.655 59.585 ;
        RECT 39.825 59.315 40.015 59.755 ;
        RECT 40.185 59.375 41.255 59.545 ;
        RECT 37.885 58.655 38.055 58.835 ;
        RECT 35.165 57.835 35.560 58.005 ;
        RECT 35.730 57.875 36.195 58.265 ;
        RECT 36.365 58.485 38.055 58.655 ;
        RECT 35.390 57.705 35.560 57.835 ;
        RECT 36.365 57.705 36.535 58.485 ;
        RECT 38.225 58.315 38.395 59.005 ;
        RECT 36.895 58.145 38.395 58.315 ;
        RECT 38.585 58.345 38.795 59.135 ;
        RECT 38.965 58.515 39.315 59.135 ;
        RECT 39.485 58.525 39.655 59.305 ;
        RECT 40.185 59.145 40.355 59.375 ;
        RECT 39.825 58.975 40.355 59.145 ;
        RECT 39.825 58.695 40.045 58.975 ;
        RECT 40.525 58.805 40.765 59.205 ;
        RECT 39.485 58.355 39.890 58.525 ;
        RECT 40.225 58.435 40.765 58.805 ;
        RECT 40.935 59.020 41.255 59.375 ;
        RECT 41.500 59.295 41.805 59.755 ;
        RECT 41.975 59.045 42.230 59.575 ;
        RECT 40.935 58.845 41.260 59.020 ;
        RECT 40.935 58.545 41.850 58.845 ;
        RECT 41.110 58.515 41.850 58.545 ;
        RECT 38.585 58.185 39.260 58.345 ;
        RECT 39.720 58.265 39.890 58.355 ;
        RECT 38.585 58.175 39.550 58.185 ;
        RECT 38.225 58.005 38.395 58.145 ;
        RECT 34.970 57.205 35.220 57.665 ;
        RECT 35.390 57.375 35.640 57.705 ;
        RECT 35.855 57.375 36.535 57.705 ;
        RECT 36.705 57.805 37.780 57.975 ;
        RECT 38.225 57.835 38.785 58.005 ;
        RECT 39.090 57.885 39.550 58.175 ;
        RECT 39.720 58.095 40.940 58.265 ;
        RECT 36.705 57.465 36.875 57.805 ;
        RECT 37.110 57.205 37.440 57.635 ;
        RECT 37.610 57.465 37.780 57.805 ;
        RECT 38.075 57.205 38.445 57.665 ;
        RECT 38.615 57.375 38.785 57.835 ;
        RECT 39.720 57.715 39.890 58.095 ;
        RECT 41.110 57.925 41.280 58.515 ;
        RECT 42.020 58.395 42.230 59.045 ;
        RECT 42.405 58.985 45.915 59.755 ;
        RECT 47.005 59.080 47.265 59.585 ;
        RECT 47.445 59.375 47.775 59.755 ;
        RECT 47.955 59.205 48.125 59.585 ;
        RECT 48.385 59.210 53.730 59.755 ;
        RECT 42.405 58.465 44.055 58.985 ;
        RECT 39.020 57.375 39.890 57.715 ;
        RECT 40.480 57.755 41.280 57.925 ;
        RECT 40.060 57.205 40.310 57.665 ;
        RECT 40.480 57.465 40.650 57.755 ;
        RECT 40.830 57.205 41.160 57.585 ;
        RECT 41.500 57.205 41.805 58.345 ;
        RECT 41.975 57.515 42.230 58.395 ;
        RECT 44.225 58.295 45.915 58.815 ;
        RECT 42.405 57.205 45.915 58.295 ;
        RECT 47.005 58.280 47.175 59.080 ;
        RECT 47.460 59.035 48.125 59.205 ;
        RECT 47.460 58.780 47.630 59.035 ;
        RECT 47.345 58.450 47.630 58.780 ;
        RECT 47.865 58.485 48.195 58.855 ;
        RECT 47.460 58.305 47.630 58.450 ;
        RECT 49.970 58.380 50.310 59.210 ;
        RECT 53.905 58.985 56.495 59.755 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 57.585 58.985 61.095 59.755 ;
        RECT 61.265 59.005 62.475 59.755 ;
        RECT 62.645 59.255 62.945 59.585 ;
        RECT 63.115 59.275 63.390 59.755 ;
        RECT 47.005 57.375 47.275 58.280 ;
        RECT 47.460 58.135 48.125 58.305 ;
        RECT 47.445 57.205 47.775 57.965 ;
        RECT 47.955 57.375 48.125 58.135 ;
        RECT 51.790 57.640 52.140 58.890 ;
        RECT 53.905 58.465 55.115 58.985 ;
        RECT 55.285 58.295 56.495 58.815 ;
        RECT 57.585 58.465 59.235 58.985 ;
        RECT 48.385 57.205 53.730 57.640 ;
        RECT 53.905 57.205 56.495 58.295 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 59.405 58.295 61.095 58.815 ;
        RECT 61.265 58.465 61.785 59.005 ;
        RECT 61.955 58.295 62.475 58.835 ;
        RECT 57.585 57.205 61.095 58.295 ;
        RECT 61.265 57.205 62.475 58.295 ;
        RECT 62.645 58.345 62.815 59.255 ;
        RECT 63.570 59.105 63.865 59.495 ;
        RECT 64.035 59.275 64.290 59.755 ;
        RECT 64.465 59.105 64.725 59.495 ;
        RECT 64.895 59.275 65.175 59.755 ;
        RECT 65.405 59.210 70.750 59.755 ;
        RECT 62.985 58.515 63.335 59.085 ;
        RECT 63.570 58.935 65.220 59.105 ;
        RECT 63.505 58.595 64.645 58.765 ;
        RECT 63.505 58.345 63.675 58.595 ;
        RECT 64.815 58.425 65.220 58.935 ;
        RECT 62.645 58.175 63.675 58.345 ;
        RECT 64.465 58.255 65.220 58.425 ;
        RECT 66.990 58.380 67.330 59.210 ;
        RECT 71.015 59.105 71.185 59.585 ;
        RECT 71.365 59.275 71.605 59.755 ;
        RECT 71.855 59.105 72.025 59.585 ;
        RECT 72.195 59.275 72.525 59.755 ;
        RECT 72.695 59.105 72.865 59.585 ;
        RECT 71.015 58.935 71.650 59.105 ;
        RECT 71.855 58.935 72.865 59.105 ;
        RECT 73.035 58.955 73.365 59.755 ;
        RECT 73.685 59.210 79.030 59.755 ;
        RECT 62.645 57.375 62.955 58.175 ;
        RECT 64.465 58.005 64.725 58.255 ;
        RECT 63.125 57.205 63.435 58.005 ;
        RECT 63.605 57.835 64.725 58.005 ;
        RECT 63.605 57.375 63.865 57.835 ;
        RECT 64.035 57.205 64.290 57.665 ;
        RECT 64.465 57.375 64.725 57.835 ;
        RECT 64.895 57.205 65.180 58.075 ;
        RECT 68.810 57.640 69.160 58.890 ;
        RECT 71.480 58.765 71.650 58.935 ;
        RECT 72.365 58.905 72.865 58.935 ;
        RECT 70.930 58.525 71.310 58.765 ;
        RECT 71.480 58.595 71.980 58.765 ;
        RECT 71.480 58.355 71.650 58.595 ;
        RECT 72.370 58.395 72.865 58.905 ;
        RECT 70.935 58.185 71.650 58.355 ;
        RECT 71.855 58.225 72.865 58.395 ;
        RECT 75.270 58.380 75.610 59.210 ;
        RECT 79.205 58.985 80.875 59.755 ;
        RECT 81.520 59.230 81.815 59.755 ;
        RECT 81.985 59.115 82.210 59.560 ;
        RECT 82.380 59.285 82.710 59.755 ;
        RECT 65.405 57.205 70.750 57.640 ;
        RECT 70.935 57.375 71.265 58.185 ;
        RECT 71.435 57.205 71.675 58.005 ;
        RECT 71.855 57.375 72.025 58.225 ;
        RECT 72.195 57.205 72.525 58.005 ;
        RECT 72.695 57.375 72.865 58.225 ;
        RECT 73.035 57.205 73.365 58.355 ;
        RECT 77.090 57.640 77.440 58.890 ;
        RECT 79.205 58.465 79.955 58.985 ;
        RECT 81.985 58.945 82.715 59.115 ;
        RECT 82.885 59.030 83.175 59.755 ;
        RECT 83.435 59.275 83.735 59.755 ;
        RECT 83.905 59.105 84.165 59.560 ;
        RECT 84.335 59.275 84.595 59.755 ;
        RECT 84.775 59.105 85.035 59.560 ;
        RECT 85.205 59.275 85.455 59.755 ;
        RECT 85.635 59.105 85.895 59.560 ;
        RECT 86.065 59.275 86.315 59.755 ;
        RECT 86.495 59.105 86.755 59.560 ;
        RECT 86.925 59.275 87.170 59.755 ;
        RECT 87.340 59.105 87.615 59.560 ;
        RECT 87.785 59.275 88.030 59.755 ;
        RECT 88.200 59.105 88.460 59.560 ;
        RECT 88.630 59.275 88.890 59.755 ;
        RECT 89.060 59.105 89.320 59.560 ;
        RECT 89.490 59.275 89.750 59.755 ;
        RECT 89.920 59.105 90.180 59.560 ;
        RECT 90.350 59.195 90.610 59.755 ;
        RECT 80.125 58.295 80.875 58.815 ;
        RECT 81.045 58.550 82.265 58.775 ;
        RECT 82.435 58.380 82.715 58.945 ;
        RECT 83.435 58.935 90.180 59.105 ;
        RECT 83.435 58.395 84.600 58.935 ;
        RECT 90.780 58.765 91.030 59.575 ;
        RECT 91.210 59.230 91.470 59.755 ;
        RECT 91.640 58.765 91.890 59.575 ;
        RECT 92.070 59.245 92.375 59.755 ;
        RECT 92.545 59.210 97.890 59.755 ;
        RECT 84.770 58.515 91.890 58.765 ;
        RECT 92.060 58.515 92.375 59.075 ;
        RECT 73.685 57.205 79.030 57.640 ;
        RECT 79.205 57.205 80.875 58.295 ;
        RECT 81.115 58.210 82.715 58.380 ;
        RECT 81.115 57.405 81.370 58.210 ;
        RECT 81.540 57.205 81.800 58.040 ;
        RECT 81.970 57.405 82.230 58.210 ;
        RECT 82.400 57.205 82.655 58.040 ;
        RECT 82.885 57.205 83.175 58.370 ;
        RECT 83.405 58.345 84.600 58.395 ;
        RECT 83.405 58.225 90.180 58.345 ;
        RECT 83.435 58.120 90.180 58.225 ;
        RECT 83.435 57.205 83.705 57.950 ;
        RECT 83.875 57.380 84.165 58.120 ;
        RECT 84.775 58.105 90.180 58.120 ;
        RECT 84.335 57.210 84.590 57.935 ;
        RECT 84.775 57.380 85.035 58.105 ;
        RECT 85.205 57.210 85.450 57.935 ;
        RECT 85.635 57.380 85.895 58.105 ;
        RECT 86.065 57.210 86.310 57.935 ;
        RECT 86.495 57.380 86.755 58.105 ;
        RECT 86.925 57.210 87.170 57.935 ;
        RECT 87.340 57.380 87.600 58.105 ;
        RECT 87.770 57.210 88.030 57.935 ;
        RECT 88.200 57.380 88.460 58.105 ;
        RECT 88.630 57.210 88.890 57.935 ;
        RECT 89.060 57.380 89.320 58.105 ;
        RECT 89.490 57.210 89.750 57.935 ;
        RECT 89.920 57.380 90.180 58.105 ;
        RECT 90.350 57.210 90.610 58.005 ;
        RECT 90.780 57.380 91.030 58.515 ;
        RECT 84.335 57.205 90.610 57.210 ;
        RECT 91.210 57.205 91.470 58.015 ;
        RECT 91.645 57.375 91.890 58.515 ;
        RECT 94.130 58.380 94.470 59.210 ;
        RECT 98.065 58.985 100.655 59.755 ;
        RECT 101.295 59.265 101.625 59.755 ;
        RECT 101.795 59.160 102.415 59.585 ;
        RECT 92.070 57.205 92.365 58.015 ;
        RECT 95.950 57.640 96.300 58.890 ;
        RECT 98.065 58.465 99.275 58.985 ;
        RECT 99.445 58.295 100.655 58.815 ;
        RECT 101.285 58.515 101.625 59.095 ;
        RECT 101.795 58.825 102.155 59.160 ;
        RECT 102.875 59.065 103.205 59.755 ;
        RECT 104.250 58.975 104.750 59.585 ;
        RECT 101.795 58.545 103.215 58.825 ;
        RECT 92.545 57.205 97.890 57.640 ;
        RECT 98.065 57.205 100.655 58.295 ;
        RECT 101.295 57.205 101.625 58.345 ;
        RECT 101.795 57.375 102.155 58.545 ;
        RECT 102.355 57.205 102.685 58.375 ;
        RECT 102.885 57.375 103.215 58.545 ;
        RECT 104.045 58.515 104.395 58.765 ;
        RECT 103.415 57.205 103.745 58.375 ;
        RECT 104.580 58.345 104.750 58.975 ;
        RECT 105.380 59.105 105.710 59.585 ;
        RECT 105.880 59.295 106.105 59.755 ;
        RECT 106.275 59.105 106.605 59.585 ;
        RECT 105.380 58.935 106.605 59.105 ;
        RECT 106.795 58.955 107.045 59.755 ;
        RECT 107.215 58.955 107.555 59.585 ;
        RECT 108.645 59.030 108.935 59.755 ;
        RECT 104.920 58.565 105.250 58.765 ;
        RECT 105.420 58.565 105.750 58.765 ;
        RECT 105.920 58.565 106.340 58.765 ;
        RECT 106.515 58.595 107.210 58.765 ;
        RECT 106.515 58.345 106.685 58.595 ;
        RECT 107.380 58.345 107.555 58.955 ;
        RECT 109.105 59.005 110.315 59.755 ;
        RECT 109.105 58.465 109.625 59.005 ;
        RECT 110.545 58.935 110.755 59.755 ;
        RECT 110.925 58.955 111.255 59.585 ;
        RECT 104.250 58.175 106.685 58.345 ;
        RECT 104.250 57.375 104.580 58.175 ;
        RECT 104.750 57.205 105.080 58.005 ;
        RECT 105.380 57.375 105.710 58.175 ;
        RECT 106.355 57.205 106.605 58.005 ;
        RECT 106.875 57.205 107.045 58.345 ;
        RECT 107.215 57.375 107.555 58.345 ;
        RECT 108.645 57.205 108.935 58.370 ;
        RECT 109.795 58.295 110.315 58.835 ;
        RECT 110.925 58.355 111.175 58.955 ;
        RECT 111.425 58.935 111.655 59.755 ;
        RECT 111.865 59.210 117.210 59.755 ;
        RECT 117.385 59.210 122.730 59.755 ;
        RECT 111.345 58.515 111.675 58.765 ;
        RECT 113.450 58.380 113.790 59.210 ;
        RECT 109.105 57.205 110.315 58.295 ;
        RECT 110.545 57.205 110.755 58.345 ;
        RECT 110.925 57.375 111.255 58.355 ;
        RECT 111.425 57.205 111.655 58.345 ;
        RECT 115.270 57.640 115.620 58.890 ;
        RECT 118.970 58.380 119.310 59.210 ;
        RECT 122.905 59.005 124.115 59.755 ;
        RECT 124.285 59.005 125.495 59.755 ;
        RECT 120.790 57.640 121.140 58.890 ;
        RECT 122.905 58.465 123.425 59.005 ;
        RECT 123.595 58.295 124.115 58.835 ;
        RECT 111.865 57.205 117.210 57.640 ;
        RECT 117.385 57.205 122.730 57.640 ;
        RECT 122.905 57.205 124.115 58.295 ;
        RECT 124.285 58.295 124.805 58.835 ;
        RECT 124.975 58.465 125.495 59.005 ;
        RECT 124.285 57.205 125.495 58.295 ;
        RECT 5.520 57.035 125.580 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 6.985 55.945 8.195 57.035 ;
        RECT 8.370 56.365 8.625 56.865 ;
        RECT 8.795 56.535 9.125 57.035 ;
        RECT 8.370 56.195 9.120 56.365 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 6.985 55.235 7.505 55.775 ;
        RECT 7.675 55.405 8.195 55.945 ;
        RECT 8.370 55.375 8.720 56.025 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 6.985 54.485 8.195 55.235 ;
        RECT 8.890 55.205 9.120 56.195 ;
        RECT 8.370 55.035 9.120 55.205 ;
        RECT 8.370 54.745 8.625 55.035 ;
        RECT 8.795 54.485 9.125 54.865 ;
        RECT 9.295 54.745 9.465 56.865 ;
        RECT 9.635 56.065 9.960 56.850 ;
        RECT 10.130 56.575 10.380 57.035 ;
        RECT 10.550 56.535 10.800 56.865 ;
        RECT 11.015 56.535 11.695 56.865 ;
        RECT 10.550 56.405 10.720 56.535 ;
        RECT 10.325 56.235 10.720 56.405 ;
        RECT 9.695 55.015 10.155 56.065 ;
        RECT 10.325 54.875 10.495 56.235 ;
        RECT 10.890 55.975 11.355 56.365 ;
        RECT 10.665 55.165 11.015 55.785 ;
        RECT 11.185 55.385 11.355 55.975 ;
        RECT 11.525 55.755 11.695 56.535 ;
        RECT 11.865 56.435 12.035 56.775 ;
        RECT 12.270 56.605 12.600 57.035 ;
        RECT 12.770 56.435 12.940 56.775 ;
        RECT 13.235 56.575 13.605 57.035 ;
        RECT 11.865 56.265 12.940 56.435 ;
        RECT 13.775 56.405 13.945 56.865 ;
        RECT 14.180 56.525 15.050 56.865 ;
        RECT 15.220 56.575 15.470 57.035 ;
        RECT 13.385 56.235 13.945 56.405 ;
        RECT 13.385 56.095 13.555 56.235 ;
        RECT 12.055 55.925 13.555 56.095 ;
        RECT 14.250 56.065 14.710 56.355 ;
        RECT 11.525 55.585 13.215 55.755 ;
        RECT 11.185 55.165 11.540 55.385 ;
        RECT 11.710 54.875 11.880 55.585 ;
        RECT 12.085 55.165 12.875 55.415 ;
        RECT 13.045 55.405 13.215 55.585 ;
        RECT 13.385 55.235 13.555 55.925 ;
        RECT 9.825 54.485 10.155 54.845 ;
        RECT 10.325 54.705 10.820 54.875 ;
        RECT 11.025 54.705 11.880 54.875 ;
        RECT 12.755 54.485 13.085 54.945 ;
        RECT 13.295 54.845 13.555 55.235 ;
        RECT 13.745 56.055 14.710 56.065 ;
        RECT 14.880 56.145 15.050 56.525 ;
        RECT 15.640 56.485 15.810 56.775 ;
        RECT 15.990 56.655 16.320 57.035 ;
        RECT 15.640 56.315 16.440 56.485 ;
        RECT 13.745 55.895 14.420 56.055 ;
        RECT 14.880 55.975 16.100 56.145 ;
        RECT 13.745 55.105 13.955 55.895 ;
        RECT 14.880 55.885 15.050 55.975 ;
        RECT 14.125 55.105 14.475 55.725 ;
        RECT 14.645 55.715 15.050 55.885 ;
        RECT 14.645 54.935 14.815 55.715 ;
        RECT 14.985 55.265 15.205 55.545 ;
        RECT 15.385 55.435 15.925 55.805 ;
        RECT 16.270 55.725 16.440 56.315 ;
        RECT 16.660 55.895 16.965 57.035 ;
        RECT 17.135 55.845 17.390 56.725 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 19.520 56.405 19.805 56.865 ;
        RECT 19.975 56.575 20.245 57.035 ;
        RECT 19.520 56.185 20.475 56.405 ;
        RECT 16.270 55.695 17.010 55.725 ;
        RECT 14.985 55.095 15.515 55.265 ;
        RECT 13.295 54.675 13.645 54.845 ;
        RECT 13.865 54.655 14.815 54.935 ;
        RECT 14.985 54.485 15.175 54.925 ;
        RECT 15.345 54.865 15.515 55.095 ;
        RECT 15.685 55.035 15.925 55.435 ;
        RECT 16.095 55.395 17.010 55.695 ;
        RECT 16.095 55.220 16.420 55.395 ;
        RECT 16.095 54.865 16.415 55.220 ;
        RECT 17.180 55.195 17.390 55.845 ;
        RECT 19.405 55.455 20.095 56.015 ;
        RECT 20.265 55.285 20.475 56.185 ;
        RECT 15.345 54.695 16.415 54.865 ;
        RECT 16.660 54.485 16.965 54.945 ;
        RECT 17.135 54.665 17.390 55.195 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 19.520 55.115 20.475 55.285 ;
        RECT 20.645 56.015 21.045 56.865 ;
        RECT 21.235 56.405 21.515 56.865 ;
        RECT 22.035 56.575 22.360 57.035 ;
        RECT 21.235 56.185 22.360 56.405 ;
        RECT 20.645 55.455 21.740 56.015 ;
        RECT 21.910 55.725 22.360 56.185 ;
        RECT 22.530 55.895 22.915 56.865 ;
        RECT 23.290 56.065 23.620 56.865 ;
        RECT 23.790 56.235 24.120 57.035 ;
        RECT 24.420 56.065 24.750 56.865 ;
        RECT 25.395 56.235 25.645 57.035 ;
        RECT 23.290 55.895 25.725 56.065 ;
        RECT 25.915 55.895 26.085 57.035 ;
        RECT 26.255 55.895 26.595 56.865 ;
        RECT 26.765 56.600 32.110 57.035 ;
        RECT 19.520 54.655 19.805 55.115 ;
        RECT 19.975 54.485 20.245 54.945 ;
        RECT 20.645 54.655 21.045 55.455 ;
        RECT 21.910 55.395 22.465 55.725 ;
        RECT 21.910 55.285 22.360 55.395 ;
        RECT 21.235 55.115 22.360 55.285 ;
        RECT 22.635 55.225 22.915 55.895 ;
        RECT 23.085 55.475 23.435 55.725 ;
        RECT 23.620 55.265 23.790 55.895 ;
        RECT 23.960 55.475 24.290 55.675 ;
        RECT 24.460 55.475 24.790 55.675 ;
        RECT 24.960 55.475 25.380 55.675 ;
        RECT 25.555 55.645 25.725 55.895 ;
        RECT 25.555 55.475 26.250 55.645 ;
        RECT 21.235 54.655 21.515 55.115 ;
        RECT 22.035 54.485 22.360 54.945 ;
        RECT 22.530 54.655 22.915 55.225 ;
        RECT 23.290 54.655 23.790 55.265 ;
        RECT 24.420 55.135 25.645 55.305 ;
        RECT 26.420 55.285 26.595 55.895 ;
        RECT 24.420 54.655 24.750 55.135 ;
        RECT 24.920 54.485 25.145 54.945 ;
        RECT 25.315 54.655 25.645 55.135 ;
        RECT 25.835 54.485 26.085 55.285 ;
        RECT 26.255 54.655 26.595 55.285 ;
        RECT 28.350 55.030 28.690 55.860 ;
        RECT 30.170 55.350 30.520 56.600 ;
        RECT 32.285 55.945 35.795 57.035 ;
        RECT 32.285 55.255 33.935 55.775 ;
        RECT 34.105 55.425 35.795 55.945 ;
        RECT 35.965 55.960 36.235 56.865 ;
        RECT 36.405 56.275 36.735 57.035 ;
        RECT 36.915 56.105 37.085 56.865 ;
        RECT 26.765 54.485 32.110 55.030 ;
        RECT 32.285 54.485 35.795 55.255 ;
        RECT 35.965 55.160 36.135 55.960 ;
        RECT 36.420 55.935 37.085 56.105 ;
        RECT 36.420 55.790 36.590 55.935 ;
        RECT 38.305 55.895 38.535 57.035 ;
        RECT 38.705 55.885 39.035 56.865 ;
        RECT 39.205 55.895 39.415 57.035 ;
        RECT 40.175 56.030 40.430 56.835 ;
        RECT 40.600 56.200 40.860 57.035 ;
        RECT 41.030 56.030 41.290 56.835 ;
        RECT 41.460 56.200 41.715 57.035 ;
        RECT 36.305 55.460 36.590 55.790 ;
        RECT 36.420 55.205 36.590 55.460 ;
        RECT 36.825 55.385 37.155 55.755 ;
        RECT 38.285 55.475 38.615 55.725 ;
        RECT 35.965 54.655 36.225 55.160 ;
        RECT 36.420 55.035 37.085 55.205 ;
        RECT 36.405 54.485 36.735 54.865 ;
        RECT 36.915 54.655 37.085 55.035 ;
        RECT 38.305 54.485 38.535 55.305 ;
        RECT 38.785 55.285 39.035 55.885 ;
        RECT 40.175 55.860 41.775 56.030 ;
        RECT 41.945 55.945 43.615 57.035 ;
        RECT 40.105 55.465 41.325 55.690 ;
        RECT 38.705 54.655 39.035 55.285 ;
        RECT 39.205 54.485 39.415 55.305 ;
        RECT 41.495 55.295 41.775 55.860 ;
        RECT 41.045 55.125 41.775 55.295 ;
        RECT 41.945 55.255 42.695 55.775 ;
        RECT 42.865 55.425 43.615 55.945 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 44.705 55.945 46.375 57.035 ;
        RECT 44.705 55.255 45.455 55.775 ;
        RECT 45.625 55.425 46.375 55.945 ;
        RECT 47.155 55.885 47.485 57.035 ;
        RECT 47.655 56.015 47.825 56.865 ;
        RECT 47.995 56.235 48.325 57.035 ;
        RECT 48.495 56.015 48.665 56.865 ;
        RECT 48.845 56.235 49.085 57.035 ;
        RECT 49.255 56.055 49.585 56.865 ;
        RECT 49.820 56.165 50.105 57.035 ;
        RECT 50.275 56.405 50.535 56.865 ;
        RECT 50.710 56.575 50.965 57.035 ;
        RECT 51.135 56.405 51.395 56.865 ;
        RECT 50.275 56.235 51.395 56.405 ;
        RECT 51.565 56.235 51.875 57.035 ;
        RECT 47.655 55.845 48.665 56.015 ;
        RECT 48.870 55.885 49.585 56.055 ;
        RECT 50.275 55.985 50.535 56.235 ;
        RECT 52.045 56.065 52.355 56.865 ;
        RECT 52.525 56.600 57.870 57.035 ;
        RECT 47.655 55.335 48.150 55.845 ;
        RECT 48.870 55.645 49.040 55.885 ;
        RECT 49.780 55.815 50.535 55.985 ;
        RECT 51.325 55.895 52.355 56.065 ;
        RECT 48.540 55.475 49.040 55.645 ;
        RECT 49.210 55.475 49.590 55.715 ;
        RECT 47.655 55.305 48.155 55.335 ;
        RECT 48.870 55.305 49.040 55.475 ;
        RECT 49.780 55.305 50.185 55.815 ;
        RECT 51.325 55.645 51.495 55.895 ;
        RECT 50.355 55.475 51.495 55.645 ;
        RECT 40.580 54.485 40.875 55.010 ;
        RECT 41.045 54.680 41.270 55.125 ;
        RECT 41.440 54.485 41.770 54.955 ;
        RECT 41.945 54.485 43.615 55.255 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 44.705 54.485 46.375 55.255 ;
        RECT 47.155 54.485 47.485 55.285 ;
        RECT 47.655 55.135 48.665 55.305 ;
        RECT 48.870 55.135 49.505 55.305 ;
        RECT 49.780 55.135 51.430 55.305 ;
        RECT 51.665 55.155 52.015 55.725 ;
        RECT 47.655 54.655 47.825 55.135 ;
        RECT 47.995 54.485 48.325 54.965 ;
        RECT 48.495 54.655 48.665 55.135 ;
        RECT 48.915 54.485 49.155 54.965 ;
        RECT 49.335 54.655 49.505 55.135 ;
        RECT 49.825 54.485 50.105 54.965 ;
        RECT 50.275 54.745 50.535 55.135 ;
        RECT 50.710 54.485 50.965 54.965 ;
        RECT 51.135 54.745 51.430 55.135 ;
        RECT 52.185 54.985 52.355 55.895 ;
        RECT 54.110 55.030 54.450 55.860 ;
        RECT 55.930 55.350 56.280 56.600 ;
        RECT 58.045 55.945 61.555 57.035 ;
        RECT 58.045 55.255 59.695 55.775 ;
        RECT 59.865 55.425 61.555 55.945 ;
        RECT 62.185 56.445 62.885 56.865 ;
        RECT 63.085 56.675 63.415 57.035 ;
        RECT 63.585 56.445 63.915 56.845 ;
        RECT 62.185 56.215 63.915 56.445 ;
        RECT 62.185 55.335 62.390 56.215 ;
        RECT 62.560 55.475 62.890 56.015 ;
        RECT 63.065 55.725 63.390 56.015 ;
        RECT 63.585 55.995 63.915 56.215 ;
        RECT 64.085 55.725 64.255 56.650 ;
        RECT 64.435 55.975 64.765 57.035 ;
        RECT 65.410 55.885 65.670 57.035 ;
        RECT 65.845 55.960 66.100 56.865 ;
        RECT 66.270 56.275 66.600 57.035 ;
        RECT 66.815 56.105 66.985 56.865 ;
        RECT 63.065 55.395 63.560 55.725 ;
        RECT 63.880 55.395 64.255 55.725 ;
        RECT 64.465 55.395 64.775 55.725 ;
        RECT 51.610 54.485 51.885 54.965 ;
        RECT 52.055 54.655 52.355 54.985 ;
        RECT 52.525 54.485 57.870 55.030 ;
        RECT 58.045 54.485 61.555 55.255 ;
        RECT 62.185 55.245 62.415 55.335 ;
        RECT 62.185 54.655 62.895 55.245 ;
        RECT 63.405 55.015 64.765 55.225 ;
        RECT 63.405 54.655 63.735 55.015 ;
        RECT 63.935 54.485 64.265 54.845 ;
        RECT 64.435 54.655 64.765 55.015 ;
        RECT 65.410 54.485 65.670 55.325 ;
        RECT 65.845 55.230 66.015 55.960 ;
        RECT 66.270 55.935 66.985 56.105 ;
        RECT 67.335 56.105 67.505 56.865 ;
        RECT 67.720 56.275 68.050 57.035 ;
        RECT 67.335 55.935 68.050 56.105 ;
        RECT 68.220 55.960 68.475 56.865 ;
        RECT 66.270 55.725 66.440 55.935 ;
        RECT 66.185 55.395 66.440 55.725 ;
        RECT 65.845 54.655 66.100 55.230 ;
        RECT 66.270 55.205 66.440 55.395 ;
        RECT 66.720 55.385 67.075 55.755 ;
        RECT 67.245 55.385 67.600 55.755 ;
        RECT 67.880 55.725 68.050 55.935 ;
        RECT 67.880 55.395 68.135 55.725 ;
        RECT 67.880 55.205 68.050 55.395 ;
        RECT 68.305 55.230 68.475 55.960 ;
        RECT 68.650 55.885 68.910 57.035 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 70.465 56.600 75.810 57.035 ;
        RECT 75.985 56.600 81.330 57.035 ;
        RECT 81.505 56.600 86.850 57.035 ;
        RECT 66.270 55.035 66.985 55.205 ;
        RECT 66.270 54.485 66.600 54.865 ;
        RECT 66.815 54.655 66.985 55.035 ;
        RECT 67.335 55.035 68.050 55.205 ;
        RECT 67.335 54.655 67.505 55.035 ;
        RECT 67.720 54.485 68.050 54.865 ;
        RECT 68.220 54.655 68.475 55.230 ;
        RECT 68.650 54.485 68.910 55.325 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 72.050 55.030 72.390 55.860 ;
        RECT 73.870 55.350 74.220 56.600 ;
        RECT 77.570 55.030 77.910 55.860 ;
        RECT 79.390 55.350 79.740 56.600 ;
        RECT 83.090 55.030 83.430 55.860 ;
        RECT 84.910 55.350 85.260 56.600 ;
        RECT 87.025 55.945 89.615 57.035 ;
        RECT 87.025 55.255 88.235 55.775 ;
        RECT 88.405 55.425 89.615 55.945 ;
        RECT 89.990 56.065 90.320 56.865 ;
        RECT 90.490 56.235 90.820 57.035 ;
        RECT 91.120 56.065 91.450 56.865 ;
        RECT 92.095 56.235 92.345 57.035 ;
        RECT 89.990 55.895 92.425 56.065 ;
        RECT 92.615 55.895 92.785 57.035 ;
        RECT 92.955 55.895 93.295 56.865 ;
        RECT 93.465 55.945 95.135 57.035 ;
        RECT 89.785 55.475 90.135 55.725 ;
        RECT 90.320 55.265 90.490 55.895 ;
        RECT 90.660 55.475 90.990 55.675 ;
        RECT 91.160 55.475 91.490 55.675 ;
        RECT 91.660 55.475 92.080 55.675 ;
        RECT 92.255 55.645 92.425 55.895 ;
        RECT 92.255 55.475 92.950 55.645 ;
        RECT 70.465 54.485 75.810 55.030 ;
        RECT 75.985 54.485 81.330 55.030 ;
        RECT 81.505 54.485 86.850 55.030 ;
        RECT 87.025 54.485 89.615 55.255 ;
        RECT 89.990 54.655 90.490 55.265 ;
        RECT 91.120 55.135 92.345 55.305 ;
        RECT 93.120 55.285 93.295 55.895 ;
        RECT 91.120 54.655 91.450 55.135 ;
        RECT 91.620 54.485 91.845 54.945 ;
        RECT 92.015 54.655 92.345 55.135 ;
        RECT 92.535 54.485 92.785 55.285 ;
        RECT 92.955 54.655 93.295 55.285 ;
        RECT 93.465 55.255 94.215 55.775 ;
        RECT 94.385 55.425 95.135 55.945 ;
        RECT 95.765 55.870 96.055 57.035 ;
        RECT 96.225 55.945 97.895 57.035 ;
        RECT 96.225 55.255 96.975 55.775 ;
        RECT 97.145 55.425 97.895 55.945 ;
        RECT 98.730 56.065 99.060 56.865 ;
        RECT 99.230 56.235 99.560 57.035 ;
        RECT 99.860 56.065 100.190 56.865 ;
        RECT 100.835 56.235 101.085 57.035 ;
        RECT 98.730 55.895 101.165 56.065 ;
        RECT 101.355 55.895 101.525 57.035 ;
        RECT 101.695 55.895 102.035 56.865 ;
        RECT 102.215 56.225 102.510 57.035 ;
        RECT 98.525 55.475 98.875 55.725 ;
        RECT 99.060 55.265 99.230 55.895 ;
        RECT 99.400 55.475 99.730 55.675 ;
        RECT 99.900 55.475 100.230 55.675 ;
        RECT 100.400 55.475 100.820 55.675 ;
        RECT 100.995 55.645 101.165 55.895 ;
        RECT 100.995 55.475 101.690 55.645 ;
        RECT 93.465 54.485 95.135 55.255 ;
        RECT 95.765 54.485 96.055 55.210 ;
        RECT 96.225 54.485 97.895 55.255 ;
        RECT 98.730 54.655 99.230 55.265 ;
        RECT 99.860 55.135 101.085 55.305 ;
        RECT 101.860 55.285 102.035 55.895 ;
        RECT 102.690 55.725 102.935 56.865 ;
        RECT 103.110 56.225 103.370 57.035 ;
        RECT 103.970 57.030 110.245 57.035 ;
        RECT 103.550 55.725 103.800 56.860 ;
        RECT 103.970 56.235 104.230 57.030 ;
        RECT 104.400 56.135 104.660 56.860 ;
        RECT 104.830 56.305 105.090 57.030 ;
        RECT 105.260 56.135 105.520 56.860 ;
        RECT 105.690 56.305 105.950 57.030 ;
        RECT 106.120 56.135 106.380 56.860 ;
        RECT 106.550 56.305 106.810 57.030 ;
        RECT 106.980 56.135 107.240 56.860 ;
        RECT 107.410 56.305 107.655 57.030 ;
        RECT 107.825 56.135 108.085 56.860 ;
        RECT 108.270 56.305 108.515 57.030 ;
        RECT 108.685 56.135 108.945 56.860 ;
        RECT 109.130 56.305 109.375 57.030 ;
        RECT 109.545 56.135 109.805 56.860 ;
        RECT 109.990 56.305 110.245 57.030 ;
        RECT 104.400 56.120 109.805 56.135 ;
        RECT 110.415 56.120 110.705 56.860 ;
        RECT 110.875 56.290 111.145 57.035 ;
        RECT 104.400 56.015 111.145 56.120 ;
        RECT 104.400 55.895 111.175 56.015 ;
        RECT 111.465 55.895 111.675 57.035 ;
        RECT 109.980 55.845 111.175 55.895 ;
        RECT 111.845 55.885 112.175 56.865 ;
        RECT 112.345 55.895 112.575 57.035 ;
        RECT 112.785 56.600 118.130 57.035 ;
        RECT 99.860 54.655 100.190 55.135 ;
        RECT 100.360 54.485 100.585 54.945 ;
        RECT 100.755 54.655 101.085 55.135 ;
        RECT 101.275 54.485 101.525 55.285 ;
        RECT 101.695 54.655 102.035 55.285 ;
        RECT 102.205 55.165 102.520 55.725 ;
        RECT 102.690 55.475 109.810 55.725 ;
        RECT 102.205 54.485 102.510 54.995 ;
        RECT 102.690 54.665 102.940 55.475 ;
        RECT 103.110 54.485 103.370 55.010 ;
        RECT 103.550 54.665 103.800 55.475 ;
        RECT 109.980 55.305 111.145 55.845 ;
        RECT 104.400 55.135 111.145 55.305 ;
        RECT 103.970 54.485 104.230 55.045 ;
        RECT 104.400 54.680 104.660 55.135 ;
        RECT 104.830 54.485 105.090 54.965 ;
        RECT 105.260 54.680 105.520 55.135 ;
        RECT 105.690 54.485 105.950 54.965 ;
        RECT 106.120 54.680 106.380 55.135 ;
        RECT 106.550 54.485 106.795 54.965 ;
        RECT 106.965 54.680 107.240 55.135 ;
        RECT 107.410 54.485 107.655 54.965 ;
        RECT 107.825 54.680 108.085 55.135 ;
        RECT 108.265 54.485 108.515 54.965 ;
        RECT 108.685 54.680 108.945 55.135 ;
        RECT 109.125 54.485 109.375 54.965 ;
        RECT 109.545 54.680 109.805 55.135 ;
        RECT 109.985 54.485 110.245 54.965 ;
        RECT 110.415 54.680 110.675 55.135 ;
        RECT 110.845 54.485 111.145 54.965 ;
        RECT 111.465 54.485 111.675 55.305 ;
        RECT 111.845 55.285 112.095 55.885 ;
        RECT 112.265 55.475 112.595 55.725 ;
        RECT 111.845 54.655 112.175 55.285 ;
        RECT 112.345 54.485 112.575 55.305 ;
        RECT 114.370 55.030 114.710 55.860 ;
        RECT 116.190 55.350 116.540 56.600 ;
        RECT 118.305 55.945 120.895 57.035 ;
        RECT 118.305 55.255 119.515 55.775 ;
        RECT 119.685 55.425 120.895 55.945 ;
        RECT 121.525 55.870 121.815 57.035 ;
        RECT 121.985 55.945 123.655 57.035 ;
        RECT 121.985 55.255 122.735 55.775 ;
        RECT 122.905 55.425 123.655 55.945 ;
        RECT 124.285 55.945 125.495 57.035 ;
        RECT 124.285 55.405 124.805 55.945 ;
        RECT 112.785 54.485 118.130 55.030 ;
        RECT 118.305 54.485 120.895 55.255 ;
        RECT 121.525 54.485 121.815 55.210 ;
        RECT 121.985 54.485 123.655 55.255 ;
        RECT 124.975 55.235 125.495 55.775 ;
        RECT 124.285 54.485 125.495 55.235 ;
        RECT 5.520 54.315 125.580 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.985 53.545 9.575 54.315 ;
        RECT 10.205 53.815 10.465 54.145 ;
        RECT 10.675 53.835 10.950 54.315 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 6.985 53.025 8.195 53.545 ;
        RECT 8.365 52.855 9.575 53.375 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 6.985 51.765 9.575 52.855 ;
        RECT 10.205 52.905 10.375 53.815 ;
        RECT 11.160 53.745 11.365 54.145 ;
        RECT 11.535 53.915 11.870 54.315 ;
        RECT 10.545 53.075 10.905 53.655 ;
        RECT 11.160 53.575 11.845 53.745 ;
        RECT 11.085 52.905 11.335 53.405 ;
        RECT 10.205 52.735 11.335 52.905 ;
        RECT 10.205 51.965 10.475 52.735 ;
        RECT 11.505 52.545 11.845 53.575 ;
        RECT 12.045 53.545 13.715 54.315 ;
        RECT 12.045 53.025 12.795 53.545 ;
        RECT 14.405 53.495 14.615 54.315 ;
        RECT 14.785 53.515 15.115 54.145 ;
        RECT 12.965 52.855 13.715 53.375 ;
        RECT 14.785 52.915 15.035 53.515 ;
        RECT 15.285 53.495 15.515 54.315 ;
        RECT 15.725 53.545 19.235 54.315 ;
        RECT 15.205 53.075 15.535 53.325 ;
        RECT 15.725 53.025 17.375 53.545 ;
        RECT 19.610 53.535 20.110 54.145 ;
        RECT 10.645 51.765 10.975 52.545 ;
        RECT 11.180 52.370 11.845 52.545 ;
        RECT 11.180 51.965 11.365 52.370 ;
        RECT 11.535 51.765 11.870 52.190 ;
        RECT 12.045 51.765 13.715 52.855 ;
        RECT 14.405 51.765 14.615 52.905 ;
        RECT 14.785 51.935 15.115 52.915 ;
        RECT 15.285 51.765 15.515 52.905 ;
        RECT 17.545 52.855 19.235 53.375 ;
        RECT 19.405 53.075 19.755 53.325 ;
        RECT 19.940 52.905 20.110 53.535 ;
        RECT 20.740 53.665 21.070 54.145 ;
        RECT 21.240 53.855 21.465 54.315 ;
        RECT 21.635 53.665 21.965 54.145 ;
        RECT 20.740 53.495 21.965 53.665 ;
        RECT 22.155 53.515 22.405 54.315 ;
        RECT 22.575 53.515 22.915 54.145 ;
        RECT 23.290 53.535 23.790 54.145 ;
        RECT 20.280 53.125 20.610 53.325 ;
        RECT 20.780 53.125 21.110 53.325 ;
        RECT 21.280 53.125 21.700 53.325 ;
        RECT 21.875 53.155 22.570 53.325 ;
        RECT 21.875 52.905 22.045 53.155 ;
        RECT 22.740 52.905 22.915 53.515 ;
        RECT 23.085 53.075 23.435 53.325 ;
        RECT 23.620 52.905 23.790 53.535 ;
        RECT 24.420 53.665 24.750 54.145 ;
        RECT 24.920 53.855 25.145 54.315 ;
        RECT 25.315 53.665 25.645 54.145 ;
        RECT 24.420 53.495 25.645 53.665 ;
        RECT 25.835 53.515 26.085 54.315 ;
        RECT 26.255 53.515 26.595 54.145 ;
        RECT 26.970 53.535 27.470 54.145 ;
        RECT 23.960 53.125 24.290 53.325 ;
        RECT 24.460 53.125 24.790 53.325 ;
        RECT 24.960 53.125 25.380 53.325 ;
        RECT 25.555 53.155 26.250 53.325 ;
        RECT 25.555 52.905 25.725 53.155 ;
        RECT 26.420 52.905 26.595 53.515 ;
        RECT 26.765 53.075 27.115 53.325 ;
        RECT 27.300 52.905 27.470 53.535 ;
        RECT 28.100 53.665 28.430 54.145 ;
        RECT 28.600 53.855 28.825 54.315 ;
        RECT 28.995 53.665 29.325 54.145 ;
        RECT 28.100 53.495 29.325 53.665 ;
        RECT 29.515 53.515 29.765 54.315 ;
        RECT 29.935 53.515 30.275 54.145 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 27.640 53.125 27.970 53.325 ;
        RECT 28.140 53.125 28.470 53.325 ;
        RECT 28.640 53.125 29.060 53.325 ;
        RECT 29.235 53.155 29.930 53.325 ;
        RECT 29.235 52.905 29.405 53.155 ;
        RECT 30.100 52.905 30.275 53.515 ;
        RECT 31.825 53.565 33.035 54.315 ;
        RECT 31.825 53.025 32.345 53.565 ;
        RECT 33.410 53.535 33.910 54.145 ;
        RECT 15.725 51.765 19.235 52.855 ;
        RECT 19.610 52.735 22.045 52.905 ;
        RECT 19.610 51.935 19.940 52.735 ;
        RECT 20.110 51.765 20.440 52.565 ;
        RECT 20.740 51.935 21.070 52.735 ;
        RECT 21.715 51.765 21.965 52.565 ;
        RECT 22.235 51.765 22.405 52.905 ;
        RECT 22.575 51.935 22.915 52.905 ;
        RECT 23.290 52.735 25.725 52.905 ;
        RECT 23.290 51.935 23.620 52.735 ;
        RECT 23.790 51.765 24.120 52.565 ;
        RECT 24.420 51.935 24.750 52.735 ;
        RECT 25.395 51.765 25.645 52.565 ;
        RECT 25.915 51.765 26.085 52.905 ;
        RECT 26.255 51.935 26.595 52.905 ;
        RECT 26.970 52.735 29.405 52.905 ;
        RECT 26.970 51.935 27.300 52.735 ;
        RECT 27.470 51.765 27.800 52.565 ;
        RECT 28.100 51.935 28.430 52.735 ;
        RECT 29.075 51.765 29.325 52.565 ;
        RECT 29.595 51.765 29.765 52.905 ;
        RECT 29.935 51.935 30.275 52.905 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 32.515 52.855 33.035 53.395 ;
        RECT 33.205 53.075 33.555 53.325 ;
        RECT 33.740 52.905 33.910 53.535 ;
        RECT 34.540 53.665 34.870 54.145 ;
        RECT 35.040 53.855 35.265 54.315 ;
        RECT 35.435 53.665 35.765 54.145 ;
        RECT 34.540 53.495 35.765 53.665 ;
        RECT 35.955 53.515 36.205 54.315 ;
        RECT 36.375 53.515 36.715 54.145 ;
        RECT 34.080 53.125 34.410 53.325 ;
        RECT 34.580 53.125 34.910 53.325 ;
        RECT 35.080 53.125 35.500 53.325 ;
        RECT 35.675 53.155 36.370 53.325 ;
        RECT 35.675 52.905 35.845 53.155 ;
        RECT 36.540 52.905 36.715 53.515 ;
        RECT 36.885 53.545 39.475 54.315 ;
        RECT 40.195 53.835 40.495 54.315 ;
        RECT 40.665 53.665 40.925 54.120 ;
        RECT 41.095 53.835 41.355 54.315 ;
        RECT 41.535 53.665 41.795 54.120 ;
        RECT 41.965 53.835 42.215 54.315 ;
        RECT 42.395 53.665 42.655 54.120 ;
        RECT 42.825 53.835 43.075 54.315 ;
        RECT 43.255 53.665 43.515 54.120 ;
        RECT 43.685 53.835 43.930 54.315 ;
        RECT 44.100 53.665 44.375 54.120 ;
        RECT 44.545 53.835 44.790 54.315 ;
        RECT 44.960 53.665 45.220 54.120 ;
        RECT 45.390 53.835 45.650 54.315 ;
        RECT 45.820 53.665 46.080 54.120 ;
        RECT 46.250 53.835 46.510 54.315 ;
        RECT 46.680 53.665 46.940 54.120 ;
        RECT 47.110 53.755 47.370 54.315 ;
        RECT 36.885 53.025 38.095 53.545 ;
        RECT 40.195 53.495 46.940 53.665 ;
        RECT 31.825 51.765 33.035 52.855 ;
        RECT 33.410 52.735 35.845 52.905 ;
        RECT 33.410 51.935 33.740 52.735 ;
        RECT 33.910 51.765 34.240 52.565 ;
        RECT 34.540 51.935 34.870 52.735 ;
        RECT 35.515 51.765 35.765 52.565 ;
        RECT 36.035 51.765 36.205 52.905 ;
        RECT 36.375 51.935 36.715 52.905 ;
        RECT 38.265 52.855 39.475 53.375 ;
        RECT 36.885 51.765 39.475 52.855 ;
        RECT 40.195 52.905 41.360 53.495 ;
        RECT 47.540 53.325 47.790 54.135 ;
        RECT 47.970 53.790 48.230 54.315 ;
        RECT 48.400 53.325 48.650 54.135 ;
        RECT 48.830 53.805 49.135 54.315 ;
        RECT 41.530 53.075 48.650 53.325 ;
        RECT 48.820 53.075 49.135 53.635 ;
        RECT 49.305 53.545 50.975 54.315 ;
        RECT 40.195 52.680 46.940 52.905 ;
        RECT 40.195 51.765 40.465 52.510 ;
        RECT 40.635 51.940 40.925 52.680 ;
        RECT 41.535 52.665 46.940 52.680 ;
        RECT 41.095 51.770 41.350 52.495 ;
        RECT 41.535 51.940 41.795 52.665 ;
        RECT 41.965 51.770 42.210 52.495 ;
        RECT 42.395 51.940 42.655 52.665 ;
        RECT 42.825 51.770 43.070 52.495 ;
        RECT 43.255 51.940 43.515 52.665 ;
        RECT 43.685 51.770 43.930 52.495 ;
        RECT 44.100 51.940 44.360 52.665 ;
        RECT 44.530 51.770 44.790 52.495 ;
        RECT 44.960 51.940 45.220 52.665 ;
        RECT 45.390 51.770 45.650 52.495 ;
        RECT 45.820 51.940 46.080 52.665 ;
        RECT 46.250 51.770 46.510 52.495 ;
        RECT 46.680 51.940 46.940 52.665 ;
        RECT 47.110 51.770 47.370 52.565 ;
        RECT 47.540 51.940 47.790 53.075 ;
        RECT 41.095 51.765 47.370 51.770 ;
        RECT 47.970 51.765 48.230 52.575 ;
        RECT 48.405 51.935 48.650 53.075 ;
        RECT 49.305 53.025 50.055 53.545 ;
        RECT 51.810 53.535 52.310 54.145 ;
        RECT 50.225 52.855 50.975 53.375 ;
        RECT 51.605 53.075 51.955 53.325 ;
        RECT 52.140 52.905 52.310 53.535 ;
        RECT 52.940 53.665 53.270 54.145 ;
        RECT 53.440 53.855 53.665 54.315 ;
        RECT 53.835 53.665 54.165 54.145 ;
        RECT 52.940 53.495 54.165 53.665 ;
        RECT 54.355 53.515 54.605 54.315 ;
        RECT 54.775 53.515 55.115 54.145 ;
        RECT 52.480 53.125 52.810 53.325 ;
        RECT 52.980 53.125 53.310 53.325 ;
        RECT 53.480 53.125 53.900 53.325 ;
        RECT 54.075 53.155 54.770 53.325 ;
        RECT 54.075 52.905 54.245 53.155 ;
        RECT 54.940 52.905 55.115 53.515 ;
        RECT 55.285 53.545 56.955 54.315 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 55.285 53.025 56.035 53.545 ;
        RECT 58.510 53.475 58.770 54.315 ;
        RECT 58.945 53.570 59.200 54.145 ;
        RECT 59.370 53.935 59.700 54.315 ;
        RECT 59.915 53.765 60.085 54.145 ;
        RECT 59.370 53.595 60.085 53.765 ;
        RECT 48.830 51.765 49.125 52.575 ;
        RECT 49.305 51.765 50.975 52.855 ;
        RECT 51.810 52.735 54.245 52.905 ;
        RECT 51.810 51.935 52.140 52.735 ;
        RECT 52.310 51.765 52.640 52.565 ;
        RECT 52.940 51.935 53.270 52.735 ;
        RECT 53.915 51.765 54.165 52.565 ;
        RECT 54.435 51.765 54.605 52.905 ;
        RECT 54.775 51.935 55.115 52.905 ;
        RECT 56.205 52.855 56.955 53.375 ;
        RECT 55.285 51.765 56.955 52.855 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 58.510 51.765 58.770 52.915 ;
        RECT 58.945 52.840 59.115 53.570 ;
        RECT 59.370 53.405 59.540 53.595 ;
        RECT 60.350 53.475 60.610 54.315 ;
        RECT 60.785 53.570 61.040 54.145 ;
        RECT 61.210 53.935 61.540 54.315 ;
        RECT 61.755 53.765 61.925 54.145 ;
        RECT 61.210 53.595 61.925 53.765 ;
        RECT 62.185 53.815 62.445 54.145 ;
        RECT 62.755 53.935 63.085 54.315 ;
        RECT 63.265 53.975 64.745 54.145 ;
        RECT 59.285 53.075 59.540 53.405 ;
        RECT 59.370 52.865 59.540 53.075 ;
        RECT 59.820 53.045 60.175 53.415 ;
        RECT 58.945 51.935 59.200 52.840 ;
        RECT 59.370 52.695 60.085 52.865 ;
        RECT 59.370 51.765 59.700 52.525 ;
        RECT 59.915 51.935 60.085 52.695 ;
        RECT 60.350 51.765 60.610 52.915 ;
        RECT 60.785 52.840 60.955 53.570 ;
        RECT 61.210 53.405 61.380 53.595 ;
        RECT 61.125 53.075 61.380 53.405 ;
        RECT 61.210 52.865 61.380 53.075 ;
        RECT 61.660 53.045 62.015 53.415 ;
        RECT 62.185 53.115 62.355 53.815 ;
        RECT 63.265 53.645 63.665 53.975 ;
        RECT 62.705 53.455 62.915 53.635 ;
        RECT 62.705 53.285 63.325 53.455 ;
        RECT 63.495 53.165 63.665 53.645 ;
        RECT 63.855 53.475 64.405 53.805 ;
        RECT 62.185 52.945 63.315 53.115 ;
        RECT 63.495 52.995 64.065 53.165 ;
        RECT 60.785 51.935 61.040 52.840 ;
        RECT 61.210 52.695 61.925 52.865 ;
        RECT 61.210 51.765 61.540 52.525 ;
        RECT 61.755 51.935 61.925 52.695 ;
        RECT 62.185 52.265 62.355 52.945 ;
        RECT 63.145 52.825 63.315 52.945 ;
        RECT 62.525 52.445 62.875 52.775 ;
        RECT 63.145 52.655 63.725 52.825 ;
        RECT 63.895 52.485 64.065 52.995 ;
        RECT 63.325 52.315 64.065 52.485 ;
        RECT 64.235 52.485 64.405 53.475 ;
        RECT 64.575 53.075 64.745 53.975 ;
        RECT 64.995 53.405 65.180 53.985 ;
        RECT 65.450 53.405 65.645 53.980 ;
        RECT 65.855 53.935 66.185 54.315 ;
        RECT 64.995 53.075 65.225 53.405 ;
        RECT 65.450 53.075 65.705 53.405 ;
        RECT 64.995 52.765 65.180 53.075 ;
        RECT 65.450 52.765 65.645 53.075 ;
        RECT 66.015 52.485 66.185 53.405 ;
        RECT 64.235 52.315 66.185 52.485 ;
        RECT 62.185 51.935 62.445 52.265 ;
        RECT 62.755 51.765 63.085 52.145 ;
        RECT 63.325 51.935 63.515 52.315 ;
        RECT 63.765 51.765 64.095 52.145 ;
        RECT 64.305 51.935 64.475 52.315 ;
        RECT 64.670 51.765 65.000 52.145 ;
        RECT 65.260 51.935 65.430 52.315 ;
        RECT 65.855 51.765 66.185 52.145 ;
        RECT 66.355 51.935 66.615 54.145 ;
        RECT 67.090 53.745 67.260 53.995 ;
        RECT 66.785 53.575 67.260 53.745 ;
        RECT 67.495 53.575 67.825 54.315 ;
        RECT 67.995 53.745 68.195 54.090 ;
        RECT 68.365 53.915 68.695 54.315 ;
        RECT 68.865 53.745 69.065 54.100 ;
        RECT 69.235 53.920 69.565 54.315 ;
        RECT 70.095 53.765 70.265 54.145 ;
        RECT 70.480 53.935 70.810 54.315 ;
        RECT 67.995 53.575 69.835 53.745 ;
        RECT 70.095 53.595 70.810 53.765 ;
        RECT 66.785 52.605 66.955 53.575 ;
        RECT 67.125 52.785 67.475 53.405 ;
        RECT 67.645 52.785 67.965 53.405 ;
        RECT 68.135 52.785 68.465 53.405 ;
        RECT 68.635 52.785 68.935 53.405 ;
        RECT 69.175 52.605 69.395 53.405 ;
        RECT 66.785 52.395 69.395 52.605 ;
        RECT 67.495 51.765 67.825 52.215 ;
        RECT 69.575 51.950 69.835 53.575 ;
        RECT 70.005 53.045 70.360 53.415 ;
        RECT 70.640 53.405 70.810 53.595 ;
        RECT 70.980 53.570 71.235 54.145 ;
        RECT 70.640 53.075 70.895 53.405 ;
        RECT 70.640 52.865 70.810 53.075 ;
        RECT 70.095 52.695 70.810 52.865 ;
        RECT 71.065 52.840 71.235 53.570 ;
        RECT 71.410 53.475 71.670 54.315 ;
        RECT 71.845 53.770 77.190 54.315 ;
        RECT 77.365 53.770 82.710 54.315 ;
        RECT 73.430 52.940 73.770 53.770 ;
        RECT 70.095 51.935 70.265 52.695 ;
        RECT 70.480 51.765 70.810 52.525 ;
        RECT 70.980 51.935 71.235 52.840 ;
        RECT 71.410 51.765 71.670 52.915 ;
        RECT 75.250 52.200 75.600 53.450 ;
        RECT 78.950 52.940 79.290 53.770 ;
        RECT 82.885 53.590 83.175 54.315 ;
        RECT 83.345 53.565 84.555 54.315 ;
        RECT 80.770 52.200 81.120 53.450 ;
        RECT 83.345 53.025 83.865 53.565 ;
        RECT 84.930 53.535 85.430 54.145 ;
        RECT 71.845 51.765 77.190 52.200 ;
        RECT 77.365 51.765 82.710 52.200 ;
        RECT 82.885 51.765 83.175 52.930 ;
        RECT 84.035 52.855 84.555 53.395 ;
        RECT 84.725 53.075 85.075 53.325 ;
        RECT 85.260 52.905 85.430 53.535 ;
        RECT 86.060 53.665 86.390 54.145 ;
        RECT 86.560 53.855 86.785 54.315 ;
        RECT 86.955 53.665 87.285 54.145 ;
        RECT 86.060 53.495 87.285 53.665 ;
        RECT 87.475 53.515 87.725 54.315 ;
        RECT 87.895 53.515 88.235 54.145 ;
        RECT 85.600 53.125 85.930 53.325 ;
        RECT 86.100 53.125 86.430 53.325 ;
        RECT 86.600 53.125 87.020 53.325 ;
        RECT 87.195 53.155 87.890 53.325 ;
        RECT 87.195 52.905 87.365 53.155 ;
        RECT 88.060 52.905 88.235 53.515 ;
        RECT 83.345 51.765 84.555 52.855 ;
        RECT 84.930 52.735 87.365 52.905 ;
        RECT 84.930 51.935 85.260 52.735 ;
        RECT 85.430 51.765 85.760 52.565 ;
        RECT 86.060 51.935 86.390 52.735 ;
        RECT 87.035 51.765 87.285 52.565 ;
        RECT 87.555 51.765 87.725 52.905 ;
        RECT 87.895 51.935 88.235 52.905 ;
        RECT 88.405 53.515 88.745 54.145 ;
        RECT 88.915 53.515 89.165 54.315 ;
        RECT 89.355 53.665 89.685 54.145 ;
        RECT 89.855 53.855 90.080 54.315 ;
        RECT 90.250 53.665 90.580 54.145 ;
        RECT 88.405 52.905 88.580 53.515 ;
        RECT 89.355 53.495 90.580 53.665 ;
        RECT 91.210 53.535 91.710 54.145 ;
        RECT 92.290 53.535 92.790 54.145 ;
        RECT 88.750 53.155 89.445 53.325 ;
        RECT 89.275 52.905 89.445 53.155 ;
        RECT 89.620 53.125 90.040 53.325 ;
        RECT 90.210 53.125 90.540 53.325 ;
        RECT 90.710 53.125 91.040 53.325 ;
        RECT 91.210 52.905 91.380 53.535 ;
        RECT 91.565 53.075 91.915 53.325 ;
        RECT 92.085 53.075 92.435 53.325 ;
        RECT 92.620 52.905 92.790 53.535 ;
        RECT 93.420 53.665 93.750 54.145 ;
        RECT 93.920 53.855 94.145 54.315 ;
        RECT 94.315 53.665 94.645 54.145 ;
        RECT 93.420 53.495 94.645 53.665 ;
        RECT 94.835 53.515 95.085 54.315 ;
        RECT 95.255 53.515 95.595 54.145 ;
        RECT 95.880 53.685 96.165 54.145 ;
        RECT 96.335 53.855 96.605 54.315 ;
        RECT 95.880 53.515 96.835 53.685 ;
        RECT 92.960 53.125 93.290 53.325 ;
        RECT 93.460 53.125 93.790 53.325 ;
        RECT 93.960 53.125 94.380 53.325 ;
        RECT 94.555 53.155 95.250 53.325 ;
        RECT 94.555 52.905 94.725 53.155 ;
        RECT 95.420 52.905 95.595 53.515 ;
        RECT 88.405 51.935 88.745 52.905 ;
        RECT 88.915 51.765 89.085 52.905 ;
        RECT 89.275 52.735 91.710 52.905 ;
        RECT 89.355 51.765 89.605 52.565 ;
        RECT 90.250 51.935 90.580 52.735 ;
        RECT 90.880 51.765 91.210 52.565 ;
        RECT 91.380 51.935 91.710 52.735 ;
        RECT 92.290 52.735 94.725 52.905 ;
        RECT 92.290 51.935 92.620 52.735 ;
        RECT 92.790 51.765 93.120 52.565 ;
        RECT 93.420 51.935 93.750 52.735 ;
        RECT 94.395 51.765 94.645 52.565 ;
        RECT 94.915 51.765 95.085 52.905 ;
        RECT 95.255 51.935 95.595 52.905 ;
        RECT 95.765 52.785 96.455 53.345 ;
        RECT 96.625 52.615 96.835 53.515 ;
        RECT 95.880 52.395 96.835 52.615 ;
        RECT 97.005 53.345 97.405 54.145 ;
        RECT 97.595 53.685 97.875 54.145 ;
        RECT 98.395 53.855 98.720 54.315 ;
        RECT 97.595 53.515 98.720 53.685 ;
        RECT 98.890 53.575 99.275 54.145 ;
        RECT 99.450 53.765 99.705 54.055 ;
        RECT 99.875 53.935 100.205 54.315 ;
        RECT 99.450 53.595 100.200 53.765 ;
        RECT 98.270 53.405 98.720 53.515 ;
        RECT 97.005 52.785 98.100 53.345 ;
        RECT 98.270 53.075 98.825 53.405 ;
        RECT 95.880 51.935 96.165 52.395 ;
        RECT 96.335 51.765 96.605 52.225 ;
        RECT 97.005 51.935 97.405 52.785 ;
        RECT 98.270 52.615 98.720 53.075 ;
        RECT 98.995 52.905 99.275 53.575 ;
        RECT 97.595 52.395 98.720 52.615 ;
        RECT 97.595 51.935 97.875 52.395 ;
        RECT 98.395 51.765 98.720 52.225 ;
        RECT 98.890 51.935 99.275 52.905 ;
        RECT 99.450 52.775 99.800 53.425 ;
        RECT 99.970 52.605 100.200 53.595 ;
        RECT 99.450 52.435 100.200 52.605 ;
        RECT 99.450 51.935 99.705 52.435 ;
        RECT 99.875 51.765 100.205 52.265 ;
        RECT 100.375 51.935 100.545 54.055 ;
        RECT 100.905 53.955 101.235 54.315 ;
        RECT 101.405 53.925 101.900 54.095 ;
        RECT 102.105 53.925 102.960 54.095 ;
        RECT 100.775 52.735 101.235 53.785 ;
        RECT 100.715 51.950 101.040 52.735 ;
        RECT 101.405 52.565 101.575 53.925 ;
        RECT 101.745 53.015 102.095 53.635 ;
        RECT 102.265 53.415 102.620 53.635 ;
        RECT 102.265 52.825 102.435 53.415 ;
        RECT 102.790 53.215 102.960 53.925 ;
        RECT 103.835 53.855 104.165 54.315 ;
        RECT 104.375 53.955 104.725 54.125 ;
        RECT 103.165 53.385 103.955 53.635 ;
        RECT 104.375 53.565 104.635 53.955 ;
        RECT 104.945 53.865 105.895 54.145 ;
        RECT 106.065 53.875 106.255 54.315 ;
        RECT 106.425 53.935 107.495 54.105 ;
        RECT 104.125 53.215 104.295 53.395 ;
        RECT 101.405 52.395 101.800 52.565 ;
        RECT 101.970 52.435 102.435 52.825 ;
        RECT 102.605 53.045 104.295 53.215 ;
        RECT 101.630 52.265 101.800 52.395 ;
        RECT 102.605 52.265 102.775 53.045 ;
        RECT 104.465 52.875 104.635 53.565 ;
        RECT 103.135 52.705 104.635 52.875 ;
        RECT 104.825 52.905 105.035 53.695 ;
        RECT 105.205 53.075 105.555 53.695 ;
        RECT 105.725 53.085 105.895 53.865 ;
        RECT 106.425 53.705 106.595 53.935 ;
        RECT 106.065 53.535 106.595 53.705 ;
        RECT 106.065 53.255 106.285 53.535 ;
        RECT 106.765 53.365 107.005 53.765 ;
        RECT 105.725 52.915 106.130 53.085 ;
        RECT 106.465 52.995 107.005 53.365 ;
        RECT 107.175 53.580 107.495 53.935 ;
        RECT 107.740 53.855 108.045 54.315 ;
        RECT 108.215 53.605 108.470 54.135 ;
        RECT 107.175 53.405 107.500 53.580 ;
        RECT 107.175 53.105 108.090 53.405 ;
        RECT 107.350 53.075 108.090 53.105 ;
        RECT 104.825 52.745 105.500 52.905 ;
        RECT 105.960 52.825 106.130 52.915 ;
        RECT 104.825 52.735 105.790 52.745 ;
        RECT 104.465 52.565 104.635 52.705 ;
        RECT 101.210 51.765 101.460 52.225 ;
        RECT 101.630 51.935 101.880 52.265 ;
        RECT 102.095 51.935 102.775 52.265 ;
        RECT 102.945 52.365 104.020 52.535 ;
        RECT 104.465 52.395 105.025 52.565 ;
        RECT 105.330 52.445 105.790 52.735 ;
        RECT 105.960 52.655 107.180 52.825 ;
        RECT 102.945 52.025 103.115 52.365 ;
        RECT 103.350 51.765 103.680 52.195 ;
        RECT 103.850 52.025 104.020 52.365 ;
        RECT 104.315 51.765 104.685 52.225 ;
        RECT 104.855 51.935 105.025 52.395 ;
        RECT 105.960 52.275 106.130 52.655 ;
        RECT 107.350 52.485 107.520 53.075 ;
        RECT 108.260 52.955 108.470 53.605 ;
        RECT 108.645 53.590 108.935 54.315 ;
        RECT 105.260 51.935 106.130 52.275 ;
        RECT 106.720 52.315 107.520 52.485 ;
        RECT 106.300 51.765 106.550 52.225 ;
        RECT 106.720 52.025 106.890 52.315 ;
        RECT 107.070 51.765 107.400 52.145 ;
        RECT 107.740 51.765 108.045 52.905 ;
        RECT 108.215 52.075 108.470 52.955 ;
        RECT 109.105 53.575 109.490 54.145 ;
        RECT 109.660 53.855 109.985 54.315 ;
        RECT 110.505 53.685 110.785 54.145 ;
        RECT 108.645 51.765 108.935 52.930 ;
        RECT 109.105 52.905 109.385 53.575 ;
        RECT 109.660 53.515 110.785 53.685 ;
        RECT 109.660 53.405 110.110 53.515 ;
        RECT 109.555 53.075 110.110 53.405 ;
        RECT 110.975 53.345 111.375 54.145 ;
        RECT 111.775 53.855 112.045 54.315 ;
        RECT 112.215 53.685 112.500 54.145 ;
        RECT 109.105 51.935 109.490 52.905 ;
        RECT 109.660 52.615 110.110 53.075 ;
        RECT 110.280 52.785 111.375 53.345 ;
        RECT 109.660 52.395 110.785 52.615 ;
        RECT 109.660 51.765 109.985 52.225 ;
        RECT 110.505 51.935 110.785 52.395 ;
        RECT 110.975 51.935 111.375 52.785 ;
        RECT 111.545 53.515 112.500 53.685 ;
        RECT 112.785 53.515 113.125 54.145 ;
        RECT 113.295 53.515 113.545 54.315 ;
        RECT 113.735 53.665 114.065 54.145 ;
        RECT 114.235 53.855 114.460 54.315 ;
        RECT 114.630 53.665 114.960 54.145 ;
        RECT 111.545 52.615 111.755 53.515 ;
        RECT 111.925 52.785 112.615 53.345 ;
        RECT 112.785 52.905 112.960 53.515 ;
        RECT 113.735 53.495 114.960 53.665 ;
        RECT 115.590 53.535 116.090 54.145 ;
        RECT 116.465 53.770 121.810 54.315 ;
        RECT 113.130 53.155 113.825 53.325 ;
        RECT 113.655 52.905 113.825 53.155 ;
        RECT 114.000 53.125 114.420 53.325 ;
        RECT 114.590 53.125 114.920 53.325 ;
        RECT 115.090 53.125 115.420 53.325 ;
        RECT 115.590 52.905 115.760 53.535 ;
        RECT 115.945 53.075 116.295 53.325 ;
        RECT 118.050 52.940 118.390 53.770 ;
        RECT 121.985 53.545 123.655 54.315 ;
        RECT 124.285 53.565 125.495 54.315 ;
        RECT 111.545 52.395 112.500 52.615 ;
        RECT 111.775 51.765 112.045 52.225 ;
        RECT 112.215 51.935 112.500 52.395 ;
        RECT 112.785 51.935 113.125 52.905 ;
        RECT 113.295 51.765 113.465 52.905 ;
        RECT 113.655 52.735 116.090 52.905 ;
        RECT 113.735 51.765 113.985 52.565 ;
        RECT 114.630 51.935 114.960 52.735 ;
        RECT 115.260 51.765 115.590 52.565 ;
        RECT 115.760 51.935 116.090 52.735 ;
        RECT 119.870 52.200 120.220 53.450 ;
        RECT 121.985 53.025 122.735 53.545 ;
        RECT 122.905 52.855 123.655 53.375 ;
        RECT 116.465 51.765 121.810 52.200 ;
        RECT 121.985 51.765 123.655 52.855 ;
        RECT 124.285 52.855 124.805 53.395 ;
        RECT 124.975 53.025 125.495 53.565 ;
        RECT 124.285 51.765 125.495 52.855 ;
        RECT 5.520 51.595 125.580 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 6.985 51.160 12.330 51.595 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 8.570 49.590 8.910 50.420 ;
        RECT 10.390 49.910 10.740 51.160 ;
        RECT 12.965 50.520 13.235 51.425 ;
        RECT 13.405 50.835 13.735 51.595 ;
        RECT 13.915 50.665 14.085 51.425 ;
        RECT 12.965 49.720 13.135 50.520 ;
        RECT 13.420 50.495 14.085 50.665 ;
        RECT 14.345 50.520 14.615 51.425 ;
        RECT 14.785 50.835 15.115 51.595 ;
        RECT 15.295 50.665 15.465 51.425 ;
        RECT 13.420 50.350 13.590 50.495 ;
        RECT 13.305 50.020 13.590 50.350 ;
        RECT 13.420 49.765 13.590 50.020 ;
        RECT 13.825 49.945 14.155 50.315 ;
        RECT 6.985 49.045 12.330 49.590 ;
        RECT 12.965 49.215 13.225 49.720 ;
        RECT 13.420 49.595 14.085 49.765 ;
        RECT 13.405 49.045 13.735 49.425 ;
        RECT 13.915 49.215 14.085 49.595 ;
        RECT 14.345 49.720 14.515 50.520 ;
        RECT 14.800 50.495 15.465 50.665 ;
        RECT 15.725 50.505 18.315 51.595 ;
        RECT 14.800 50.350 14.970 50.495 ;
        RECT 14.685 50.020 14.970 50.350 ;
        RECT 14.800 49.765 14.970 50.020 ;
        RECT 15.205 49.945 15.535 50.315 ;
        RECT 15.725 49.815 16.935 50.335 ;
        RECT 17.105 49.985 18.315 50.505 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 18.945 50.505 21.535 51.595 ;
        RECT 22.280 50.965 22.565 51.425 ;
        RECT 22.735 51.135 23.005 51.595 ;
        RECT 22.280 50.745 23.235 50.965 ;
        RECT 18.945 49.815 20.155 50.335 ;
        RECT 20.325 49.985 21.535 50.505 ;
        RECT 22.165 50.015 22.855 50.575 ;
        RECT 23.025 49.845 23.235 50.745 ;
        RECT 14.345 49.215 14.605 49.720 ;
        RECT 14.800 49.595 15.465 49.765 ;
        RECT 14.785 49.045 15.115 49.425 ;
        RECT 15.295 49.215 15.465 49.595 ;
        RECT 15.725 49.045 18.315 49.815 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 18.945 49.045 21.535 49.815 ;
        RECT 22.280 49.675 23.235 49.845 ;
        RECT 23.405 50.575 23.805 51.425 ;
        RECT 23.995 50.965 24.275 51.425 ;
        RECT 24.795 51.135 25.120 51.595 ;
        RECT 23.995 50.745 25.120 50.965 ;
        RECT 23.405 50.015 24.500 50.575 ;
        RECT 24.670 50.285 25.120 50.745 ;
        RECT 25.290 50.455 25.675 51.425 ;
        RECT 26.050 50.625 26.380 51.425 ;
        RECT 26.550 50.795 26.880 51.595 ;
        RECT 27.180 50.625 27.510 51.425 ;
        RECT 28.155 50.795 28.405 51.595 ;
        RECT 26.050 50.455 28.485 50.625 ;
        RECT 28.675 50.455 28.845 51.595 ;
        RECT 29.015 50.455 29.355 51.425 ;
        RECT 22.280 49.215 22.565 49.675 ;
        RECT 22.735 49.045 23.005 49.505 ;
        RECT 23.405 49.215 23.805 50.015 ;
        RECT 24.670 49.955 25.225 50.285 ;
        RECT 24.670 49.845 25.120 49.955 ;
        RECT 23.995 49.675 25.120 49.845 ;
        RECT 25.395 49.785 25.675 50.455 ;
        RECT 25.845 50.035 26.195 50.285 ;
        RECT 26.380 49.825 26.550 50.455 ;
        RECT 26.720 50.035 27.050 50.235 ;
        RECT 27.220 50.035 27.550 50.235 ;
        RECT 27.720 50.035 28.140 50.235 ;
        RECT 28.315 50.205 28.485 50.455 ;
        RECT 28.315 50.035 29.010 50.205 ;
        RECT 23.995 49.215 24.275 49.675 ;
        RECT 24.795 49.045 25.120 49.505 ;
        RECT 25.290 49.215 25.675 49.785 ;
        RECT 26.050 49.215 26.550 49.825 ;
        RECT 27.180 49.695 28.405 49.865 ;
        RECT 29.180 49.845 29.355 50.455 ;
        RECT 27.180 49.215 27.510 49.695 ;
        RECT 27.680 49.045 27.905 49.505 ;
        RECT 28.075 49.215 28.405 49.695 ;
        RECT 28.595 49.045 28.845 49.845 ;
        RECT 29.015 49.215 29.355 49.845 ;
        RECT 29.525 50.455 29.910 51.425 ;
        RECT 30.080 51.135 30.405 51.595 ;
        RECT 30.925 50.965 31.205 51.425 ;
        RECT 30.080 50.745 31.205 50.965 ;
        RECT 29.525 49.785 29.805 50.455 ;
        RECT 30.080 50.285 30.530 50.745 ;
        RECT 31.395 50.575 31.795 51.425 ;
        RECT 32.195 51.135 32.465 51.595 ;
        RECT 32.635 50.965 32.920 51.425 ;
        RECT 29.975 49.955 30.530 50.285 ;
        RECT 30.700 50.015 31.795 50.575 ;
        RECT 30.080 49.845 30.530 49.955 ;
        RECT 29.525 49.215 29.910 49.785 ;
        RECT 30.080 49.675 31.205 49.845 ;
        RECT 30.080 49.045 30.405 49.505 ;
        RECT 30.925 49.215 31.205 49.675 ;
        RECT 31.395 49.215 31.795 50.015 ;
        RECT 31.965 50.745 32.920 50.965 ;
        RECT 31.965 49.845 32.175 50.745 ;
        RECT 32.345 50.015 33.035 50.575 ;
        RECT 33.205 50.505 34.415 51.595 ;
        RECT 31.965 49.675 32.920 49.845 ;
        RECT 32.195 49.045 32.465 49.505 ;
        RECT 32.635 49.215 32.920 49.675 ;
        RECT 33.205 49.795 33.725 50.335 ;
        RECT 33.895 49.965 34.415 50.505 ;
        RECT 34.585 50.835 35.100 51.245 ;
        RECT 35.335 50.835 35.505 51.595 ;
        RECT 35.675 51.255 37.705 51.425 ;
        RECT 34.585 50.025 34.925 50.835 ;
        RECT 35.675 50.590 35.845 51.255 ;
        RECT 36.240 50.915 37.365 51.085 ;
        RECT 35.095 50.400 35.845 50.590 ;
        RECT 36.015 50.575 37.025 50.745 ;
        RECT 34.585 49.855 35.815 50.025 ;
        RECT 33.205 49.045 34.415 49.795 ;
        RECT 34.860 49.250 35.105 49.855 ;
        RECT 35.325 49.045 35.835 49.580 ;
        RECT 36.015 49.215 36.205 50.575 ;
        RECT 36.375 49.555 36.650 50.375 ;
        RECT 36.855 49.775 37.025 50.575 ;
        RECT 37.195 49.785 37.365 50.915 ;
        RECT 37.535 50.285 37.705 51.255 ;
        RECT 37.875 50.455 38.045 51.595 ;
        RECT 38.215 50.455 38.550 51.425 ;
        RECT 37.535 49.955 37.730 50.285 ;
        RECT 37.955 49.955 38.210 50.285 ;
        RECT 37.955 49.785 38.125 49.955 ;
        RECT 38.380 49.785 38.550 50.455 ;
        RECT 37.195 49.615 38.125 49.785 ;
        RECT 37.195 49.580 37.370 49.615 ;
        RECT 36.375 49.385 36.655 49.555 ;
        RECT 36.375 49.215 36.650 49.385 ;
        RECT 36.840 49.215 37.370 49.580 ;
        RECT 37.795 49.045 38.125 49.445 ;
        RECT 38.295 49.215 38.550 49.785 ;
        RECT 38.725 50.455 39.110 51.425 ;
        RECT 39.280 51.135 39.605 51.595 ;
        RECT 40.125 50.965 40.405 51.425 ;
        RECT 39.280 50.745 40.405 50.965 ;
        RECT 38.725 49.785 39.005 50.455 ;
        RECT 39.280 50.285 39.730 50.745 ;
        RECT 40.595 50.575 40.995 51.425 ;
        RECT 41.395 51.135 41.665 51.595 ;
        RECT 41.835 50.965 42.120 51.425 ;
        RECT 39.175 49.955 39.730 50.285 ;
        RECT 39.900 50.015 40.995 50.575 ;
        RECT 39.280 49.845 39.730 49.955 ;
        RECT 38.725 49.215 39.110 49.785 ;
        RECT 39.280 49.675 40.405 49.845 ;
        RECT 39.280 49.045 39.605 49.505 ;
        RECT 40.125 49.215 40.405 49.675 ;
        RECT 40.595 49.215 40.995 50.015 ;
        RECT 41.165 50.745 42.120 50.965 ;
        RECT 41.165 49.845 41.375 50.745 ;
        RECT 42.955 50.665 43.125 51.425 ;
        RECT 43.305 50.835 43.635 51.595 ;
        RECT 41.545 50.015 42.235 50.575 ;
        RECT 42.955 50.495 43.620 50.665 ;
        RECT 43.805 50.520 44.075 51.425 ;
        RECT 43.450 50.350 43.620 50.495 ;
        RECT 42.885 49.945 43.215 50.315 ;
        RECT 43.450 50.020 43.735 50.350 ;
        RECT 41.165 49.675 42.120 49.845 ;
        RECT 43.450 49.765 43.620 50.020 ;
        RECT 41.395 49.045 41.665 49.505 ;
        RECT 41.835 49.215 42.120 49.675 ;
        RECT 42.955 49.595 43.620 49.765 ;
        RECT 43.905 49.720 44.075 50.520 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 45.625 50.455 46.010 51.425 ;
        RECT 46.180 51.135 46.505 51.595 ;
        RECT 47.025 50.965 47.305 51.425 ;
        RECT 46.180 50.745 47.305 50.965 ;
        RECT 45.625 49.785 45.905 50.455 ;
        RECT 46.180 50.285 46.630 50.745 ;
        RECT 47.495 50.575 47.895 51.425 ;
        RECT 48.295 51.135 48.565 51.595 ;
        RECT 48.735 50.965 49.020 51.425 ;
        RECT 46.075 49.955 46.630 50.285 ;
        RECT 46.800 50.015 47.895 50.575 ;
        RECT 46.180 49.845 46.630 49.955 ;
        RECT 42.955 49.215 43.125 49.595 ;
        RECT 43.305 49.045 43.635 49.425 ;
        RECT 43.815 49.215 44.075 49.720 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 45.625 49.215 46.010 49.785 ;
        RECT 46.180 49.675 47.305 49.845 ;
        RECT 46.180 49.045 46.505 49.505 ;
        RECT 47.025 49.215 47.305 49.675 ;
        RECT 47.495 49.215 47.895 50.015 ;
        RECT 48.065 50.745 49.020 50.965 ;
        RECT 48.065 49.845 48.275 50.745 ;
        RECT 48.445 50.015 49.135 50.575 ;
        RECT 49.455 50.445 49.785 51.595 ;
        RECT 49.955 50.575 50.125 51.425 ;
        RECT 50.295 50.795 50.625 51.595 ;
        RECT 50.795 50.575 50.965 51.425 ;
        RECT 51.145 50.795 51.385 51.595 ;
        RECT 51.555 50.615 51.885 51.425 ;
        RECT 49.955 50.405 50.965 50.575 ;
        RECT 51.170 50.445 51.885 50.615 ;
        RECT 52.730 50.625 53.060 51.425 ;
        RECT 53.230 50.795 53.560 51.595 ;
        RECT 53.860 50.625 54.190 51.425 ;
        RECT 54.835 50.795 55.085 51.595 ;
        RECT 52.730 50.455 55.165 50.625 ;
        RECT 55.355 50.455 55.525 51.595 ;
        RECT 55.695 50.455 56.035 51.425 ;
        RECT 49.955 49.895 50.450 50.405 ;
        RECT 51.170 50.205 51.340 50.445 ;
        RECT 50.840 50.035 51.340 50.205 ;
        RECT 51.510 50.035 51.890 50.275 ;
        RECT 52.525 50.035 52.875 50.285 ;
        RECT 49.955 49.865 50.455 49.895 ;
        RECT 51.170 49.865 51.340 50.035 ;
        RECT 48.065 49.675 49.020 49.845 ;
        RECT 48.295 49.045 48.565 49.505 ;
        RECT 48.735 49.215 49.020 49.675 ;
        RECT 49.455 49.045 49.785 49.845 ;
        RECT 49.955 49.695 50.965 49.865 ;
        RECT 51.170 49.695 51.805 49.865 ;
        RECT 53.060 49.825 53.230 50.455 ;
        RECT 53.400 50.035 53.730 50.235 ;
        RECT 53.900 50.035 54.230 50.235 ;
        RECT 54.400 50.035 54.820 50.235 ;
        RECT 54.995 50.205 55.165 50.455 ;
        RECT 54.995 50.035 55.690 50.205 ;
        RECT 49.955 49.215 50.125 49.695 ;
        RECT 50.295 49.045 50.625 49.525 ;
        RECT 50.795 49.215 50.965 49.695 ;
        RECT 51.215 49.045 51.455 49.525 ;
        RECT 51.635 49.215 51.805 49.695 ;
        RECT 52.730 49.215 53.230 49.825 ;
        RECT 53.860 49.695 55.085 49.865 ;
        RECT 55.860 49.845 56.035 50.455 ;
        RECT 53.860 49.215 54.190 49.695 ;
        RECT 54.360 49.045 54.585 49.505 ;
        RECT 54.755 49.215 55.085 49.695 ;
        RECT 55.275 49.045 55.525 49.845 ;
        RECT 55.695 49.215 56.035 49.845 ;
        RECT 56.205 50.455 56.545 51.425 ;
        RECT 56.715 50.455 56.885 51.595 ;
        RECT 57.155 50.795 57.405 51.595 ;
        RECT 58.050 50.625 58.380 51.425 ;
        RECT 58.680 50.795 59.010 51.595 ;
        RECT 59.180 50.625 59.510 51.425 ;
        RECT 57.075 50.455 59.510 50.625 ;
        RECT 59.885 50.505 61.555 51.595 ;
        RECT 62.435 51.145 62.765 51.595 ;
        RECT 56.205 49.845 56.380 50.455 ;
        RECT 57.075 50.205 57.245 50.455 ;
        RECT 56.550 50.035 57.245 50.205 ;
        RECT 57.420 50.035 57.840 50.235 ;
        RECT 58.010 50.035 58.340 50.235 ;
        RECT 58.510 50.035 58.840 50.235 ;
        RECT 56.205 49.215 56.545 49.845 ;
        RECT 56.715 49.045 56.965 49.845 ;
        RECT 57.155 49.695 58.380 49.865 ;
        RECT 57.155 49.215 57.485 49.695 ;
        RECT 57.655 49.045 57.880 49.505 ;
        RECT 58.050 49.215 58.380 49.695 ;
        RECT 59.010 49.825 59.180 50.455 ;
        RECT 59.365 50.035 59.715 50.285 ;
        RECT 59.010 49.215 59.510 49.825 ;
        RECT 59.885 49.815 60.635 50.335 ;
        RECT 60.805 49.985 61.555 50.505 ;
        RECT 61.725 50.755 64.335 50.965 ;
        RECT 59.885 49.045 61.555 49.815 ;
        RECT 61.725 49.785 61.895 50.755 ;
        RECT 62.065 49.955 62.415 50.575 ;
        RECT 62.585 49.955 62.905 50.575 ;
        RECT 63.075 49.955 63.405 50.575 ;
        RECT 63.575 49.955 63.875 50.575 ;
        RECT 64.115 49.955 64.335 50.755 ;
        RECT 64.515 49.785 64.775 51.410 ;
        RECT 65.655 51.145 65.985 51.595 ;
        RECT 61.725 49.615 62.200 49.785 ;
        RECT 62.030 49.365 62.200 49.615 ;
        RECT 62.435 49.045 62.765 49.785 ;
        RECT 62.935 49.615 64.775 49.785 ;
        RECT 64.945 50.755 67.555 50.965 ;
        RECT 64.945 49.785 65.115 50.755 ;
        RECT 65.285 49.955 65.635 50.575 ;
        RECT 65.805 49.955 66.125 50.575 ;
        RECT 66.295 49.955 66.625 50.575 ;
        RECT 66.795 49.955 67.095 50.575 ;
        RECT 67.335 49.955 67.555 50.755 ;
        RECT 67.735 49.785 67.995 51.410 ;
        RECT 68.225 50.455 68.435 51.595 ;
        RECT 68.605 50.445 68.935 51.425 ;
        RECT 69.105 50.455 69.335 51.595 ;
        RECT 64.945 49.615 65.420 49.785 ;
        RECT 62.935 49.270 63.135 49.615 ;
        RECT 63.305 49.045 63.635 49.445 ;
        RECT 63.805 49.260 64.005 49.615 ;
        RECT 64.175 49.045 64.505 49.440 ;
        RECT 65.250 49.365 65.420 49.615 ;
        RECT 65.655 49.045 65.985 49.785 ;
        RECT 66.155 49.615 67.995 49.785 ;
        RECT 66.155 49.270 66.355 49.615 ;
        RECT 66.525 49.045 66.855 49.445 ;
        RECT 67.025 49.260 67.225 49.615 ;
        RECT 67.395 49.045 67.725 49.440 ;
        RECT 68.225 49.045 68.435 49.865 ;
        RECT 68.605 49.845 68.855 50.445 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 70.465 50.505 73.975 51.595 ;
        RECT 69.025 50.035 69.355 50.285 ;
        RECT 68.605 49.215 68.935 49.845 ;
        RECT 69.105 49.045 69.335 49.865 ;
        RECT 70.465 49.815 72.115 50.335 ;
        RECT 72.285 49.985 73.975 50.505 ;
        RECT 74.145 50.625 74.455 51.425 ;
        RECT 74.625 50.795 74.935 51.595 ;
        RECT 75.105 50.965 75.365 51.425 ;
        RECT 75.535 51.135 75.790 51.595 ;
        RECT 75.965 50.965 76.225 51.425 ;
        RECT 75.105 50.795 76.225 50.965 ;
        RECT 74.145 50.455 75.175 50.625 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 70.465 49.045 73.975 49.815 ;
        RECT 74.145 49.545 74.315 50.455 ;
        RECT 74.485 49.715 74.835 50.285 ;
        RECT 75.005 50.205 75.175 50.455 ;
        RECT 75.965 50.545 76.225 50.795 ;
        RECT 76.395 50.725 76.680 51.595 ;
        RECT 77.110 50.625 77.440 51.425 ;
        RECT 77.610 50.795 77.940 51.595 ;
        RECT 78.240 50.625 78.570 51.425 ;
        RECT 79.215 50.795 79.465 51.595 ;
        RECT 75.965 50.375 76.720 50.545 ;
        RECT 77.110 50.455 79.545 50.625 ;
        RECT 79.735 50.455 79.905 51.595 ;
        RECT 80.075 50.455 80.415 51.425 ;
        RECT 75.005 50.035 76.145 50.205 ;
        RECT 76.315 49.865 76.720 50.375 ;
        RECT 76.905 50.035 77.255 50.285 ;
        RECT 75.070 49.695 76.720 49.865 ;
        RECT 77.440 49.825 77.610 50.455 ;
        RECT 77.780 50.035 78.110 50.235 ;
        RECT 78.280 50.035 78.610 50.235 ;
        RECT 78.780 50.065 79.205 50.235 ;
        RECT 79.375 50.205 79.545 50.455 ;
        RECT 78.780 50.035 79.200 50.065 ;
        RECT 79.375 50.035 80.070 50.205 ;
        RECT 74.145 49.215 74.445 49.545 ;
        RECT 74.615 49.045 74.890 49.525 ;
        RECT 75.070 49.305 75.365 49.695 ;
        RECT 75.535 49.045 75.790 49.525 ;
        RECT 75.965 49.305 76.225 49.695 ;
        RECT 76.395 49.045 76.675 49.525 ;
        RECT 77.110 49.215 77.610 49.825 ;
        RECT 78.240 49.695 79.465 49.865 ;
        RECT 80.240 49.845 80.415 50.455 ;
        RECT 78.240 49.215 78.570 49.695 ;
        RECT 78.740 49.045 78.965 49.505 ;
        RECT 79.135 49.215 79.465 49.695 ;
        RECT 79.655 49.045 79.905 49.845 ;
        RECT 80.075 49.215 80.415 49.845 ;
        RECT 80.585 50.455 80.970 51.425 ;
        RECT 81.140 51.135 81.465 51.595 ;
        RECT 81.985 50.965 82.265 51.425 ;
        RECT 81.140 50.745 82.265 50.965 ;
        RECT 80.585 49.785 80.865 50.455 ;
        RECT 81.140 50.285 81.590 50.745 ;
        RECT 82.455 50.575 82.855 51.425 ;
        RECT 83.255 51.135 83.525 51.595 ;
        RECT 83.695 50.965 83.980 51.425 ;
        RECT 81.035 49.955 81.590 50.285 ;
        RECT 81.760 50.015 82.855 50.575 ;
        RECT 81.140 49.845 81.590 49.955 ;
        RECT 80.585 49.215 80.970 49.785 ;
        RECT 81.140 49.675 82.265 49.845 ;
        RECT 81.140 49.045 81.465 49.505 ;
        RECT 81.985 49.215 82.265 49.675 ;
        RECT 82.455 49.215 82.855 50.015 ;
        RECT 83.025 50.745 83.980 50.965 ;
        RECT 83.025 49.845 83.235 50.745 ;
        RECT 85.275 50.665 85.445 51.425 ;
        RECT 85.625 50.835 85.955 51.595 ;
        RECT 83.405 50.015 84.095 50.575 ;
        RECT 85.275 50.495 85.940 50.665 ;
        RECT 86.125 50.520 86.395 51.425 ;
        RECT 86.570 50.925 86.825 51.425 ;
        RECT 86.995 51.095 87.325 51.595 ;
        RECT 86.570 50.755 87.320 50.925 ;
        RECT 85.770 50.350 85.940 50.495 ;
        RECT 85.205 49.945 85.535 50.315 ;
        RECT 85.770 50.020 86.055 50.350 ;
        RECT 83.025 49.675 83.980 49.845 ;
        RECT 85.770 49.765 85.940 50.020 ;
        RECT 83.255 49.045 83.525 49.505 ;
        RECT 83.695 49.215 83.980 49.675 ;
        RECT 85.275 49.595 85.940 49.765 ;
        RECT 86.225 49.720 86.395 50.520 ;
        RECT 86.570 49.935 86.920 50.585 ;
        RECT 87.090 49.765 87.320 50.755 ;
        RECT 85.275 49.215 85.445 49.595 ;
        RECT 85.625 49.045 85.955 49.425 ;
        RECT 86.135 49.215 86.395 49.720 ;
        RECT 86.570 49.595 87.320 49.765 ;
        RECT 86.570 49.305 86.825 49.595 ;
        RECT 86.995 49.045 87.325 49.425 ;
        RECT 87.495 49.305 87.665 51.425 ;
        RECT 87.835 50.625 88.160 51.410 ;
        RECT 88.330 51.135 88.580 51.595 ;
        RECT 88.750 51.095 89.000 51.425 ;
        RECT 89.215 51.095 89.895 51.425 ;
        RECT 88.750 50.965 88.920 51.095 ;
        RECT 88.525 50.795 88.920 50.965 ;
        RECT 87.895 49.575 88.355 50.625 ;
        RECT 88.525 49.435 88.695 50.795 ;
        RECT 89.090 50.535 89.555 50.925 ;
        RECT 88.865 49.725 89.215 50.345 ;
        RECT 89.385 49.945 89.555 50.535 ;
        RECT 89.725 50.315 89.895 51.095 ;
        RECT 90.065 50.995 90.235 51.335 ;
        RECT 90.470 51.165 90.800 51.595 ;
        RECT 90.970 50.995 91.140 51.335 ;
        RECT 91.435 51.135 91.805 51.595 ;
        RECT 90.065 50.825 91.140 50.995 ;
        RECT 91.975 50.965 92.145 51.425 ;
        RECT 92.380 51.085 93.250 51.425 ;
        RECT 93.420 51.135 93.670 51.595 ;
        RECT 91.585 50.795 92.145 50.965 ;
        RECT 91.585 50.655 91.755 50.795 ;
        RECT 90.255 50.485 91.755 50.655 ;
        RECT 92.450 50.625 92.910 50.915 ;
        RECT 89.725 50.145 91.415 50.315 ;
        RECT 89.385 49.725 89.740 49.945 ;
        RECT 89.910 49.435 90.080 50.145 ;
        RECT 90.285 49.725 91.075 49.975 ;
        RECT 91.245 49.965 91.415 50.145 ;
        RECT 91.585 49.795 91.755 50.485 ;
        RECT 88.025 49.045 88.355 49.405 ;
        RECT 88.525 49.265 89.020 49.435 ;
        RECT 89.225 49.265 90.080 49.435 ;
        RECT 90.955 49.045 91.285 49.505 ;
        RECT 91.495 49.405 91.755 49.795 ;
        RECT 91.945 50.615 92.910 50.625 ;
        RECT 93.080 50.705 93.250 51.085 ;
        RECT 93.840 51.045 94.010 51.335 ;
        RECT 94.190 51.215 94.520 51.595 ;
        RECT 93.840 50.875 94.640 51.045 ;
        RECT 91.945 50.455 92.620 50.615 ;
        RECT 93.080 50.535 94.300 50.705 ;
        RECT 91.945 49.665 92.155 50.455 ;
        RECT 93.080 50.445 93.250 50.535 ;
        RECT 92.325 49.665 92.675 50.285 ;
        RECT 92.845 50.275 93.250 50.445 ;
        RECT 92.845 49.495 93.015 50.275 ;
        RECT 93.185 49.825 93.405 50.105 ;
        RECT 93.585 49.995 94.125 50.365 ;
        RECT 94.470 50.285 94.640 50.875 ;
        RECT 94.860 50.455 95.165 51.595 ;
        RECT 95.335 50.405 95.590 51.285 ;
        RECT 95.765 50.430 96.055 51.595 ;
        RECT 96.285 50.455 96.495 51.595 ;
        RECT 96.665 50.445 96.995 51.425 ;
        RECT 97.165 50.455 97.395 51.595 ;
        RECT 98.070 50.455 98.405 51.425 ;
        RECT 98.575 50.455 98.745 51.595 ;
        RECT 98.915 51.255 100.945 51.425 ;
        RECT 94.470 50.255 95.210 50.285 ;
        RECT 93.185 49.655 93.715 49.825 ;
        RECT 91.495 49.235 91.845 49.405 ;
        RECT 92.065 49.215 93.015 49.495 ;
        RECT 93.185 49.045 93.375 49.485 ;
        RECT 93.545 49.425 93.715 49.655 ;
        RECT 93.885 49.595 94.125 49.995 ;
        RECT 94.295 49.955 95.210 50.255 ;
        RECT 94.295 49.780 94.620 49.955 ;
        RECT 94.295 49.425 94.615 49.780 ;
        RECT 95.380 49.755 95.590 50.405 ;
        RECT 93.545 49.255 94.615 49.425 ;
        RECT 94.860 49.045 95.165 49.505 ;
        RECT 95.335 49.225 95.590 49.755 ;
        RECT 95.765 49.045 96.055 49.770 ;
        RECT 96.285 49.045 96.495 49.865 ;
        RECT 96.665 49.845 96.915 50.445 ;
        RECT 97.085 50.035 97.415 50.285 ;
        RECT 96.665 49.215 96.995 49.845 ;
        RECT 97.165 49.045 97.395 49.865 ;
        RECT 98.070 49.785 98.240 50.455 ;
        RECT 98.915 50.285 99.085 51.255 ;
        RECT 98.410 49.955 98.665 50.285 ;
        RECT 98.890 49.955 99.085 50.285 ;
        RECT 99.255 50.915 100.380 51.085 ;
        RECT 98.495 49.785 98.665 49.955 ;
        RECT 99.255 49.785 99.425 50.915 ;
        RECT 98.070 49.215 98.325 49.785 ;
        RECT 98.495 49.615 99.425 49.785 ;
        RECT 99.595 50.575 100.605 50.745 ;
        RECT 99.595 49.775 99.765 50.575 ;
        RECT 99.250 49.580 99.425 49.615 ;
        RECT 98.495 49.045 98.825 49.445 ;
        RECT 99.250 49.215 99.780 49.580 ;
        RECT 99.970 49.555 100.245 50.375 ;
        RECT 99.965 49.385 100.245 49.555 ;
        RECT 99.970 49.215 100.245 49.385 ;
        RECT 100.415 49.215 100.605 50.575 ;
        RECT 100.775 50.590 100.945 51.255 ;
        RECT 101.115 50.835 101.285 51.595 ;
        RECT 101.520 50.835 102.035 51.245 ;
        RECT 100.775 50.400 101.525 50.590 ;
        RECT 101.695 50.025 102.035 50.835 ;
        RECT 100.805 49.855 102.035 50.025 ;
        RECT 102.205 50.520 102.475 51.425 ;
        RECT 102.645 50.835 102.975 51.595 ;
        RECT 103.155 50.665 103.325 51.425 ;
        RECT 100.785 49.045 101.295 49.580 ;
        RECT 101.515 49.250 101.760 49.855 ;
        RECT 102.205 49.720 102.375 50.520 ;
        RECT 102.660 50.495 103.325 50.665 ;
        RECT 103.585 50.835 104.100 51.245 ;
        RECT 104.335 50.835 104.505 51.595 ;
        RECT 104.675 51.255 106.705 51.425 ;
        RECT 102.660 50.350 102.830 50.495 ;
        RECT 102.545 50.020 102.830 50.350 ;
        RECT 102.660 49.765 102.830 50.020 ;
        RECT 103.065 49.945 103.395 50.315 ;
        RECT 103.585 50.025 103.925 50.835 ;
        RECT 104.675 50.590 104.845 51.255 ;
        RECT 105.240 50.915 106.365 51.085 ;
        RECT 104.095 50.400 104.845 50.590 ;
        RECT 105.015 50.575 106.025 50.745 ;
        RECT 103.585 49.855 104.815 50.025 ;
        RECT 102.205 49.215 102.465 49.720 ;
        RECT 102.660 49.595 103.325 49.765 ;
        RECT 102.645 49.045 102.975 49.425 ;
        RECT 103.155 49.215 103.325 49.595 ;
        RECT 103.860 49.250 104.105 49.855 ;
        RECT 104.325 49.045 104.835 49.580 ;
        RECT 105.015 49.215 105.205 50.575 ;
        RECT 105.375 50.235 105.650 50.375 ;
        RECT 105.375 50.065 105.655 50.235 ;
        RECT 105.375 49.215 105.650 50.065 ;
        RECT 105.855 49.775 106.025 50.575 ;
        RECT 106.195 49.785 106.365 50.915 ;
        RECT 106.535 50.285 106.705 51.255 ;
        RECT 106.875 50.455 107.045 51.595 ;
        RECT 107.215 50.455 107.550 51.425 ;
        RECT 107.730 50.925 107.985 51.425 ;
        RECT 108.155 51.095 108.485 51.595 ;
        RECT 107.730 50.755 108.480 50.925 ;
        RECT 106.535 49.955 106.730 50.285 ;
        RECT 106.955 49.955 107.210 50.285 ;
        RECT 106.955 49.785 107.125 49.955 ;
        RECT 107.380 49.785 107.550 50.455 ;
        RECT 107.730 49.935 108.080 50.585 ;
        RECT 106.195 49.615 107.125 49.785 ;
        RECT 106.195 49.580 106.370 49.615 ;
        RECT 105.840 49.215 106.370 49.580 ;
        RECT 106.795 49.045 107.125 49.445 ;
        RECT 107.295 49.215 107.550 49.785 ;
        RECT 108.250 49.765 108.480 50.755 ;
        RECT 107.730 49.595 108.480 49.765 ;
        RECT 107.730 49.305 107.985 49.595 ;
        RECT 108.155 49.045 108.485 49.425 ;
        RECT 108.655 49.305 108.825 51.425 ;
        RECT 108.995 50.625 109.320 51.410 ;
        RECT 109.490 51.135 109.740 51.595 ;
        RECT 109.910 51.095 110.160 51.425 ;
        RECT 110.375 51.095 111.055 51.425 ;
        RECT 109.910 50.965 110.080 51.095 ;
        RECT 109.685 50.795 110.080 50.965 ;
        RECT 109.055 49.575 109.515 50.625 ;
        RECT 109.685 49.435 109.855 50.795 ;
        RECT 110.250 50.535 110.715 50.925 ;
        RECT 110.025 49.725 110.375 50.345 ;
        RECT 110.545 49.945 110.715 50.535 ;
        RECT 110.885 50.315 111.055 51.095 ;
        RECT 111.225 50.995 111.395 51.335 ;
        RECT 111.630 51.165 111.960 51.595 ;
        RECT 112.130 50.995 112.300 51.335 ;
        RECT 112.595 51.135 112.965 51.595 ;
        RECT 111.225 50.825 112.300 50.995 ;
        RECT 113.135 50.965 113.305 51.425 ;
        RECT 113.540 51.085 114.410 51.425 ;
        RECT 114.580 51.135 114.830 51.595 ;
        RECT 112.745 50.795 113.305 50.965 ;
        RECT 112.745 50.655 112.915 50.795 ;
        RECT 111.415 50.485 112.915 50.655 ;
        RECT 113.610 50.625 114.070 50.915 ;
        RECT 110.885 50.145 112.575 50.315 ;
        RECT 110.545 49.725 110.900 49.945 ;
        RECT 111.070 49.435 111.240 50.145 ;
        RECT 111.445 49.725 112.235 49.975 ;
        RECT 112.405 49.965 112.575 50.145 ;
        RECT 112.745 49.795 112.915 50.485 ;
        RECT 109.185 49.045 109.515 49.405 ;
        RECT 109.685 49.265 110.180 49.435 ;
        RECT 110.385 49.265 111.240 49.435 ;
        RECT 112.115 49.045 112.445 49.505 ;
        RECT 112.655 49.405 112.915 49.795 ;
        RECT 113.105 50.615 114.070 50.625 ;
        RECT 114.240 50.705 114.410 51.085 ;
        RECT 115.000 51.045 115.170 51.335 ;
        RECT 115.350 51.215 115.680 51.595 ;
        RECT 115.000 50.875 115.800 51.045 ;
        RECT 113.105 50.455 113.780 50.615 ;
        RECT 114.240 50.535 115.460 50.705 ;
        RECT 113.105 49.665 113.315 50.455 ;
        RECT 114.240 50.445 114.410 50.535 ;
        RECT 113.485 49.665 113.835 50.285 ;
        RECT 114.005 50.275 114.410 50.445 ;
        RECT 114.005 49.495 114.175 50.275 ;
        RECT 114.345 49.825 114.565 50.105 ;
        RECT 114.745 49.995 115.285 50.365 ;
        RECT 115.630 50.285 115.800 50.875 ;
        RECT 116.020 50.455 116.325 51.595 ;
        RECT 116.495 50.405 116.750 51.285 ;
        RECT 116.925 50.505 120.435 51.595 ;
        RECT 115.630 50.255 116.370 50.285 ;
        RECT 114.345 49.655 114.875 49.825 ;
        RECT 112.655 49.235 113.005 49.405 ;
        RECT 113.225 49.215 114.175 49.495 ;
        RECT 114.345 49.045 114.535 49.485 ;
        RECT 114.705 49.425 114.875 49.655 ;
        RECT 115.045 49.595 115.285 49.995 ;
        RECT 115.455 49.955 116.370 50.255 ;
        RECT 115.455 49.780 115.780 49.955 ;
        RECT 115.455 49.425 115.775 49.780 ;
        RECT 116.540 49.755 116.750 50.405 ;
        RECT 114.705 49.255 115.775 49.425 ;
        RECT 116.020 49.045 116.325 49.505 ;
        RECT 116.495 49.225 116.750 49.755 ;
        RECT 116.925 49.815 118.575 50.335 ;
        RECT 118.745 49.985 120.435 50.505 ;
        RECT 121.525 50.430 121.815 51.595 ;
        RECT 121.985 50.505 123.655 51.595 ;
        RECT 121.985 49.815 122.735 50.335 ;
        RECT 122.905 49.985 123.655 50.505 ;
        RECT 124.285 50.505 125.495 51.595 ;
        RECT 124.285 49.965 124.805 50.505 ;
        RECT 116.925 49.045 120.435 49.815 ;
        RECT 121.525 49.045 121.815 49.770 ;
        RECT 121.985 49.045 123.655 49.815 ;
        RECT 124.975 49.795 125.495 50.335 ;
        RECT 124.285 49.045 125.495 49.795 ;
        RECT 5.520 48.875 125.580 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.985 48.105 10.495 48.875 ;
        RECT 11.590 48.325 11.845 48.615 ;
        RECT 12.015 48.495 12.345 48.875 ;
        RECT 11.590 48.155 12.340 48.325 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 6.985 47.585 8.635 48.105 ;
        RECT 8.805 47.415 10.495 47.935 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 6.985 46.325 10.495 47.415 ;
        RECT 11.590 47.335 11.940 47.985 ;
        RECT 12.110 47.165 12.340 48.155 ;
        RECT 11.590 46.995 12.340 47.165 ;
        RECT 11.590 46.495 11.845 46.995 ;
        RECT 12.015 46.325 12.345 46.825 ;
        RECT 12.515 46.495 12.685 48.615 ;
        RECT 13.045 48.515 13.375 48.875 ;
        RECT 13.545 48.485 14.040 48.655 ;
        RECT 14.245 48.485 15.100 48.655 ;
        RECT 12.915 47.295 13.375 48.345 ;
        RECT 12.855 46.510 13.180 47.295 ;
        RECT 13.545 47.125 13.715 48.485 ;
        RECT 13.885 47.575 14.235 48.195 ;
        RECT 14.405 47.975 14.760 48.195 ;
        RECT 14.405 47.385 14.575 47.975 ;
        RECT 14.930 47.775 15.100 48.485 ;
        RECT 15.975 48.415 16.305 48.875 ;
        RECT 16.515 48.515 16.865 48.685 ;
        RECT 15.305 47.945 16.095 48.195 ;
        RECT 16.515 48.125 16.775 48.515 ;
        RECT 17.085 48.425 18.035 48.705 ;
        RECT 18.205 48.435 18.395 48.875 ;
        RECT 18.565 48.495 19.635 48.665 ;
        RECT 16.265 47.775 16.435 47.955 ;
        RECT 13.545 46.955 13.940 47.125 ;
        RECT 14.110 46.995 14.575 47.385 ;
        RECT 14.745 47.605 16.435 47.775 ;
        RECT 13.770 46.825 13.940 46.955 ;
        RECT 14.745 46.825 14.915 47.605 ;
        RECT 16.605 47.435 16.775 48.125 ;
        RECT 15.275 47.265 16.775 47.435 ;
        RECT 16.965 47.465 17.175 48.255 ;
        RECT 17.345 47.635 17.695 48.255 ;
        RECT 17.865 47.645 18.035 48.425 ;
        RECT 18.565 48.265 18.735 48.495 ;
        RECT 18.205 48.095 18.735 48.265 ;
        RECT 18.205 47.815 18.425 48.095 ;
        RECT 18.905 47.925 19.145 48.325 ;
        RECT 17.865 47.475 18.270 47.645 ;
        RECT 18.605 47.555 19.145 47.925 ;
        RECT 19.315 48.140 19.635 48.495 ;
        RECT 19.880 48.415 20.185 48.875 ;
        RECT 20.355 48.165 20.610 48.695 ;
        RECT 19.315 47.965 19.640 48.140 ;
        RECT 19.315 47.665 20.230 47.965 ;
        RECT 19.490 47.635 20.230 47.665 ;
        RECT 16.965 47.305 17.640 47.465 ;
        RECT 18.100 47.385 18.270 47.475 ;
        RECT 16.965 47.295 17.930 47.305 ;
        RECT 16.605 47.125 16.775 47.265 ;
        RECT 13.350 46.325 13.600 46.785 ;
        RECT 13.770 46.495 14.020 46.825 ;
        RECT 14.235 46.495 14.915 46.825 ;
        RECT 15.085 46.925 16.160 47.095 ;
        RECT 16.605 46.955 17.165 47.125 ;
        RECT 17.470 47.005 17.930 47.295 ;
        RECT 18.100 47.215 19.320 47.385 ;
        RECT 15.085 46.585 15.255 46.925 ;
        RECT 15.490 46.325 15.820 46.755 ;
        RECT 15.990 46.585 16.160 46.925 ;
        RECT 16.455 46.325 16.825 46.785 ;
        RECT 16.995 46.495 17.165 46.955 ;
        RECT 18.100 46.835 18.270 47.215 ;
        RECT 19.490 47.045 19.660 47.635 ;
        RECT 20.400 47.515 20.610 48.165 ;
        RECT 17.400 46.495 18.270 46.835 ;
        RECT 18.860 46.875 19.660 47.045 ;
        RECT 18.440 46.325 18.690 46.785 ;
        RECT 18.860 46.585 19.030 46.875 ;
        RECT 19.210 46.325 19.540 46.705 ;
        RECT 19.880 46.325 20.185 47.465 ;
        RECT 20.355 46.635 20.610 47.515 ;
        RECT 20.790 48.135 21.045 48.705 ;
        RECT 21.215 48.475 21.545 48.875 ;
        RECT 21.970 48.340 22.500 48.705 ;
        RECT 21.970 48.305 22.145 48.340 ;
        RECT 21.215 48.135 22.145 48.305 ;
        RECT 20.790 47.465 20.960 48.135 ;
        RECT 21.215 47.965 21.385 48.135 ;
        RECT 21.130 47.635 21.385 47.965 ;
        RECT 21.610 47.635 21.805 47.965 ;
        RECT 20.790 46.495 21.125 47.465 ;
        RECT 21.295 46.325 21.465 47.465 ;
        RECT 21.635 46.665 21.805 47.635 ;
        RECT 21.975 47.005 22.145 48.135 ;
        RECT 22.315 47.345 22.485 48.145 ;
        RECT 22.690 47.855 22.965 48.705 ;
        RECT 22.685 47.685 22.965 47.855 ;
        RECT 22.690 47.545 22.965 47.685 ;
        RECT 23.135 47.345 23.325 48.705 ;
        RECT 23.505 48.340 24.015 48.875 ;
        RECT 24.235 48.065 24.480 48.670 ;
        RECT 24.925 48.105 26.595 48.875 ;
        RECT 23.525 47.895 24.755 48.065 ;
        RECT 22.315 47.175 23.325 47.345 ;
        RECT 23.495 47.330 24.245 47.520 ;
        RECT 21.975 46.835 23.100 47.005 ;
        RECT 23.495 46.665 23.665 47.330 ;
        RECT 24.415 47.085 24.755 47.895 ;
        RECT 24.925 47.585 25.675 48.105 ;
        RECT 27.040 48.065 27.285 48.670 ;
        RECT 27.505 48.340 28.015 48.875 ;
        RECT 25.845 47.415 26.595 47.935 ;
        RECT 21.635 46.495 23.665 46.665 ;
        RECT 23.835 46.325 24.005 47.085 ;
        RECT 24.240 46.675 24.755 47.085 ;
        RECT 24.925 46.325 26.595 47.415 ;
        RECT 26.765 47.895 27.995 48.065 ;
        RECT 26.765 47.085 27.105 47.895 ;
        RECT 27.275 47.330 28.025 47.520 ;
        RECT 26.765 46.675 27.280 47.085 ;
        RECT 27.515 46.325 27.685 47.085 ;
        RECT 27.855 46.665 28.025 47.330 ;
        RECT 28.195 47.345 28.385 48.705 ;
        RECT 28.555 48.195 28.830 48.705 ;
        RECT 29.020 48.340 29.550 48.705 ;
        RECT 29.975 48.475 30.305 48.875 ;
        RECT 29.375 48.305 29.550 48.340 ;
        RECT 28.555 48.025 28.835 48.195 ;
        RECT 28.555 47.545 28.830 48.025 ;
        RECT 29.035 47.345 29.205 48.145 ;
        RECT 28.195 47.175 29.205 47.345 ;
        RECT 29.375 48.135 30.305 48.305 ;
        RECT 30.475 48.135 30.730 48.705 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 32.750 48.325 33.005 48.615 ;
        RECT 33.175 48.495 33.505 48.875 ;
        RECT 32.750 48.155 33.500 48.325 ;
        RECT 29.375 47.005 29.545 48.135 ;
        RECT 30.135 47.965 30.305 48.135 ;
        RECT 28.420 46.835 29.545 47.005 ;
        RECT 29.715 47.635 29.910 47.965 ;
        RECT 30.135 47.635 30.390 47.965 ;
        RECT 29.715 46.665 29.885 47.635 ;
        RECT 30.560 47.465 30.730 48.135 ;
        RECT 27.855 46.495 29.885 46.665 ;
        RECT 30.055 46.325 30.225 47.465 ;
        RECT 30.395 46.495 30.730 47.465 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 32.750 47.335 33.100 47.985 ;
        RECT 33.270 47.165 33.500 48.155 ;
        RECT 32.750 46.995 33.500 47.165 ;
        RECT 32.750 46.495 33.005 46.995 ;
        RECT 33.175 46.325 33.505 46.825 ;
        RECT 33.675 46.495 33.845 48.615 ;
        RECT 34.205 48.515 34.535 48.875 ;
        RECT 34.705 48.485 35.200 48.655 ;
        RECT 35.405 48.485 36.260 48.655 ;
        RECT 34.075 47.295 34.535 48.345 ;
        RECT 34.015 46.510 34.340 47.295 ;
        RECT 34.705 47.125 34.875 48.485 ;
        RECT 35.045 47.575 35.395 48.195 ;
        RECT 35.565 47.975 35.920 48.195 ;
        RECT 35.565 47.385 35.735 47.975 ;
        RECT 36.090 47.775 36.260 48.485 ;
        RECT 37.135 48.415 37.465 48.875 ;
        RECT 37.675 48.515 38.025 48.685 ;
        RECT 36.465 47.945 37.255 48.195 ;
        RECT 37.675 48.125 37.935 48.515 ;
        RECT 38.245 48.425 39.195 48.705 ;
        RECT 39.365 48.435 39.555 48.875 ;
        RECT 39.725 48.495 40.795 48.665 ;
        RECT 37.425 47.775 37.595 47.955 ;
        RECT 34.705 46.955 35.100 47.125 ;
        RECT 35.270 46.995 35.735 47.385 ;
        RECT 35.905 47.605 37.595 47.775 ;
        RECT 34.930 46.825 35.100 46.955 ;
        RECT 35.905 46.825 36.075 47.605 ;
        RECT 37.765 47.435 37.935 48.125 ;
        RECT 36.435 47.265 37.935 47.435 ;
        RECT 38.125 47.465 38.335 48.255 ;
        RECT 38.505 47.635 38.855 48.255 ;
        RECT 39.025 47.645 39.195 48.425 ;
        RECT 39.725 48.265 39.895 48.495 ;
        RECT 39.365 48.095 39.895 48.265 ;
        RECT 39.365 47.815 39.585 48.095 ;
        RECT 40.065 47.925 40.305 48.325 ;
        RECT 39.025 47.475 39.430 47.645 ;
        RECT 39.765 47.555 40.305 47.925 ;
        RECT 40.475 48.140 40.795 48.495 ;
        RECT 41.040 48.415 41.345 48.875 ;
        RECT 41.515 48.165 41.770 48.695 ;
        RECT 40.475 47.965 40.800 48.140 ;
        RECT 40.475 47.665 41.390 47.965 ;
        RECT 40.650 47.635 41.390 47.665 ;
        RECT 38.125 47.305 38.800 47.465 ;
        RECT 39.260 47.385 39.430 47.475 ;
        RECT 38.125 47.295 39.090 47.305 ;
        RECT 37.765 47.125 37.935 47.265 ;
        RECT 34.510 46.325 34.760 46.785 ;
        RECT 34.930 46.495 35.180 46.825 ;
        RECT 35.395 46.495 36.075 46.825 ;
        RECT 36.245 46.925 37.320 47.095 ;
        RECT 37.765 46.955 38.325 47.125 ;
        RECT 38.630 47.005 39.090 47.295 ;
        RECT 39.260 47.215 40.480 47.385 ;
        RECT 36.245 46.585 36.415 46.925 ;
        RECT 36.650 46.325 36.980 46.755 ;
        RECT 37.150 46.585 37.320 46.925 ;
        RECT 37.615 46.325 37.985 46.785 ;
        RECT 38.155 46.495 38.325 46.955 ;
        RECT 39.260 46.835 39.430 47.215 ;
        RECT 40.650 47.045 40.820 47.635 ;
        RECT 41.560 47.515 41.770 48.165 ;
        RECT 42.870 48.325 43.125 48.615 ;
        RECT 43.295 48.495 43.625 48.875 ;
        RECT 42.870 48.155 43.620 48.325 ;
        RECT 38.560 46.495 39.430 46.835 ;
        RECT 40.020 46.875 40.820 47.045 ;
        RECT 39.600 46.325 39.850 46.785 ;
        RECT 40.020 46.585 40.190 46.875 ;
        RECT 40.370 46.325 40.700 46.705 ;
        RECT 41.040 46.325 41.345 47.465 ;
        RECT 41.515 46.635 41.770 47.515 ;
        RECT 42.870 47.335 43.220 47.985 ;
        RECT 43.390 47.165 43.620 48.155 ;
        RECT 42.870 46.995 43.620 47.165 ;
        RECT 42.870 46.495 43.125 46.995 ;
        RECT 43.295 46.325 43.625 46.825 ;
        RECT 43.795 46.495 43.965 48.615 ;
        RECT 44.325 48.515 44.655 48.875 ;
        RECT 44.825 48.485 45.320 48.655 ;
        RECT 45.525 48.485 46.380 48.655 ;
        RECT 44.195 47.295 44.655 48.345 ;
        RECT 44.135 46.510 44.460 47.295 ;
        RECT 44.825 47.125 44.995 48.485 ;
        RECT 45.165 47.575 45.515 48.195 ;
        RECT 45.685 47.975 46.040 48.195 ;
        RECT 45.685 47.385 45.855 47.975 ;
        RECT 46.210 47.775 46.380 48.485 ;
        RECT 47.255 48.415 47.585 48.875 ;
        RECT 47.795 48.515 48.145 48.685 ;
        RECT 46.585 47.945 47.375 48.195 ;
        RECT 47.795 48.125 48.055 48.515 ;
        RECT 48.365 48.425 49.315 48.705 ;
        RECT 49.485 48.435 49.675 48.875 ;
        RECT 49.845 48.495 50.915 48.665 ;
        RECT 47.545 47.775 47.715 47.955 ;
        RECT 44.825 46.955 45.220 47.125 ;
        RECT 45.390 46.995 45.855 47.385 ;
        RECT 46.025 47.605 47.715 47.775 ;
        RECT 45.050 46.825 45.220 46.955 ;
        RECT 46.025 46.825 46.195 47.605 ;
        RECT 47.885 47.435 48.055 48.125 ;
        RECT 46.555 47.265 48.055 47.435 ;
        RECT 48.245 47.465 48.455 48.255 ;
        RECT 48.625 47.635 48.975 48.255 ;
        RECT 49.145 47.645 49.315 48.425 ;
        RECT 49.845 48.265 50.015 48.495 ;
        RECT 49.485 48.095 50.015 48.265 ;
        RECT 49.485 47.815 49.705 48.095 ;
        RECT 50.185 47.925 50.425 48.325 ;
        RECT 49.145 47.475 49.550 47.645 ;
        RECT 49.885 47.555 50.425 47.925 ;
        RECT 50.595 48.140 50.915 48.495 ;
        RECT 51.160 48.415 51.465 48.875 ;
        RECT 51.635 48.165 51.890 48.695 ;
        RECT 50.595 47.965 50.920 48.140 ;
        RECT 50.595 47.665 51.510 47.965 ;
        RECT 50.770 47.635 51.510 47.665 ;
        RECT 48.245 47.305 48.920 47.465 ;
        RECT 49.380 47.385 49.550 47.475 ;
        RECT 48.245 47.295 49.210 47.305 ;
        RECT 47.885 47.125 48.055 47.265 ;
        RECT 44.630 46.325 44.880 46.785 ;
        RECT 45.050 46.495 45.300 46.825 ;
        RECT 45.515 46.495 46.195 46.825 ;
        RECT 46.365 46.925 47.440 47.095 ;
        RECT 47.885 46.955 48.445 47.125 ;
        RECT 48.750 47.005 49.210 47.295 ;
        RECT 49.380 47.215 50.600 47.385 ;
        RECT 46.365 46.585 46.535 46.925 ;
        RECT 46.770 46.325 47.100 46.755 ;
        RECT 47.270 46.585 47.440 46.925 ;
        RECT 47.735 46.325 48.105 46.785 ;
        RECT 48.275 46.495 48.445 46.955 ;
        RECT 49.380 46.835 49.550 47.215 ;
        RECT 50.770 47.045 50.940 47.635 ;
        RECT 51.680 47.515 51.890 48.165 ;
        RECT 52.270 48.095 52.770 48.705 ;
        RECT 52.065 47.635 52.415 47.885 ;
        RECT 48.680 46.495 49.550 46.835 ;
        RECT 50.140 46.875 50.940 47.045 ;
        RECT 49.720 46.325 49.970 46.785 ;
        RECT 50.140 46.585 50.310 46.875 ;
        RECT 50.490 46.325 50.820 46.705 ;
        RECT 51.160 46.325 51.465 47.465 ;
        RECT 51.635 46.635 51.890 47.515 ;
        RECT 52.600 47.465 52.770 48.095 ;
        RECT 53.400 48.225 53.730 48.705 ;
        RECT 53.900 48.415 54.125 48.875 ;
        RECT 54.295 48.225 54.625 48.705 ;
        RECT 53.400 48.055 54.625 48.225 ;
        RECT 54.815 48.075 55.065 48.875 ;
        RECT 55.235 48.075 55.575 48.705 ;
        RECT 55.345 48.025 55.575 48.075 ;
        RECT 55.785 48.055 56.015 48.875 ;
        RECT 56.185 48.075 56.515 48.705 ;
        RECT 52.940 47.685 53.270 47.885 ;
        RECT 53.440 47.685 53.770 47.885 ;
        RECT 53.940 47.685 54.360 47.885 ;
        RECT 54.535 47.715 55.230 47.885 ;
        RECT 54.535 47.465 54.705 47.715 ;
        RECT 55.400 47.465 55.575 48.025 ;
        RECT 55.765 47.635 56.095 47.885 ;
        RECT 56.265 47.475 56.515 48.075 ;
        RECT 56.685 48.055 56.895 48.875 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 57.585 48.105 61.095 48.875 ;
        RECT 62.490 48.305 62.660 48.555 ;
        RECT 62.185 48.135 62.660 48.305 ;
        RECT 62.895 48.135 63.225 48.875 ;
        RECT 63.395 48.305 63.595 48.650 ;
        RECT 63.765 48.475 64.095 48.875 ;
        RECT 64.265 48.305 64.465 48.660 ;
        RECT 64.635 48.480 64.965 48.875 ;
        RECT 65.405 48.330 70.750 48.875 ;
        RECT 63.395 48.135 65.235 48.305 ;
        RECT 57.585 47.585 59.235 48.105 ;
        RECT 52.270 47.295 54.705 47.465 ;
        RECT 52.270 46.495 52.600 47.295 ;
        RECT 52.770 46.325 53.100 47.125 ;
        RECT 53.400 46.495 53.730 47.295 ;
        RECT 54.375 46.325 54.625 47.125 ;
        RECT 54.895 46.325 55.065 47.465 ;
        RECT 55.235 46.495 55.575 47.465 ;
        RECT 55.785 46.325 56.015 47.465 ;
        RECT 56.185 46.495 56.515 47.475 ;
        RECT 56.685 46.325 56.895 47.465 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 59.405 47.415 61.095 47.935 ;
        RECT 57.585 46.325 61.095 47.415 ;
        RECT 62.185 47.165 62.355 48.135 ;
        RECT 62.525 47.345 62.875 47.965 ;
        RECT 63.045 47.345 63.365 47.965 ;
        RECT 63.535 47.345 63.865 47.965 ;
        RECT 64.035 47.345 64.335 47.965 ;
        RECT 64.575 47.165 64.795 47.965 ;
        RECT 62.185 46.955 64.795 47.165 ;
        RECT 62.895 46.325 63.225 46.775 ;
        RECT 64.975 46.510 65.235 48.135 ;
        RECT 66.990 47.500 67.330 48.330 ;
        RECT 70.925 48.105 74.435 48.875 ;
        RECT 75.525 48.200 75.785 48.705 ;
        RECT 75.965 48.495 76.295 48.875 ;
        RECT 76.475 48.325 76.645 48.705 ;
        RECT 68.810 46.760 69.160 48.010 ;
        RECT 70.925 47.585 72.575 48.105 ;
        RECT 72.745 47.415 74.435 47.935 ;
        RECT 65.405 46.325 70.750 46.760 ;
        RECT 70.925 46.325 74.435 47.415 ;
        RECT 75.525 47.400 75.695 48.200 ;
        RECT 75.980 48.155 76.645 48.325 ;
        RECT 75.980 47.900 76.150 48.155 ;
        RECT 77.180 48.065 77.425 48.670 ;
        RECT 77.645 48.340 78.155 48.875 ;
        RECT 75.865 47.570 76.150 47.900 ;
        RECT 76.385 47.605 76.715 47.975 ;
        RECT 76.905 47.895 78.135 48.065 ;
        RECT 75.980 47.425 76.150 47.570 ;
        RECT 75.525 46.495 75.795 47.400 ;
        RECT 75.980 47.255 76.645 47.425 ;
        RECT 75.965 46.325 76.295 47.085 ;
        RECT 76.475 46.495 76.645 47.255 ;
        RECT 76.905 47.085 77.245 47.895 ;
        RECT 77.415 47.330 78.165 47.520 ;
        RECT 76.905 46.675 77.420 47.085 ;
        RECT 77.655 46.325 77.825 47.085 ;
        RECT 77.995 46.665 78.165 47.330 ;
        RECT 78.335 47.345 78.525 48.705 ;
        RECT 78.695 47.855 78.970 48.705 ;
        RECT 79.160 48.340 79.690 48.705 ;
        RECT 80.115 48.475 80.445 48.875 ;
        RECT 79.515 48.305 79.690 48.340 ;
        RECT 78.695 47.685 78.975 47.855 ;
        RECT 78.695 47.545 78.970 47.685 ;
        RECT 79.175 47.345 79.345 48.145 ;
        RECT 78.335 47.175 79.345 47.345 ;
        RECT 79.515 48.135 80.445 48.305 ;
        RECT 80.615 48.135 80.870 48.705 ;
        RECT 79.515 47.005 79.685 48.135 ;
        RECT 80.275 47.965 80.445 48.135 ;
        RECT 78.560 46.835 79.685 47.005 ;
        RECT 79.855 47.635 80.050 47.965 ;
        RECT 80.275 47.635 80.530 47.965 ;
        RECT 79.855 46.665 80.025 47.635 ;
        RECT 80.700 47.465 80.870 48.135 ;
        RECT 81.045 48.105 82.715 48.875 ;
        RECT 82.885 48.150 83.175 48.875 ;
        RECT 81.045 47.585 81.795 48.105 ;
        RECT 83.345 48.075 83.685 48.705 ;
        RECT 83.855 48.075 84.105 48.875 ;
        RECT 84.295 48.225 84.625 48.705 ;
        RECT 84.795 48.415 85.020 48.875 ;
        RECT 85.190 48.225 85.520 48.705 ;
        RECT 77.995 46.495 80.025 46.665 ;
        RECT 80.195 46.325 80.365 47.465 ;
        RECT 80.535 46.495 80.870 47.465 ;
        RECT 81.965 47.415 82.715 47.935 ;
        RECT 81.045 46.325 82.715 47.415 ;
        RECT 82.885 46.325 83.175 47.490 ;
        RECT 83.345 47.465 83.520 48.075 ;
        RECT 84.295 48.055 85.520 48.225 ;
        RECT 86.150 48.095 86.650 48.705 ;
        RECT 87.025 48.105 89.615 48.875 ;
        RECT 89.790 48.135 90.045 48.705 ;
        RECT 90.215 48.475 90.545 48.875 ;
        RECT 90.970 48.340 91.500 48.705 ;
        RECT 90.970 48.305 91.145 48.340 ;
        RECT 90.215 48.135 91.145 48.305 ;
        RECT 83.690 47.715 84.385 47.885 ;
        RECT 84.215 47.465 84.385 47.715 ;
        RECT 84.560 47.685 84.980 47.885 ;
        RECT 85.150 47.685 85.480 47.885 ;
        RECT 85.650 47.685 85.980 47.885 ;
        RECT 86.150 47.465 86.320 48.095 ;
        RECT 86.505 47.635 86.855 47.885 ;
        RECT 87.025 47.585 88.235 48.105 ;
        RECT 83.345 46.495 83.685 47.465 ;
        RECT 83.855 46.325 84.025 47.465 ;
        RECT 84.215 47.295 86.650 47.465 ;
        RECT 88.405 47.415 89.615 47.935 ;
        RECT 84.295 46.325 84.545 47.125 ;
        RECT 85.190 46.495 85.520 47.295 ;
        RECT 85.820 46.325 86.150 47.125 ;
        RECT 86.320 46.495 86.650 47.295 ;
        RECT 87.025 46.325 89.615 47.415 ;
        RECT 89.790 47.465 89.960 48.135 ;
        RECT 90.215 47.965 90.385 48.135 ;
        RECT 90.130 47.635 90.385 47.965 ;
        RECT 90.610 47.635 90.805 47.965 ;
        RECT 89.790 46.495 90.125 47.465 ;
        RECT 90.295 46.325 90.465 47.465 ;
        RECT 90.635 46.665 90.805 47.635 ;
        RECT 90.975 47.005 91.145 48.135 ;
        RECT 91.315 47.345 91.485 48.145 ;
        RECT 91.690 47.855 91.965 48.705 ;
        RECT 91.685 47.685 91.965 47.855 ;
        RECT 91.690 47.545 91.965 47.685 ;
        RECT 92.135 47.345 92.325 48.705 ;
        RECT 92.505 48.340 93.015 48.875 ;
        RECT 93.235 48.065 93.480 48.670 ;
        RECT 93.925 48.105 97.435 48.875 ;
        RECT 98.180 48.245 98.465 48.705 ;
        RECT 98.635 48.415 98.905 48.875 ;
        RECT 92.525 47.895 93.755 48.065 ;
        RECT 91.315 47.175 92.325 47.345 ;
        RECT 92.495 47.330 93.245 47.520 ;
        RECT 90.975 46.835 92.100 47.005 ;
        RECT 92.495 46.665 92.665 47.330 ;
        RECT 93.415 47.085 93.755 47.895 ;
        RECT 93.925 47.585 95.575 48.105 ;
        RECT 98.180 48.075 99.135 48.245 ;
        RECT 95.745 47.415 97.435 47.935 ;
        RECT 90.635 46.495 92.665 46.665 ;
        RECT 92.835 46.325 93.005 47.085 ;
        RECT 93.240 46.675 93.755 47.085 ;
        RECT 93.925 46.325 97.435 47.415 ;
        RECT 98.065 47.345 98.755 47.905 ;
        RECT 98.925 47.175 99.135 48.075 ;
        RECT 98.180 46.955 99.135 47.175 ;
        RECT 99.305 47.905 99.705 48.705 ;
        RECT 99.895 48.245 100.175 48.705 ;
        RECT 100.695 48.415 101.020 48.875 ;
        RECT 99.895 48.075 101.020 48.245 ;
        RECT 101.190 48.135 101.575 48.705 ;
        RECT 101.745 48.330 107.090 48.875 ;
        RECT 100.570 47.965 101.020 48.075 ;
        RECT 99.305 47.345 100.400 47.905 ;
        RECT 100.570 47.635 101.125 47.965 ;
        RECT 98.180 46.495 98.465 46.955 ;
        RECT 98.635 46.325 98.905 46.785 ;
        RECT 99.305 46.495 99.705 47.345 ;
        RECT 100.570 47.175 101.020 47.635 ;
        RECT 101.295 47.465 101.575 48.135 ;
        RECT 103.330 47.500 103.670 48.330 ;
        RECT 107.355 48.325 107.525 48.705 ;
        RECT 107.705 48.495 108.035 48.875 ;
        RECT 107.355 48.155 108.020 48.325 ;
        RECT 108.215 48.200 108.475 48.705 ;
        RECT 99.895 46.955 101.020 47.175 ;
        RECT 99.895 46.495 100.175 46.955 ;
        RECT 100.695 46.325 101.020 46.785 ;
        RECT 101.190 46.495 101.575 47.465 ;
        RECT 105.150 46.760 105.500 48.010 ;
        RECT 107.285 47.605 107.615 47.975 ;
        RECT 107.850 47.900 108.020 48.155 ;
        RECT 107.850 47.570 108.135 47.900 ;
        RECT 107.850 47.425 108.020 47.570 ;
        RECT 107.355 47.255 108.020 47.425 ;
        RECT 108.305 47.400 108.475 48.200 ;
        RECT 108.645 48.150 108.935 48.875 ;
        RECT 109.105 48.135 109.490 48.705 ;
        RECT 109.660 48.415 109.985 48.875 ;
        RECT 110.505 48.245 110.785 48.705 ;
        RECT 101.745 46.325 107.090 46.760 ;
        RECT 107.355 46.495 107.525 47.255 ;
        RECT 107.705 46.325 108.035 47.085 ;
        RECT 108.205 46.495 108.475 47.400 ;
        RECT 108.645 46.325 108.935 47.490 ;
        RECT 109.105 47.465 109.385 48.135 ;
        RECT 109.660 48.075 110.785 48.245 ;
        RECT 109.660 47.965 110.110 48.075 ;
        RECT 109.555 47.635 110.110 47.965 ;
        RECT 110.975 47.905 111.375 48.705 ;
        RECT 111.775 48.415 112.045 48.875 ;
        RECT 112.215 48.245 112.500 48.705 ;
        RECT 109.105 46.495 109.490 47.465 ;
        RECT 109.660 47.175 110.110 47.635 ;
        RECT 110.280 47.345 111.375 47.905 ;
        RECT 109.660 46.955 110.785 47.175 ;
        RECT 109.660 46.325 109.985 46.785 ;
        RECT 110.505 46.495 110.785 46.955 ;
        RECT 110.975 46.495 111.375 47.345 ;
        RECT 111.545 48.075 112.500 48.245 ;
        RECT 112.785 48.135 113.170 48.705 ;
        RECT 113.340 48.415 113.665 48.875 ;
        RECT 114.185 48.245 114.465 48.705 ;
        RECT 111.545 47.175 111.755 48.075 ;
        RECT 111.925 47.345 112.615 47.905 ;
        RECT 112.785 47.465 113.065 48.135 ;
        RECT 113.340 48.075 114.465 48.245 ;
        RECT 113.340 47.965 113.790 48.075 ;
        RECT 113.235 47.635 113.790 47.965 ;
        RECT 114.655 47.905 115.055 48.705 ;
        RECT 115.455 48.415 115.725 48.875 ;
        RECT 115.895 48.245 116.180 48.705 ;
        RECT 116.465 48.330 121.810 48.875 ;
        RECT 111.545 46.955 112.500 47.175 ;
        RECT 111.775 46.325 112.045 46.785 ;
        RECT 112.215 46.495 112.500 46.955 ;
        RECT 112.785 46.495 113.170 47.465 ;
        RECT 113.340 47.175 113.790 47.635 ;
        RECT 113.960 47.345 115.055 47.905 ;
        RECT 113.340 46.955 114.465 47.175 ;
        RECT 113.340 46.325 113.665 46.785 ;
        RECT 114.185 46.495 114.465 46.955 ;
        RECT 114.655 46.495 115.055 47.345 ;
        RECT 115.225 48.075 116.180 48.245 ;
        RECT 115.225 47.175 115.435 48.075 ;
        RECT 115.605 47.345 116.295 47.905 ;
        RECT 118.050 47.500 118.390 48.330 ;
        RECT 121.985 48.105 123.655 48.875 ;
        RECT 124.285 48.125 125.495 48.875 ;
        RECT 115.225 46.955 116.180 47.175 ;
        RECT 115.455 46.325 115.725 46.785 ;
        RECT 115.895 46.495 116.180 46.955 ;
        RECT 119.870 46.760 120.220 48.010 ;
        RECT 121.985 47.585 122.735 48.105 ;
        RECT 122.905 47.415 123.655 47.935 ;
        RECT 116.465 46.325 121.810 46.760 ;
        RECT 121.985 46.325 123.655 47.415 ;
        RECT 124.285 47.415 124.805 47.955 ;
        RECT 124.975 47.585 125.495 48.125 ;
        RECT 124.285 46.325 125.495 47.415 ;
        RECT 5.520 46.155 125.580 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 6.985 45.065 8.655 46.155 ;
        RECT 9.290 45.485 9.545 45.985 ;
        RECT 9.715 45.655 10.045 46.155 ;
        RECT 9.290 45.315 10.040 45.485 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 6.985 44.375 7.735 44.895 ;
        RECT 7.905 44.545 8.655 45.065 ;
        RECT 9.290 44.495 9.640 45.145 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 6.985 43.605 8.655 44.375 ;
        RECT 9.810 44.325 10.040 45.315 ;
        RECT 9.290 44.155 10.040 44.325 ;
        RECT 9.290 43.865 9.545 44.155 ;
        RECT 9.715 43.605 10.045 43.985 ;
        RECT 10.215 43.865 10.385 45.985 ;
        RECT 10.555 45.185 10.880 45.970 ;
        RECT 11.050 45.695 11.300 46.155 ;
        RECT 11.470 45.655 11.720 45.985 ;
        RECT 11.935 45.655 12.615 45.985 ;
        RECT 11.470 45.525 11.640 45.655 ;
        RECT 11.245 45.355 11.640 45.525 ;
        RECT 10.615 44.135 11.075 45.185 ;
        RECT 11.245 43.995 11.415 45.355 ;
        RECT 11.810 45.095 12.275 45.485 ;
        RECT 11.585 44.285 11.935 44.905 ;
        RECT 12.105 44.505 12.275 45.095 ;
        RECT 12.445 44.875 12.615 45.655 ;
        RECT 12.785 45.555 12.955 45.895 ;
        RECT 13.190 45.725 13.520 46.155 ;
        RECT 13.690 45.555 13.860 45.895 ;
        RECT 14.155 45.695 14.525 46.155 ;
        RECT 12.785 45.385 13.860 45.555 ;
        RECT 14.695 45.525 14.865 45.985 ;
        RECT 15.100 45.645 15.970 45.985 ;
        RECT 16.140 45.695 16.390 46.155 ;
        RECT 14.305 45.355 14.865 45.525 ;
        RECT 14.305 45.215 14.475 45.355 ;
        RECT 12.975 45.045 14.475 45.215 ;
        RECT 15.170 45.185 15.630 45.475 ;
        RECT 12.445 44.705 14.135 44.875 ;
        RECT 12.105 44.285 12.460 44.505 ;
        RECT 12.630 43.995 12.800 44.705 ;
        RECT 13.005 44.285 13.795 44.535 ;
        RECT 13.965 44.525 14.135 44.705 ;
        RECT 14.305 44.355 14.475 45.045 ;
        RECT 10.745 43.605 11.075 43.965 ;
        RECT 11.245 43.825 11.740 43.995 ;
        RECT 11.945 43.825 12.800 43.995 ;
        RECT 13.675 43.605 14.005 44.065 ;
        RECT 14.215 43.965 14.475 44.355 ;
        RECT 14.665 45.175 15.630 45.185 ;
        RECT 15.800 45.265 15.970 45.645 ;
        RECT 16.560 45.605 16.730 45.895 ;
        RECT 16.910 45.775 17.240 46.155 ;
        RECT 16.560 45.435 17.360 45.605 ;
        RECT 14.665 45.015 15.340 45.175 ;
        RECT 15.800 45.095 17.020 45.265 ;
        RECT 14.665 44.225 14.875 45.015 ;
        RECT 15.800 45.005 15.970 45.095 ;
        RECT 15.045 44.225 15.395 44.845 ;
        RECT 15.565 44.835 15.970 45.005 ;
        RECT 15.565 44.055 15.735 44.835 ;
        RECT 15.905 44.385 16.125 44.665 ;
        RECT 16.305 44.555 16.845 44.925 ;
        RECT 17.190 44.845 17.360 45.435 ;
        RECT 17.580 45.015 17.885 46.155 ;
        RECT 18.055 44.965 18.310 45.845 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 18.950 45.015 19.285 45.985 ;
        RECT 19.455 45.015 19.625 46.155 ;
        RECT 19.795 45.815 21.825 45.985 ;
        RECT 17.190 44.815 17.930 44.845 ;
        RECT 15.905 44.215 16.435 44.385 ;
        RECT 14.215 43.795 14.565 43.965 ;
        RECT 14.785 43.775 15.735 44.055 ;
        RECT 15.905 43.605 16.095 44.045 ;
        RECT 16.265 43.985 16.435 44.215 ;
        RECT 16.605 44.155 16.845 44.555 ;
        RECT 17.015 44.515 17.930 44.815 ;
        RECT 17.015 44.340 17.340 44.515 ;
        RECT 17.015 43.985 17.335 44.340 ;
        RECT 18.100 44.315 18.310 44.965 ;
        RECT 18.950 44.345 19.120 45.015 ;
        RECT 19.795 44.845 19.965 45.815 ;
        RECT 19.290 44.515 19.545 44.845 ;
        RECT 19.770 44.515 19.965 44.845 ;
        RECT 20.135 45.475 21.260 45.645 ;
        RECT 19.375 44.345 19.545 44.515 ;
        RECT 20.135 44.345 20.305 45.475 ;
        RECT 16.265 43.815 17.335 43.985 ;
        RECT 17.580 43.605 17.885 44.065 ;
        RECT 18.055 43.785 18.310 44.315 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 18.950 43.775 19.205 44.345 ;
        RECT 19.375 44.175 20.305 44.345 ;
        RECT 20.475 45.135 21.485 45.305 ;
        RECT 20.475 44.335 20.645 45.135 ;
        RECT 20.130 44.140 20.305 44.175 ;
        RECT 19.375 43.605 19.705 44.005 ;
        RECT 20.130 43.775 20.660 44.140 ;
        RECT 20.850 44.115 21.125 44.935 ;
        RECT 20.845 43.945 21.125 44.115 ;
        RECT 20.850 43.775 21.125 43.945 ;
        RECT 21.295 43.775 21.485 45.135 ;
        RECT 21.655 45.150 21.825 45.815 ;
        RECT 21.995 45.395 22.165 46.155 ;
        RECT 22.400 45.395 22.915 45.805 ;
        RECT 21.655 44.960 22.405 45.150 ;
        RECT 22.575 44.585 22.915 45.395 ;
        RECT 23.085 45.065 24.295 46.155 ;
        RECT 21.685 44.415 22.915 44.585 ;
        RECT 21.665 43.605 22.175 44.140 ;
        RECT 22.395 43.810 22.640 44.415 ;
        RECT 23.085 44.355 23.605 44.895 ;
        RECT 23.775 44.525 24.295 45.065 ;
        RECT 24.555 45.225 24.725 45.985 ;
        RECT 24.905 45.395 25.235 46.155 ;
        RECT 24.555 45.055 25.220 45.225 ;
        RECT 25.405 45.080 25.675 45.985 ;
        RECT 25.850 45.485 26.105 45.985 ;
        RECT 26.275 45.655 26.605 46.155 ;
        RECT 25.850 45.315 26.600 45.485 ;
        RECT 25.050 44.910 25.220 45.055 ;
        RECT 24.485 44.505 24.815 44.875 ;
        RECT 25.050 44.580 25.335 44.910 ;
        RECT 23.085 43.605 24.295 44.355 ;
        RECT 25.050 44.325 25.220 44.580 ;
        RECT 24.555 44.155 25.220 44.325 ;
        RECT 25.505 44.280 25.675 45.080 ;
        RECT 25.850 44.495 26.200 45.145 ;
        RECT 26.370 44.325 26.600 45.315 ;
        RECT 24.555 43.775 24.725 44.155 ;
        RECT 24.905 43.605 25.235 43.985 ;
        RECT 25.415 43.775 25.675 44.280 ;
        RECT 25.850 44.155 26.600 44.325 ;
        RECT 25.850 43.865 26.105 44.155 ;
        RECT 26.275 43.605 26.605 43.985 ;
        RECT 26.775 43.865 26.945 45.985 ;
        RECT 27.115 45.185 27.440 45.970 ;
        RECT 27.610 45.695 27.860 46.155 ;
        RECT 28.030 45.655 28.280 45.985 ;
        RECT 28.495 45.655 29.175 45.985 ;
        RECT 28.030 45.525 28.200 45.655 ;
        RECT 27.805 45.355 28.200 45.525 ;
        RECT 27.175 44.135 27.635 45.185 ;
        RECT 27.805 43.995 27.975 45.355 ;
        RECT 28.370 45.095 28.835 45.485 ;
        RECT 28.145 44.285 28.495 44.905 ;
        RECT 28.665 44.505 28.835 45.095 ;
        RECT 29.005 44.875 29.175 45.655 ;
        RECT 29.345 45.555 29.515 45.895 ;
        RECT 29.750 45.725 30.080 46.155 ;
        RECT 30.250 45.555 30.420 45.895 ;
        RECT 30.715 45.695 31.085 46.155 ;
        RECT 29.345 45.385 30.420 45.555 ;
        RECT 31.255 45.525 31.425 45.985 ;
        RECT 31.660 45.645 32.530 45.985 ;
        RECT 32.700 45.695 32.950 46.155 ;
        RECT 30.865 45.355 31.425 45.525 ;
        RECT 30.865 45.215 31.035 45.355 ;
        RECT 29.535 45.045 31.035 45.215 ;
        RECT 31.730 45.185 32.190 45.475 ;
        RECT 29.005 44.705 30.695 44.875 ;
        RECT 28.665 44.285 29.020 44.505 ;
        RECT 29.190 43.995 29.360 44.705 ;
        RECT 29.565 44.285 30.355 44.535 ;
        RECT 30.525 44.525 30.695 44.705 ;
        RECT 30.865 44.355 31.035 45.045 ;
        RECT 27.305 43.605 27.635 43.965 ;
        RECT 27.805 43.825 28.300 43.995 ;
        RECT 28.505 43.825 29.360 43.995 ;
        RECT 30.235 43.605 30.565 44.065 ;
        RECT 30.775 43.965 31.035 44.355 ;
        RECT 31.225 45.175 32.190 45.185 ;
        RECT 32.360 45.265 32.530 45.645 ;
        RECT 33.120 45.605 33.290 45.895 ;
        RECT 33.470 45.775 33.800 46.155 ;
        RECT 33.120 45.435 33.920 45.605 ;
        RECT 31.225 45.015 31.900 45.175 ;
        RECT 32.360 45.095 33.580 45.265 ;
        RECT 31.225 44.225 31.435 45.015 ;
        RECT 32.360 45.005 32.530 45.095 ;
        RECT 31.605 44.225 31.955 44.845 ;
        RECT 32.125 44.835 32.530 45.005 ;
        RECT 32.125 44.055 32.295 44.835 ;
        RECT 32.465 44.385 32.685 44.665 ;
        RECT 32.865 44.555 33.405 44.925 ;
        RECT 33.750 44.845 33.920 45.435 ;
        RECT 34.140 45.015 34.445 46.155 ;
        RECT 34.615 44.965 34.870 45.845 ;
        RECT 36.080 45.525 36.365 45.985 ;
        RECT 36.535 45.695 36.805 46.155 ;
        RECT 36.080 45.305 37.035 45.525 ;
        RECT 33.750 44.815 34.490 44.845 ;
        RECT 32.465 44.215 32.995 44.385 ;
        RECT 30.775 43.795 31.125 43.965 ;
        RECT 31.345 43.775 32.295 44.055 ;
        RECT 32.465 43.605 32.655 44.045 ;
        RECT 32.825 43.985 32.995 44.215 ;
        RECT 33.165 44.155 33.405 44.555 ;
        RECT 33.575 44.515 34.490 44.815 ;
        RECT 33.575 44.340 33.900 44.515 ;
        RECT 33.575 43.985 33.895 44.340 ;
        RECT 34.660 44.315 34.870 44.965 ;
        RECT 35.965 44.575 36.655 45.135 ;
        RECT 36.825 44.405 37.035 45.305 ;
        RECT 32.825 43.815 33.895 43.985 ;
        RECT 34.140 43.605 34.445 44.065 ;
        RECT 34.615 43.785 34.870 44.315 ;
        RECT 36.080 44.235 37.035 44.405 ;
        RECT 37.205 45.135 37.605 45.985 ;
        RECT 37.795 45.525 38.075 45.985 ;
        RECT 38.595 45.695 38.920 46.155 ;
        RECT 37.795 45.305 38.920 45.525 ;
        RECT 37.205 44.575 38.300 45.135 ;
        RECT 38.470 44.845 38.920 45.305 ;
        RECT 39.090 45.015 39.475 45.985 ;
        RECT 39.705 45.015 39.915 46.155 ;
        RECT 36.080 43.775 36.365 44.235 ;
        RECT 36.535 43.605 36.805 44.065 ;
        RECT 37.205 43.775 37.605 44.575 ;
        RECT 38.470 44.515 39.025 44.845 ;
        RECT 38.470 44.405 38.920 44.515 ;
        RECT 37.795 44.235 38.920 44.405 ;
        RECT 39.195 44.345 39.475 45.015 ;
        RECT 40.085 45.005 40.415 45.985 ;
        RECT 40.585 45.015 40.815 46.155 ;
        RECT 41.025 45.065 43.615 46.155 ;
        RECT 37.795 43.775 38.075 44.235 ;
        RECT 38.595 43.605 38.920 44.065 ;
        RECT 39.090 43.775 39.475 44.345 ;
        RECT 39.705 43.605 39.915 44.425 ;
        RECT 40.085 44.405 40.335 45.005 ;
        RECT 40.505 44.595 40.835 44.845 ;
        RECT 40.085 43.775 40.415 44.405 ;
        RECT 40.585 43.605 40.815 44.425 ;
        RECT 41.025 44.375 42.235 44.895 ;
        RECT 42.405 44.545 43.615 45.065 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 45.630 45.015 45.965 45.985 ;
        RECT 46.135 45.015 46.305 46.155 ;
        RECT 46.475 45.815 48.505 45.985 ;
        RECT 41.025 43.605 43.615 44.375 ;
        RECT 45.630 44.345 45.800 45.015 ;
        RECT 46.475 44.845 46.645 45.815 ;
        RECT 45.970 44.515 46.225 44.845 ;
        RECT 46.450 44.515 46.645 44.845 ;
        RECT 46.815 45.475 47.940 45.645 ;
        RECT 46.055 44.345 46.225 44.515 ;
        RECT 46.815 44.345 46.985 45.475 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 45.630 43.775 45.885 44.345 ;
        RECT 46.055 44.175 46.985 44.345 ;
        RECT 47.155 45.135 48.165 45.305 ;
        RECT 47.155 44.335 47.325 45.135 ;
        RECT 47.530 44.795 47.805 44.935 ;
        RECT 47.525 44.625 47.805 44.795 ;
        RECT 46.810 44.140 46.985 44.175 ;
        RECT 46.055 43.605 46.385 44.005 ;
        RECT 46.810 43.775 47.340 44.140 ;
        RECT 47.530 43.775 47.805 44.625 ;
        RECT 47.975 43.775 48.165 45.135 ;
        RECT 48.335 45.150 48.505 45.815 ;
        RECT 48.675 45.395 48.845 46.155 ;
        RECT 49.080 45.395 49.595 45.805 ;
        RECT 48.335 44.960 49.085 45.150 ;
        RECT 49.255 44.585 49.595 45.395 ;
        RECT 48.365 44.415 49.595 44.585 ;
        RECT 49.770 45.015 50.105 45.985 ;
        RECT 50.275 45.015 50.445 46.155 ;
        RECT 50.615 45.815 52.645 45.985 ;
        RECT 48.345 43.605 48.855 44.140 ;
        RECT 49.075 43.810 49.320 44.415 ;
        RECT 49.770 44.345 49.940 45.015 ;
        RECT 50.615 44.845 50.785 45.815 ;
        RECT 50.110 44.515 50.365 44.845 ;
        RECT 50.590 44.515 50.785 44.845 ;
        RECT 50.955 45.475 52.080 45.645 ;
        RECT 50.195 44.345 50.365 44.515 ;
        RECT 50.955 44.345 51.125 45.475 ;
        RECT 49.770 43.775 50.025 44.345 ;
        RECT 50.195 44.175 51.125 44.345 ;
        RECT 51.295 45.135 52.305 45.305 ;
        RECT 51.295 44.335 51.465 45.135 ;
        RECT 51.670 44.455 51.945 44.935 ;
        RECT 51.665 44.285 51.945 44.455 ;
        RECT 50.950 44.140 51.125 44.175 ;
        RECT 50.195 43.605 50.525 44.005 ;
        RECT 50.950 43.775 51.480 44.140 ;
        RECT 51.670 43.775 51.945 44.285 ;
        RECT 52.115 43.775 52.305 45.135 ;
        RECT 52.475 45.150 52.645 45.815 ;
        RECT 52.815 45.395 52.985 46.155 ;
        RECT 53.220 45.395 53.735 45.805 ;
        RECT 52.475 44.960 53.225 45.150 ;
        RECT 53.395 44.585 53.735 45.395 ;
        RECT 52.505 44.415 53.735 44.585 ;
        RECT 53.905 45.015 54.290 45.985 ;
        RECT 54.460 45.695 54.785 46.155 ;
        RECT 55.305 45.525 55.585 45.985 ;
        RECT 54.460 45.305 55.585 45.525 ;
        RECT 52.485 43.605 52.995 44.140 ;
        RECT 53.215 43.810 53.460 44.415 ;
        RECT 53.905 44.345 54.185 45.015 ;
        RECT 54.460 44.845 54.910 45.305 ;
        RECT 55.775 45.135 56.175 45.985 ;
        RECT 56.575 45.695 56.845 46.155 ;
        RECT 57.015 45.525 57.300 45.985 ;
        RECT 57.585 45.720 62.930 46.155 ;
        RECT 63.105 45.720 68.450 46.155 ;
        RECT 54.355 44.515 54.910 44.845 ;
        RECT 55.080 44.575 56.175 45.135 ;
        RECT 54.460 44.405 54.910 44.515 ;
        RECT 53.905 43.775 54.290 44.345 ;
        RECT 54.460 44.235 55.585 44.405 ;
        RECT 54.460 43.605 54.785 44.065 ;
        RECT 55.305 43.775 55.585 44.235 ;
        RECT 55.775 43.775 56.175 44.575 ;
        RECT 56.345 45.305 57.300 45.525 ;
        RECT 56.345 44.405 56.555 45.305 ;
        RECT 56.725 44.575 57.415 45.135 ;
        RECT 56.345 44.235 57.300 44.405 ;
        RECT 56.575 43.605 56.845 44.065 ;
        RECT 57.015 43.775 57.300 44.235 ;
        RECT 59.170 44.150 59.510 44.980 ;
        RECT 60.990 44.470 61.340 45.720 ;
        RECT 64.690 44.150 65.030 44.980 ;
        RECT 66.510 44.470 66.860 45.720 ;
        RECT 68.625 45.065 69.835 46.155 ;
        RECT 68.625 44.355 69.145 44.895 ;
        RECT 69.315 44.525 69.835 45.065 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.465 45.065 73.055 46.155 ;
        RECT 73.690 45.485 73.945 45.985 ;
        RECT 74.115 45.655 74.445 46.155 ;
        RECT 73.690 45.315 74.440 45.485 ;
        RECT 70.465 44.375 71.675 44.895 ;
        RECT 71.845 44.545 73.055 45.065 ;
        RECT 73.690 44.495 74.040 45.145 ;
        RECT 57.585 43.605 62.930 44.150 ;
        RECT 63.105 43.605 68.450 44.150 ;
        RECT 68.625 43.605 69.835 44.355 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 70.465 43.605 73.055 44.375 ;
        RECT 74.210 44.325 74.440 45.315 ;
        RECT 73.690 44.155 74.440 44.325 ;
        RECT 73.690 43.865 73.945 44.155 ;
        RECT 74.115 43.605 74.445 43.985 ;
        RECT 74.615 43.865 74.785 45.985 ;
        RECT 74.955 45.185 75.280 45.970 ;
        RECT 75.450 45.695 75.700 46.155 ;
        RECT 75.870 45.655 76.120 45.985 ;
        RECT 76.335 45.655 77.015 45.985 ;
        RECT 75.870 45.525 76.040 45.655 ;
        RECT 75.645 45.355 76.040 45.525 ;
        RECT 75.015 44.135 75.475 45.185 ;
        RECT 75.645 43.995 75.815 45.355 ;
        RECT 76.210 45.095 76.675 45.485 ;
        RECT 75.985 44.285 76.335 44.905 ;
        RECT 76.505 44.505 76.675 45.095 ;
        RECT 76.845 44.875 77.015 45.655 ;
        RECT 77.185 45.555 77.355 45.895 ;
        RECT 77.590 45.725 77.920 46.155 ;
        RECT 78.090 45.555 78.260 45.895 ;
        RECT 78.555 45.695 78.925 46.155 ;
        RECT 77.185 45.385 78.260 45.555 ;
        RECT 79.095 45.525 79.265 45.985 ;
        RECT 79.500 45.645 80.370 45.985 ;
        RECT 80.540 45.695 80.790 46.155 ;
        RECT 78.705 45.355 79.265 45.525 ;
        RECT 78.705 45.215 78.875 45.355 ;
        RECT 77.375 45.045 78.875 45.215 ;
        RECT 79.570 45.185 80.030 45.475 ;
        RECT 76.845 44.705 78.535 44.875 ;
        RECT 76.505 44.285 76.860 44.505 ;
        RECT 77.030 43.995 77.200 44.705 ;
        RECT 77.405 44.285 78.195 44.535 ;
        RECT 78.365 44.525 78.535 44.705 ;
        RECT 78.705 44.355 78.875 45.045 ;
        RECT 75.145 43.605 75.475 43.965 ;
        RECT 75.645 43.825 76.140 43.995 ;
        RECT 76.345 43.825 77.200 43.995 ;
        RECT 78.075 43.605 78.405 44.065 ;
        RECT 78.615 43.965 78.875 44.355 ;
        RECT 79.065 45.175 80.030 45.185 ;
        RECT 80.200 45.265 80.370 45.645 ;
        RECT 80.960 45.605 81.130 45.895 ;
        RECT 81.310 45.775 81.640 46.155 ;
        RECT 80.960 45.435 81.760 45.605 ;
        RECT 79.065 45.015 79.740 45.175 ;
        RECT 80.200 45.095 81.420 45.265 ;
        RECT 79.065 44.225 79.275 45.015 ;
        RECT 80.200 45.005 80.370 45.095 ;
        RECT 79.445 44.225 79.795 44.845 ;
        RECT 79.965 44.835 80.370 45.005 ;
        RECT 79.965 44.055 80.135 44.835 ;
        RECT 80.305 44.385 80.525 44.665 ;
        RECT 80.705 44.555 81.245 44.925 ;
        RECT 81.590 44.845 81.760 45.435 ;
        RECT 81.980 45.015 82.285 46.155 ;
        RECT 82.455 44.965 82.710 45.845 ;
        RECT 81.590 44.815 82.330 44.845 ;
        RECT 80.305 44.215 80.835 44.385 ;
        RECT 78.615 43.795 78.965 43.965 ;
        RECT 79.185 43.775 80.135 44.055 ;
        RECT 80.305 43.605 80.495 44.045 ;
        RECT 80.665 43.985 80.835 44.215 ;
        RECT 81.005 44.155 81.245 44.555 ;
        RECT 81.415 44.515 82.330 44.815 ;
        RECT 81.415 44.340 81.740 44.515 ;
        RECT 81.415 43.985 81.735 44.340 ;
        RECT 82.500 44.315 82.710 44.965 ;
        RECT 80.665 43.815 81.735 43.985 ;
        RECT 81.980 43.605 82.285 44.065 ;
        RECT 82.455 43.785 82.710 44.315 ;
        RECT 82.885 45.015 83.270 45.985 ;
        RECT 83.440 45.695 83.765 46.155 ;
        RECT 84.285 45.525 84.565 45.985 ;
        RECT 83.440 45.305 84.565 45.525 ;
        RECT 82.885 44.345 83.165 45.015 ;
        RECT 83.440 44.845 83.890 45.305 ;
        RECT 84.755 45.135 85.155 45.985 ;
        RECT 85.555 45.695 85.825 46.155 ;
        RECT 85.995 45.525 86.280 45.985 ;
        RECT 83.335 44.515 83.890 44.845 ;
        RECT 84.060 44.575 85.155 45.135 ;
        RECT 83.440 44.405 83.890 44.515 ;
        RECT 82.885 43.775 83.270 44.345 ;
        RECT 83.440 44.235 84.565 44.405 ;
        RECT 83.440 43.605 83.765 44.065 ;
        RECT 84.285 43.775 84.565 44.235 ;
        RECT 84.755 43.775 85.155 44.575 ;
        RECT 85.325 45.305 86.280 45.525 ;
        RECT 85.325 44.405 85.535 45.305 ;
        RECT 85.705 44.575 86.395 45.135 ;
        RECT 86.565 45.015 86.905 45.985 ;
        RECT 87.075 45.015 87.245 46.155 ;
        RECT 87.515 45.355 87.765 46.155 ;
        RECT 88.410 45.185 88.740 45.985 ;
        RECT 89.040 45.355 89.370 46.155 ;
        RECT 89.540 45.185 89.870 45.985 ;
        RECT 87.435 45.015 89.870 45.185 ;
        RECT 90.245 45.015 90.630 45.985 ;
        RECT 90.800 45.695 91.125 46.155 ;
        RECT 91.645 45.525 91.925 45.985 ;
        RECT 90.800 45.305 91.925 45.525 ;
        RECT 86.565 44.405 86.740 45.015 ;
        RECT 87.435 44.765 87.605 45.015 ;
        RECT 86.910 44.595 87.605 44.765 ;
        RECT 87.780 44.595 88.200 44.795 ;
        RECT 88.370 44.595 88.700 44.795 ;
        RECT 88.870 44.595 89.200 44.795 ;
        RECT 85.325 44.235 86.280 44.405 ;
        RECT 85.555 43.605 85.825 44.065 ;
        RECT 85.995 43.775 86.280 44.235 ;
        RECT 86.565 43.775 86.905 44.405 ;
        RECT 87.075 43.605 87.325 44.405 ;
        RECT 87.515 44.255 88.740 44.425 ;
        RECT 87.515 43.775 87.845 44.255 ;
        RECT 88.015 43.605 88.240 44.065 ;
        RECT 88.410 43.775 88.740 44.255 ;
        RECT 89.370 44.385 89.540 45.015 ;
        RECT 89.725 44.595 90.075 44.845 ;
        RECT 89.370 43.775 89.870 44.385 ;
        RECT 90.245 44.345 90.525 45.015 ;
        RECT 90.800 44.845 91.250 45.305 ;
        RECT 92.115 45.135 92.515 45.985 ;
        RECT 92.915 45.695 93.185 46.155 ;
        RECT 93.355 45.525 93.640 45.985 ;
        RECT 90.695 44.515 91.250 44.845 ;
        RECT 91.420 44.575 92.515 45.135 ;
        RECT 90.800 44.405 91.250 44.515 ;
        RECT 90.245 43.775 90.630 44.345 ;
        RECT 90.800 44.235 91.925 44.405 ;
        RECT 90.800 43.605 91.125 44.065 ;
        RECT 91.645 43.775 91.925 44.235 ;
        RECT 92.115 43.775 92.515 44.575 ;
        RECT 92.685 45.305 93.640 45.525 ;
        RECT 92.685 44.405 92.895 45.305 ;
        RECT 93.065 44.575 93.755 45.135 ;
        RECT 93.925 45.065 95.595 46.155 ;
        RECT 92.685 44.235 93.640 44.405 ;
        RECT 92.915 43.605 93.185 44.065 ;
        RECT 93.355 43.775 93.640 44.235 ;
        RECT 93.925 44.375 94.675 44.895 ;
        RECT 94.845 44.545 95.595 45.065 ;
        RECT 95.765 44.990 96.055 46.155 ;
        RECT 96.225 45.720 101.570 46.155 ;
        RECT 93.925 43.605 95.595 44.375 ;
        RECT 95.765 43.605 96.055 44.330 ;
        RECT 97.810 44.150 98.150 44.980 ;
        RECT 99.630 44.470 99.980 45.720 ;
        RECT 101.745 45.065 103.415 46.155 ;
        RECT 101.745 44.375 102.495 44.895 ;
        RECT 102.665 44.545 103.415 45.065 ;
        RECT 103.585 45.395 104.100 45.805 ;
        RECT 104.335 45.395 104.505 46.155 ;
        RECT 104.675 45.815 106.705 45.985 ;
        RECT 103.585 44.585 103.925 45.395 ;
        RECT 104.675 45.150 104.845 45.815 ;
        RECT 105.240 45.475 106.365 45.645 ;
        RECT 104.095 44.960 104.845 45.150 ;
        RECT 105.015 45.135 106.025 45.305 ;
        RECT 103.585 44.415 104.815 44.585 ;
        RECT 96.225 43.605 101.570 44.150 ;
        RECT 101.745 43.605 103.415 44.375 ;
        RECT 103.860 43.810 104.105 44.415 ;
        RECT 104.325 43.605 104.835 44.140 ;
        RECT 105.015 43.775 105.205 45.135 ;
        RECT 105.375 44.795 105.650 44.935 ;
        RECT 105.375 44.625 105.655 44.795 ;
        RECT 105.375 43.775 105.650 44.625 ;
        RECT 105.855 44.335 106.025 45.135 ;
        RECT 106.195 44.345 106.365 45.475 ;
        RECT 106.535 44.845 106.705 45.815 ;
        RECT 106.875 45.015 107.045 46.155 ;
        RECT 107.215 45.015 107.550 45.985 ;
        RECT 106.535 44.515 106.730 44.845 ;
        RECT 106.955 44.515 107.210 44.845 ;
        RECT 106.955 44.345 107.125 44.515 ;
        RECT 107.380 44.345 107.550 45.015 ;
        RECT 106.195 44.175 107.125 44.345 ;
        RECT 106.195 44.140 106.370 44.175 ;
        RECT 105.840 43.775 106.370 44.140 ;
        RECT 106.795 43.605 107.125 44.005 ;
        RECT 107.295 43.775 107.550 44.345 ;
        RECT 107.725 45.015 108.110 45.985 ;
        RECT 108.280 45.695 108.605 46.155 ;
        RECT 109.125 45.525 109.405 45.985 ;
        RECT 108.280 45.305 109.405 45.525 ;
        RECT 107.725 44.345 108.005 45.015 ;
        RECT 108.280 44.845 108.730 45.305 ;
        RECT 109.595 45.135 109.995 45.985 ;
        RECT 110.395 45.695 110.665 46.155 ;
        RECT 110.835 45.525 111.120 45.985 ;
        RECT 108.175 44.515 108.730 44.845 ;
        RECT 108.900 44.575 109.995 45.135 ;
        RECT 108.280 44.405 108.730 44.515 ;
        RECT 107.725 43.775 108.110 44.345 ;
        RECT 108.280 44.235 109.405 44.405 ;
        RECT 108.280 43.605 108.605 44.065 ;
        RECT 109.125 43.775 109.405 44.235 ;
        RECT 109.595 43.775 109.995 44.575 ;
        RECT 110.165 45.305 111.120 45.525 ;
        RECT 110.165 44.405 110.375 45.305 ;
        RECT 110.545 44.575 111.235 45.135 ;
        RECT 111.445 45.015 111.675 46.155 ;
        RECT 111.845 45.005 112.175 45.985 ;
        RECT 112.345 45.015 112.555 46.155 ;
        RECT 112.785 45.720 118.130 46.155 ;
        RECT 111.425 44.595 111.755 44.845 ;
        RECT 110.165 44.235 111.120 44.405 ;
        RECT 110.395 43.605 110.665 44.065 ;
        RECT 110.835 43.775 111.120 44.235 ;
        RECT 111.445 43.605 111.675 44.425 ;
        RECT 111.925 44.405 112.175 45.005 ;
        RECT 111.845 43.775 112.175 44.405 ;
        RECT 112.345 43.605 112.555 44.425 ;
        RECT 114.370 44.150 114.710 44.980 ;
        RECT 116.190 44.470 116.540 45.720 ;
        RECT 118.305 45.065 120.895 46.155 ;
        RECT 118.305 44.375 119.515 44.895 ;
        RECT 119.685 44.545 120.895 45.065 ;
        RECT 121.525 44.990 121.815 46.155 ;
        RECT 121.985 45.065 123.655 46.155 ;
        RECT 121.985 44.375 122.735 44.895 ;
        RECT 122.905 44.545 123.655 45.065 ;
        RECT 124.285 45.065 125.495 46.155 ;
        RECT 124.285 44.525 124.805 45.065 ;
        RECT 112.785 43.605 118.130 44.150 ;
        RECT 118.305 43.605 120.895 44.375 ;
        RECT 121.525 43.605 121.815 44.330 ;
        RECT 121.985 43.605 123.655 44.375 ;
        RECT 124.975 44.355 125.495 44.895 ;
        RECT 124.285 43.605 125.495 44.355 ;
        RECT 5.520 43.435 125.580 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 6.985 42.890 12.330 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 8.570 42.060 8.910 42.890 ;
        RECT 12.505 42.665 16.015 43.435 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 10.390 41.320 10.740 42.570 ;
        RECT 12.505 42.145 14.155 42.665 ;
        RECT 17.165 42.615 17.375 43.435 ;
        RECT 17.545 42.635 17.875 43.265 ;
        RECT 14.325 41.975 16.015 42.495 ;
        RECT 17.545 42.035 17.795 42.635 ;
        RECT 18.045 42.615 18.275 43.435 ;
        RECT 18.545 42.615 18.755 43.435 ;
        RECT 18.925 42.635 19.255 43.265 ;
        RECT 17.965 42.195 18.295 42.445 ;
        RECT 18.925 42.035 19.175 42.635 ;
        RECT 19.425 42.615 19.655 43.435 ;
        RECT 20.900 42.805 21.185 43.265 ;
        RECT 21.355 42.975 21.625 43.435 ;
        RECT 20.900 42.635 21.855 42.805 ;
        RECT 19.345 42.195 19.675 42.445 ;
        RECT 6.985 40.885 12.330 41.320 ;
        RECT 12.505 40.885 16.015 41.975 ;
        RECT 17.165 40.885 17.375 42.025 ;
        RECT 17.545 41.055 17.875 42.035 ;
        RECT 18.045 40.885 18.275 42.025 ;
        RECT 18.545 40.885 18.755 42.025 ;
        RECT 18.925 41.055 19.255 42.035 ;
        RECT 19.425 40.885 19.655 42.025 ;
        RECT 20.785 41.905 21.475 42.465 ;
        RECT 21.645 41.735 21.855 42.635 ;
        RECT 20.900 41.515 21.855 41.735 ;
        RECT 22.025 42.465 22.425 43.265 ;
        RECT 22.615 42.805 22.895 43.265 ;
        RECT 23.415 42.975 23.740 43.435 ;
        RECT 22.615 42.635 23.740 42.805 ;
        RECT 23.910 42.695 24.295 43.265 ;
        RECT 23.290 42.525 23.740 42.635 ;
        RECT 22.025 41.905 23.120 42.465 ;
        RECT 23.290 42.195 23.845 42.525 ;
        RECT 20.900 41.055 21.185 41.515 ;
        RECT 21.355 40.885 21.625 41.345 ;
        RECT 22.025 41.055 22.425 41.905 ;
        RECT 23.290 41.735 23.740 42.195 ;
        RECT 24.015 42.025 24.295 42.695 ;
        RECT 22.615 41.515 23.740 41.735 ;
        RECT 22.615 41.055 22.895 41.515 ;
        RECT 23.415 40.885 23.740 41.345 ;
        RECT 23.910 41.055 24.295 42.025 ;
        RECT 24.465 42.695 24.850 43.265 ;
        RECT 25.020 42.975 25.345 43.435 ;
        RECT 25.865 42.805 26.145 43.265 ;
        RECT 24.465 42.025 24.745 42.695 ;
        RECT 25.020 42.635 26.145 42.805 ;
        RECT 25.020 42.525 25.470 42.635 ;
        RECT 24.915 42.195 25.470 42.525 ;
        RECT 26.335 42.465 26.735 43.265 ;
        RECT 27.135 42.975 27.405 43.435 ;
        RECT 27.575 42.805 27.860 43.265 ;
        RECT 24.465 41.055 24.850 42.025 ;
        RECT 25.020 41.735 25.470 42.195 ;
        RECT 25.640 41.905 26.735 42.465 ;
        RECT 25.020 41.515 26.145 41.735 ;
        RECT 25.020 40.885 25.345 41.345 ;
        RECT 25.865 41.055 26.145 41.515 ;
        RECT 26.335 41.055 26.735 41.905 ;
        RECT 26.905 42.635 27.860 42.805 ;
        RECT 28.145 42.665 30.735 43.435 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 26.905 41.735 27.115 42.635 ;
        RECT 27.285 41.905 27.975 42.465 ;
        RECT 28.145 42.145 29.355 42.665 ;
        RECT 31.885 42.615 32.095 43.435 ;
        RECT 32.265 42.635 32.595 43.265 ;
        RECT 29.525 41.975 30.735 42.495 ;
        RECT 26.905 41.515 27.860 41.735 ;
        RECT 27.135 40.885 27.405 41.345 ;
        RECT 27.575 41.055 27.860 41.515 ;
        RECT 28.145 40.885 30.735 41.975 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 32.265 42.035 32.515 42.635 ;
        RECT 32.765 42.615 32.995 43.435 ;
        RECT 33.205 42.665 34.875 43.435 ;
        RECT 35.045 42.760 35.305 43.265 ;
        RECT 35.485 43.055 35.815 43.435 ;
        RECT 35.995 42.885 36.165 43.265 ;
        RECT 36.425 42.890 41.770 43.435 ;
        RECT 32.685 42.195 33.015 42.445 ;
        RECT 33.205 42.145 33.955 42.665 ;
        RECT 31.885 40.885 32.095 42.025 ;
        RECT 32.265 41.055 32.595 42.035 ;
        RECT 32.765 40.885 32.995 42.025 ;
        RECT 34.125 41.975 34.875 42.495 ;
        RECT 33.205 40.885 34.875 41.975 ;
        RECT 35.045 41.960 35.215 42.760 ;
        RECT 35.500 42.715 36.165 42.885 ;
        RECT 35.500 42.460 35.670 42.715 ;
        RECT 35.385 42.130 35.670 42.460 ;
        RECT 35.905 42.165 36.235 42.535 ;
        RECT 35.500 41.985 35.670 42.130 ;
        RECT 38.010 42.060 38.350 42.890 ;
        RECT 41.945 42.665 43.615 43.435 ;
        RECT 43.875 42.885 44.045 43.265 ;
        RECT 44.225 43.055 44.555 43.435 ;
        RECT 43.875 42.715 44.540 42.885 ;
        RECT 44.735 42.760 44.995 43.265 ;
        RECT 35.045 41.055 35.315 41.960 ;
        RECT 35.500 41.815 36.165 41.985 ;
        RECT 35.485 40.885 35.815 41.645 ;
        RECT 35.995 41.055 36.165 41.815 ;
        RECT 39.830 41.320 40.180 42.570 ;
        RECT 41.945 42.145 42.695 42.665 ;
        RECT 42.865 41.975 43.615 42.495 ;
        RECT 43.805 42.165 44.135 42.535 ;
        RECT 44.370 42.460 44.540 42.715 ;
        RECT 44.370 42.130 44.655 42.460 ;
        RECT 44.370 41.985 44.540 42.130 ;
        RECT 36.425 40.885 41.770 41.320 ;
        RECT 41.945 40.885 43.615 41.975 ;
        RECT 43.875 41.815 44.540 41.985 ;
        RECT 44.825 41.960 44.995 42.760 ;
        RECT 46.125 42.615 46.355 43.435 ;
        RECT 46.525 42.635 46.855 43.265 ;
        RECT 46.105 42.195 46.435 42.445 ;
        RECT 46.605 42.035 46.855 42.635 ;
        RECT 47.025 42.615 47.235 43.435 ;
        RECT 47.465 42.890 52.810 43.435 ;
        RECT 49.050 42.060 49.390 42.890 ;
        RECT 52.985 42.665 56.495 43.435 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 57.585 42.665 61.095 43.435 ;
        RECT 61.725 42.935 61.985 43.265 ;
        RECT 62.295 43.055 62.625 43.435 ;
        RECT 62.805 43.095 64.285 43.265 ;
        RECT 43.875 41.055 44.045 41.815 ;
        RECT 44.225 40.885 44.555 41.645 ;
        RECT 44.725 41.055 44.995 41.960 ;
        RECT 46.125 40.885 46.355 42.025 ;
        RECT 46.525 41.055 46.855 42.035 ;
        RECT 47.025 40.885 47.235 42.025 ;
        RECT 50.870 41.320 51.220 42.570 ;
        RECT 52.985 42.145 54.635 42.665 ;
        RECT 54.805 41.975 56.495 42.495 ;
        RECT 57.585 42.145 59.235 42.665 ;
        RECT 47.465 40.885 52.810 41.320 ;
        RECT 52.985 40.885 56.495 41.975 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 59.405 41.975 61.095 42.495 ;
        RECT 57.585 40.885 61.095 41.975 ;
        RECT 61.725 42.235 61.895 42.935 ;
        RECT 62.805 42.765 63.205 43.095 ;
        RECT 62.245 42.575 62.455 42.755 ;
        RECT 62.245 42.405 62.865 42.575 ;
        RECT 63.035 42.285 63.205 42.765 ;
        RECT 63.395 42.595 63.945 42.925 ;
        RECT 61.725 42.065 62.855 42.235 ;
        RECT 63.035 42.115 63.605 42.285 ;
        RECT 61.725 41.385 61.895 42.065 ;
        RECT 62.685 41.945 62.855 42.065 ;
        RECT 62.065 41.565 62.415 41.895 ;
        RECT 62.685 41.775 63.265 41.945 ;
        RECT 63.435 41.605 63.605 42.115 ;
        RECT 62.865 41.435 63.605 41.605 ;
        RECT 63.775 41.605 63.945 42.595 ;
        RECT 64.115 42.195 64.285 43.095 ;
        RECT 64.535 42.525 64.720 43.105 ;
        RECT 64.990 42.525 65.185 43.100 ;
        RECT 65.395 43.055 65.725 43.435 ;
        RECT 64.535 42.195 64.765 42.525 ;
        RECT 64.990 42.195 65.245 42.525 ;
        RECT 64.535 41.885 64.720 42.195 ;
        RECT 64.990 41.885 65.185 42.195 ;
        RECT 65.555 41.605 65.725 42.525 ;
        RECT 63.775 41.435 65.725 41.605 ;
        RECT 61.725 41.055 61.985 41.385 ;
        RECT 62.295 40.885 62.625 41.265 ;
        RECT 62.865 41.055 63.055 41.435 ;
        RECT 63.305 40.885 63.635 41.265 ;
        RECT 63.845 41.055 64.015 41.435 ;
        RECT 64.210 40.885 64.540 41.265 ;
        RECT 64.800 41.055 64.970 41.435 ;
        RECT 65.395 40.885 65.725 41.265 ;
        RECT 65.895 41.055 66.155 43.265 ;
        RECT 66.385 42.615 66.595 43.435 ;
        RECT 66.765 42.635 67.095 43.265 ;
        RECT 66.765 42.035 67.015 42.635 ;
        RECT 67.265 42.615 67.495 43.435 ;
        RECT 67.705 42.890 73.050 43.435 ;
        RECT 67.185 42.195 67.515 42.445 ;
        RECT 69.290 42.060 69.630 42.890 ;
        RECT 73.225 42.665 76.735 43.435 ;
        RECT 76.905 42.685 78.115 43.435 ;
        RECT 66.385 40.885 66.595 42.025 ;
        RECT 66.765 41.055 67.095 42.035 ;
        RECT 67.265 40.885 67.495 42.025 ;
        RECT 71.110 41.320 71.460 42.570 ;
        RECT 73.225 42.145 74.875 42.665 ;
        RECT 75.045 41.975 76.735 42.495 ;
        RECT 76.905 42.145 77.425 42.685 ;
        RECT 78.325 42.615 78.555 43.435 ;
        RECT 78.725 42.635 79.055 43.265 ;
        RECT 77.595 41.975 78.115 42.515 ;
        RECT 78.305 42.195 78.635 42.445 ;
        RECT 78.805 42.035 79.055 42.635 ;
        RECT 79.225 42.615 79.435 43.435 ;
        RECT 79.665 42.665 82.255 43.435 ;
        RECT 82.885 42.710 83.175 43.435 ;
        RECT 83.350 42.695 83.605 43.265 ;
        RECT 83.775 43.035 84.105 43.435 ;
        RECT 84.530 42.900 85.060 43.265 ;
        RECT 84.530 42.865 84.705 42.900 ;
        RECT 83.775 42.695 84.705 42.865 ;
        RECT 79.665 42.145 80.875 42.665 ;
        RECT 67.705 40.885 73.050 41.320 ;
        RECT 73.225 40.885 76.735 41.975 ;
        RECT 76.905 40.885 78.115 41.975 ;
        RECT 78.325 40.885 78.555 42.025 ;
        RECT 78.725 41.055 79.055 42.035 ;
        RECT 79.225 40.885 79.435 42.025 ;
        RECT 81.045 41.975 82.255 42.495 ;
        RECT 79.665 40.885 82.255 41.975 ;
        RECT 82.885 40.885 83.175 42.050 ;
        RECT 83.350 42.025 83.520 42.695 ;
        RECT 83.775 42.525 83.945 42.695 ;
        RECT 83.690 42.195 83.945 42.525 ;
        RECT 84.170 42.195 84.365 42.525 ;
        RECT 83.350 41.055 83.685 42.025 ;
        RECT 83.855 40.885 84.025 42.025 ;
        RECT 84.195 41.225 84.365 42.195 ;
        RECT 84.535 41.565 84.705 42.695 ;
        RECT 84.875 41.905 85.045 42.705 ;
        RECT 85.250 42.415 85.525 43.265 ;
        RECT 85.245 42.245 85.525 42.415 ;
        RECT 85.250 42.105 85.525 42.245 ;
        RECT 85.695 41.905 85.885 43.265 ;
        RECT 86.065 42.900 86.575 43.435 ;
        RECT 86.795 42.625 87.040 43.230 ;
        RECT 87.485 42.695 87.870 43.265 ;
        RECT 88.040 42.975 88.365 43.435 ;
        RECT 88.885 42.805 89.165 43.265 ;
        RECT 86.085 42.455 87.315 42.625 ;
        RECT 84.875 41.735 85.885 41.905 ;
        RECT 86.055 41.890 86.805 42.080 ;
        RECT 84.535 41.395 85.660 41.565 ;
        RECT 86.055 41.225 86.225 41.890 ;
        RECT 86.975 41.645 87.315 42.455 ;
        RECT 84.195 41.055 86.225 41.225 ;
        RECT 86.395 40.885 86.565 41.645 ;
        RECT 86.800 41.235 87.315 41.645 ;
        RECT 87.485 42.025 87.765 42.695 ;
        RECT 88.040 42.635 89.165 42.805 ;
        RECT 88.040 42.525 88.490 42.635 ;
        RECT 87.935 42.195 88.490 42.525 ;
        RECT 89.355 42.465 89.755 43.265 ;
        RECT 90.155 42.975 90.425 43.435 ;
        RECT 90.595 42.805 90.880 43.265 ;
        RECT 87.485 41.055 87.870 42.025 ;
        RECT 88.040 41.735 88.490 42.195 ;
        RECT 88.660 41.905 89.755 42.465 ;
        RECT 88.040 41.515 89.165 41.735 ;
        RECT 88.040 40.885 88.365 41.345 ;
        RECT 88.885 41.055 89.165 41.515 ;
        RECT 89.355 41.055 89.755 41.905 ;
        RECT 89.925 42.635 90.880 42.805 ;
        RECT 89.925 41.735 90.135 42.635 ;
        RECT 91.205 42.615 91.435 43.435 ;
        RECT 91.605 42.635 91.935 43.265 ;
        RECT 90.305 41.905 90.995 42.465 ;
        RECT 91.185 42.195 91.515 42.445 ;
        RECT 91.685 42.035 91.935 42.635 ;
        RECT 92.105 42.615 92.315 43.435 ;
        RECT 92.545 42.695 92.930 43.265 ;
        RECT 93.100 42.975 93.425 43.435 ;
        RECT 93.945 42.805 94.225 43.265 ;
        RECT 89.925 41.515 90.880 41.735 ;
        RECT 90.155 40.885 90.425 41.345 ;
        RECT 90.595 41.055 90.880 41.515 ;
        RECT 91.205 40.885 91.435 42.025 ;
        RECT 91.605 41.055 91.935 42.035 ;
        RECT 92.545 42.025 92.825 42.695 ;
        RECT 93.100 42.635 94.225 42.805 ;
        RECT 93.100 42.525 93.550 42.635 ;
        RECT 92.995 42.195 93.550 42.525 ;
        RECT 94.415 42.465 94.815 43.265 ;
        RECT 95.215 42.975 95.485 43.435 ;
        RECT 95.655 42.805 95.940 43.265 ;
        RECT 92.105 40.885 92.315 42.025 ;
        RECT 92.545 41.055 92.930 42.025 ;
        RECT 93.100 41.735 93.550 42.195 ;
        RECT 93.720 41.905 94.815 42.465 ;
        RECT 93.100 41.515 94.225 41.735 ;
        RECT 93.100 40.885 93.425 41.345 ;
        RECT 93.945 41.055 94.225 41.515 ;
        RECT 94.415 41.055 94.815 41.905 ;
        RECT 94.985 42.635 95.940 42.805 ;
        RECT 96.230 42.695 96.485 43.265 ;
        RECT 96.655 43.035 96.985 43.435 ;
        RECT 97.410 42.900 97.940 43.265 ;
        RECT 98.130 43.095 98.405 43.265 ;
        RECT 98.125 42.925 98.405 43.095 ;
        RECT 97.410 42.865 97.585 42.900 ;
        RECT 96.655 42.695 97.585 42.865 ;
        RECT 94.985 41.735 95.195 42.635 ;
        RECT 95.365 41.905 96.055 42.465 ;
        RECT 96.230 42.025 96.400 42.695 ;
        RECT 96.655 42.525 96.825 42.695 ;
        RECT 96.570 42.195 96.825 42.525 ;
        RECT 97.050 42.195 97.245 42.525 ;
        RECT 94.985 41.515 95.940 41.735 ;
        RECT 95.215 40.885 95.485 41.345 ;
        RECT 95.655 41.055 95.940 41.515 ;
        RECT 96.230 41.055 96.565 42.025 ;
        RECT 96.735 40.885 96.905 42.025 ;
        RECT 97.075 41.225 97.245 42.195 ;
        RECT 97.415 41.565 97.585 42.695 ;
        RECT 97.755 41.905 97.925 42.705 ;
        RECT 98.130 42.105 98.405 42.925 ;
        RECT 98.575 41.905 98.765 43.265 ;
        RECT 98.945 42.900 99.455 43.435 ;
        RECT 99.675 42.625 99.920 43.230 ;
        RECT 100.830 42.695 101.085 43.265 ;
        RECT 101.255 43.035 101.585 43.435 ;
        RECT 102.010 42.900 102.540 43.265 ;
        RECT 102.010 42.865 102.185 42.900 ;
        RECT 101.255 42.695 102.185 42.865 ;
        RECT 102.730 42.755 103.005 43.265 ;
        RECT 98.965 42.455 100.195 42.625 ;
        RECT 97.755 41.735 98.765 41.905 ;
        RECT 98.935 41.890 99.685 42.080 ;
        RECT 97.415 41.395 98.540 41.565 ;
        RECT 98.935 41.225 99.105 41.890 ;
        RECT 99.855 41.645 100.195 42.455 ;
        RECT 97.075 41.055 99.105 41.225 ;
        RECT 99.275 40.885 99.445 41.645 ;
        RECT 99.680 41.235 100.195 41.645 ;
        RECT 100.830 42.025 101.000 42.695 ;
        RECT 101.255 42.525 101.425 42.695 ;
        RECT 101.170 42.195 101.425 42.525 ;
        RECT 101.650 42.195 101.845 42.525 ;
        RECT 100.830 41.055 101.165 42.025 ;
        RECT 101.335 40.885 101.505 42.025 ;
        RECT 101.675 41.225 101.845 42.195 ;
        RECT 102.015 41.565 102.185 42.695 ;
        RECT 102.355 41.905 102.525 42.705 ;
        RECT 102.725 42.585 103.005 42.755 ;
        RECT 102.730 42.105 103.005 42.585 ;
        RECT 103.175 41.905 103.365 43.265 ;
        RECT 103.545 42.900 104.055 43.435 ;
        RECT 104.275 42.625 104.520 43.230 ;
        RECT 105.055 42.885 105.225 43.265 ;
        RECT 105.405 43.055 105.735 43.435 ;
        RECT 105.055 42.715 105.720 42.885 ;
        RECT 105.915 42.760 106.175 43.265 ;
        RECT 103.565 42.455 104.795 42.625 ;
        RECT 102.355 41.735 103.365 41.905 ;
        RECT 103.535 41.890 104.285 42.080 ;
        RECT 102.015 41.395 103.140 41.565 ;
        RECT 103.535 41.225 103.705 41.890 ;
        RECT 104.455 41.645 104.795 42.455 ;
        RECT 104.985 42.165 105.315 42.535 ;
        RECT 105.550 42.460 105.720 42.715 ;
        RECT 105.550 42.130 105.835 42.460 ;
        RECT 105.550 41.985 105.720 42.130 ;
        RECT 101.675 41.055 103.705 41.225 ;
        RECT 103.875 40.885 104.045 41.645 ;
        RECT 104.280 41.235 104.795 41.645 ;
        RECT 105.055 41.815 105.720 41.985 ;
        RECT 106.005 41.960 106.175 42.760 ;
        RECT 106.345 42.665 108.015 43.435 ;
        RECT 108.645 42.710 108.935 43.435 ;
        RECT 109.105 42.695 109.490 43.265 ;
        RECT 109.660 42.975 109.985 43.435 ;
        RECT 110.505 42.805 110.785 43.265 ;
        RECT 106.345 42.145 107.095 42.665 ;
        RECT 107.265 41.975 108.015 42.495 ;
        RECT 105.055 41.055 105.225 41.815 ;
        RECT 105.405 40.885 105.735 41.645 ;
        RECT 105.905 41.055 106.175 41.960 ;
        RECT 106.345 40.885 108.015 41.975 ;
        RECT 108.645 40.885 108.935 42.050 ;
        RECT 109.105 42.025 109.385 42.695 ;
        RECT 109.660 42.635 110.785 42.805 ;
        RECT 109.660 42.525 110.110 42.635 ;
        RECT 109.555 42.195 110.110 42.525 ;
        RECT 110.975 42.465 111.375 43.265 ;
        RECT 111.775 42.975 112.045 43.435 ;
        RECT 112.215 42.805 112.500 43.265 ;
        RECT 109.105 41.055 109.490 42.025 ;
        RECT 109.660 41.735 110.110 42.195 ;
        RECT 110.280 41.905 111.375 42.465 ;
        RECT 109.660 41.515 110.785 41.735 ;
        RECT 109.660 40.885 109.985 41.345 ;
        RECT 110.505 41.055 110.785 41.515 ;
        RECT 110.975 41.055 111.375 41.905 ;
        RECT 111.545 42.635 112.500 42.805 ;
        RECT 111.545 41.735 111.755 42.635 ;
        RECT 112.825 42.615 113.055 43.435 ;
        RECT 113.225 42.635 113.555 43.265 ;
        RECT 111.925 41.905 112.615 42.465 ;
        RECT 112.805 42.195 113.135 42.445 ;
        RECT 113.305 42.035 113.555 42.635 ;
        RECT 113.725 42.615 113.935 43.435 ;
        RECT 114.165 42.890 119.510 43.435 ;
        RECT 115.750 42.060 116.090 42.890 ;
        RECT 119.685 42.665 123.195 43.435 ;
        RECT 124.285 42.685 125.495 43.435 ;
        RECT 111.545 41.515 112.500 41.735 ;
        RECT 111.775 40.885 112.045 41.345 ;
        RECT 112.215 41.055 112.500 41.515 ;
        RECT 112.825 40.885 113.055 42.025 ;
        RECT 113.225 41.055 113.555 42.035 ;
        RECT 113.725 40.885 113.935 42.025 ;
        RECT 117.570 41.320 117.920 42.570 ;
        RECT 119.685 42.145 121.335 42.665 ;
        RECT 121.505 41.975 123.195 42.495 ;
        RECT 114.165 40.885 119.510 41.320 ;
        RECT 119.685 40.885 123.195 41.975 ;
        RECT 124.285 41.975 124.805 42.515 ;
        RECT 124.975 42.145 125.495 42.685 ;
        RECT 124.285 40.885 125.495 41.975 ;
        RECT 5.520 40.715 125.580 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 6.985 40.280 12.330 40.715 ;
        RECT 12.505 40.280 17.850 40.715 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 8.570 38.710 8.910 39.540 ;
        RECT 10.390 39.030 10.740 40.280 ;
        RECT 14.090 38.710 14.430 39.540 ;
        RECT 15.910 39.030 16.260 40.280 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.945 40.280 24.290 40.715 ;
        RECT 24.465 40.280 29.810 40.715 ;
        RECT 6.985 38.165 12.330 38.710 ;
        RECT 12.505 38.165 17.850 38.710 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 20.530 38.710 20.870 39.540 ;
        RECT 22.350 39.030 22.700 40.280 ;
        RECT 26.050 38.710 26.390 39.540 ;
        RECT 27.870 39.030 28.220 40.280 ;
        RECT 31.020 40.085 31.305 40.545 ;
        RECT 31.475 40.255 31.745 40.715 ;
        RECT 31.020 39.865 31.975 40.085 ;
        RECT 30.905 39.135 31.595 39.695 ;
        RECT 31.765 38.965 31.975 39.865 ;
        RECT 31.020 38.795 31.975 38.965 ;
        RECT 32.145 39.695 32.545 40.545 ;
        RECT 32.735 40.085 33.015 40.545 ;
        RECT 33.535 40.255 33.860 40.715 ;
        RECT 32.735 39.865 33.860 40.085 ;
        RECT 32.145 39.135 33.240 39.695 ;
        RECT 33.410 39.405 33.860 39.865 ;
        RECT 34.030 39.575 34.415 40.545 ;
        RECT 34.585 39.625 38.095 40.715 ;
        RECT 38.265 39.625 39.475 40.715 ;
        RECT 18.945 38.165 24.290 38.710 ;
        RECT 24.465 38.165 29.810 38.710 ;
        RECT 31.020 38.335 31.305 38.795 ;
        RECT 31.475 38.165 31.745 38.625 ;
        RECT 32.145 38.335 32.545 39.135 ;
        RECT 33.410 39.075 33.965 39.405 ;
        RECT 33.410 38.965 33.860 39.075 ;
        RECT 32.735 38.795 33.860 38.965 ;
        RECT 34.135 38.905 34.415 39.575 ;
        RECT 32.735 38.335 33.015 38.795 ;
        RECT 33.535 38.165 33.860 38.625 ;
        RECT 34.030 38.335 34.415 38.905 ;
        RECT 34.585 38.935 36.235 39.455 ;
        RECT 36.405 39.105 38.095 39.625 ;
        RECT 34.585 38.165 38.095 38.935 ;
        RECT 38.265 38.915 38.785 39.455 ;
        RECT 38.955 39.085 39.475 39.625 ;
        RECT 39.645 39.640 39.915 40.545 ;
        RECT 40.085 39.955 40.415 40.715 ;
        RECT 40.595 39.785 40.765 40.545 ;
        RECT 38.265 38.165 39.475 38.915 ;
        RECT 39.645 38.840 39.815 39.640 ;
        RECT 40.100 39.615 40.765 39.785 ;
        RECT 41.025 39.625 43.615 40.715 ;
        RECT 40.100 39.470 40.270 39.615 ;
        RECT 39.985 39.140 40.270 39.470 ;
        RECT 40.100 38.885 40.270 39.140 ;
        RECT 40.505 39.065 40.835 39.435 ;
        RECT 41.025 38.935 42.235 39.455 ;
        RECT 42.405 39.105 43.615 39.625 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.795 40.045 44.965 40.545 ;
        RECT 45.135 40.215 45.465 40.715 ;
        RECT 44.795 39.875 45.460 40.045 ;
        RECT 44.710 39.055 45.060 39.705 ;
        RECT 39.645 38.335 39.905 38.840 ;
        RECT 40.100 38.715 40.765 38.885 ;
        RECT 40.085 38.165 40.415 38.545 ;
        RECT 40.595 38.335 40.765 38.715 ;
        RECT 41.025 38.165 43.615 38.935 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 45.230 38.885 45.460 39.875 ;
        RECT 44.795 38.715 45.460 38.885 ;
        RECT 44.795 38.425 44.965 38.715 ;
        RECT 45.135 38.165 45.465 38.545 ;
        RECT 45.635 38.425 45.860 40.545 ;
        RECT 46.075 40.215 46.405 40.715 ;
        RECT 46.575 40.045 46.745 40.545 ;
        RECT 46.980 40.330 47.810 40.500 ;
        RECT 48.050 40.335 48.430 40.715 ;
        RECT 46.050 39.875 46.745 40.045 ;
        RECT 46.050 38.905 46.220 39.875 ;
        RECT 46.390 39.085 46.800 39.705 ;
        RECT 46.970 39.655 47.470 40.035 ;
        RECT 46.050 38.715 46.745 38.905 ;
        RECT 46.970 38.785 47.190 39.655 ;
        RECT 47.640 39.485 47.810 40.330 ;
        RECT 48.610 40.165 48.780 40.455 ;
        RECT 48.950 40.335 49.280 40.715 ;
        RECT 49.750 40.245 50.380 40.495 ;
        RECT 50.560 40.335 50.980 40.715 ;
        RECT 50.210 40.165 50.380 40.245 ;
        RECT 51.180 40.165 51.420 40.455 ;
        RECT 47.980 39.915 49.350 40.165 ;
        RECT 47.980 39.655 48.230 39.915 ;
        RECT 48.740 39.485 48.990 39.645 ;
        RECT 47.640 39.315 48.990 39.485 ;
        RECT 47.640 39.275 48.060 39.315 ;
        RECT 47.370 38.725 47.720 39.095 ;
        RECT 46.075 38.165 46.405 38.545 ;
        RECT 46.575 38.385 46.745 38.715 ;
        RECT 47.890 38.545 48.060 39.275 ;
        RECT 49.160 39.145 49.350 39.915 ;
        RECT 48.230 38.815 48.640 39.145 ;
        RECT 48.930 38.805 49.350 39.145 ;
        RECT 49.520 39.735 50.040 40.045 ;
        RECT 50.210 39.995 51.420 40.165 ;
        RECT 51.650 40.025 51.980 40.715 ;
        RECT 49.520 38.975 49.690 39.735 ;
        RECT 49.860 39.145 50.040 39.555 ;
        RECT 50.210 39.485 50.380 39.995 ;
        RECT 52.150 39.845 52.320 40.455 ;
        RECT 52.590 39.995 52.920 40.505 ;
        RECT 52.150 39.825 52.470 39.845 ;
        RECT 50.550 39.655 52.470 39.825 ;
        RECT 50.210 39.315 52.110 39.485 ;
        RECT 50.440 38.975 50.770 39.095 ;
        RECT 49.520 38.805 50.770 38.975 ;
        RECT 47.045 38.345 48.060 38.545 ;
        RECT 48.230 38.165 48.640 38.605 ;
        RECT 48.930 38.375 49.180 38.805 ;
        RECT 49.380 38.165 49.700 38.625 ;
        RECT 50.940 38.555 51.110 39.315 ;
        RECT 51.780 39.255 52.110 39.315 ;
        RECT 51.300 39.085 51.630 39.145 ;
        RECT 51.300 38.815 51.960 39.085 ;
        RECT 52.280 38.760 52.470 39.655 ;
        RECT 50.260 38.385 51.110 38.555 ;
        RECT 51.310 38.165 51.970 38.645 ;
        RECT 52.150 38.430 52.470 38.760 ;
        RECT 52.670 39.405 52.920 39.995 ;
        RECT 53.100 39.915 53.385 40.715 ;
        RECT 53.565 40.375 53.820 40.405 ;
        RECT 53.565 40.205 53.905 40.375 ;
        RECT 53.565 39.735 53.820 40.205 ;
        RECT 52.670 39.075 53.470 39.405 ;
        RECT 52.670 38.425 52.920 39.075 ;
        RECT 53.640 38.875 53.820 39.735 ;
        RECT 54.365 39.625 57.875 40.715 ;
        RECT 58.050 40.045 58.305 40.545 ;
        RECT 58.475 40.215 58.805 40.715 ;
        RECT 58.050 39.875 58.800 40.045 ;
        RECT 53.100 38.165 53.385 38.625 ;
        RECT 53.565 38.345 53.820 38.875 ;
        RECT 54.365 38.935 56.015 39.455 ;
        RECT 56.185 39.105 57.875 39.625 ;
        RECT 58.050 39.055 58.400 39.705 ;
        RECT 54.365 38.165 57.875 38.935 ;
        RECT 58.570 38.885 58.800 39.875 ;
        RECT 58.050 38.715 58.800 38.885 ;
        RECT 58.050 38.425 58.305 38.715 ;
        RECT 58.475 38.165 58.805 38.545 ;
        RECT 58.975 38.425 59.145 40.545 ;
        RECT 59.315 39.745 59.640 40.530 ;
        RECT 59.810 40.255 60.060 40.715 ;
        RECT 60.230 40.215 60.480 40.545 ;
        RECT 60.695 40.215 61.375 40.545 ;
        RECT 60.230 40.085 60.400 40.215 ;
        RECT 60.005 39.915 60.400 40.085 ;
        RECT 59.375 38.695 59.835 39.745 ;
        RECT 60.005 38.555 60.175 39.915 ;
        RECT 60.570 39.655 61.035 40.045 ;
        RECT 60.345 38.845 60.695 39.465 ;
        RECT 60.865 39.065 61.035 39.655 ;
        RECT 61.205 39.435 61.375 40.215 ;
        RECT 61.545 40.115 61.715 40.455 ;
        RECT 61.950 40.285 62.280 40.715 ;
        RECT 62.450 40.115 62.620 40.455 ;
        RECT 62.915 40.255 63.285 40.715 ;
        RECT 61.545 39.945 62.620 40.115 ;
        RECT 63.455 40.085 63.625 40.545 ;
        RECT 63.860 40.205 64.730 40.545 ;
        RECT 64.900 40.255 65.150 40.715 ;
        RECT 63.065 39.915 63.625 40.085 ;
        RECT 63.065 39.775 63.235 39.915 ;
        RECT 61.735 39.605 63.235 39.775 ;
        RECT 63.930 39.745 64.390 40.035 ;
        RECT 61.205 39.265 62.895 39.435 ;
        RECT 60.865 38.845 61.220 39.065 ;
        RECT 61.390 38.555 61.560 39.265 ;
        RECT 61.765 38.845 62.555 39.095 ;
        RECT 62.725 39.085 62.895 39.265 ;
        RECT 63.065 38.915 63.235 39.605 ;
        RECT 59.505 38.165 59.835 38.525 ;
        RECT 60.005 38.385 60.500 38.555 ;
        RECT 60.705 38.385 61.560 38.555 ;
        RECT 62.435 38.165 62.765 38.625 ;
        RECT 62.975 38.525 63.235 38.915 ;
        RECT 63.425 39.735 64.390 39.745 ;
        RECT 64.560 39.825 64.730 40.205 ;
        RECT 65.320 40.165 65.490 40.455 ;
        RECT 65.670 40.335 66.000 40.715 ;
        RECT 65.320 39.995 66.120 40.165 ;
        RECT 63.425 39.575 64.100 39.735 ;
        RECT 64.560 39.655 65.780 39.825 ;
        RECT 63.425 38.785 63.635 39.575 ;
        RECT 64.560 39.565 64.730 39.655 ;
        RECT 63.805 38.785 64.155 39.405 ;
        RECT 64.325 39.395 64.730 39.565 ;
        RECT 64.325 38.615 64.495 39.395 ;
        RECT 64.665 38.945 64.885 39.225 ;
        RECT 65.065 39.115 65.605 39.485 ;
        RECT 65.950 39.405 66.120 39.995 ;
        RECT 66.340 39.575 66.645 40.715 ;
        RECT 66.815 39.525 67.070 40.405 ;
        RECT 67.250 39.565 67.510 40.715 ;
        RECT 67.685 39.640 67.940 40.545 ;
        RECT 68.110 39.955 68.440 40.715 ;
        RECT 68.655 39.785 68.825 40.545 ;
        RECT 65.950 39.375 66.690 39.405 ;
        RECT 64.665 38.775 65.195 38.945 ;
        RECT 62.975 38.355 63.325 38.525 ;
        RECT 63.545 38.335 64.495 38.615 ;
        RECT 64.665 38.165 64.855 38.605 ;
        RECT 65.025 38.545 65.195 38.775 ;
        RECT 65.365 38.715 65.605 39.115 ;
        RECT 65.775 39.075 66.690 39.375 ;
        RECT 65.775 38.900 66.100 39.075 ;
        RECT 65.775 38.545 66.095 38.900 ;
        RECT 66.860 38.875 67.070 39.525 ;
        RECT 65.025 38.375 66.095 38.545 ;
        RECT 66.340 38.165 66.645 38.625 ;
        RECT 66.815 38.345 67.070 38.875 ;
        RECT 67.250 38.165 67.510 39.005 ;
        RECT 67.685 38.910 67.855 39.640 ;
        RECT 68.110 39.615 68.825 39.785 ;
        RECT 68.110 39.405 68.280 39.615 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.930 40.045 71.185 40.545 ;
        RECT 71.355 40.215 71.685 40.715 ;
        RECT 70.930 39.875 71.680 40.045 ;
        RECT 68.025 39.075 68.280 39.405 ;
        RECT 67.685 38.335 67.940 38.910 ;
        RECT 68.110 38.885 68.280 39.075 ;
        RECT 68.560 39.065 68.915 39.435 ;
        RECT 70.930 39.055 71.280 39.705 ;
        RECT 68.110 38.715 68.825 38.885 ;
        RECT 68.110 38.165 68.440 38.545 ;
        RECT 68.655 38.335 68.825 38.715 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 71.450 38.885 71.680 39.875 ;
        RECT 70.930 38.715 71.680 38.885 ;
        RECT 70.930 38.425 71.185 38.715 ;
        RECT 71.355 38.165 71.685 38.545 ;
        RECT 71.855 38.425 72.025 40.545 ;
        RECT 72.195 39.745 72.520 40.530 ;
        RECT 72.690 40.255 72.940 40.715 ;
        RECT 73.110 40.215 73.360 40.545 ;
        RECT 73.575 40.215 74.255 40.545 ;
        RECT 73.110 40.085 73.280 40.215 ;
        RECT 72.885 39.915 73.280 40.085 ;
        RECT 72.255 38.695 72.715 39.745 ;
        RECT 72.885 38.555 73.055 39.915 ;
        RECT 73.450 39.655 73.915 40.045 ;
        RECT 73.225 38.845 73.575 39.465 ;
        RECT 73.745 39.065 73.915 39.655 ;
        RECT 74.085 39.435 74.255 40.215 ;
        RECT 74.425 40.115 74.595 40.455 ;
        RECT 74.830 40.285 75.160 40.715 ;
        RECT 75.330 40.115 75.500 40.455 ;
        RECT 75.795 40.255 76.165 40.715 ;
        RECT 74.425 39.945 75.500 40.115 ;
        RECT 76.335 40.085 76.505 40.545 ;
        RECT 76.740 40.205 77.610 40.545 ;
        RECT 77.780 40.255 78.030 40.715 ;
        RECT 75.945 39.915 76.505 40.085 ;
        RECT 75.945 39.775 76.115 39.915 ;
        RECT 74.615 39.605 76.115 39.775 ;
        RECT 76.810 39.745 77.270 40.035 ;
        RECT 74.085 39.265 75.775 39.435 ;
        RECT 73.745 38.845 74.100 39.065 ;
        RECT 74.270 38.555 74.440 39.265 ;
        RECT 74.645 38.845 75.435 39.095 ;
        RECT 75.605 39.085 75.775 39.265 ;
        RECT 75.945 38.915 76.115 39.605 ;
        RECT 72.385 38.165 72.715 38.525 ;
        RECT 72.885 38.385 73.380 38.555 ;
        RECT 73.585 38.385 74.440 38.555 ;
        RECT 75.315 38.165 75.645 38.625 ;
        RECT 75.855 38.525 76.115 38.915 ;
        RECT 76.305 39.735 77.270 39.745 ;
        RECT 77.440 39.825 77.610 40.205 ;
        RECT 78.200 40.165 78.370 40.455 ;
        RECT 78.550 40.335 78.880 40.715 ;
        RECT 78.200 39.995 79.000 40.165 ;
        RECT 76.305 39.575 76.980 39.735 ;
        RECT 77.440 39.655 78.660 39.825 ;
        RECT 76.305 38.785 76.515 39.575 ;
        RECT 77.440 39.565 77.610 39.655 ;
        RECT 76.685 38.785 77.035 39.405 ;
        RECT 77.205 39.395 77.610 39.565 ;
        RECT 77.205 38.615 77.375 39.395 ;
        RECT 77.545 38.945 77.765 39.225 ;
        RECT 77.945 39.115 78.485 39.485 ;
        RECT 78.830 39.405 79.000 39.995 ;
        RECT 79.220 39.575 79.525 40.715 ;
        RECT 79.695 39.525 79.950 40.405 ;
        RECT 81.135 39.785 81.305 40.545 ;
        RECT 81.485 39.955 81.815 40.715 ;
        RECT 81.135 39.615 81.800 39.785 ;
        RECT 81.985 39.640 82.255 40.545 ;
        RECT 78.830 39.375 79.570 39.405 ;
        RECT 77.545 38.775 78.075 38.945 ;
        RECT 75.855 38.355 76.205 38.525 ;
        RECT 76.425 38.335 77.375 38.615 ;
        RECT 77.545 38.165 77.735 38.605 ;
        RECT 77.905 38.545 78.075 38.775 ;
        RECT 78.245 38.715 78.485 39.115 ;
        RECT 78.655 39.075 79.570 39.375 ;
        RECT 78.655 38.900 78.980 39.075 ;
        RECT 78.655 38.545 78.975 38.900 ;
        RECT 79.740 38.875 79.950 39.525 ;
        RECT 81.630 39.470 81.800 39.615 ;
        RECT 81.065 39.065 81.395 39.435 ;
        RECT 81.630 39.140 81.915 39.470 ;
        RECT 81.630 38.885 81.800 39.140 ;
        RECT 77.905 38.375 78.975 38.545 ;
        RECT 79.220 38.165 79.525 38.625 ;
        RECT 79.695 38.345 79.950 38.875 ;
        RECT 81.135 38.715 81.800 38.885 ;
        RECT 82.085 38.840 82.255 39.640 ;
        RECT 81.135 38.335 81.305 38.715 ;
        RECT 81.485 38.165 81.815 38.545 ;
        RECT 81.995 38.335 82.255 38.840 ;
        RECT 82.425 39.575 82.810 40.545 ;
        RECT 82.980 40.255 83.305 40.715 ;
        RECT 83.825 40.085 84.105 40.545 ;
        RECT 82.980 39.865 84.105 40.085 ;
        RECT 82.425 38.905 82.705 39.575 ;
        RECT 82.980 39.405 83.430 39.865 ;
        RECT 84.295 39.695 84.695 40.545 ;
        RECT 85.095 40.255 85.365 40.715 ;
        RECT 85.535 40.085 85.820 40.545 ;
        RECT 82.875 39.075 83.430 39.405 ;
        RECT 83.600 39.135 84.695 39.695 ;
        RECT 82.980 38.965 83.430 39.075 ;
        RECT 82.425 38.335 82.810 38.905 ;
        RECT 82.980 38.795 84.105 38.965 ;
        RECT 82.980 38.165 83.305 38.625 ;
        RECT 83.825 38.335 84.105 38.795 ;
        RECT 84.295 38.335 84.695 39.135 ;
        RECT 84.865 39.865 85.820 40.085 ;
        RECT 86.105 39.955 86.620 40.365 ;
        RECT 86.855 39.955 87.025 40.715 ;
        RECT 87.195 40.375 89.225 40.545 ;
        RECT 84.865 38.965 85.075 39.865 ;
        RECT 85.245 39.135 85.935 39.695 ;
        RECT 86.105 39.145 86.445 39.955 ;
        RECT 87.195 39.710 87.365 40.375 ;
        RECT 87.760 40.035 88.885 40.205 ;
        RECT 86.615 39.520 87.365 39.710 ;
        RECT 87.535 39.695 88.545 39.865 ;
        RECT 86.105 38.975 87.335 39.145 ;
        RECT 84.865 38.795 85.820 38.965 ;
        RECT 85.095 38.165 85.365 38.625 ;
        RECT 85.535 38.335 85.820 38.795 ;
        RECT 86.380 38.370 86.625 38.975 ;
        RECT 86.845 38.165 87.355 38.700 ;
        RECT 87.535 38.335 87.725 39.695 ;
        RECT 87.895 39.355 88.170 39.495 ;
        RECT 87.895 39.185 88.175 39.355 ;
        RECT 87.895 38.335 88.170 39.185 ;
        RECT 88.375 38.895 88.545 39.695 ;
        RECT 88.715 38.905 88.885 40.035 ;
        RECT 89.055 39.405 89.225 40.375 ;
        RECT 89.395 39.575 89.565 40.715 ;
        RECT 89.735 39.575 90.070 40.545 ;
        RECT 90.360 40.085 90.645 40.545 ;
        RECT 90.815 40.255 91.085 40.715 ;
        RECT 90.360 39.865 91.315 40.085 ;
        RECT 89.055 39.075 89.250 39.405 ;
        RECT 89.475 39.075 89.730 39.405 ;
        RECT 89.475 38.905 89.645 39.075 ;
        RECT 89.900 38.905 90.070 39.575 ;
        RECT 90.245 39.135 90.935 39.695 ;
        RECT 91.105 38.965 91.315 39.865 ;
        RECT 88.715 38.735 89.645 38.905 ;
        RECT 88.715 38.700 88.890 38.735 ;
        RECT 88.360 38.335 88.890 38.700 ;
        RECT 89.315 38.165 89.645 38.565 ;
        RECT 89.815 38.335 90.070 38.905 ;
        RECT 90.360 38.795 91.315 38.965 ;
        RECT 91.485 39.695 91.885 40.545 ;
        RECT 92.075 40.085 92.355 40.545 ;
        RECT 92.875 40.255 93.200 40.715 ;
        RECT 92.075 39.865 93.200 40.085 ;
        RECT 91.485 39.135 92.580 39.695 ;
        RECT 92.750 39.405 93.200 39.865 ;
        RECT 93.370 39.575 93.755 40.545 ;
        RECT 90.360 38.335 90.645 38.795 ;
        RECT 90.815 38.165 91.085 38.625 ;
        RECT 91.485 38.335 91.885 39.135 ;
        RECT 92.750 39.075 93.305 39.405 ;
        RECT 92.750 38.965 93.200 39.075 ;
        RECT 92.075 38.795 93.200 38.965 ;
        RECT 93.475 38.905 93.755 39.575 ;
        RECT 92.075 38.335 92.355 38.795 ;
        RECT 92.875 38.165 93.200 38.625 ;
        RECT 93.370 38.335 93.755 38.905 ;
        RECT 93.925 39.640 94.195 40.545 ;
        RECT 94.365 39.955 94.695 40.715 ;
        RECT 94.875 39.785 95.045 40.545 ;
        RECT 93.925 38.840 94.095 39.640 ;
        RECT 94.380 39.615 95.045 39.785 ;
        RECT 94.380 39.470 94.550 39.615 ;
        RECT 95.765 39.550 96.055 40.715 ;
        RECT 96.265 39.575 96.495 40.715 ;
        RECT 96.665 39.565 96.995 40.545 ;
        RECT 97.165 39.575 97.375 40.715 ;
        RECT 98.615 40.045 98.785 40.545 ;
        RECT 98.955 40.215 99.285 40.715 ;
        RECT 98.615 39.875 99.280 40.045 ;
        RECT 94.265 39.140 94.550 39.470 ;
        RECT 94.380 38.885 94.550 39.140 ;
        RECT 94.785 39.065 95.115 39.435 ;
        RECT 96.245 39.155 96.575 39.405 ;
        RECT 93.925 38.335 94.185 38.840 ;
        RECT 94.380 38.715 95.045 38.885 ;
        RECT 94.365 38.165 94.695 38.545 ;
        RECT 94.875 38.335 95.045 38.715 ;
        RECT 95.765 38.165 96.055 38.890 ;
        RECT 96.265 38.165 96.495 38.985 ;
        RECT 96.745 38.965 96.995 39.565 ;
        RECT 98.530 39.055 98.880 39.705 ;
        RECT 96.665 38.335 96.995 38.965 ;
        RECT 97.165 38.165 97.375 38.985 ;
        RECT 99.050 38.885 99.280 39.875 ;
        RECT 98.615 38.715 99.280 38.885 ;
        RECT 98.615 38.425 98.785 38.715 ;
        RECT 98.955 38.165 99.285 38.545 ;
        RECT 99.455 38.425 99.680 40.545 ;
        RECT 99.895 40.215 100.225 40.715 ;
        RECT 100.395 40.045 100.565 40.545 ;
        RECT 100.800 40.330 101.630 40.500 ;
        RECT 101.870 40.335 102.250 40.715 ;
        RECT 99.870 39.875 100.565 40.045 ;
        RECT 99.870 38.905 100.040 39.875 ;
        RECT 100.210 39.085 100.620 39.705 ;
        RECT 100.790 39.655 101.290 40.035 ;
        RECT 99.870 38.715 100.565 38.905 ;
        RECT 100.790 38.785 101.010 39.655 ;
        RECT 101.460 39.485 101.630 40.330 ;
        RECT 102.430 40.165 102.600 40.455 ;
        RECT 102.770 40.335 103.100 40.715 ;
        RECT 103.570 40.245 104.200 40.495 ;
        RECT 104.380 40.335 104.800 40.715 ;
        RECT 104.030 40.165 104.200 40.245 ;
        RECT 105.000 40.165 105.240 40.455 ;
        RECT 101.800 39.915 103.170 40.165 ;
        RECT 101.800 39.655 102.050 39.915 ;
        RECT 102.560 39.485 102.810 39.645 ;
        RECT 101.460 39.315 102.810 39.485 ;
        RECT 101.460 39.275 101.880 39.315 ;
        RECT 101.190 38.725 101.540 39.095 ;
        RECT 99.895 38.165 100.225 38.545 ;
        RECT 100.395 38.385 100.565 38.715 ;
        RECT 101.710 38.545 101.880 39.275 ;
        RECT 102.980 39.145 103.170 39.915 ;
        RECT 102.050 38.815 102.460 39.145 ;
        RECT 102.750 38.805 103.170 39.145 ;
        RECT 103.340 39.735 103.860 40.045 ;
        RECT 104.030 39.995 105.240 40.165 ;
        RECT 105.470 40.025 105.800 40.715 ;
        RECT 103.340 38.975 103.510 39.735 ;
        RECT 103.680 39.145 103.860 39.555 ;
        RECT 104.030 39.485 104.200 39.995 ;
        RECT 105.970 39.845 106.140 40.455 ;
        RECT 106.410 39.995 106.740 40.505 ;
        RECT 105.970 39.825 106.290 39.845 ;
        RECT 104.370 39.655 106.290 39.825 ;
        RECT 104.030 39.315 105.930 39.485 ;
        RECT 104.260 38.975 104.590 39.095 ;
        RECT 103.340 38.805 104.590 38.975 ;
        RECT 100.865 38.345 101.880 38.545 ;
        RECT 102.050 38.165 102.460 38.605 ;
        RECT 102.750 38.375 103.000 38.805 ;
        RECT 103.200 38.165 103.520 38.625 ;
        RECT 104.760 38.555 104.930 39.315 ;
        RECT 105.600 39.255 105.930 39.315 ;
        RECT 105.120 39.085 105.450 39.145 ;
        RECT 105.120 38.815 105.780 39.085 ;
        RECT 106.100 38.760 106.290 39.655 ;
        RECT 104.080 38.385 104.930 38.555 ;
        RECT 105.130 38.165 105.790 38.645 ;
        RECT 105.970 38.430 106.290 38.760 ;
        RECT 106.490 39.405 106.740 39.995 ;
        RECT 106.920 39.915 107.205 40.715 ;
        RECT 107.385 40.375 107.640 40.405 ;
        RECT 107.385 40.205 107.725 40.375 ;
        RECT 107.385 39.735 107.640 40.205 ;
        RECT 108.190 40.045 108.445 40.545 ;
        RECT 108.615 40.215 108.945 40.715 ;
        RECT 108.190 39.875 108.940 40.045 ;
        RECT 106.490 39.075 107.290 39.405 ;
        RECT 106.490 38.425 106.740 39.075 ;
        RECT 107.460 38.875 107.640 39.735 ;
        RECT 108.190 39.055 108.540 39.705 ;
        RECT 108.710 38.885 108.940 39.875 ;
        RECT 106.920 38.165 107.205 38.625 ;
        RECT 107.385 38.345 107.640 38.875 ;
        RECT 108.190 38.715 108.940 38.885 ;
        RECT 108.190 38.425 108.445 38.715 ;
        RECT 108.615 38.165 108.945 38.545 ;
        RECT 109.115 38.425 109.285 40.545 ;
        RECT 109.455 39.745 109.780 40.530 ;
        RECT 109.950 40.255 110.200 40.715 ;
        RECT 110.370 40.215 110.620 40.545 ;
        RECT 110.835 40.215 111.515 40.545 ;
        RECT 110.370 40.085 110.540 40.215 ;
        RECT 110.145 39.915 110.540 40.085 ;
        RECT 109.515 38.695 109.975 39.745 ;
        RECT 110.145 38.555 110.315 39.915 ;
        RECT 110.710 39.655 111.175 40.045 ;
        RECT 110.485 38.845 110.835 39.465 ;
        RECT 111.005 39.065 111.175 39.655 ;
        RECT 111.345 39.435 111.515 40.215 ;
        RECT 111.685 40.115 111.855 40.455 ;
        RECT 112.090 40.285 112.420 40.715 ;
        RECT 112.590 40.115 112.760 40.455 ;
        RECT 113.055 40.255 113.425 40.715 ;
        RECT 111.685 39.945 112.760 40.115 ;
        RECT 113.595 40.085 113.765 40.545 ;
        RECT 114.000 40.205 114.870 40.545 ;
        RECT 115.040 40.255 115.290 40.715 ;
        RECT 113.205 39.915 113.765 40.085 ;
        RECT 113.205 39.775 113.375 39.915 ;
        RECT 111.875 39.605 113.375 39.775 ;
        RECT 114.070 39.745 114.530 40.035 ;
        RECT 111.345 39.265 113.035 39.435 ;
        RECT 111.005 38.845 111.360 39.065 ;
        RECT 111.530 38.555 111.700 39.265 ;
        RECT 111.905 38.845 112.695 39.095 ;
        RECT 112.865 39.085 113.035 39.265 ;
        RECT 113.205 38.915 113.375 39.605 ;
        RECT 109.645 38.165 109.975 38.525 ;
        RECT 110.145 38.385 110.640 38.555 ;
        RECT 110.845 38.385 111.700 38.555 ;
        RECT 112.575 38.165 112.905 38.625 ;
        RECT 113.115 38.525 113.375 38.915 ;
        RECT 113.565 39.735 114.530 39.745 ;
        RECT 114.700 39.825 114.870 40.205 ;
        RECT 115.460 40.165 115.630 40.455 ;
        RECT 115.810 40.335 116.140 40.715 ;
        RECT 115.460 39.995 116.260 40.165 ;
        RECT 113.565 39.575 114.240 39.735 ;
        RECT 114.700 39.655 115.920 39.825 ;
        RECT 113.565 38.785 113.775 39.575 ;
        RECT 114.700 39.565 114.870 39.655 ;
        RECT 113.945 38.785 114.295 39.405 ;
        RECT 114.465 39.395 114.870 39.565 ;
        RECT 114.465 38.615 114.635 39.395 ;
        RECT 114.805 38.945 115.025 39.225 ;
        RECT 115.205 39.115 115.745 39.485 ;
        RECT 116.090 39.405 116.260 39.995 ;
        RECT 116.480 39.575 116.785 40.715 ;
        RECT 116.955 39.525 117.210 40.405 ;
        RECT 117.385 39.625 120.895 40.715 ;
        RECT 116.090 39.375 116.830 39.405 ;
        RECT 114.805 38.775 115.335 38.945 ;
        RECT 113.115 38.355 113.465 38.525 ;
        RECT 113.685 38.335 114.635 38.615 ;
        RECT 114.805 38.165 114.995 38.605 ;
        RECT 115.165 38.545 115.335 38.775 ;
        RECT 115.505 38.715 115.745 39.115 ;
        RECT 115.915 39.075 116.830 39.375 ;
        RECT 115.915 38.900 116.240 39.075 ;
        RECT 115.915 38.545 116.235 38.900 ;
        RECT 117.000 38.875 117.210 39.525 ;
        RECT 115.165 38.375 116.235 38.545 ;
        RECT 116.480 38.165 116.785 38.625 ;
        RECT 116.955 38.345 117.210 38.875 ;
        RECT 117.385 38.935 119.035 39.455 ;
        RECT 119.205 39.105 120.895 39.625 ;
        RECT 121.525 39.550 121.815 40.715 ;
        RECT 121.985 39.625 123.655 40.715 ;
        RECT 121.985 38.935 122.735 39.455 ;
        RECT 122.905 39.105 123.655 39.625 ;
        RECT 124.285 39.625 125.495 40.715 ;
        RECT 124.285 39.085 124.805 39.625 ;
        RECT 117.385 38.165 120.895 38.935 ;
        RECT 121.525 38.165 121.815 38.890 ;
        RECT 121.985 38.165 123.655 38.935 ;
        RECT 124.975 38.915 125.495 39.455 ;
        RECT 124.285 38.165 125.495 38.915 ;
        RECT 5.520 37.995 125.580 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 6.985 37.450 12.330 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 8.570 36.620 8.910 37.450 ;
        RECT 12.505 37.225 14.175 37.995 ;
        RECT 14.350 37.445 14.605 37.735 ;
        RECT 14.775 37.615 15.105 37.995 ;
        RECT 14.350 37.275 15.100 37.445 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 10.390 35.880 10.740 37.130 ;
        RECT 12.505 36.705 13.255 37.225 ;
        RECT 13.425 36.535 14.175 37.055 ;
        RECT 6.985 35.445 12.330 35.880 ;
        RECT 12.505 35.445 14.175 36.535 ;
        RECT 14.350 36.455 14.700 37.105 ;
        RECT 14.870 36.285 15.100 37.275 ;
        RECT 14.350 36.115 15.100 36.285 ;
        RECT 14.350 35.615 14.605 36.115 ;
        RECT 14.775 35.445 15.105 35.945 ;
        RECT 15.275 35.615 15.445 37.735 ;
        RECT 15.805 37.635 16.135 37.995 ;
        RECT 16.305 37.605 16.800 37.775 ;
        RECT 17.005 37.605 17.860 37.775 ;
        RECT 15.675 36.415 16.135 37.465 ;
        RECT 15.615 35.630 15.940 36.415 ;
        RECT 16.305 36.245 16.475 37.605 ;
        RECT 16.645 36.695 16.995 37.315 ;
        RECT 17.165 37.095 17.520 37.315 ;
        RECT 17.165 36.505 17.335 37.095 ;
        RECT 17.690 36.895 17.860 37.605 ;
        RECT 18.735 37.535 19.065 37.995 ;
        RECT 19.275 37.635 19.625 37.805 ;
        RECT 18.065 37.065 18.855 37.315 ;
        RECT 19.275 37.245 19.535 37.635 ;
        RECT 19.845 37.545 20.795 37.825 ;
        RECT 20.965 37.555 21.155 37.995 ;
        RECT 21.325 37.615 22.395 37.785 ;
        RECT 19.025 36.895 19.195 37.075 ;
        RECT 16.305 36.075 16.700 36.245 ;
        RECT 16.870 36.115 17.335 36.505 ;
        RECT 17.505 36.725 19.195 36.895 ;
        RECT 16.530 35.945 16.700 36.075 ;
        RECT 17.505 35.945 17.675 36.725 ;
        RECT 19.365 36.555 19.535 37.245 ;
        RECT 18.035 36.385 19.535 36.555 ;
        RECT 19.725 36.585 19.935 37.375 ;
        RECT 20.105 36.755 20.455 37.375 ;
        RECT 20.625 36.765 20.795 37.545 ;
        RECT 21.325 37.385 21.495 37.615 ;
        RECT 20.965 37.215 21.495 37.385 ;
        RECT 20.965 36.935 21.185 37.215 ;
        RECT 21.665 37.045 21.905 37.445 ;
        RECT 20.625 36.595 21.030 36.765 ;
        RECT 21.365 36.675 21.905 37.045 ;
        RECT 22.075 37.260 22.395 37.615 ;
        RECT 22.640 37.535 22.945 37.995 ;
        RECT 23.115 37.285 23.370 37.815 ;
        RECT 22.075 37.085 22.400 37.260 ;
        RECT 22.075 36.785 22.990 37.085 ;
        RECT 22.250 36.755 22.990 36.785 ;
        RECT 19.725 36.425 20.400 36.585 ;
        RECT 20.860 36.505 21.030 36.595 ;
        RECT 19.725 36.415 20.690 36.425 ;
        RECT 19.365 36.245 19.535 36.385 ;
        RECT 16.110 35.445 16.360 35.905 ;
        RECT 16.530 35.615 16.780 35.945 ;
        RECT 16.995 35.615 17.675 35.945 ;
        RECT 17.845 36.045 18.920 36.215 ;
        RECT 19.365 36.075 19.925 36.245 ;
        RECT 20.230 36.125 20.690 36.415 ;
        RECT 20.860 36.335 22.080 36.505 ;
        RECT 17.845 35.705 18.015 36.045 ;
        RECT 18.250 35.445 18.580 35.875 ;
        RECT 18.750 35.705 18.920 36.045 ;
        RECT 19.215 35.445 19.585 35.905 ;
        RECT 19.755 35.615 19.925 36.075 ;
        RECT 20.860 35.955 21.030 36.335 ;
        RECT 22.250 36.165 22.420 36.755 ;
        RECT 23.160 36.635 23.370 37.285 ;
        RECT 20.160 35.615 21.030 35.955 ;
        RECT 21.620 35.995 22.420 36.165 ;
        RECT 21.200 35.445 21.450 35.905 ;
        RECT 21.620 35.705 21.790 35.995 ;
        RECT 21.970 35.445 22.300 35.825 ;
        RECT 22.640 35.445 22.945 36.585 ;
        RECT 23.115 35.755 23.370 36.635 ;
        RECT 23.550 37.255 23.805 37.825 ;
        RECT 23.975 37.595 24.305 37.995 ;
        RECT 24.730 37.460 25.260 37.825 ;
        RECT 25.450 37.655 25.725 37.825 ;
        RECT 25.445 37.485 25.725 37.655 ;
        RECT 24.730 37.425 24.905 37.460 ;
        RECT 23.975 37.255 24.905 37.425 ;
        RECT 23.550 36.585 23.720 37.255 ;
        RECT 23.975 37.085 24.145 37.255 ;
        RECT 23.890 36.755 24.145 37.085 ;
        RECT 24.370 36.755 24.565 37.085 ;
        RECT 23.550 35.615 23.885 36.585 ;
        RECT 24.055 35.445 24.225 36.585 ;
        RECT 24.395 35.785 24.565 36.755 ;
        RECT 24.735 36.125 24.905 37.255 ;
        RECT 25.075 36.465 25.245 37.265 ;
        RECT 25.450 36.665 25.725 37.485 ;
        RECT 25.895 36.465 26.085 37.825 ;
        RECT 26.265 37.460 26.775 37.995 ;
        RECT 26.995 37.185 27.240 37.790 ;
        RECT 27.685 37.225 31.195 37.995 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 26.285 37.015 27.515 37.185 ;
        RECT 25.075 36.295 26.085 36.465 ;
        RECT 26.255 36.450 27.005 36.640 ;
        RECT 24.735 35.955 25.860 36.125 ;
        RECT 26.255 35.785 26.425 36.450 ;
        RECT 27.175 36.205 27.515 37.015 ;
        RECT 27.685 36.705 29.335 37.225 ;
        RECT 32.100 37.185 32.345 37.790 ;
        RECT 32.565 37.460 33.075 37.995 ;
        RECT 29.505 36.535 31.195 37.055 ;
        RECT 31.825 37.015 33.055 37.185 ;
        RECT 24.395 35.615 26.425 35.785 ;
        RECT 26.595 35.445 26.765 36.205 ;
        RECT 27.000 35.795 27.515 36.205 ;
        RECT 27.685 35.445 31.195 36.535 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 31.825 36.205 32.165 37.015 ;
        RECT 32.335 36.450 33.085 36.640 ;
        RECT 31.825 35.795 32.340 36.205 ;
        RECT 32.575 35.445 32.745 36.205 ;
        RECT 32.915 35.785 33.085 36.450 ;
        RECT 33.255 36.465 33.445 37.825 ;
        RECT 33.615 36.975 33.890 37.825 ;
        RECT 34.080 37.460 34.610 37.825 ;
        RECT 35.035 37.595 35.365 37.995 ;
        RECT 34.435 37.425 34.610 37.460 ;
        RECT 33.615 36.805 33.895 36.975 ;
        RECT 33.615 36.665 33.890 36.805 ;
        RECT 34.095 36.465 34.265 37.265 ;
        RECT 33.255 36.295 34.265 36.465 ;
        RECT 34.435 37.255 35.365 37.425 ;
        RECT 35.535 37.255 35.790 37.825 ;
        RECT 36.515 37.445 36.685 37.735 ;
        RECT 36.855 37.615 37.185 37.995 ;
        RECT 36.515 37.275 37.180 37.445 ;
        RECT 34.435 36.125 34.605 37.255 ;
        RECT 35.195 37.085 35.365 37.255 ;
        RECT 33.480 35.955 34.605 36.125 ;
        RECT 34.775 36.755 34.970 37.085 ;
        RECT 35.195 36.755 35.450 37.085 ;
        RECT 34.775 35.785 34.945 36.755 ;
        RECT 35.620 36.585 35.790 37.255 ;
        RECT 32.915 35.615 34.945 35.785 ;
        RECT 35.115 35.445 35.285 36.585 ;
        RECT 35.455 35.615 35.790 36.585 ;
        RECT 36.430 36.455 36.780 37.105 ;
        RECT 36.950 36.285 37.180 37.275 ;
        RECT 36.515 36.115 37.180 36.285 ;
        RECT 36.515 35.615 36.685 36.115 ;
        RECT 36.855 35.445 37.185 35.945 ;
        RECT 37.355 35.615 37.580 37.735 ;
        RECT 37.795 37.615 38.125 37.995 ;
        RECT 38.295 37.445 38.465 37.775 ;
        RECT 38.765 37.615 39.780 37.815 ;
        RECT 37.770 37.255 38.465 37.445 ;
        RECT 37.770 36.285 37.940 37.255 ;
        RECT 38.110 36.455 38.520 37.075 ;
        RECT 38.690 36.505 38.910 37.375 ;
        RECT 39.090 37.065 39.440 37.435 ;
        RECT 39.610 36.885 39.780 37.615 ;
        RECT 39.950 37.555 40.360 37.995 ;
        RECT 40.650 37.355 40.900 37.785 ;
        RECT 41.100 37.535 41.420 37.995 ;
        RECT 41.980 37.605 42.830 37.775 ;
        RECT 39.950 37.015 40.360 37.345 ;
        RECT 40.650 37.015 41.070 37.355 ;
        RECT 39.360 36.845 39.780 36.885 ;
        RECT 39.360 36.675 40.710 36.845 ;
        RECT 37.770 36.115 38.465 36.285 ;
        RECT 38.690 36.125 39.190 36.505 ;
        RECT 37.795 35.445 38.125 35.945 ;
        RECT 38.295 35.615 38.465 36.115 ;
        RECT 39.360 35.830 39.530 36.675 ;
        RECT 40.460 36.515 40.710 36.675 ;
        RECT 39.700 36.245 39.950 36.505 ;
        RECT 40.880 36.245 41.070 37.015 ;
        RECT 39.700 35.995 41.070 36.245 ;
        RECT 41.240 37.185 42.490 37.355 ;
        RECT 41.240 36.425 41.410 37.185 ;
        RECT 42.160 37.065 42.490 37.185 ;
        RECT 41.580 36.605 41.760 37.015 ;
        RECT 42.660 36.845 42.830 37.605 ;
        RECT 43.030 37.515 43.690 37.995 ;
        RECT 43.870 37.400 44.190 37.730 ;
        RECT 43.020 37.075 43.680 37.345 ;
        RECT 43.020 37.015 43.350 37.075 ;
        RECT 43.500 36.845 43.830 36.905 ;
        RECT 41.930 36.675 43.830 36.845 ;
        RECT 41.240 36.115 41.760 36.425 ;
        RECT 41.930 36.165 42.100 36.675 ;
        RECT 44.000 36.505 44.190 37.400 ;
        RECT 42.270 36.335 44.190 36.505 ;
        RECT 43.870 36.315 44.190 36.335 ;
        RECT 44.390 37.085 44.640 37.735 ;
        RECT 44.820 37.535 45.105 37.995 ;
        RECT 45.285 37.285 45.540 37.815 ;
        RECT 44.390 36.755 45.190 37.085 ;
        RECT 41.930 35.995 43.140 36.165 ;
        RECT 38.700 35.660 39.530 35.830 ;
        RECT 39.770 35.445 40.150 35.825 ;
        RECT 40.330 35.705 40.500 35.995 ;
        RECT 41.930 35.915 42.100 35.995 ;
        RECT 40.670 35.445 41.000 35.825 ;
        RECT 41.470 35.665 42.100 35.915 ;
        RECT 42.280 35.445 42.700 35.825 ;
        RECT 42.900 35.705 43.140 35.995 ;
        RECT 43.370 35.445 43.700 36.135 ;
        RECT 43.870 35.705 44.040 36.315 ;
        RECT 44.390 36.165 44.640 36.755 ;
        RECT 45.360 36.425 45.540 37.285 ;
        RECT 44.310 35.655 44.640 36.165 ;
        RECT 44.820 35.445 45.105 36.245 ;
        RECT 45.285 35.955 45.540 36.425 ;
        RECT 46.090 37.255 46.345 37.825 ;
        RECT 46.515 37.595 46.845 37.995 ;
        RECT 47.270 37.460 47.800 37.825 ;
        RECT 47.990 37.655 48.265 37.825 ;
        RECT 47.985 37.485 48.265 37.655 ;
        RECT 47.270 37.425 47.445 37.460 ;
        RECT 46.515 37.255 47.445 37.425 ;
        RECT 46.090 36.585 46.260 37.255 ;
        RECT 46.515 37.085 46.685 37.255 ;
        RECT 46.430 36.755 46.685 37.085 ;
        RECT 46.910 36.755 47.105 37.085 ;
        RECT 45.285 35.785 45.625 35.955 ;
        RECT 45.285 35.755 45.540 35.785 ;
        RECT 46.090 35.615 46.425 36.585 ;
        RECT 46.595 35.445 46.765 36.585 ;
        RECT 46.935 35.785 47.105 36.755 ;
        RECT 47.275 36.125 47.445 37.255 ;
        RECT 47.615 36.465 47.785 37.265 ;
        RECT 47.990 36.665 48.265 37.485 ;
        RECT 48.435 36.465 48.625 37.825 ;
        RECT 48.805 37.460 49.315 37.995 ;
        RECT 49.535 37.185 49.780 37.790 ;
        RECT 50.225 37.450 55.570 37.995 ;
        RECT 48.825 37.015 50.055 37.185 ;
        RECT 47.615 36.295 48.625 36.465 ;
        RECT 48.795 36.450 49.545 36.640 ;
        RECT 47.275 35.955 48.400 36.125 ;
        RECT 48.795 35.785 48.965 36.450 ;
        RECT 49.715 36.205 50.055 37.015 ;
        RECT 51.810 36.620 52.150 37.450 ;
        RECT 55.745 37.245 56.955 37.995 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 46.935 35.615 48.965 35.785 ;
        RECT 49.135 35.445 49.305 36.205 ;
        RECT 49.540 35.795 50.055 36.205 ;
        RECT 53.630 35.880 53.980 37.130 ;
        RECT 55.745 36.705 56.265 37.245 ;
        RECT 57.645 37.175 57.855 37.995 ;
        RECT 58.025 37.195 58.355 37.825 ;
        RECT 56.435 36.535 56.955 37.075 ;
        RECT 50.225 35.445 55.570 35.880 ;
        RECT 55.745 35.445 56.955 36.535 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 58.025 36.595 58.275 37.195 ;
        RECT 58.525 37.175 58.755 37.995 ;
        RECT 59.485 37.175 59.695 37.995 ;
        RECT 59.865 37.195 60.195 37.825 ;
        RECT 58.445 36.755 58.775 37.005 ;
        RECT 59.865 36.595 60.115 37.195 ;
        RECT 60.365 37.175 60.595 37.995 ;
        RECT 61.350 37.425 61.525 37.825 ;
        RECT 61.695 37.615 62.025 37.995 ;
        RECT 62.270 37.495 62.500 37.825 ;
        RECT 61.350 37.255 61.980 37.425 ;
        RECT 61.810 37.085 61.980 37.255 ;
        RECT 60.285 36.755 60.615 37.005 ;
        RECT 57.645 35.445 57.855 36.585 ;
        RECT 58.025 35.615 58.355 36.595 ;
        RECT 58.525 35.445 58.755 36.585 ;
        RECT 59.485 35.445 59.695 36.585 ;
        RECT 59.865 35.615 60.195 36.595 ;
        RECT 60.365 35.445 60.595 36.585 ;
        RECT 61.265 36.405 61.630 37.085 ;
        RECT 61.810 36.755 62.160 37.085 ;
        RECT 61.810 36.235 61.980 36.755 ;
        RECT 61.350 36.065 61.980 36.235 ;
        RECT 62.330 36.205 62.500 37.495 ;
        RECT 62.700 36.385 62.980 37.660 ;
        RECT 63.205 37.315 63.475 37.660 ;
        RECT 63.935 37.615 64.265 37.995 ;
        RECT 64.435 37.740 64.770 37.785 ;
        RECT 63.165 37.145 63.475 37.315 ;
        RECT 63.205 36.385 63.475 37.145 ;
        RECT 63.665 36.385 64.005 37.415 ;
        RECT 64.435 37.275 64.775 37.740 ;
        RECT 64.175 36.755 64.435 37.085 ;
        RECT 64.175 36.205 64.345 36.755 ;
        RECT 64.605 36.585 64.775 37.275 ;
        RECT 61.350 35.615 61.525 36.065 ;
        RECT 62.330 36.035 64.345 36.205 ;
        RECT 61.695 35.445 62.025 35.885 ;
        RECT 62.330 35.615 62.500 36.035 ;
        RECT 62.735 35.445 63.405 35.855 ;
        RECT 63.620 35.615 63.790 36.035 ;
        RECT 63.990 35.445 64.320 35.855 ;
        RECT 64.515 35.615 64.775 36.585 ;
        RECT 64.945 37.495 65.205 37.825 ;
        RECT 65.415 37.515 65.690 37.995 ;
        RECT 64.945 36.585 65.115 37.495 ;
        RECT 65.900 37.425 66.105 37.825 ;
        RECT 66.275 37.595 66.610 37.995 ;
        RECT 65.285 36.755 65.645 37.335 ;
        RECT 65.900 37.255 66.585 37.425 ;
        RECT 65.825 36.585 66.075 37.085 ;
        RECT 64.945 36.415 66.075 36.585 ;
        RECT 64.945 35.645 65.215 36.415 ;
        RECT 66.245 36.225 66.585 37.255 ;
        RECT 67.360 37.365 67.645 37.825 ;
        RECT 67.815 37.535 68.085 37.995 ;
        RECT 67.360 37.195 68.315 37.365 ;
        RECT 67.245 36.465 67.935 37.025 ;
        RECT 68.105 36.295 68.315 37.195 ;
        RECT 65.385 35.445 65.715 36.225 ;
        RECT 65.920 36.050 66.585 36.225 ;
        RECT 67.360 36.075 68.315 36.295 ;
        RECT 68.485 37.025 68.885 37.825 ;
        RECT 69.075 37.365 69.355 37.825 ;
        RECT 69.875 37.535 70.200 37.995 ;
        RECT 69.075 37.195 70.200 37.365 ;
        RECT 70.370 37.255 70.755 37.825 ;
        RECT 69.750 37.085 70.200 37.195 ;
        RECT 68.485 36.465 69.580 37.025 ;
        RECT 69.750 36.755 70.305 37.085 ;
        RECT 65.920 35.645 66.105 36.050 ;
        RECT 66.275 35.445 66.610 35.870 ;
        RECT 67.360 35.615 67.645 36.075 ;
        RECT 67.815 35.445 68.085 35.905 ;
        RECT 68.485 35.615 68.885 36.465 ;
        RECT 69.750 36.295 70.200 36.755 ;
        RECT 70.475 36.585 70.755 37.255 ;
        RECT 70.925 37.225 73.515 37.995 ;
        RECT 73.685 37.320 73.945 37.825 ;
        RECT 74.125 37.615 74.455 37.995 ;
        RECT 74.635 37.445 74.805 37.825 ;
        RECT 70.925 36.705 72.135 37.225 ;
        RECT 69.075 36.075 70.200 36.295 ;
        RECT 69.075 35.615 69.355 36.075 ;
        RECT 69.875 35.445 70.200 35.905 ;
        RECT 70.370 35.615 70.755 36.585 ;
        RECT 72.305 36.535 73.515 37.055 ;
        RECT 70.925 35.445 73.515 36.535 ;
        RECT 73.685 36.520 73.855 37.320 ;
        RECT 74.140 37.275 74.805 37.445 ;
        RECT 74.140 37.020 74.310 37.275 ;
        RECT 75.530 37.255 75.785 37.825 ;
        RECT 75.955 37.595 76.285 37.995 ;
        RECT 76.710 37.460 77.240 37.825 ;
        RECT 76.710 37.425 76.885 37.460 ;
        RECT 75.955 37.255 76.885 37.425 ;
        RECT 77.430 37.315 77.705 37.825 ;
        RECT 74.025 36.690 74.310 37.020 ;
        RECT 74.545 36.725 74.875 37.095 ;
        RECT 74.140 36.545 74.310 36.690 ;
        RECT 75.530 36.585 75.700 37.255 ;
        RECT 75.955 37.085 76.125 37.255 ;
        RECT 75.870 36.755 76.125 37.085 ;
        RECT 76.350 36.755 76.545 37.085 ;
        RECT 73.685 35.615 73.955 36.520 ;
        RECT 74.140 36.375 74.805 36.545 ;
        RECT 74.125 35.445 74.455 36.205 ;
        RECT 74.635 35.615 74.805 36.375 ;
        RECT 75.530 35.615 75.865 36.585 ;
        RECT 76.035 35.445 76.205 36.585 ;
        RECT 76.375 35.785 76.545 36.755 ;
        RECT 76.715 36.125 76.885 37.255 ;
        RECT 77.055 36.465 77.225 37.265 ;
        RECT 77.425 37.145 77.705 37.315 ;
        RECT 77.430 36.665 77.705 37.145 ;
        RECT 77.875 36.465 78.065 37.825 ;
        RECT 78.245 37.460 78.755 37.995 ;
        RECT 78.975 37.185 79.220 37.790 ;
        RECT 78.265 37.015 79.495 37.185 ;
        RECT 79.725 37.175 79.935 37.995 ;
        RECT 80.105 37.195 80.435 37.825 ;
        RECT 77.055 36.295 78.065 36.465 ;
        RECT 78.235 36.450 78.985 36.640 ;
        RECT 76.715 35.955 77.840 36.125 ;
        RECT 78.235 35.785 78.405 36.450 ;
        RECT 79.155 36.205 79.495 37.015 ;
        RECT 80.105 36.595 80.355 37.195 ;
        RECT 80.605 37.175 80.835 37.995 ;
        RECT 81.545 37.175 81.775 37.995 ;
        RECT 81.945 37.195 82.275 37.825 ;
        RECT 80.525 36.755 80.855 37.005 ;
        RECT 81.525 36.755 81.855 37.005 ;
        RECT 82.025 36.595 82.275 37.195 ;
        RECT 82.445 37.175 82.655 37.995 ;
        RECT 82.885 37.270 83.175 37.995 ;
        RECT 83.350 37.445 83.605 37.735 ;
        RECT 83.775 37.615 84.105 37.995 ;
        RECT 83.350 37.275 84.100 37.445 ;
        RECT 76.375 35.615 78.405 35.785 ;
        RECT 78.575 35.445 78.745 36.205 ;
        RECT 78.980 35.795 79.495 36.205 ;
        RECT 79.725 35.445 79.935 36.585 ;
        RECT 80.105 35.615 80.435 36.595 ;
        RECT 80.605 35.445 80.835 36.585 ;
        RECT 81.545 35.445 81.775 36.585 ;
        RECT 81.945 35.615 82.275 36.595 ;
        RECT 82.445 35.445 82.655 36.585 ;
        RECT 82.885 35.445 83.175 36.610 ;
        RECT 83.350 36.455 83.700 37.105 ;
        RECT 83.870 36.285 84.100 37.275 ;
        RECT 83.350 36.115 84.100 36.285 ;
        RECT 83.350 35.615 83.605 36.115 ;
        RECT 83.775 35.445 84.105 35.945 ;
        RECT 84.275 35.615 84.445 37.735 ;
        RECT 84.805 37.635 85.135 37.995 ;
        RECT 85.305 37.605 85.800 37.775 ;
        RECT 86.005 37.605 86.860 37.775 ;
        RECT 84.675 36.415 85.135 37.465 ;
        RECT 84.615 35.630 84.940 36.415 ;
        RECT 85.305 36.245 85.475 37.605 ;
        RECT 85.645 36.695 85.995 37.315 ;
        RECT 86.165 37.095 86.520 37.315 ;
        RECT 86.165 36.505 86.335 37.095 ;
        RECT 86.690 36.895 86.860 37.605 ;
        RECT 87.735 37.535 88.065 37.995 ;
        RECT 88.275 37.635 88.625 37.805 ;
        RECT 87.065 37.065 87.855 37.315 ;
        RECT 88.275 37.245 88.535 37.635 ;
        RECT 88.845 37.545 89.795 37.825 ;
        RECT 89.965 37.555 90.155 37.995 ;
        RECT 90.325 37.615 91.395 37.785 ;
        RECT 88.025 36.895 88.195 37.075 ;
        RECT 85.305 36.075 85.700 36.245 ;
        RECT 85.870 36.115 86.335 36.505 ;
        RECT 86.505 36.725 88.195 36.895 ;
        RECT 85.530 35.945 85.700 36.075 ;
        RECT 86.505 35.945 86.675 36.725 ;
        RECT 88.365 36.555 88.535 37.245 ;
        RECT 87.035 36.385 88.535 36.555 ;
        RECT 88.725 36.585 88.935 37.375 ;
        RECT 89.105 36.755 89.455 37.375 ;
        RECT 89.625 36.765 89.795 37.545 ;
        RECT 90.325 37.385 90.495 37.615 ;
        RECT 89.965 37.215 90.495 37.385 ;
        RECT 89.965 36.935 90.185 37.215 ;
        RECT 90.665 37.045 90.905 37.445 ;
        RECT 89.625 36.595 90.030 36.765 ;
        RECT 90.365 36.675 90.905 37.045 ;
        RECT 91.075 37.260 91.395 37.615 ;
        RECT 91.640 37.535 91.945 37.995 ;
        RECT 92.115 37.285 92.370 37.815 ;
        RECT 91.075 37.085 91.400 37.260 ;
        RECT 91.075 36.785 91.990 37.085 ;
        RECT 91.250 36.755 91.990 36.785 ;
        RECT 88.725 36.425 89.400 36.585 ;
        RECT 89.860 36.505 90.030 36.595 ;
        RECT 88.725 36.415 89.690 36.425 ;
        RECT 88.365 36.245 88.535 36.385 ;
        RECT 85.110 35.445 85.360 35.905 ;
        RECT 85.530 35.615 85.780 35.945 ;
        RECT 85.995 35.615 86.675 35.945 ;
        RECT 86.845 36.045 87.920 36.215 ;
        RECT 88.365 36.075 88.925 36.245 ;
        RECT 89.230 36.125 89.690 36.415 ;
        RECT 89.860 36.335 91.080 36.505 ;
        RECT 86.845 35.705 87.015 36.045 ;
        RECT 87.250 35.445 87.580 35.875 ;
        RECT 87.750 35.705 87.920 36.045 ;
        RECT 88.215 35.445 88.585 35.905 ;
        RECT 88.755 35.615 88.925 36.075 ;
        RECT 89.860 35.955 90.030 36.335 ;
        RECT 91.250 36.165 91.420 36.755 ;
        RECT 92.160 36.635 92.370 37.285 ;
        RECT 89.160 35.615 90.030 35.955 ;
        RECT 90.620 35.995 91.420 36.165 ;
        RECT 90.200 35.445 90.450 35.905 ;
        RECT 90.620 35.705 90.790 35.995 ;
        RECT 90.970 35.445 91.300 35.825 ;
        RECT 91.640 35.445 91.945 36.585 ;
        RECT 92.115 35.755 92.370 36.635 ;
        RECT 92.550 37.285 92.805 37.815 ;
        RECT 92.975 37.535 93.280 37.995 ;
        RECT 93.525 37.615 94.595 37.785 ;
        RECT 92.550 36.635 92.760 37.285 ;
        RECT 93.525 37.260 93.845 37.615 ;
        RECT 93.520 37.085 93.845 37.260 ;
        RECT 92.930 36.785 93.845 37.085 ;
        RECT 94.015 37.045 94.255 37.445 ;
        RECT 94.425 37.385 94.595 37.615 ;
        RECT 94.765 37.555 94.955 37.995 ;
        RECT 95.125 37.545 96.075 37.825 ;
        RECT 96.295 37.635 96.645 37.805 ;
        RECT 94.425 37.215 94.955 37.385 ;
        RECT 92.930 36.755 93.670 36.785 ;
        RECT 92.550 35.755 92.805 36.635 ;
        RECT 92.975 35.445 93.280 36.585 ;
        RECT 93.500 36.165 93.670 36.755 ;
        RECT 94.015 36.675 94.555 37.045 ;
        RECT 94.735 36.935 94.955 37.215 ;
        RECT 95.125 36.765 95.295 37.545 ;
        RECT 94.890 36.595 95.295 36.765 ;
        RECT 95.465 36.755 95.815 37.375 ;
        RECT 94.890 36.505 95.060 36.595 ;
        RECT 95.985 36.585 96.195 37.375 ;
        RECT 93.840 36.335 95.060 36.505 ;
        RECT 95.520 36.425 96.195 36.585 ;
        RECT 93.500 35.995 94.300 36.165 ;
        RECT 93.620 35.445 93.950 35.825 ;
        RECT 94.130 35.705 94.300 35.995 ;
        RECT 94.890 35.955 95.060 36.335 ;
        RECT 95.230 36.415 96.195 36.425 ;
        RECT 96.385 37.245 96.645 37.635 ;
        RECT 96.855 37.535 97.185 37.995 ;
        RECT 98.060 37.605 98.915 37.775 ;
        RECT 99.120 37.605 99.615 37.775 ;
        RECT 99.785 37.635 100.115 37.995 ;
        RECT 96.385 36.555 96.555 37.245 ;
        RECT 96.725 36.895 96.895 37.075 ;
        RECT 97.065 37.065 97.855 37.315 ;
        RECT 98.060 36.895 98.230 37.605 ;
        RECT 98.400 37.095 98.755 37.315 ;
        RECT 96.725 36.725 98.415 36.895 ;
        RECT 95.230 36.125 95.690 36.415 ;
        RECT 96.385 36.385 97.885 36.555 ;
        RECT 96.385 36.245 96.555 36.385 ;
        RECT 95.995 36.075 96.555 36.245 ;
        RECT 94.470 35.445 94.720 35.905 ;
        RECT 94.890 35.615 95.760 35.955 ;
        RECT 95.995 35.615 96.165 36.075 ;
        RECT 97.000 36.045 98.075 36.215 ;
        RECT 96.335 35.445 96.705 35.905 ;
        RECT 97.000 35.705 97.170 36.045 ;
        RECT 97.340 35.445 97.670 35.875 ;
        RECT 97.905 35.705 98.075 36.045 ;
        RECT 98.245 35.945 98.415 36.725 ;
        RECT 98.585 36.505 98.755 37.095 ;
        RECT 98.925 36.695 99.275 37.315 ;
        RECT 98.585 36.115 99.050 36.505 ;
        RECT 99.445 36.245 99.615 37.605 ;
        RECT 99.785 36.415 100.245 37.465 ;
        RECT 99.220 36.075 99.615 36.245 ;
        RECT 99.220 35.945 99.390 36.075 ;
        RECT 98.245 35.615 98.925 35.945 ;
        RECT 99.140 35.615 99.390 35.945 ;
        RECT 99.560 35.445 99.810 35.905 ;
        RECT 99.980 35.630 100.305 36.415 ;
        RECT 100.475 35.615 100.645 37.735 ;
        RECT 100.815 37.615 101.145 37.995 ;
        RECT 101.315 37.445 101.570 37.735 ;
        RECT 100.820 37.275 101.570 37.445 ;
        RECT 100.820 36.285 101.050 37.275 ;
        RECT 101.745 37.225 103.415 37.995 ;
        RECT 101.220 36.455 101.570 37.105 ;
        RECT 101.745 36.705 102.495 37.225 ;
        RECT 104.105 37.175 104.315 37.995 ;
        RECT 104.485 37.195 104.815 37.825 ;
        RECT 102.665 36.535 103.415 37.055 ;
        RECT 104.485 36.595 104.735 37.195 ;
        RECT 104.985 37.175 105.215 37.995 ;
        RECT 105.425 37.225 108.015 37.995 ;
        RECT 108.645 37.270 108.935 37.995 ;
        RECT 109.105 37.450 114.450 37.995 ;
        RECT 114.625 37.450 119.970 37.995 ;
        RECT 104.905 36.755 105.235 37.005 ;
        RECT 105.425 36.705 106.635 37.225 ;
        RECT 100.820 36.115 101.570 36.285 ;
        RECT 100.815 35.445 101.145 35.945 ;
        RECT 101.315 35.615 101.570 36.115 ;
        RECT 101.745 35.445 103.415 36.535 ;
        RECT 104.105 35.445 104.315 36.585 ;
        RECT 104.485 35.615 104.815 36.595 ;
        RECT 104.985 35.445 105.215 36.585 ;
        RECT 106.805 36.535 108.015 37.055 ;
        RECT 110.690 36.620 111.030 37.450 ;
        RECT 105.425 35.445 108.015 36.535 ;
        RECT 108.645 35.445 108.935 36.610 ;
        RECT 112.510 35.880 112.860 37.130 ;
        RECT 116.210 36.620 116.550 37.450 ;
        RECT 120.145 37.225 123.655 37.995 ;
        RECT 124.285 37.245 125.495 37.995 ;
        RECT 118.030 35.880 118.380 37.130 ;
        RECT 120.145 36.705 121.795 37.225 ;
        RECT 121.965 36.535 123.655 37.055 ;
        RECT 109.105 35.445 114.450 35.880 ;
        RECT 114.625 35.445 119.970 35.880 ;
        RECT 120.145 35.445 123.655 36.535 ;
        RECT 124.285 36.535 124.805 37.075 ;
        RECT 124.975 36.705 125.495 37.245 ;
        RECT 124.285 35.445 125.495 36.535 ;
        RECT 5.520 35.275 125.580 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.840 12.330 35.275 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 8.570 33.270 8.910 34.100 ;
        RECT 10.390 33.590 10.740 34.840 ;
        RECT 13.515 34.345 13.685 35.105 ;
        RECT 13.865 34.515 14.195 35.275 ;
        RECT 13.515 34.175 14.180 34.345 ;
        RECT 14.365 34.200 14.635 35.105 ;
        RECT 14.010 34.030 14.180 34.175 ;
        RECT 13.445 33.625 13.775 33.995 ;
        RECT 14.010 33.700 14.295 34.030 ;
        RECT 14.010 33.445 14.180 33.700 ;
        RECT 13.515 33.275 14.180 33.445 ;
        RECT 14.465 33.400 14.635 34.200 ;
        RECT 6.985 32.725 12.330 33.270 ;
        RECT 13.515 32.895 13.685 33.275 ;
        RECT 13.865 32.725 14.195 33.105 ;
        RECT 14.375 32.895 14.635 33.400 ;
        RECT 14.805 34.135 15.190 35.105 ;
        RECT 15.360 34.815 15.685 35.275 ;
        RECT 16.205 34.645 16.485 35.105 ;
        RECT 15.360 34.425 16.485 34.645 ;
        RECT 14.805 33.465 15.085 34.135 ;
        RECT 15.360 33.965 15.810 34.425 ;
        RECT 16.675 34.255 17.075 35.105 ;
        RECT 17.475 34.815 17.745 35.275 ;
        RECT 17.915 34.645 18.200 35.105 ;
        RECT 15.255 33.635 15.810 33.965 ;
        RECT 15.980 33.695 17.075 34.255 ;
        RECT 15.360 33.525 15.810 33.635 ;
        RECT 14.805 32.895 15.190 33.465 ;
        RECT 15.360 33.355 16.485 33.525 ;
        RECT 15.360 32.725 15.685 33.185 ;
        RECT 16.205 32.895 16.485 33.355 ;
        RECT 16.675 32.895 17.075 33.695 ;
        RECT 17.245 34.425 18.200 34.645 ;
        RECT 17.245 33.525 17.455 34.425 ;
        RECT 17.625 33.695 18.315 34.255 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 19.870 34.135 20.205 35.105 ;
        RECT 20.375 34.135 20.545 35.275 ;
        RECT 20.715 34.935 22.745 35.105 ;
        RECT 17.245 33.355 18.200 33.525 ;
        RECT 19.870 33.465 20.040 34.135 ;
        RECT 20.715 33.965 20.885 34.935 ;
        RECT 20.210 33.635 20.465 33.965 ;
        RECT 20.690 33.635 20.885 33.965 ;
        RECT 21.055 34.595 22.180 34.765 ;
        RECT 20.295 33.465 20.465 33.635 ;
        RECT 21.055 33.465 21.225 34.595 ;
        RECT 17.475 32.725 17.745 33.185 ;
        RECT 17.915 32.895 18.200 33.355 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 19.870 32.895 20.125 33.465 ;
        RECT 20.295 33.295 21.225 33.465 ;
        RECT 21.395 34.255 22.405 34.425 ;
        RECT 21.395 33.455 21.565 34.255 ;
        RECT 21.770 33.575 22.045 34.055 ;
        RECT 21.765 33.405 22.045 33.575 ;
        RECT 21.050 33.260 21.225 33.295 ;
        RECT 20.295 32.725 20.625 33.125 ;
        RECT 21.050 32.895 21.580 33.260 ;
        RECT 21.770 32.895 22.045 33.405 ;
        RECT 22.215 32.895 22.405 34.255 ;
        RECT 22.575 34.270 22.745 34.935 ;
        RECT 22.915 34.515 23.085 35.275 ;
        RECT 23.320 34.515 23.835 34.925 ;
        RECT 22.575 34.080 23.325 34.270 ;
        RECT 23.495 33.705 23.835 34.515 ;
        RECT 22.605 33.535 23.835 33.705 ;
        RECT 24.005 34.200 24.275 35.105 ;
        RECT 24.445 34.515 24.775 35.275 ;
        RECT 24.955 34.345 25.125 35.105 ;
        RECT 22.585 32.725 23.095 33.260 ;
        RECT 23.315 32.930 23.560 33.535 ;
        RECT 24.005 33.400 24.175 34.200 ;
        RECT 24.460 34.175 25.125 34.345 ;
        RECT 25.385 34.185 27.055 35.275 ;
        RECT 24.460 34.030 24.630 34.175 ;
        RECT 24.345 33.700 24.630 34.030 ;
        RECT 24.460 33.445 24.630 33.700 ;
        RECT 24.865 33.625 25.195 33.995 ;
        RECT 25.385 33.495 26.135 34.015 ;
        RECT 26.305 33.665 27.055 34.185 ;
        RECT 27.230 34.085 27.485 34.965 ;
        RECT 27.655 34.135 27.960 35.275 ;
        RECT 28.300 34.895 28.630 35.275 ;
        RECT 28.810 34.725 28.980 35.015 ;
        RECT 29.150 34.815 29.400 35.275 ;
        RECT 28.180 34.555 28.980 34.725 ;
        RECT 29.570 34.765 30.440 35.105 ;
        RECT 24.005 32.895 24.265 33.400 ;
        RECT 24.460 33.275 25.125 33.445 ;
        RECT 24.445 32.725 24.775 33.105 ;
        RECT 24.955 32.895 25.125 33.275 ;
        RECT 25.385 32.725 27.055 33.495 ;
        RECT 27.230 33.435 27.440 34.085 ;
        RECT 28.180 33.965 28.350 34.555 ;
        RECT 29.570 34.385 29.740 34.765 ;
        RECT 30.675 34.645 30.845 35.105 ;
        RECT 31.015 34.815 31.385 35.275 ;
        RECT 31.680 34.675 31.850 35.015 ;
        RECT 32.020 34.845 32.350 35.275 ;
        RECT 32.585 34.675 32.755 35.015 ;
        RECT 28.520 34.215 29.740 34.385 ;
        RECT 29.910 34.305 30.370 34.595 ;
        RECT 30.675 34.475 31.235 34.645 ;
        RECT 31.680 34.505 32.755 34.675 ;
        RECT 32.925 34.775 33.605 35.105 ;
        RECT 33.820 34.775 34.070 35.105 ;
        RECT 34.240 34.815 34.490 35.275 ;
        RECT 31.065 34.335 31.235 34.475 ;
        RECT 29.910 34.295 30.875 34.305 ;
        RECT 29.570 34.125 29.740 34.215 ;
        RECT 30.200 34.135 30.875 34.295 ;
        RECT 27.610 33.935 28.350 33.965 ;
        RECT 27.610 33.635 28.525 33.935 ;
        RECT 28.200 33.460 28.525 33.635 ;
        RECT 27.230 32.905 27.485 33.435 ;
        RECT 27.655 32.725 27.960 33.185 ;
        RECT 28.205 33.105 28.525 33.460 ;
        RECT 28.695 33.675 29.235 34.045 ;
        RECT 29.570 33.955 29.975 34.125 ;
        RECT 28.695 33.275 28.935 33.675 ;
        RECT 29.415 33.505 29.635 33.785 ;
        RECT 29.105 33.335 29.635 33.505 ;
        RECT 29.105 33.105 29.275 33.335 ;
        RECT 29.805 33.175 29.975 33.955 ;
        RECT 30.145 33.345 30.495 33.965 ;
        RECT 30.665 33.345 30.875 34.135 ;
        RECT 31.065 34.165 32.565 34.335 ;
        RECT 31.065 33.475 31.235 34.165 ;
        RECT 32.925 33.995 33.095 34.775 ;
        RECT 33.900 34.645 34.070 34.775 ;
        RECT 31.405 33.825 33.095 33.995 ;
        RECT 33.265 34.215 33.730 34.605 ;
        RECT 33.900 34.475 34.295 34.645 ;
        RECT 31.405 33.645 31.575 33.825 ;
        RECT 28.205 32.935 29.275 33.105 ;
        RECT 29.445 32.725 29.635 33.165 ;
        RECT 29.805 32.895 30.755 33.175 ;
        RECT 31.065 33.085 31.325 33.475 ;
        RECT 31.745 33.405 32.535 33.655 ;
        RECT 30.975 32.915 31.325 33.085 ;
        RECT 31.535 32.725 31.865 33.185 ;
        RECT 32.740 33.115 32.910 33.825 ;
        RECT 33.265 33.625 33.435 34.215 ;
        RECT 33.080 33.405 33.435 33.625 ;
        RECT 33.605 33.405 33.955 34.025 ;
        RECT 34.125 33.115 34.295 34.475 ;
        RECT 34.660 34.305 34.985 35.090 ;
        RECT 34.465 33.255 34.925 34.305 ;
        RECT 32.740 32.945 33.595 33.115 ;
        RECT 33.800 32.945 34.295 33.115 ;
        RECT 34.465 32.725 34.795 33.085 ;
        RECT 35.155 32.985 35.325 35.105 ;
        RECT 35.495 34.775 35.825 35.275 ;
        RECT 35.995 34.605 36.250 35.105 ;
        RECT 35.500 34.435 36.250 34.605 ;
        RECT 35.500 33.445 35.730 34.435 ;
        RECT 35.900 33.615 36.250 34.265 ;
        RECT 36.425 34.185 39.935 35.275 ;
        RECT 36.425 33.495 38.075 34.015 ;
        RECT 38.245 33.665 39.935 34.185 ;
        RECT 40.605 34.135 40.835 35.275 ;
        RECT 41.005 34.125 41.335 35.105 ;
        RECT 41.505 34.135 41.715 35.275 ;
        RECT 41.945 34.185 43.615 35.275 ;
        RECT 40.585 33.715 40.915 33.965 ;
        RECT 35.500 33.275 36.250 33.445 ;
        RECT 35.495 32.725 35.825 33.105 ;
        RECT 35.995 32.985 36.250 33.275 ;
        RECT 36.425 32.725 39.935 33.495 ;
        RECT 40.605 32.725 40.835 33.545 ;
        RECT 41.085 33.525 41.335 34.125 ;
        RECT 41.005 32.895 41.335 33.525 ;
        RECT 41.505 32.725 41.715 33.545 ;
        RECT 41.945 33.495 42.695 34.015 ;
        RECT 42.865 33.665 43.615 34.185 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 44.705 34.840 50.050 35.275 ;
        RECT 41.945 32.725 43.615 33.495 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 46.290 33.270 46.630 34.100 ;
        RECT 48.110 33.590 48.460 34.840 ;
        RECT 50.225 34.185 51.895 35.275 ;
        RECT 52.070 34.605 52.325 35.105 ;
        RECT 52.495 34.775 52.825 35.275 ;
        RECT 52.070 34.435 52.820 34.605 ;
        RECT 50.225 33.495 50.975 34.015 ;
        RECT 51.145 33.665 51.895 34.185 ;
        RECT 52.070 33.615 52.420 34.265 ;
        RECT 44.705 32.725 50.050 33.270 ;
        RECT 50.225 32.725 51.895 33.495 ;
        RECT 52.590 33.445 52.820 34.435 ;
        RECT 52.070 33.275 52.820 33.445 ;
        RECT 52.070 32.985 52.325 33.275 ;
        RECT 52.495 32.725 52.825 33.105 ;
        RECT 52.995 32.985 53.165 35.105 ;
        RECT 53.335 34.305 53.660 35.090 ;
        RECT 53.830 34.815 54.080 35.275 ;
        RECT 54.250 34.775 54.500 35.105 ;
        RECT 54.715 34.775 55.395 35.105 ;
        RECT 54.250 34.645 54.420 34.775 ;
        RECT 54.025 34.475 54.420 34.645 ;
        RECT 53.395 33.255 53.855 34.305 ;
        RECT 54.025 33.115 54.195 34.475 ;
        RECT 54.590 34.215 55.055 34.605 ;
        RECT 54.365 33.405 54.715 34.025 ;
        RECT 54.885 33.625 55.055 34.215 ;
        RECT 55.225 33.995 55.395 34.775 ;
        RECT 55.565 34.675 55.735 35.015 ;
        RECT 55.970 34.845 56.300 35.275 ;
        RECT 56.470 34.675 56.640 35.015 ;
        RECT 56.935 34.815 57.305 35.275 ;
        RECT 55.565 34.505 56.640 34.675 ;
        RECT 57.475 34.645 57.645 35.105 ;
        RECT 57.880 34.765 58.750 35.105 ;
        RECT 58.920 34.815 59.170 35.275 ;
        RECT 57.085 34.475 57.645 34.645 ;
        RECT 57.085 34.335 57.255 34.475 ;
        RECT 55.755 34.165 57.255 34.335 ;
        RECT 57.950 34.305 58.410 34.595 ;
        RECT 55.225 33.825 56.915 33.995 ;
        RECT 54.885 33.405 55.240 33.625 ;
        RECT 55.410 33.115 55.580 33.825 ;
        RECT 55.785 33.405 56.575 33.655 ;
        RECT 56.745 33.645 56.915 33.825 ;
        RECT 57.085 33.475 57.255 34.165 ;
        RECT 53.525 32.725 53.855 33.085 ;
        RECT 54.025 32.945 54.520 33.115 ;
        RECT 54.725 32.945 55.580 33.115 ;
        RECT 56.455 32.725 56.785 33.185 ;
        RECT 56.995 33.085 57.255 33.475 ;
        RECT 57.445 34.295 58.410 34.305 ;
        RECT 58.580 34.385 58.750 34.765 ;
        RECT 59.340 34.725 59.510 35.015 ;
        RECT 59.690 34.895 60.020 35.275 ;
        RECT 59.340 34.555 60.140 34.725 ;
        RECT 57.445 34.135 58.120 34.295 ;
        RECT 58.580 34.215 59.800 34.385 ;
        RECT 57.445 33.345 57.655 34.135 ;
        RECT 58.580 34.125 58.750 34.215 ;
        RECT 57.825 33.345 58.175 33.965 ;
        RECT 58.345 33.955 58.750 34.125 ;
        RECT 58.345 33.175 58.515 33.955 ;
        RECT 58.685 33.505 58.905 33.785 ;
        RECT 59.085 33.675 59.625 34.045 ;
        RECT 59.970 33.965 60.140 34.555 ;
        RECT 60.360 34.135 60.665 35.275 ;
        RECT 60.835 34.085 61.090 34.965 ;
        RECT 61.355 34.345 61.525 35.105 ;
        RECT 61.740 34.515 62.070 35.275 ;
        RECT 61.355 34.175 62.070 34.345 ;
        RECT 62.240 34.200 62.495 35.105 ;
        RECT 59.970 33.935 60.710 33.965 ;
        RECT 58.685 33.335 59.215 33.505 ;
        RECT 56.995 32.915 57.345 33.085 ;
        RECT 57.565 32.895 58.515 33.175 ;
        RECT 58.685 32.725 58.875 33.165 ;
        RECT 59.045 33.105 59.215 33.335 ;
        RECT 59.385 33.275 59.625 33.675 ;
        RECT 59.795 33.635 60.710 33.935 ;
        RECT 59.795 33.460 60.120 33.635 ;
        RECT 59.795 33.105 60.115 33.460 ;
        RECT 60.880 33.435 61.090 34.085 ;
        RECT 61.265 33.625 61.620 33.995 ;
        RECT 61.900 33.965 62.070 34.175 ;
        RECT 61.900 33.635 62.155 33.965 ;
        RECT 61.900 33.445 62.070 33.635 ;
        RECT 62.325 33.470 62.495 34.200 ;
        RECT 62.670 34.125 62.930 35.275 ;
        RECT 63.105 34.840 68.450 35.275 ;
        RECT 59.045 32.935 60.115 33.105 ;
        RECT 60.360 32.725 60.665 33.185 ;
        RECT 60.835 32.905 61.090 33.435 ;
        RECT 61.355 33.275 62.070 33.445 ;
        RECT 61.355 32.895 61.525 33.275 ;
        RECT 61.740 32.725 62.070 33.105 ;
        RECT 62.240 32.895 62.495 33.470 ;
        RECT 62.670 32.725 62.930 33.565 ;
        RECT 64.690 33.270 65.030 34.100 ;
        RECT 66.510 33.590 66.860 34.840 ;
        RECT 68.625 34.185 69.835 35.275 ;
        RECT 68.625 33.475 69.145 34.015 ;
        RECT 69.315 33.645 69.835 34.185 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 70.465 34.840 75.810 35.275 ;
        RECT 75.985 34.840 81.330 35.275 ;
        RECT 63.105 32.725 68.450 33.270 ;
        RECT 68.625 32.725 69.835 33.475 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 72.050 33.270 72.390 34.100 ;
        RECT 73.870 33.590 74.220 34.840 ;
        RECT 77.570 33.270 77.910 34.100 ;
        RECT 79.390 33.590 79.740 34.840 ;
        RECT 81.505 34.185 84.095 35.275 ;
        RECT 84.270 34.605 84.525 35.105 ;
        RECT 84.695 34.775 85.025 35.275 ;
        RECT 84.270 34.435 85.020 34.605 ;
        RECT 81.505 33.495 82.715 34.015 ;
        RECT 82.885 33.665 84.095 34.185 ;
        RECT 84.270 33.615 84.620 34.265 ;
        RECT 70.465 32.725 75.810 33.270 ;
        RECT 75.985 32.725 81.330 33.270 ;
        RECT 81.505 32.725 84.095 33.495 ;
        RECT 84.790 33.445 85.020 34.435 ;
        RECT 84.270 33.275 85.020 33.445 ;
        RECT 84.270 32.985 84.525 33.275 ;
        RECT 84.695 32.725 85.025 33.105 ;
        RECT 85.195 32.985 85.365 35.105 ;
        RECT 85.535 34.305 85.860 35.090 ;
        RECT 86.030 34.815 86.280 35.275 ;
        RECT 86.450 34.775 86.700 35.105 ;
        RECT 86.915 34.775 87.595 35.105 ;
        RECT 86.450 34.645 86.620 34.775 ;
        RECT 86.225 34.475 86.620 34.645 ;
        RECT 85.595 33.255 86.055 34.305 ;
        RECT 86.225 33.115 86.395 34.475 ;
        RECT 86.790 34.215 87.255 34.605 ;
        RECT 86.565 33.405 86.915 34.025 ;
        RECT 87.085 33.625 87.255 34.215 ;
        RECT 87.425 33.995 87.595 34.775 ;
        RECT 87.765 34.675 87.935 35.015 ;
        RECT 88.170 34.845 88.500 35.275 ;
        RECT 88.670 34.675 88.840 35.015 ;
        RECT 89.135 34.815 89.505 35.275 ;
        RECT 87.765 34.505 88.840 34.675 ;
        RECT 89.675 34.645 89.845 35.105 ;
        RECT 90.080 34.765 90.950 35.105 ;
        RECT 91.120 34.815 91.370 35.275 ;
        RECT 89.285 34.475 89.845 34.645 ;
        RECT 89.285 34.335 89.455 34.475 ;
        RECT 87.955 34.165 89.455 34.335 ;
        RECT 90.150 34.305 90.610 34.595 ;
        RECT 87.425 33.825 89.115 33.995 ;
        RECT 87.085 33.405 87.440 33.625 ;
        RECT 87.610 33.115 87.780 33.825 ;
        RECT 87.985 33.405 88.775 33.655 ;
        RECT 88.945 33.645 89.115 33.825 ;
        RECT 89.285 33.475 89.455 34.165 ;
        RECT 85.725 32.725 86.055 33.085 ;
        RECT 86.225 32.945 86.720 33.115 ;
        RECT 86.925 32.945 87.780 33.115 ;
        RECT 88.655 32.725 88.985 33.185 ;
        RECT 89.195 33.085 89.455 33.475 ;
        RECT 89.645 34.295 90.610 34.305 ;
        RECT 90.780 34.385 90.950 34.765 ;
        RECT 91.540 34.725 91.710 35.015 ;
        RECT 91.890 34.895 92.220 35.275 ;
        RECT 91.540 34.555 92.340 34.725 ;
        RECT 89.645 34.135 90.320 34.295 ;
        RECT 90.780 34.215 92.000 34.385 ;
        RECT 89.645 33.345 89.855 34.135 ;
        RECT 90.780 34.125 90.950 34.215 ;
        RECT 90.025 33.345 90.375 33.965 ;
        RECT 90.545 33.955 90.950 34.125 ;
        RECT 90.545 33.175 90.715 33.955 ;
        RECT 90.885 33.505 91.105 33.785 ;
        RECT 91.285 33.675 91.825 34.045 ;
        RECT 92.170 33.965 92.340 34.555 ;
        RECT 92.560 34.135 92.865 35.275 ;
        RECT 93.035 34.085 93.290 34.965 ;
        RECT 94.015 34.345 94.185 35.105 ;
        RECT 94.365 34.515 94.695 35.275 ;
        RECT 94.015 34.175 94.680 34.345 ;
        RECT 94.865 34.200 95.135 35.105 ;
        RECT 92.170 33.935 92.910 33.965 ;
        RECT 90.885 33.335 91.415 33.505 ;
        RECT 89.195 32.915 89.545 33.085 ;
        RECT 89.765 32.895 90.715 33.175 ;
        RECT 90.885 32.725 91.075 33.165 ;
        RECT 91.245 33.105 91.415 33.335 ;
        RECT 91.585 33.275 91.825 33.675 ;
        RECT 91.995 33.635 92.910 33.935 ;
        RECT 91.995 33.460 92.320 33.635 ;
        RECT 91.995 33.105 92.315 33.460 ;
        RECT 93.080 33.435 93.290 34.085 ;
        RECT 94.510 34.030 94.680 34.175 ;
        RECT 93.945 33.625 94.275 33.995 ;
        RECT 94.510 33.700 94.795 34.030 ;
        RECT 94.510 33.445 94.680 33.700 ;
        RECT 91.245 32.935 92.315 33.105 ;
        RECT 92.560 32.725 92.865 33.185 ;
        RECT 93.035 32.905 93.290 33.435 ;
        RECT 94.015 33.275 94.680 33.445 ;
        RECT 94.965 33.400 95.135 34.200 ;
        RECT 95.765 34.110 96.055 35.275 ;
        RECT 97.235 34.345 97.405 35.105 ;
        RECT 97.585 34.515 97.915 35.275 ;
        RECT 97.235 34.175 97.900 34.345 ;
        RECT 98.085 34.200 98.355 35.105 ;
        RECT 98.525 34.840 103.870 35.275 ;
        RECT 104.045 34.840 109.390 35.275 ;
        RECT 109.565 34.840 114.910 35.275 ;
        RECT 115.085 34.840 120.430 35.275 ;
        RECT 97.730 34.030 97.900 34.175 ;
        RECT 97.165 33.625 97.495 33.995 ;
        RECT 97.730 33.700 98.015 34.030 ;
        RECT 94.015 32.895 94.185 33.275 ;
        RECT 94.365 32.725 94.695 33.105 ;
        RECT 94.875 32.895 95.135 33.400 ;
        RECT 95.765 32.725 96.055 33.450 ;
        RECT 97.730 33.445 97.900 33.700 ;
        RECT 97.235 33.275 97.900 33.445 ;
        RECT 98.185 33.400 98.355 34.200 ;
        RECT 97.235 32.895 97.405 33.275 ;
        RECT 97.585 32.725 97.915 33.105 ;
        RECT 98.095 32.895 98.355 33.400 ;
        RECT 100.110 33.270 100.450 34.100 ;
        RECT 101.930 33.590 102.280 34.840 ;
        RECT 105.630 33.270 105.970 34.100 ;
        RECT 107.450 33.590 107.800 34.840 ;
        RECT 111.150 33.270 111.490 34.100 ;
        RECT 112.970 33.590 113.320 34.840 ;
        RECT 116.670 33.270 117.010 34.100 ;
        RECT 118.490 33.590 118.840 34.840 ;
        RECT 121.525 34.110 121.815 35.275 ;
        RECT 121.985 34.185 123.655 35.275 ;
        RECT 121.985 33.495 122.735 34.015 ;
        RECT 122.905 33.665 123.655 34.185 ;
        RECT 124.285 34.185 125.495 35.275 ;
        RECT 124.285 33.645 124.805 34.185 ;
        RECT 98.525 32.725 103.870 33.270 ;
        RECT 104.045 32.725 109.390 33.270 ;
        RECT 109.565 32.725 114.910 33.270 ;
        RECT 115.085 32.725 120.430 33.270 ;
        RECT 121.525 32.725 121.815 33.450 ;
        RECT 121.985 32.725 123.655 33.495 ;
        RECT 124.975 33.475 125.495 34.015 ;
        RECT 124.285 32.725 125.495 33.475 ;
        RECT 5.520 32.555 125.580 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 6.985 32.010 12.330 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 8.570 31.180 8.910 32.010 ;
        RECT 12.505 31.785 16.015 32.555 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 10.390 30.440 10.740 31.690 ;
        RECT 12.505 31.265 14.155 31.785 ;
        RECT 17.165 31.735 17.375 32.555 ;
        RECT 17.545 31.755 17.875 32.385 ;
        RECT 14.325 31.095 16.015 31.615 ;
        RECT 17.545 31.155 17.795 31.755 ;
        RECT 18.045 31.735 18.275 32.555 ;
        RECT 18.490 32.005 18.745 32.295 ;
        RECT 18.915 32.175 19.245 32.555 ;
        RECT 18.490 31.835 19.240 32.005 ;
        RECT 17.965 31.315 18.295 31.565 ;
        RECT 6.985 30.005 12.330 30.440 ;
        RECT 12.505 30.005 16.015 31.095 ;
        RECT 17.165 30.005 17.375 31.145 ;
        RECT 17.545 30.175 17.875 31.155 ;
        RECT 18.045 30.005 18.275 31.145 ;
        RECT 18.490 31.015 18.840 31.665 ;
        RECT 19.010 30.845 19.240 31.835 ;
        RECT 18.490 30.675 19.240 30.845 ;
        RECT 18.490 30.175 18.745 30.675 ;
        RECT 18.915 30.005 19.245 30.505 ;
        RECT 19.415 30.175 19.585 32.295 ;
        RECT 19.945 32.195 20.275 32.555 ;
        RECT 20.445 32.165 20.940 32.335 ;
        RECT 21.145 32.165 22.000 32.335 ;
        RECT 19.815 30.975 20.275 32.025 ;
        RECT 19.755 30.190 20.080 30.975 ;
        RECT 20.445 30.805 20.615 32.165 ;
        RECT 20.785 31.255 21.135 31.875 ;
        RECT 21.305 31.655 21.660 31.875 ;
        RECT 21.305 31.065 21.475 31.655 ;
        RECT 21.830 31.455 22.000 32.165 ;
        RECT 22.875 32.095 23.205 32.555 ;
        RECT 23.415 32.195 23.765 32.365 ;
        RECT 22.205 31.625 22.995 31.875 ;
        RECT 23.415 31.805 23.675 32.195 ;
        RECT 23.985 32.105 24.935 32.385 ;
        RECT 25.105 32.115 25.295 32.555 ;
        RECT 25.465 32.175 26.535 32.345 ;
        RECT 23.165 31.455 23.335 31.635 ;
        RECT 20.445 30.635 20.840 30.805 ;
        RECT 21.010 30.675 21.475 31.065 ;
        RECT 21.645 31.285 23.335 31.455 ;
        RECT 20.670 30.505 20.840 30.635 ;
        RECT 21.645 30.505 21.815 31.285 ;
        RECT 23.505 31.115 23.675 31.805 ;
        RECT 22.175 30.945 23.675 31.115 ;
        RECT 23.865 31.145 24.075 31.935 ;
        RECT 24.245 31.315 24.595 31.935 ;
        RECT 24.765 31.325 24.935 32.105 ;
        RECT 25.465 31.945 25.635 32.175 ;
        RECT 25.105 31.775 25.635 31.945 ;
        RECT 25.105 31.495 25.325 31.775 ;
        RECT 25.805 31.605 26.045 32.005 ;
        RECT 24.765 31.155 25.170 31.325 ;
        RECT 25.505 31.235 26.045 31.605 ;
        RECT 26.215 31.820 26.535 32.175 ;
        RECT 26.780 32.095 27.085 32.555 ;
        RECT 27.255 31.845 27.510 32.375 ;
        RECT 26.215 31.645 26.540 31.820 ;
        RECT 26.215 31.345 27.130 31.645 ;
        RECT 26.390 31.315 27.130 31.345 ;
        RECT 23.865 30.985 24.540 31.145 ;
        RECT 25.000 31.065 25.170 31.155 ;
        RECT 23.865 30.975 24.830 30.985 ;
        RECT 23.505 30.805 23.675 30.945 ;
        RECT 20.250 30.005 20.500 30.465 ;
        RECT 20.670 30.175 20.920 30.505 ;
        RECT 21.135 30.175 21.815 30.505 ;
        RECT 21.985 30.605 23.060 30.775 ;
        RECT 23.505 30.635 24.065 30.805 ;
        RECT 24.370 30.685 24.830 30.975 ;
        RECT 25.000 30.895 26.220 31.065 ;
        RECT 21.985 30.265 22.155 30.605 ;
        RECT 22.390 30.005 22.720 30.435 ;
        RECT 22.890 30.265 23.060 30.605 ;
        RECT 23.355 30.005 23.725 30.465 ;
        RECT 23.895 30.175 24.065 30.635 ;
        RECT 25.000 30.515 25.170 30.895 ;
        RECT 26.390 30.725 26.560 31.315 ;
        RECT 27.300 31.195 27.510 31.845 ;
        RECT 24.300 30.175 25.170 30.515 ;
        RECT 25.760 30.555 26.560 30.725 ;
        RECT 25.340 30.005 25.590 30.465 ;
        RECT 25.760 30.265 25.930 30.555 ;
        RECT 26.110 30.005 26.440 30.385 ;
        RECT 26.780 30.005 27.085 31.145 ;
        RECT 27.255 30.315 27.510 31.195 ;
        RECT 27.685 31.815 28.070 32.385 ;
        RECT 28.240 32.095 28.565 32.555 ;
        RECT 29.085 31.925 29.365 32.385 ;
        RECT 27.685 31.145 27.965 31.815 ;
        RECT 28.240 31.755 29.365 31.925 ;
        RECT 28.240 31.645 28.690 31.755 ;
        RECT 28.135 31.315 28.690 31.645 ;
        RECT 29.555 31.585 29.955 32.385 ;
        RECT 30.355 32.095 30.625 32.555 ;
        RECT 30.795 31.925 31.080 32.385 ;
        RECT 27.685 30.175 28.070 31.145 ;
        RECT 28.240 30.855 28.690 31.315 ;
        RECT 28.860 31.025 29.955 31.585 ;
        RECT 28.240 30.635 29.365 30.855 ;
        RECT 28.240 30.005 28.565 30.465 ;
        RECT 29.085 30.175 29.365 30.635 ;
        RECT 29.555 30.175 29.955 31.025 ;
        RECT 30.125 31.755 31.080 31.925 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 30.125 30.855 30.335 31.755 ;
        RECT 31.885 31.735 32.095 32.555 ;
        RECT 32.265 31.755 32.595 32.385 ;
        RECT 30.505 31.025 31.195 31.585 ;
        RECT 30.125 30.635 31.080 30.855 ;
        RECT 30.355 30.005 30.625 30.465 ;
        RECT 30.795 30.175 31.080 30.635 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 32.265 31.155 32.515 31.755 ;
        RECT 32.765 31.735 32.995 32.555 ;
        RECT 33.295 32.005 33.465 32.385 ;
        RECT 33.645 32.175 33.975 32.555 ;
        RECT 33.295 31.835 33.960 32.005 ;
        RECT 34.155 31.880 34.415 32.385 ;
        RECT 34.585 32.010 39.930 32.555 ;
        RECT 40.105 32.010 45.450 32.555 ;
        RECT 45.625 32.010 50.970 32.555 ;
        RECT 32.685 31.315 33.015 31.565 ;
        RECT 33.225 31.285 33.555 31.655 ;
        RECT 33.790 31.580 33.960 31.835 ;
        RECT 33.790 31.250 34.075 31.580 ;
        RECT 31.885 30.005 32.095 31.145 ;
        RECT 32.265 30.175 32.595 31.155 ;
        RECT 32.765 30.005 32.995 31.145 ;
        RECT 33.790 31.105 33.960 31.250 ;
        RECT 33.295 30.935 33.960 31.105 ;
        RECT 34.245 31.080 34.415 31.880 ;
        RECT 36.170 31.180 36.510 32.010 ;
        RECT 33.295 30.175 33.465 30.935 ;
        RECT 33.645 30.005 33.975 30.765 ;
        RECT 34.145 30.175 34.415 31.080 ;
        RECT 37.990 30.440 38.340 31.690 ;
        RECT 41.690 31.180 42.030 32.010 ;
        RECT 43.510 30.440 43.860 31.690 ;
        RECT 47.210 31.180 47.550 32.010 ;
        RECT 51.145 31.785 52.815 32.555 ;
        RECT 49.030 30.440 49.380 31.690 ;
        RECT 51.145 31.265 51.895 31.785 ;
        RECT 53.485 31.735 53.715 32.555 ;
        RECT 53.885 31.755 54.215 32.385 ;
        RECT 52.065 31.095 52.815 31.615 ;
        RECT 53.465 31.315 53.795 31.565 ;
        RECT 53.965 31.155 54.215 31.755 ;
        RECT 54.385 31.735 54.595 32.555 ;
        RECT 55.285 31.880 55.545 32.385 ;
        RECT 55.725 32.175 56.055 32.555 ;
        RECT 56.235 32.005 56.405 32.385 ;
        RECT 34.585 30.005 39.930 30.440 ;
        RECT 40.105 30.005 45.450 30.440 ;
        RECT 45.625 30.005 50.970 30.440 ;
        RECT 51.145 30.005 52.815 31.095 ;
        RECT 53.485 30.005 53.715 31.145 ;
        RECT 53.885 30.175 54.215 31.155 ;
        RECT 54.385 30.005 54.595 31.145 ;
        RECT 55.285 31.080 55.455 31.880 ;
        RECT 55.740 31.835 56.405 32.005 ;
        RECT 55.740 31.580 55.910 31.835 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 57.585 31.905 57.845 32.385 ;
        RECT 58.015 32.015 58.265 32.555 ;
        RECT 55.625 31.250 55.910 31.580 ;
        RECT 56.145 31.285 56.475 31.655 ;
        RECT 55.740 31.105 55.910 31.250 ;
        RECT 55.285 30.175 55.555 31.080 ;
        RECT 55.740 30.935 56.405 31.105 ;
        RECT 55.725 30.005 56.055 30.765 ;
        RECT 56.235 30.175 56.405 30.935 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 57.585 30.875 57.755 31.905 ;
        RECT 58.435 31.850 58.655 32.335 ;
        RECT 57.925 31.255 58.155 31.650 ;
        RECT 58.325 31.425 58.655 31.850 ;
        RECT 58.825 32.175 59.715 32.345 ;
        RECT 60.805 32.175 61.695 32.345 ;
        RECT 58.825 31.450 58.995 32.175 ;
        RECT 59.165 31.620 59.715 32.005 ;
        RECT 60.805 31.620 61.355 32.005 ;
        RECT 61.525 31.450 61.695 32.175 ;
        RECT 58.825 31.380 59.715 31.450 ;
        RECT 58.820 31.355 59.715 31.380 ;
        RECT 58.810 31.340 59.715 31.355 ;
        RECT 58.805 31.325 59.715 31.340 ;
        RECT 58.795 31.320 59.715 31.325 ;
        RECT 58.790 31.310 59.715 31.320 ;
        RECT 58.785 31.300 59.715 31.310 ;
        RECT 58.775 31.295 59.715 31.300 ;
        RECT 58.765 31.285 59.715 31.295 ;
        RECT 58.755 31.280 59.715 31.285 ;
        RECT 58.755 31.275 59.090 31.280 ;
        RECT 58.740 31.270 59.090 31.275 ;
        RECT 58.725 31.260 59.090 31.270 ;
        RECT 58.700 31.255 59.090 31.260 ;
        RECT 57.925 31.250 59.090 31.255 ;
        RECT 57.925 31.215 59.060 31.250 ;
        RECT 57.925 31.190 59.025 31.215 ;
        RECT 57.925 31.160 58.995 31.190 ;
        RECT 57.925 31.130 58.975 31.160 ;
        RECT 57.925 31.100 58.955 31.130 ;
        RECT 57.925 31.090 58.885 31.100 ;
        RECT 57.925 31.080 58.860 31.090 ;
        RECT 57.925 31.065 58.840 31.080 ;
        RECT 57.925 31.050 58.820 31.065 ;
        RECT 58.030 31.040 58.815 31.050 ;
        RECT 58.030 31.005 58.800 31.040 ;
        RECT 57.585 30.175 57.860 30.875 ;
        RECT 58.030 30.755 58.785 31.005 ;
        RECT 58.955 30.685 59.285 30.930 ;
        RECT 59.455 30.830 59.715 31.280 ;
        RECT 60.805 31.380 61.695 31.450 ;
        RECT 61.865 31.850 62.085 32.335 ;
        RECT 62.255 32.015 62.505 32.555 ;
        RECT 62.675 31.905 62.935 32.385 ;
        RECT 61.865 31.425 62.195 31.850 ;
        RECT 60.805 31.355 61.700 31.380 ;
        RECT 60.805 31.340 61.710 31.355 ;
        RECT 60.805 31.325 61.715 31.340 ;
        RECT 60.805 31.320 61.725 31.325 ;
        RECT 60.805 31.310 61.730 31.320 ;
        RECT 60.805 31.300 61.735 31.310 ;
        RECT 60.805 31.295 61.745 31.300 ;
        RECT 60.805 31.285 61.755 31.295 ;
        RECT 60.805 31.280 61.765 31.285 ;
        RECT 60.805 30.830 61.065 31.280 ;
        RECT 61.430 31.275 61.765 31.280 ;
        RECT 61.430 31.270 61.780 31.275 ;
        RECT 61.430 31.260 61.795 31.270 ;
        RECT 61.430 31.255 61.820 31.260 ;
        RECT 62.365 31.255 62.595 31.650 ;
        RECT 61.430 31.250 62.595 31.255 ;
        RECT 61.460 31.215 62.595 31.250 ;
        RECT 61.495 31.190 62.595 31.215 ;
        RECT 61.525 31.160 62.595 31.190 ;
        RECT 61.545 31.130 62.595 31.160 ;
        RECT 61.565 31.100 62.595 31.130 ;
        RECT 61.635 31.090 62.595 31.100 ;
        RECT 61.660 31.080 62.595 31.090 ;
        RECT 61.680 31.065 62.595 31.080 ;
        RECT 61.700 31.050 62.595 31.065 ;
        RECT 61.705 31.040 62.490 31.050 ;
        RECT 61.720 31.005 62.490 31.040 ;
        RECT 59.100 30.660 59.285 30.685 ;
        RECT 61.235 30.685 61.565 30.930 ;
        RECT 61.735 30.755 62.490 31.005 ;
        RECT 62.765 30.875 62.935 31.905 ;
        RECT 61.235 30.660 61.420 30.685 ;
        RECT 59.100 30.560 59.715 30.660 ;
        RECT 58.030 30.005 58.285 30.550 ;
        RECT 58.455 30.175 58.935 30.515 ;
        RECT 59.110 30.005 59.715 30.560 ;
        RECT 60.805 30.560 61.420 30.660 ;
        RECT 60.805 30.005 61.410 30.560 ;
        RECT 61.585 30.175 62.065 30.515 ;
        RECT 62.235 30.005 62.490 30.550 ;
        RECT 62.660 30.175 62.935 30.875 ;
        RECT 63.115 31.830 63.445 32.340 ;
        RECT 63.615 32.155 63.945 32.555 ;
        RECT 64.995 31.985 65.325 32.325 ;
        RECT 65.495 32.155 65.825 32.555 ;
        RECT 63.115 31.065 63.305 31.830 ;
        RECT 63.615 31.815 65.980 31.985 ;
        RECT 63.615 31.645 63.785 31.815 ;
        RECT 63.475 31.315 63.785 31.645 ;
        RECT 63.955 31.315 64.260 31.645 ;
        RECT 63.115 30.215 63.445 31.065 ;
        RECT 63.615 30.005 63.865 31.145 ;
        RECT 64.045 30.985 64.260 31.315 ;
        RECT 64.435 30.985 64.720 31.645 ;
        RECT 64.915 30.985 65.180 31.645 ;
        RECT 65.395 30.985 65.640 31.645 ;
        RECT 65.810 30.815 65.980 31.815 ;
        RECT 66.325 31.785 68.915 32.555 ;
        RECT 69.085 31.815 69.470 32.385 ;
        RECT 69.640 32.095 69.965 32.555 ;
        RECT 70.485 31.925 70.765 32.385 ;
        RECT 66.325 31.265 67.535 31.785 ;
        RECT 67.705 31.095 68.915 31.615 ;
        RECT 64.055 30.645 65.345 30.815 ;
        RECT 64.055 30.225 64.305 30.645 ;
        RECT 64.535 30.005 64.865 30.475 ;
        RECT 65.095 30.225 65.345 30.645 ;
        RECT 65.525 30.645 65.980 30.815 ;
        RECT 65.525 30.215 65.855 30.645 ;
        RECT 66.325 30.005 68.915 31.095 ;
        RECT 69.085 31.145 69.365 31.815 ;
        RECT 69.640 31.755 70.765 31.925 ;
        RECT 69.640 31.645 70.090 31.755 ;
        RECT 69.535 31.315 70.090 31.645 ;
        RECT 70.955 31.585 71.355 32.385 ;
        RECT 71.755 32.095 72.025 32.555 ;
        RECT 72.195 31.925 72.480 32.385 ;
        RECT 69.085 30.175 69.470 31.145 ;
        RECT 69.640 30.855 70.090 31.315 ;
        RECT 70.260 31.025 71.355 31.585 ;
        RECT 69.640 30.635 70.765 30.855 ;
        RECT 69.640 30.005 69.965 30.465 ;
        RECT 70.485 30.175 70.765 30.635 ;
        RECT 70.955 30.175 71.355 31.025 ;
        RECT 71.525 31.755 72.480 31.925 ;
        RECT 71.525 30.855 71.735 31.755 ;
        RECT 72.805 31.735 73.035 32.555 ;
        RECT 73.205 31.755 73.535 32.385 ;
        RECT 71.905 31.025 72.595 31.585 ;
        RECT 72.785 31.315 73.115 31.565 ;
        RECT 73.285 31.155 73.535 31.755 ;
        RECT 73.705 31.735 73.915 32.555 ;
        RECT 74.145 32.010 79.490 32.555 ;
        RECT 75.730 31.180 76.070 32.010 ;
        RECT 79.665 31.785 82.255 32.555 ;
        RECT 82.885 31.830 83.175 32.555 ;
        RECT 83.345 32.010 88.690 32.555 ;
        RECT 88.865 32.010 94.210 32.555 ;
        RECT 94.385 32.010 99.730 32.555 ;
        RECT 99.905 32.010 105.250 32.555 ;
        RECT 71.525 30.635 72.480 30.855 ;
        RECT 71.755 30.005 72.025 30.465 ;
        RECT 72.195 30.175 72.480 30.635 ;
        RECT 72.805 30.005 73.035 31.145 ;
        RECT 73.205 30.175 73.535 31.155 ;
        RECT 73.705 30.005 73.915 31.145 ;
        RECT 77.550 30.440 77.900 31.690 ;
        RECT 79.665 31.265 80.875 31.785 ;
        RECT 81.045 31.095 82.255 31.615 ;
        RECT 84.930 31.180 85.270 32.010 ;
        RECT 74.145 30.005 79.490 30.440 ;
        RECT 79.665 30.005 82.255 31.095 ;
        RECT 82.885 30.005 83.175 31.170 ;
        RECT 86.750 30.440 87.100 31.690 ;
        RECT 90.450 31.180 90.790 32.010 ;
        RECT 92.270 30.440 92.620 31.690 ;
        RECT 95.970 31.180 96.310 32.010 ;
        RECT 97.790 30.440 98.140 31.690 ;
        RECT 101.490 31.180 101.830 32.010 ;
        RECT 105.425 31.785 108.015 32.555 ;
        RECT 108.645 31.830 108.935 32.555 ;
        RECT 109.105 32.010 114.450 32.555 ;
        RECT 114.625 32.010 119.970 32.555 ;
        RECT 103.310 30.440 103.660 31.690 ;
        RECT 105.425 31.265 106.635 31.785 ;
        RECT 106.805 31.095 108.015 31.615 ;
        RECT 110.690 31.180 111.030 32.010 ;
        RECT 83.345 30.005 88.690 30.440 ;
        RECT 88.865 30.005 94.210 30.440 ;
        RECT 94.385 30.005 99.730 30.440 ;
        RECT 99.905 30.005 105.250 30.440 ;
        RECT 105.425 30.005 108.015 31.095 ;
        RECT 108.645 30.005 108.935 31.170 ;
        RECT 112.510 30.440 112.860 31.690 ;
        RECT 116.210 31.180 116.550 32.010 ;
        RECT 120.145 31.785 123.655 32.555 ;
        RECT 124.285 31.805 125.495 32.555 ;
        RECT 118.030 30.440 118.380 31.690 ;
        RECT 120.145 31.265 121.795 31.785 ;
        RECT 121.965 31.095 123.655 31.615 ;
        RECT 109.105 30.005 114.450 30.440 ;
        RECT 114.625 30.005 119.970 30.440 ;
        RECT 120.145 30.005 123.655 31.095 ;
        RECT 124.285 31.095 124.805 31.635 ;
        RECT 124.975 31.265 125.495 31.805 ;
        RECT 124.285 30.005 125.495 31.095 ;
        RECT 5.520 29.835 125.580 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 6.985 29.400 12.330 29.835 ;
        RECT 12.505 29.400 17.850 29.835 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 8.570 27.830 8.910 28.660 ;
        RECT 10.390 28.150 10.740 29.400 ;
        RECT 14.090 27.830 14.430 28.660 ;
        RECT 15.910 28.150 16.260 29.400 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.945 29.400 24.290 29.835 ;
        RECT 6.985 27.285 12.330 27.830 ;
        RECT 12.505 27.285 17.850 27.830 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 20.530 27.830 20.870 28.660 ;
        RECT 22.350 28.150 22.700 29.400 ;
        RECT 24.465 28.745 27.055 29.835 ;
        RECT 24.465 28.055 25.675 28.575 ;
        RECT 25.845 28.225 27.055 28.745 ;
        RECT 27.745 28.695 27.955 29.835 ;
        RECT 28.125 28.685 28.455 29.665 ;
        RECT 28.625 28.695 28.855 29.835 ;
        RECT 29.065 29.400 34.410 29.835 ;
        RECT 34.585 29.400 39.930 29.835 ;
        RECT 18.945 27.285 24.290 27.830 ;
        RECT 24.465 27.285 27.055 28.055 ;
        RECT 27.745 27.285 27.955 28.105 ;
        RECT 28.125 28.085 28.375 28.685 ;
        RECT 28.545 28.275 28.875 28.525 ;
        RECT 28.125 27.455 28.455 28.085 ;
        RECT 28.625 27.285 28.855 28.105 ;
        RECT 30.650 27.830 30.990 28.660 ;
        RECT 32.470 28.150 32.820 29.400 ;
        RECT 36.170 27.830 36.510 28.660 ;
        RECT 37.990 28.150 38.340 29.400 ;
        RECT 40.105 28.745 43.615 29.835 ;
        RECT 40.105 28.055 41.755 28.575 ;
        RECT 41.925 28.225 43.615 28.745 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.705 28.745 48.215 29.835 ;
        RECT 49.310 29.165 49.565 29.665 ;
        RECT 49.735 29.335 50.065 29.835 ;
        RECT 49.310 28.995 50.060 29.165 ;
        RECT 44.705 28.055 46.355 28.575 ;
        RECT 46.525 28.225 48.215 28.745 ;
        RECT 49.310 28.175 49.660 28.825 ;
        RECT 29.065 27.285 34.410 27.830 ;
        RECT 34.585 27.285 39.930 27.830 ;
        RECT 40.105 27.285 43.615 28.055 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 44.705 27.285 48.215 28.055 ;
        RECT 49.830 28.005 50.060 28.995 ;
        RECT 49.310 27.835 50.060 28.005 ;
        RECT 49.310 27.545 49.565 27.835 ;
        RECT 49.735 27.285 50.065 27.665 ;
        RECT 50.235 27.545 50.405 29.665 ;
        RECT 50.575 28.865 50.900 29.650 ;
        RECT 51.070 29.375 51.320 29.835 ;
        RECT 51.490 29.335 51.740 29.665 ;
        RECT 51.955 29.335 52.635 29.665 ;
        RECT 51.490 29.205 51.660 29.335 ;
        RECT 51.265 29.035 51.660 29.205 ;
        RECT 50.635 27.815 51.095 28.865 ;
        RECT 51.265 27.675 51.435 29.035 ;
        RECT 51.830 28.775 52.295 29.165 ;
        RECT 51.605 27.965 51.955 28.585 ;
        RECT 52.125 28.185 52.295 28.775 ;
        RECT 52.465 28.555 52.635 29.335 ;
        RECT 52.805 29.235 52.975 29.575 ;
        RECT 53.210 29.405 53.540 29.835 ;
        RECT 53.710 29.235 53.880 29.575 ;
        RECT 54.175 29.375 54.545 29.835 ;
        RECT 52.805 29.065 53.880 29.235 ;
        RECT 54.715 29.205 54.885 29.665 ;
        RECT 55.120 29.325 55.990 29.665 ;
        RECT 56.160 29.375 56.410 29.835 ;
        RECT 54.325 29.035 54.885 29.205 ;
        RECT 54.325 28.895 54.495 29.035 ;
        RECT 52.995 28.725 54.495 28.895 ;
        RECT 55.190 28.865 55.650 29.155 ;
        RECT 52.465 28.385 54.155 28.555 ;
        RECT 52.125 27.965 52.480 28.185 ;
        RECT 52.650 27.675 52.820 28.385 ;
        RECT 53.025 27.965 53.815 28.215 ;
        RECT 53.985 28.205 54.155 28.385 ;
        RECT 54.325 28.035 54.495 28.725 ;
        RECT 50.765 27.285 51.095 27.645 ;
        RECT 51.265 27.505 51.760 27.675 ;
        RECT 51.965 27.505 52.820 27.675 ;
        RECT 53.695 27.285 54.025 27.745 ;
        RECT 54.235 27.645 54.495 28.035 ;
        RECT 54.685 28.855 55.650 28.865 ;
        RECT 55.820 28.945 55.990 29.325 ;
        RECT 56.580 29.285 56.750 29.575 ;
        RECT 56.930 29.455 57.260 29.835 ;
        RECT 56.580 29.115 57.380 29.285 ;
        RECT 54.685 28.695 55.360 28.855 ;
        RECT 55.820 28.775 57.040 28.945 ;
        RECT 54.685 27.905 54.895 28.695 ;
        RECT 55.820 28.685 55.990 28.775 ;
        RECT 55.065 27.905 55.415 28.525 ;
        RECT 55.585 28.515 55.990 28.685 ;
        RECT 55.585 27.735 55.755 28.515 ;
        RECT 55.925 28.065 56.145 28.345 ;
        RECT 56.325 28.235 56.865 28.605 ;
        RECT 57.210 28.525 57.380 29.115 ;
        RECT 57.600 28.695 57.905 29.835 ;
        RECT 58.075 28.645 58.330 29.525 ;
        RECT 58.505 28.695 58.765 29.835 ;
        RECT 58.935 28.685 59.265 29.665 ;
        RECT 59.435 28.695 59.715 29.835 ;
        RECT 60.365 29.035 60.645 29.835 ;
        RECT 60.845 28.865 61.175 29.665 ;
        RECT 61.375 29.035 61.545 29.835 ;
        RECT 61.715 28.865 62.045 29.665 ;
        RECT 57.210 28.495 57.950 28.525 ;
        RECT 55.925 27.895 56.455 28.065 ;
        RECT 54.235 27.475 54.585 27.645 ;
        RECT 54.805 27.455 55.755 27.735 ;
        RECT 55.925 27.285 56.115 27.725 ;
        RECT 56.285 27.665 56.455 27.895 ;
        RECT 56.625 27.835 56.865 28.235 ;
        RECT 57.035 28.195 57.950 28.495 ;
        RECT 57.035 28.020 57.360 28.195 ;
        RECT 57.035 27.665 57.355 28.020 ;
        RECT 58.120 27.995 58.330 28.645 ;
        RECT 58.525 28.275 58.860 28.525 ;
        RECT 59.030 28.085 59.200 28.685 ;
        RECT 59.370 28.255 59.705 28.525 ;
        RECT 60.345 28.195 60.585 28.865 ;
        RECT 60.765 28.695 62.045 28.865 ;
        RECT 62.215 28.695 62.475 29.835 ;
        RECT 62.645 28.695 62.920 29.665 ;
        RECT 63.130 29.035 63.410 29.835 ;
        RECT 63.580 29.325 65.195 29.655 ;
        RECT 63.580 28.985 64.755 29.155 ;
        RECT 63.580 28.865 63.750 28.985 ;
        RECT 63.090 28.695 63.750 28.865 ;
        RECT 56.285 27.495 57.355 27.665 ;
        RECT 57.600 27.285 57.905 27.745 ;
        RECT 58.075 27.465 58.330 27.995 ;
        RECT 58.505 27.455 59.200 28.085 ;
        RECT 59.405 27.285 59.715 28.085 ;
        RECT 60.765 28.025 60.935 28.695 ;
        RECT 61.105 28.195 61.415 28.525 ;
        RECT 61.585 28.195 61.965 28.525 ;
        RECT 62.165 28.195 62.450 28.525 ;
        RECT 61.210 28.025 61.415 28.195 ;
        RECT 60.345 27.455 61.040 28.025 ;
        RECT 61.210 27.500 61.560 28.025 ;
        RECT 61.750 27.500 61.965 28.195 ;
        RECT 62.135 27.285 62.470 28.025 ;
        RECT 62.645 27.960 62.815 28.695 ;
        RECT 63.090 28.525 63.260 28.695 ;
        RECT 64.010 28.525 64.255 28.815 ;
        RECT 64.425 28.695 64.755 28.985 ;
        RECT 65.015 28.525 65.185 29.085 ;
        RECT 65.435 28.695 65.695 29.835 ;
        RECT 65.865 29.325 66.165 29.835 ;
        RECT 66.335 29.155 66.665 29.665 ;
        RECT 66.835 29.325 67.465 29.835 ;
        RECT 68.045 29.325 68.425 29.495 ;
        RECT 68.595 29.325 68.895 29.835 ;
        RECT 68.255 29.155 68.425 29.325 ;
        RECT 65.865 28.985 68.085 29.155 ;
        RECT 62.985 28.195 63.260 28.525 ;
        RECT 63.430 28.195 64.255 28.525 ;
        RECT 64.470 28.195 65.185 28.525 ;
        RECT 65.355 28.275 65.690 28.525 ;
        RECT 63.090 28.025 63.260 28.195 ;
        RECT 64.935 28.105 65.185 28.195 ;
        RECT 62.645 27.615 62.920 27.960 ;
        RECT 63.090 27.855 64.755 28.025 ;
        RECT 63.110 27.285 63.485 27.685 ;
        RECT 63.655 27.505 63.825 27.855 ;
        RECT 63.995 27.285 64.325 27.685 ;
        RECT 64.495 27.455 64.755 27.855 ;
        RECT 64.935 27.685 65.265 28.105 ;
        RECT 65.435 27.285 65.695 28.105 ;
        RECT 65.865 28.025 66.035 28.985 ;
        RECT 66.205 28.645 67.745 28.815 ;
        RECT 66.205 28.195 66.450 28.645 ;
        RECT 66.710 28.275 67.405 28.475 ;
        RECT 67.575 28.445 67.745 28.645 ;
        RECT 67.915 28.785 68.085 28.985 ;
        RECT 68.255 28.955 68.915 29.155 ;
        RECT 67.915 28.615 68.575 28.785 ;
        RECT 67.575 28.275 68.175 28.445 ;
        RECT 68.405 28.195 68.575 28.615 ;
        RECT 65.865 27.480 66.330 28.025 ;
        RECT 66.835 27.285 67.005 28.105 ;
        RECT 67.175 28.025 68.085 28.105 ;
        RECT 68.745 28.025 68.915 28.955 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 70.515 28.695 70.765 29.835 ;
        RECT 70.935 28.645 71.185 29.525 ;
        RECT 71.355 28.695 71.660 29.835 ;
        RECT 72.000 29.455 72.330 29.835 ;
        RECT 72.510 29.285 72.680 29.575 ;
        RECT 72.850 29.375 73.100 29.835 ;
        RECT 71.880 29.115 72.680 29.285 ;
        RECT 73.270 29.325 74.140 29.665 ;
        RECT 67.175 27.935 68.425 28.025 ;
        RECT 67.175 27.455 67.505 27.935 ;
        RECT 67.915 27.855 68.425 27.935 ;
        RECT 67.675 27.285 68.025 27.675 ;
        RECT 68.195 27.455 68.425 27.855 ;
        RECT 68.595 27.545 68.915 28.025 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 70.515 27.285 70.765 28.040 ;
        RECT 70.935 27.995 71.140 28.645 ;
        RECT 71.880 28.525 72.050 29.115 ;
        RECT 73.270 28.945 73.440 29.325 ;
        RECT 74.375 29.205 74.545 29.665 ;
        RECT 74.715 29.375 75.085 29.835 ;
        RECT 75.380 29.235 75.550 29.575 ;
        RECT 75.720 29.405 76.050 29.835 ;
        RECT 76.285 29.235 76.455 29.575 ;
        RECT 72.220 28.775 73.440 28.945 ;
        RECT 73.610 28.865 74.070 29.155 ;
        RECT 74.375 29.035 74.935 29.205 ;
        RECT 75.380 29.065 76.455 29.235 ;
        RECT 76.625 29.335 77.305 29.665 ;
        RECT 77.520 29.335 77.770 29.665 ;
        RECT 77.940 29.375 78.190 29.835 ;
        RECT 74.765 28.895 74.935 29.035 ;
        RECT 73.610 28.855 74.575 28.865 ;
        RECT 73.270 28.685 73.440 28.775 ;
        RECT 73.900 28.695 74.575 28.855 ;
        RECT 71.310 28.495 72.050 28.525 ;
        RECT 71.310 28.195 72.225 28.495 ;
        RECT 71.900 28.020 72.225 28.195 ;
        RECT 70.935 27.465 71.185 27.995 ;
        RECT 71.355 27.285 71.660 27.745 ;
        RECT 71.905 27.665 72.225 28.020 ;
        RECT 72.395 28.235 72.935 28.605 ;
        RECT 73.270 28.515 73.675 28.685 ;
        RECT 72.395 27.835 72.635 28.235 ;
        RECT 73.115 28.065 73.335 28.345 ;
        RECT 72.805 27.895 73.335 28.065 ;
        RECT 72.805 27.665 72.975 27.895 ;
        RECT 73.505 27.735 73.675 28.515 ;
        RECT 73.845 27.905 74.195 28.525 ;
        RECT 74.365 27.905 74.575 28.695 ;
        RECT 74.765 28.725 76.265 28.895 ;
        RECT 74.765 28.035 74.935 28.725 ;
        RECT 76.625 28.555 76.795 29.335 ;
        RECT 77.600 29.205 77.770 29.335 ;
        RECT 75.105 28.385 76.795 28.555 ;
        RECT 76.965 28.775 77.430 29.165 ;
        RECT 77.600 29.035 77.995 29.205 ;
        RECT 75.105 28.205 75.275 28.385 ;
        RECT 71.905 27.495 72.975 27.665 ;
        RECT 73.145 27.285 73.335 27.725 ;
        RECT 73.505 27.455 74.455 27.735 ;
        RECT 74.765 27.645 75.025 28.035 ;
        RECT 75.445 27.965 76.235 28.215 ;
        RECT 74.675 27.475 75.025 27.645 ;
        RECT 75.235 27.285 75.565 27.745 ;
        RECT 76.440 27.675 76.610 28.385 ;
        RECT 76.965 28.185 77.135 28.775 ;
        RECT 76.780 27.965 77.135 28.185 ;
        RECT 77.305 27.965 77.655 28.585 ;
        RECT 77.825 27.675 77.995 29.035 ;
        RECT 78.360 28.865 78.685 29.650 ;
        RECT 78.165 27.815 78.625 28.865 ;
        RECT 76.440 27.505 77.295 27.675 ;
        RECT 77.500 27.505 77.995 27.675 ;
        RECT 78.165 27.285 78.495 27.645 ;
        RECT 78.855 27.545 79.025 29.665 ;
        RECT 79.195 29.335 79.525 29.835 ;
        RECT 79.695 29.165 79.950 29.665 ;
        RECT 80.125 29.400 85.470 29.835 ;
        RECT 85.645 29.400 90.990 29.835 ;
        RECT 79.200 28.995 79.950 29.165 ;
        RECT 79.200 28.005 79.430 28.995 ;
        RECT 79.600 28.175 79.950 28.825 ;
        RECT 79.200 27.835 79.950 28.005 ;
        RECT 79.195 27.285 79.525 27.665 ;
        RECT 79.695 27.545 79.950 27.835 ;
        RECT 81.710 27.830 82.050 28.660 ;
        RECT 83.530 28.150 83.880 29.400 ;
        RECT 87.230 27.830 87.570 28.660 ;
        RECT 89.050 28.150 89.400 29.400 ;
        RECT 91.165 28.745 94.675 29.835 ;
        RECT 91.165 28.055 92.815 28.575 ;
        RECT 92.985 28.225 94.675 28.745 ;
        RECT 95.765 28.670 96.055 29.835 ;
        RECT 96.225 29.400 101.570 29.835 ;
        RECT 101.745 29.400 107.090 29.835 ;
        RECT 107.265 29.400 112.610 29.835 ;
        RECT 112.785 29.400 118.130 29.835 ;
        RECT 80.125 27.285 85.470 27.830 ;
        RECT 85.645 27.285 90.990 27.830 ;
        RECT 91.165 27.285 94.675 28.055 ;
        RECT 95.765 27.285 96.055 28.010 ;
        RECT 97.810 27.830 98.150 28.660 ;
        RECT 99.630 28.150 99.980 29.400 ;
        RECT 103.330 27.830 103.670 28.660 ;
        RECT 105.150 28.150 105.500 29.400 ;
        RECT 108.850 27.830 109.190 28.660 ;
        RECT 110.670 28.150 111.020 29.400 ;
        RECT 114.370 27.830 114.710 28.660 ;
        RECT 116.190 28.150 116.540 29.400 ;
        RECT 118.305 28.745 120.895 29.835 ;
        RECT 118.305 28.055 119.515 28.575 ;
        RECT 119.685 28.225 120.895 28.745 ;
        RECT 121.525 28.670 121.815 29.835 ;
        RECT 121.985 28.745 123.655 29.835 ;
        RECT 121.985 28.055 122.735 28.575 ;
        RECT 122.905 28.225 123.655 28.745 ;
        RECT 124.285 28.745 125.495 29.835 ;
        RECT 124.285 28.205 124.805 28.745 ;
        RECT 96.225 27.285 101.570 27.830 ;
        RECT 101.745 27.285 107.090 27.830 ;
        RECT 107.265 27.285 112.610 27.830 ;
        RECT 112.785 27.285 118.130 27.830 ;
        RECT 118.305 27.285 120.895 28.055 ;
        RECT 121.525 27.285 121.815 28.010 ;
        RECT 121.985 27.285 123.655 28.055 ;
        RECT 124.975 28.035 125.495 28.575 ;
        RECT 124.285 27.285 125.495 28.035 ;
        RECT 5.520 27.115 125.580 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 6.985 26.570 12.330 27.115 ;
        RECT 12.505 26.570 17.850 27.115 ;
        RECT 18.025 26.570 23.370 27.115 ;
        RECT 23.545 26.570 28.890 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 8.570 25.740 8.910 26.570 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 10.390 25.000 10.740 26.250 ;
        RECT 14.090 25.740 14.430 26.570 ;
        RECT 15.910 25.000 16.260 26.250 ;
        RECT 19.610 25.740 19.950 26.570 ;
        RECT 21.430 25.000 21.780 26.250 ;
        RECT 25.130 25.740 25.470 26.570 ;
        RECT 29.065 26.345 30.735 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.825 26.570 37.170 27.115 ;
        RECT 37.345 26.570 42.690 27.115 ;
        RECT 42.865 26.570 48.210 27.115 ;
        RECT 26.950 25.000 27.300 26.250 ;
        RECT 29.065 25.825 29.815 26.345 ;
        RECT 29.985 25.655 30.735 26.175 ;
        RECT 33.410 25.740 33.750 26.570 ;
        RECT 6.985 24.565 12.330 25.000 ;
        RECT 12.505 24.565 17.850 25.000 ;
        RECT 18.025 24.565 23.370 25.000 ;
        RECT 23.545 24.565 28.890 25.000 ;
        RECT 29.065 24.565 30.735 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 35.230 25.000 35.580 26.250 ;
        RECT 38.930 25.740 39.270 26.570 ;
        RECT 40.750 25.000 41.100 26.250 ;
        RECT 44.450 25.740 44.790 26.570 ;
        RECT 48.385 26.345 51.895 27.115 ;
        RECT 52.525 26.375 52.845 26.855 ;
        RECT 53.015 26.545 53.245 26.945 ;
        RECT 53.415 26.725 53.765 27.115 ;
        RECT 53.015 26.465 53.525 26.545 ;
        RECT 53.935 26.465 54.265 26.945 ;
        RECT 53.015 26.375 54.265 26.465 ;
        RECT 46.270 25.000 46.620 26.250 ;
        RECT 48.385 25.825 50.035 26.345 ;
        RECT 50.205 25.655 51.895 26.175 ;
        RECT 31.825 24.565 37.170 25.000 ;
        RECT 37.345 24.565 42.690 25.000 ;
        RECT 42.865 24.565 48.210 25.000 ;
        RECT 48.385 24.565 51.895 25.655 ;
        RECT 52.525 25.445 52.695 26.375 ;
        RECT 53.355 26.295 54.265 26.375 ;
        RECT 54.435 26.295 54.605 27.115 ;
        RECT 55.110 26.375 55.575 26.920 ;
        RECT 52.865 25.785 53.035 26.205 ;
        RECT 53.265 25.955 53.865 26.125 ;
        RECT 52.865 25.615 53.525 25.785 ;
        RECT 52.525 25.245 53.185 25.445 ;
        RECT 53.355 25.415 53.525 25.615 ;
        RECT 53.695 25.755 53.865 25.955 ;
        RECT 54.035 25.925 54.730 26.125 ;
        RECT 54.990 25.755 55.235 26.205 ;
        RECT 53.695 25.585 55.235 25.755 ;
        RECT 55.405 25.415 55.575 26.375 ;
        RECT 55.745 26.365 56.955 27.115 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 58.540 26.375 59.155 26.945 ;
        RECT 59.325 26.605 59.540 27.115 ;
        RECT 59.770 26.605 60.050 26.935 ;
        RECT 60.230 26.605 60.470 27.115 ;
        RECT 55.745 25.825 56.265 26.365 ;
        RECT 56.435 25.655 56.955 26.195 ;
        RECT 53.355 25.245 55.575 25.415 ;
        RECT 53.015 25.075 53.185 25.245 ;
        RECT 52.545 24.565 52.845 25.075 ;
        RECT 53.015 24.905 53.395 25.075 ;
        RECT 53.975 24.565 54.605 25.075 ;
        RECT 54.775 24.735 55.105 25.245 ;
        RECT 55.275 24.565 55.575 25.075 ;
        RECT 55.745 24.565 56.955 25.655 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 58.540 25.355 58.855 26.375 ;
        RECT 59.025 25.705 59.195 26.205 ;
        RECT 59.445 25.875 59.710 26.435 ;
        RECT 59.880 25.705 60.050 26.605 ;
        RECT 61.265 26.440 61.540 26.785 ;
        RECT 61.730 26.715 62.105 27.115 ;
        RECT 62.275 26.545 62.445 26.895 ;
        RECT 62.615 26.715 62.945 27.115 ;
        RECT 63.115 26.545 63.375 26.945 ;
        RECT 60.220 25.875 60.575 26.435 ;
        RECT 61.265 25.705 61.435 26.440 ;
        RECT 61.710 26.375 63.375 26.545 ;
        RECT 61.710 26.205 61.880 26.375 ;
        RECT 63.555 26.295 63.885 26.715 ;
        RECT 64.055 26.295 64.315 27.115 ;
        RECT 64.490 26.565 64.745 26.855 ;
        RECT 64.915 26.735 65.245 27.115 ;
        RECT 64.490 26.395 65.240 26.565 ;
        RECT 63.555 26.205 63.805 26.295 ;
        RECT 61.605 25.875 61.880 26.205 ;
        RECT 62.050 25.875 62.875 26.205 ;
        RECT 63.090 25.875 63.805 26.205 ;
        RECT 63.975 25.875 64.310 26.125 ;
        RECT 61.710 25.705 61.880 25.875 ;
        RECT 59.025 25.535 60.450 25.705 ;
        RECT 58.540 24.735 59.075 25.355 ;
        RECT 59.245 24.565 59.575 25.365 ;
        RECT 60.060 25.360 60.450 25.535 ;
        RECT 61.265 24.735 61.540 25.705 ;
        RECT 61.710 25.535 62.370 25.705 ;
        RECT 62.630 25.585 62.875 25.875 ;
        RECT 62.200 25.415 62.370 25.535 ;
        RECT 63.045 25.415 63.375 25.705 ;
        RECT 61.750 24.565 62.030 25.365 ;
        RECT 62.200 25.245 63.375 25.415 ;
        RECT 63.635 25.315 63.805 25.875 ;
        RECT 62.200 24.745 63.815 25.075 ;
        RECT 64.055 24.565 64.315 25.705 ;
        RECT 64.490 25.575 64.840 26.225 ;
        RECT 65.010 25.405 65.240 26.395 ;
        RECT 64.490 25.235 65.240 25.405 ;
        RECT 64.490 24.735 64.745 25.235 ;
        RECT 64.915 24.565 65.245 25.065 ;
        RECT 65.415 24.735 65.585 26.855 ;
        RECT 65.945 26.755 66.275 27.115 ;
        RECT 66.445 26.725 66.940 26.895 ;
        RECT 67.145 26.725 68.000 26.895 ;
        RECT 65.815 25.535 66.275 26.585 ;
        RECT 65.755 24.750 66.080 25.535 ;
        RECT 66.445 25.365 66.615 26.725 ;
        RECT 66.785 25.815 67.135 26.435 ;
        RECT 67.305 26.215 67.660 26.435 ;
        RECT 67.305 25.625 67.475 26.215 ;
        RECT 67.830 26.015 68.000 26.725 ;
        RECT 68.875 26.655 69.205 27.115 ;
        RECT 69.415 26.755 69.765 26.925 ;
        RECT 68.205 26.185 68.995 26.435 ;
        RECT 69.415 26.365 69.675 26.755 ;
        RECT 69.985 26.665 70.935 26.945 ;
        RECT 71.105 26.675 71.295 27.115 ;
        RECT 71.465 26.735 72.535 26.905 ;
        RECT 69.165 26.015 69.335 26.195 ;
        RECT 66.445 25.195 66.840 25.365 ;
        RECT 67.010 25.235 67.475 25.625 ;
        RECT 67.645 25.845 69.335 26.015 ;
        RECT 66.670 25.065 66.840 25.195 ;
        RECT 67.645 25.065 67.815 25.845 ;
        RECT 69.505 25.675 69.675 26.365 ;
        RECT 68.175 25.505 69.675 25.675 ;
        RECT 69.865 25.705 70.075 26.495 ;
        RECT 70.245 25.875 70.595 26.495 ;
        RECT 70.765 25.885 70.935 26.665 ;
        RECT 71.465 26.505 71.635 26.735 ;
        RECT 71.105 26.335 71.635 26.505 ;
        RECT 71.105 26.055 71.325 26.335 ;
        RECT 71.805 26.165 72.045 26.565 ;
        RECT 70.765 25.715 71.170 25.885 ;
        RECT 71.505 25.795 72.045 26.165 ;
        RECT 72.215 26.380 72.535 26.735 ;
        RECT 72.215 26.125 72.540 26.380 ;
        RECT 72.735 26.305 72.905 27.115 ;
        RECT 73.075 26.465 73.405 26.945 ;
        RECT 73.575 26.645 73.745 27.115 ;
        RECT 73.915 26.465 74.245 26.945 ;
        RECT 74.415 26.645 74.585 27.115 ;
        RECT 75.065 26.570 80.410 27.115 ;
        RECT 73.075 26.295 74.840 26.465 ;
        RECT 72.215 25.915 74.245 26.125 ;
        RECT 72.215 25.905 72.560 25.915 ;
        RECT 69.865 25.545 70.540 25.705 ;
        RECT 71.000 25.625 71.170 25.715 ;
        RECT 69.865 25.535 70.830 25.545 ;
        RECT 69.505 25.365 69.675 25.505 ;
        RECT 66.250 24.565 66.500 25.025 ;
        RECT 66.670 24.735 66.920 25.065 ;
        RECT 67.135 24.735 67.815 25.065 ;
        RECT 67.985 25.165 69.060 25.335 ;
        RECT 69.505 25.195 70.065 25.365 ;
        RECT 70.370 25.245 70.830 25.535 ;
        RECT 71.000 25.455 72.220 25.625 ;
        RECT 67.985 24.825 68.155 25.165 ;
        RECT 68.390 24.565 68.720 24.995 ;
        RECT 68.890 24.825 69.060 25.165 ;
        RECT 69.355 24.565 69.725 25.025 ;
        RECT 69.895 24.735 70.065 25.195 ;
        RECT 71.000 25.075 71.170 25.455 ;
        RECT 72.390 25.285 72.560 25.905 ;
        RECT 74.430 25.745 74.840 26.295 ;
        RECT 70.300 24.735 71.170 25.075 ;
        RECT 71.760 25.115 72.560 25.285 ;
        RECT 71.340 24.565 71.590 25.025 ;
        RECT 71.760 24.825 71.930 25.115 ;
        RECT 72.110 24.565 72.440 24.945 ;
        RECT 72.735 24.565 72.905 25.625 ;
        RECT 73.115 25.575 74.840 25.745 ;
        RECT 76.650 25.740 76.990 26.570 ;
        RECT 80.585 26.345 82.255 27.115 ;
        RECT 82.885 26.390 83.175 27.115 ;
        RECT 83.345 26.570 88.690 27.115 ;
        RECT 88.865 26.570 94.210 27.115 ;
        RECT 94.385 26.570 99.730 27.115 ;
        RECT 99.905 26.570 105.250 27.115 ;
        RECT 73.115 24.735 73.405 25.575 ;
        RECT 73.575 24.565 73.745 25.405 ;
        RECT 73.955 24.735 74.205 25.575 ;
        RECT 74.415 24.565 74.585 25.405 ;
        RECT 78.470 25.000 78.820 26.250 ;
        RECT 80.585 25.825 81.335 26.345 ;
        RECT 81.505 25.655 82.255 26.175 ;
        RECT 84.930 25.740 85.270 26.570 ;
        RECT 75.065 24.565 80.410 25.000 ;
        RECT 80.585 24.565 82.255 25.655 ;
        RECT 82.885 24.565 83.175 25.730 ;
        RECT 86.750 25.000 87.100 26.250 ;
        RECT 90.450 25.740 90.790 26.570 ;
        RECT 92.270 25.000 92.620 26.250 ;
        RECT 95.970 25.740 96.310 26.570 ;
        RECT 97.790 25.000 98.140 26.250 ;
        RECT 101.490 25.740 101.830 26.570 ;
        RECT 105.425 26.345 108.015 27.115 ;
        RECT 108.645 26.390 108.935 27.115 ;
        RECT 109.105 26.570 114.450 27.115 ;
        RECT 114.625 26.570 119.970 27.115 ;
        RECT 103.310 25.000 103.660 26.250 ;
        RECT 105.425 25.825 106.635 26.345 ;
        RECT 106.805 25.655 108.015 26.175 ;
        RECT 110.690 25.740 111.030 26.570 ;
        RECT 83.345 24.565 88.690 25.000 ;
        RECT 88.865 24.565 94.210 25.000 ;
        RECT 94.385 24.565 99.730 25.000 ;
        RECT 99.905 24.565 105.250 25.000 ;
        RECT 105.425 24.565 108.015 25.655 ;
        RECT 108.645 24.565 108.935 25.730 ;
        RECT 112.510 25.000 112.860 26.250 ;
        RECT 116.210 25.740 116.550 26.570 ;
        RECT 120.145 26.345 123.655 27.115 ;
        RECT 124.285 26.365 125.495 27.115 ;
        RECT 118.030 25.000 118.380 26.250 ;
        RECT 120.145 25.825 121.795 26.345 ;
        RECT 121.965 25.655 123.655 26.175 ;
        RECT 109.105 24.565 114.450 25.000 ;
        RECT 114.625 24.565 119.970 25.000 ;
        RECT 120.145 24.565 123.655 25.655 ;
        RECT 124.285 25.655 124.805 26.195 ;
        RECT 124.975 25.825 125.495 26.365 ;
        RECT 124.285 24.565 125.495 25.655 ;
        RECT 5.520 24.395 125.580 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 6.985 23.960 12.330 24.395 ;
        RECT 12.505 23.960 17.850 24.395 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 8.570 22.390 8.910 23.220 ;
        RECT 10.390 22.710 10.740 23.960 ;
        RECT 14.090 22.390 14.430 23.220 ;
        RECT 15.910 22.710 16.260 23.960 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.960 24.290 24.395 ;
        RECT 24.465 23.960 29.810 24.395 ;
        RECT 29.985 23.960 35.330 24.395 ;
        RECT 35.505 23.960 40.850 24.395 ;
        RECT 6.985 21.845 12.330 22.390 ;
        RECT 12.505 21.845 17.850 22.390 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 20.530 22.390 20.870 23.220 ;
        RECT 22.350 22.710 22.700 23.960 ;
        RECT 26.050 22.390 26.390 23.220 ;
        RECT 27.870 22.710 28.220 23.960 ;
        RECT 31.570 22.390 31.910 23.220 ;
        RECT 33.390 22.710 33.740 23.960 ;
        RECT 37.090 22.390 37.430 23.220 ;
        RECT 38.910 22.710 39.260 23.960 ;
        RECT 41.025 23.305 43.615 24.395 ;
        RECT 41.025 22.615 42.235 23.135 ;
        RECT 42.405 22.785 43.615 23.305 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.705 23.960 50.050 24.395 ;
        RECT 50.225 23.960 55.570 24.395 ;
        RECT 55.745 23.960 61.090 24.395 ;
        RECT 61.265 23.960 66.610 24.395 ;
        RECT 18.945 21.845 24.290 22.390 ;
        RECT 24.465 21.845 29.810 22.390 ;
        RECT 29.985 21.845 35.330 22.390 ;
        RECT 35.505 21.845 40.850 22.390 ;
        RECT 41.025 21.845 43.615 22.615 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 46.290 22.390 46.630 23.220 ;
        RECT 48.110 22.710 48.460 23.960 ;
        RECT 51.810 22.390 52.150 23.220 ;
        RECT 53.630 22.710 53.980 23.960 ;
        RECT 57.330 22.390 57.670 23.220 ;
        RECT 59.150 22.710 59.500 23.960 ;
        RECT 62.850 22.390 63.190 23.220 ;
        RECT 64.670 22.710 65.020 23.960 ;
        RECT 67.245 23.320 67.515 24.225 ;
        RECT 67.685 23.635 68.015 24.395 ;
        RECT 68.195 23.465 68.365 24.225 ;
        RECT 67.245 22.520 67.415 23.320 ;
        RECT 67.700 23.295 68.365 23.465 ;
        RECT 68.625 23.305 69.835 24.395 ;
        RECT 67.700 23.150 67.870 23.295 ;
        RECT 67.585 22.820 67.870 23.150 ;
        RECT 67.700 22.565 67.870 22.820 ;
        RECT 68.105 22.745 68.435 23.115 ;
        RECT 68.625 22.595 69.145 23.135 ;
        RECT 69.315 22.765 69.835 23.305 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.525 23.255 70.735 24.395 ;
        RECT 70.905 23.245 71.235 24.225 ;
        RECT 71.405 23.255 71.635 24.395 ;
        RECT 71.845 23.960 77.190 24.395 ;
        RECT 77.365 23.960 82.710 24.395 ;
        RECT 82.885 23.960 88.230 24.395 ;
        RECT 88.405 23.960 93.750 24.395 ;
        RECT 44.705 21.845 50.050 22.390 ;
        RECT 50.225 21.845 55.570 22.390 ;
        RECT 55.745 21.845 61.090 22.390 ;
        RECT 61.265 21.845 66.610 22.390 ;
        RECT 67.245 22.015 67.505 22.520 ;
        RECT 67.700 22.395 68.365 22.565 ;
        RECT 67.685 21.845 68.015 22.225 ;
        RECT 68.195 22.015 68.365 22.395 ;
        RECT 68.625 21.845 69.835 22.595 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 70.525 21.845 70.735 22.665 ;
        RECT 70.905 22.645 71.155 23.245 ;
        RECT 71.325 22.835 71.655 23.085 ;
        RECT 70.905 22.015 71.235 22.645 ;
        RECT 71.405 21.845 71.635 22.665 ;
        RECT 73.430 22.390 73.770 23.220 ;
        RECT 75.250 22.710 75.600 23.960 ;
        RECT 78.950 22.390 79.290 23.220 ;
        RECT 80.770 22.710 81.120 23.960 ;
        RECT 84.470 22.390 84.810 23.220 ;
        RECT 86.290 22.710 86.640 23.960 ;
        RECT 89.990 22.390 90.330 23.220 ;
        RECT 91.810 22.710 92.160 23.960 ;
        RECT 93.925 23.305 95.595 24.395 ;
        RECT 93.925 22.615 94.675 23.135 ;
        RECT 94.845 22.785 95.595 23.305 ;
        RECT 95.765 23.230 96.055 24.395 ;
        RECT 96.225 23.960 101.570 24.395 ;
        RECT 101.745 23.960 107.090 24.395 ;
        RECT 107.265 23.960 112.610 24.395 ;
        RECT 112.785 23.960 118.130 24.395 ;
        RECT 71.845 21.845 77.190 22.390 ;
        RECT 77.365 21.845 82.710 22.390 ;
        RECT 82.885 21.845 88.230 22.390 ;
        RECT 88.405 21.845 93.750 22.390 ;
        RECT 93.925 21.845 95.595 22.615 ;
        RECT 95.765 21.845 96.055 22.570 ;
        RECT 97.810 22.390 98.150 23.220 ;
        RECT 99.630 22.710 99.980 23.960 ;
        RECT 103.330 22.390 103.670 23.220 ;
        RECT 105.150 22.710 105.500 23.960 ;
        RECT 108.850 22.390 109.190 23.220 ;
        RECT 110.670 22.710 111.020 23.960 ;
        RECT 114.370 22.390 114.710 23.220 ;
        RECT 116.190 22.710 116.540 23.960 ;
        RECT 118.305 23.305 120.895 24.395 ;
        RECT 118.305 22.615 119.515 23.135 ;
        RECT 119.685 22.785 120.895 23.305 ;
        RECT 121.525 23.230 121.815 24.395 ;
        RECT 121.985 23.305 123.655 24.395 ;
        RECT 121.985 22.615 122.735 23.135 ;
        RECT 122.905 22.785 123.655 23.305 ;
        RECT 124.285 23.305 125.495 24.395 ;
        RECT 124.285 22.765 124.805 23.305 ;
        RECT 96.225 21.845 101.570 22.390 ;
        RECT 101.745 21.845 107.090 22.390 ;
        RECT 107.265 21.845 112.610 22.390 ;
        RECT 112.785 21.845 118.130 22.390 ;
        RECT 118.305 21.845 120.895 22.615 ;
        RECT 121.525 21.845 121.815 22.570 ;
        RECT 121.985 21.845 123.655 22.615 ;
        RECT 124.975 22.595 125.495 23.135 ;
        RECT 124.285 21.845 125.495 22.595 ;
        RECT 5.520 21.675 125.580 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 6.985 21.130 12.330 21.675 ;
        RECT 12.505 21.130 17.850 21.675 ;
        RECT 18.025 21.130 23.370 21.675 ;
        RECT 23.545 21.130 28.890 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 8.570 20.300 8.910 21.130 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 10.390 19.560 10.740 20.810 ;
        RECT 14.090 20.300 14.430 21.130 ;
        RECT 15.910 19.560 16.260 20.810 ;
        RECT 19.610 20.300 19.950 21.130 ;
        RECT 21.430 19.560 21.780 20.810 ;
        RECT 25.130 20.300 25.470 21.130 ;
        RECT 29.065 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 37.345 21.130 42.690 21.675 ;
        RECT 42.865 21.130 48.210 21.675 ;
        RECT 48.385 21.130 53.730 21.675 ;
        RECT 26.950 19.560 27.300 20.810 ;
        RECT 29.065 20.385 29.815 20.905 ;
        RECT 29.985 20.215 30.735 20.735 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 6.985 19.125 12.330 19.560 ;
        RECT 12.505 19.125 17.850 19.560 ;
        RECT 18.025 19.125 23.370 19.560 ;
        RECT 23.545 19.125 28.890 19.560 ;
        RECT 29.065 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 38.930 20.300 39.270 21.130 ;
        RECT 40.750 19.560 41.100 20.810 ;
        RECT 44.450 20.300 44.790 21.130 ;
        RECT 46.270 19.560 46.620 20.810 ;
        RECT 49.970 20.300 50.310 21.130 ;
        RECT 53.905 20.905 56.495 21.675 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 57.585 21.130 62.930 21.675 ;
        RECT 63.105 21.130 68.450 21.675 ;
        RECT 68.625 21.130 73.970 21.675 ;
        RECT 74.145 21.130 79.490 21.675 ;
        RECT 51.790 19.560 52.140 20.810 ;
        RECT 53.905 20.385 55.115 20.905 ;
        RECT 55.285 20.215 56.495 20.735 ;
        RECT 59.170 20.300 59.510 21.130 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.345 19.125 42.690 19.560 ;
        RECT 42.865 19.125 48.210 19.560 ;
        RECT 48.385 19.125 53.730 19.560 ;
        RECT 53.905 19.125 56.495 20.215 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 60.990 19.560 61.340 20.810 ;
        RECT 64.690 20.300 65.030 21.130 ;
        RECT 66.510 19.560 66.860 20.810 ;
        RECT 70.210 20.300 70.550 21.130 ;
        RECT 72.030 19.560 72.380 20.810 ;
        RECT 75.730 20.300 76.070 21.130 ;
        RECT 79.665 20.905 82.255 21.675 ;
        RECT 82.885 20.950 83.175 21.675 ;
        RECT 83.345 21.130 88.690 21.675 ;
        RECT 88.865 21.130 94.210 21.675 ;
        RECT 94.385 21.130 99.730 21.675 ;
        RECT 99.905 21.130 105.250 21.675 ;
        RECT 77.550 19.560 77.900 20.810 ;
        RECT 79.665 20.385 80.875 20.905 ;
        RECT 81.045 20.215 82.255 20.735 ;
        RECT 84.930 20.300 85.270 21.130 ;
        RECT 57.585 19.125 62.930 19.560 ;
        RECT 63.105 19.125 68.450 19.560 ;
        RECT 68.625 19.125 73.970 19.560 ;
        RECT 74.145 19.125 79.490 19.560 ;
        RECT 79.665 19.125 82.255 20.215 ;
        RECT 82.885 19.125 83.175 20.290 ;
        RECT 86.750 19.560 87.100 20.810 ;
        RECT 90.450 20.300 90.790 21.130 ;
        RECT 92.270 19.560 92.620 20.810 ;
        RECT 95.970 20.300 96.310 21.130 ;
        RECT 97.790 19.560 98.140 20.810 ;
        RECT 101.490 20.300 101.830 21.130 ;
        RECT 105.425 20.905 108.015 21.675 ;
        RECT 108.645 20.950 108.935 21.675 ;
        RECT 109.105 21.130 114.450 21.675 ;
        RECT 114.625 21.130 119.970 21.675 ;
        RECT 103.310 19.560 103.660 20.810 ;
        RECT 105.425 20.385 106.635 20.905 ;
        RECT 106.805 20.215 108.015 20.735 ;
        RECT 110.690 20.300 111.030 21.130 ;
        RECT 83.345 19.125 88.690 19.560 ;
        RECT 88.865 19.125 94.210 19.560 ;
        RECT 94.385 19.125 99.730 19.560 ;
        RECT 99.905 19.125 105.250 19.560 ;
        RECT 105.425 19.125 108.015 20.215 ;
        RECT 108.645 19.125 108.935 20.290 ;
        RECT 112.510 19.560 112.860 20.810 ;
        RECT 116.210 20.300 116.550 21.130 ;
        RECT 120.145 20.905 123.655 21.675 ;
        RECT 124.285 20.925 125.495 21.675 ;
        RECT 118.030 19.560 118.380 20.810 ;
        RECT 120.145 20.385 121.795 20.905 ;
        RECT 121.965 20.215 123.655 20.735 ;
        RECT 109.105 19.125 114.450 19.560 ;
        RECT 114.625 19.125 119.970 19.560 ;
        RECT 120.145 19.125 123.655 20.215 ;
        RECT 124.285 20.215 124.805 20.755 ;
        RECT 124.975 20.385 125.495 20.925 ;
        RECT 124.285 19.125 125.495 20.215 ;
        RECT 5.520 18.955 125.580 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 6.985 18.520 12.330 18.955 ;
        RECT 12.505 18.520 17.850 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 8.570 16.950 8.910 17.780 ;
        RECT 10.390 17.270 10.740 18.520 ;
        RECT 14.090 16.950 14.430 17.780 ;
        RECT 15.910 17.270 16.260 18.520 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 18.520 24.290 18.955 ;
        RECT 24.465 18.520 29.810 18.955 ;
        RECT 29.985 18.520 35.330 18.955 ;
        RECT 35.505 18.520 40.850 18.955 ;
        RECT 6.985 16.405 12.330 16.950 ;
        RECT 12.505 16.405 17.850 16.950 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 20.530 16.950 20.870 17.780 ;
        RECT 22.350 17.270 22.700 18.520 ;
        RECT 26.050 16.950 26.390 17.780 ;
        RECT 27.870 17.270 28.220 18.520 ;
        RECT 31.570 16.950 31.910 17.780 ;
        RECT 33.390 17.270 33.740 18.520 ;
        RECT 37.090 16.950 37.430 17.780 ;
        RECT 38.910 17.270 39.260 18.520 ;
        RECT 41.025 17.865 43.615 18.955 ;
        RECT 41.025 17.175 42.235 17.695 ;
        RECT 42.405 17.345 43.615 17.865 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 44.705 18.520 50.050 18.955 ;
        RECT 50.225 18.520 55.570 18.955 ;
        RECT 55.745 18.520 61.090 18.955 ;
        RECT 61.265 18.520 66.610 18.955 ;
        RECT 18.945 16.405 24.290 16.950 ;
        RECT 24.465 16.405 29.810 16.950 ;
        RECT 29.985 16.405 35.330 16.950 ;
        RECT 35.505 16.405 40.850 16.950 ;
        RECT 41.025 16.405 43.615 17.175 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 46.290 16.950 46.630 17.780 ;
        RECT 48.110 17.270 48.460 18.520 ;
        RECT 51.810 16.950 52.150 17.780 ;
        RECT 53.630 17.270 53.980 18.520 ;
        RECT 57.330 16.950 57.670 17.780 ;
        RECT 59.150 17.270 59.500 18.520 ;
        RECT 62.850 16.950 63.190 17.780 ;
        RECT 64.670 17.270 65.020 18.520 ;
        RECT 66.785 17.865 69.375 18.955 ;
        RECT 66.785 17.175 67.995 17.695 ;
        RECT 68.165 17.345 69.375 17.865 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 70.465 18.520 75.810 18.955 ;
        RECT 75.985 18.520 81.330 18.955 ;
        RECT 81.505 18.520 86.850 18.955 ;
        RECT 87.025 18.520 92.370 18.955 ;
        RECT 44.705 16.405 50.050 16.950 ;
        RECT 50.225 16.405 55.570 16.950 ;
        RECT 55.745 16.405 61.090 16.950 ;
        RECT 61.265 16.405 66.610 16.950 ;
        RECT 66.785 16.405 69.375 17.175 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 72.050 16.950 72.390 17.780 ;
        RECT 73.870 17.270 74.220 18.520 ;
        RECT 77.570 16.950 77.910 17.780 ;
        RECT 79.390 17.270 79.740 18.520 ;
        RECT 83.090 16.950 83.430 17.780 ;
        RECT 84.910 17.270 85.260 18.520 ;
        RECT 88.610 16.950 88.950 17.780 ;
        RECT 90.430 17.270 90.780 18.520 ;
        RECT 92.545 17.865 95.135 18.955 ;
        RECT 92.545 17.175 93.755 17.695 ;
        RECT 93.925 17.345 95.135 17.865 ;
        RECT 95.765 17.790 96.055 18.955 ;
        RECT 96.225 18.520 101.570 18.955 ;
        RECT 101.745 18.520 107.090 18.955 ;
        RECT 107.265 18.520 112.610 18.955 ;
        RECT 112.785 18.520 118.130 18.955 ;
        RECT 70.465 16.405 75.810 16.950 ;
        RECT 75.985 16.405 81.330 16.950 ;
        RECT 81.505 16.405 86.850 16.950 ;
        RECT 87.025 16.405 92.370 16.950 ;
        RECT 92.545 16.405 95.135 17.175 ;
        RECT 95.765 16.405 96.055 17.130 ;
        RECT 97.810 16.950 98.150 17.780 ;
        RECT 99.630 17.270 99.980 18.520 ;
        RECT 103.330 16.950 103.670 17.780 ;
        RECT 105.150 17.270 105.500 18.520 ;
        RECT 108.850 16.950 109.190 17.780 ;
        RECT 110.670 17.270 111.020 18.520 ;
        RECT 114.370 16.950 114.710 17.780 ;
        RECT 116.190 17.270 116.540 18.520 ;
        RECT 118.305 17.865 120.895 18.955 ;
        RECT 118.305 17.175 119.515 17.695 ;
        RECT 119.685 17.345 120.895 17.865 ;
        RECT 121.525 17.790 121.815 18.955 ;
        RECT 121.985 17.865 123.655 18.955 ;
        RECT 121.985 17.175 122.735 17.695 ;
        RECT 122.905 17.345 123.655 17.865 ;
        RECT 124.285 17.865 125.495 18.955 ;
        RECT 124.285 17.325 124.805 17.865 ;
        RECT 96.225 16.405 101.570 16.950 ;
        RECT 101.745 16.405 107.090 16.950 ;
        RECT 107.265 16.405 112.610 16.950 ;
        RECT 112.785 16.405 118.130 16.950 ;
        RECT 118.305 16.405 120.895 17.175 ;
        RECT 121.525 16.405 121.815 17.130 ;
        RECT 121.985 16.405 123.655 17.175 ;
        RECT 124.975 17.155 125.495 17.695 ;
        RECT 124.285 16.405 125.495 17.155 ;
        RECT 5.520 16.235 125.580 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 18.025 15.690 23.370 16.235 ;
        RECT 23.545 15.690 28.890 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 19.610 14.860 19.950 15.690 ;
        RECT 21.430 14.120 21.780 15.370 ;
        RECT 25.130 14.860 25.470 15.690 ;
        RECT 29.065 15.465 30.735 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.690 37.170 16.235 ;
        RECT 37.345 15.690 42.690 16.235 ;
        RECT 42.865 15.690 48.210 16.235 ;
        RECT 48.385 15.690 53.730 16.235 ;
        RECT 26.950 14.120 27.300 15.370 ;
        RECT 29.065 14.945 29.815 15.465 ;
        RECT 29.985 14.775 30.735 15.295 ;
        RECT 33.410 14.860 33.750 15.690 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 23.370 14.120 ;
        RECT 23.545 13.685 28.890 14.120 ;
        RECT 29.065 13.685 30.735 14.775 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 35.230 14.120 35.580 15.370 ;
        RECT 38.930 14.860 39.270 15.690 ;
        RECT 40.750 14.120 41.100 15.370 ;
        RECT 44.450 14.860 44.790 15.690 ;
        RECT 46.270 14.120 46.620 15.370 ;
        RECT 49.970 14.860 50.310 15.690 ;
        RECT 53.905 15.465 56.495 16.235 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 57.585 15.690 62.930 16.235 ;
        RECT 63.105 15.690 68.450 16.235 ;
        RECT 68.625 15.690 73.970 16.235 ;
        RECT 74.145 15.690 79.490 16.235 ;
        RECT 51.790 14.120 52.140 15.370 ;
        RECT 53.905 14.945 55.115 15.465 ;
        RECT 55.285 14.775 56.495 15.295 ;
        RECT 59.170 14.860 59.510 15.690 ;
        RECT 31.825 13.685 37.170 14.120 ;
        RECT 37.345 13.685 42.690 14.120 ;
        RECT 42.865 13.685 48.210 14.120 ;
        RECT 48.385 13.685 53.730 14.120 ;
        RECT 53.905 13.685 56.495 14.775 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 60.990 14.120 61.340 15.370 ;
        RECT 64.690 14.860 65.030 15.690 ;
        RECT 66.510 14.120 66.860 15.370 ;
        RECT 70.210 14.860 70.550 15.690 ;
        RECT 72.030 14.120 72.380 15.370 ;
        RECT 75.730 14.860 76.070 15.690 ;
        RECT 79.665 15.465 82.255 16.235 ;
        RECT 82.885 15.510 83.175 16.235 ;
        RECT 83.345 15.690 88.690 16.235 ;
        RECT 88.865 15.690 94.210 16.235 ;
        RECT 94.385 15.690 99.730 16.235 ;
        RECT 99.905 15.690 105.250 16.235 ;
        RECT 77.550 14.120 77.900 15.370 ;
        RECT 79.665 14.945 80.875 15.465 ;
        RECT 81.045 14.775 82.255 15.295 ;
        RECT 84.930 14.860 85.270 15.690 ;
        RECT 57.585 13.685 62.930 14.120 ;
        RECT 63.105 13.685 68.450 14.120 ;
        RECT 68.625 13.685 73.970 14.120 ;
        RECT 74.145 13.685 79.490 14.120 ;
        RECT 79.665 13.685 82.255 14.775 ;
        RECT 82.885 13.685 83.175 14.850 ;
        RECT 86.750 14.120 87.100 15.370 ;
        RECT 90.450 14.860 90.790 15.690 ;
        RECT 92.270 14.120 92.620 15.370 ;
        RECT 95.970 14.860 96.310 15.690 ;
        RECT 97.790 14.120 98.140 15.370 ;
        RECT 101.490 14.860 101.830 15.690 ;
        RECT 105.425 15.465 108.015 16.235 ;
        RECT 108.645 15.510 108.935 16.235 ;
        RECT 109.105 15.690 114.450 16.235 ;
        RECT 114.625 15.690 119.970 16.235 ;
        RECT 103.310 14.120 103.660 15.370 ;
        RECT 105.425 14.945 106.635 15.465 ;
        RECT 106.805 14.775 108.015 15.295 ;
        RECT 110.690 14.860 111.030 15.690 ;
        RECT 83.345 13.685 88.690 14.120 ;
        RECT 88.865 13.685 94.210 14.120 ;
        RECT 94.385 13.685 99.730 14.120 ;
        RECT 99.905 13.685 105.250 14.120 ;
        RECT 105.425 13.685 108.015 14.775 ;
        RECT 108.645 13.685 108.935 14.850 ;
        RECT 112.510 14.120 112.860 15.370 ;
        RECT 116.210 14.860 116.550 15.690 ;
        RECT 120.145 15.465 123.655 16.235 ;
        RECT 124.285 15.485 125.495 16.235 ;
        RECT 118.030 14.120 118.380 15.370 ;
        RECT 120.145 14.945 121.795 15.465 ;
        RECT 121.965 14.775 123.655 15.295 ;
        RECT 109.105 13.685 114.450 14.120 ;
        RECT 114.625 13.685 119.970 14.120 ;
        RECT 120.145 13.685 123.655 14.775 ;
        RECT 124.285 14.775 124.805 15.315 ;
        RECT 124.975 14.945 125.495 15.485 ;
        RECT 124.285 13.685 125.495 14.775 ;
        RECT 5.520 13.515 125.580 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 12.505 13.080 17.850 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 14.090 11.510 14.430 12.340 ;
        RECT 15.910 11.830 16.260 13.080 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 13.080 24.290 13.515 ;
        RECT 24.465 13.080 29.810 13.515 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 12.505 10.965 17.850 11.510 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 20.530 11.510 20.870 12.340 ;
        RECT 22.350 11.830 22.700 13.080 ;
        RECT 26.050 11.510 26.390 12.340 ;
        RECT 27.870 11.830 28.220 13.080 ;
        RECT 29.985 12.425 31.195 13.515 ;
        RECT 29.985 11.715 30.505 12.255 ;
        RECT 30.675 11.885 31.195 12.425 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 31.825 13.080 37.170 13.515 ;
        RECT 37.345 13.080 42.690 13.515 ;
        RECT 18.945 10.965 24.290 11.510 ;
        RECT 24.465 10.965 29.810 11.510 ;
        RECT 29.985 10.965 31.195 11.715 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 33.410 11.510 33.750 12.340 ;
        RECT 35.230 11.830 35.580 13.080 ;
        RECT 38.930 11.510 39.270 12.340 ;
        RECT 40.750 11.830 41.100 13.080 ;
        RECT 42.865 12.425 44.075 13.515 ;
        RECT 42.865 11.715 43.385 12.255 ;
        RECT 43.555 11.885 44.075 12.425 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 44.705 13.080 50.050 13.515 ;
        RECT 50.225 13.080 55.570 13.515 ;
        RECT 31.825 10.965 37.170 11.510 ;
        RECT 37.345 10.965 42.690 11.510 ;
        RECT 42.865 10.965 44.075 11.715 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 46.290 11.510 46.630 12.340 ;
        RECT 48.110 11.830 48.460 13.080 ;
        RECT 51.810 11.510 52.150 12.340 ;
        RECT 53.630 11.830 53.980 13.080 ;
        RECT 55.745 12.425 56.955 13.515 ;
        RECT 55.745 11.715 56.265 12.255 ;
        RECT 56.435 11.885 56.955 12.425 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 57.585 13.080 62.930 13.515 ;
        RECT 63.105 13.080 68.450 13.515 ;
        RECT 44.705 10.965 50.050 11.510 ;
        RECT 50.225 10.965 55.570 11.510 ;
        RECT 55.745 10.965 56.955 11.715 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 59.170 11.510 59.510 12.340 ;
        RECT 60.990 11.830 61.340 13.080 ;
        RECT 64.690 11.510 65.030 12.340 ;
        RECT 66.510 11.830 66.860 13.080 ;
        RECT 68.625 12.425 69.835 13.515 ;
        RECT 68.625 11.715 69.145 12.255 ;
        RECT 69.315 11.885 69.835 12.425 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 70.465 13.080 75.810 13.515 ;
        RECT 75.985 13.080 81.330 13.515 ;
        RECT 57.585 10.965 62.930 11.510 ;
        RECT 63.105 10.965 68.450 11.510 ;
        RECT 68.625 10.965 69.835 11.715 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 72.050 11.510 72.390 12.340 ;
        RECT 73.870 11.830 74.220 13.080 ;
        RECT 77.570 11.510 77.910 12.340 ;
        RECT 79.390 11.830 79.740 13.080 ;
        RECT 81.505 12.425 82.715 13.515 ;
        RECT 81.505 11.715 82.025 12.255 ;
        RECT 82.195 11.885 82.715 12.425 ;
        RECT 82.885 12.350 83.175 13.515 ;
        RECT 83.345 13.080 88.690 13.515 ;
        RECT 88.865 13.080 94.210 13.515 ;
        RECT 70.465 10.965 75.810 11.510 ;
        RECT 75.985 10.965 81.330 11.510 ;
        RECT 81.505 10.965 82.715 11.715 ;
        RECT 82.885 10.965 83.175 11.690 ;
        RECT 84.930 11.510 85.270 12.340 ;
        RECT 86.750 11.830 87.100 13.080 ;
        RECT 90.450 11.510 90.790 12.340 ;
        RECT 92.270 11.830 92.620 13.080 ;
        RECT 94.385 12.425 95.595 13.515 ;
        RECT 94.385 11.715 94.905 12.255 ;
        RECT 95.075 11.885 95.595 12.425 ;
        RECT 95.765 12.350 96.055 13.515 ;
        RECT 96.225 13.080 101.570 13.515 ;
        RECT 101.745 13.080 107.090 13.515 ;
        RECT 83.345 10.965 88.690 11.510 ;
        RECT 88.865 10.965 94.210 11.510 ;
        RECT 94.385 10.965 95.595 11.715 ;
        RECT 95.765 10.965 96.055 11.690 ;
        RECT 97.810 11.510 98.150 12.340 ;
        RECT 99.630 11.830 99.980 13.080 ;
        RECT 103.330 11.510 103.670 12.340 ;
        RECT 105.150 11.830 105.500 13.080 ;
        RECT 107.265 12.425 108.475 13.515 ;
        RECT 107.265 11.715 107.785 12.255 ;
        RECT 107.955 11.885 108.475 12.425 ;
        RECT 108.645 12.350 108.935 13.515 ;
        RECT 109.105 13.080 114.450 13.515 ;
        RECT 114.625 13.080 119.970 13.515 ;
        RECT 96.225 10.965 101.570 11.510 ;
        RECT 101.745 10.965 107.090 11.510 ;
        RECT 107.265 10.965 108.475 11.715 ;
        RECT 108.645 10.965 108.935 11.690 ;
        RECT 110.690 11.510 111.030 12.340 ;
        RECT 112.510 11.830 112.860 13.080 ;
        RECT 116.210 11.510 116.550 12.340 ;
        RECT 118.030 11.830 118.380 13.080 ;
        RECT 120.145 12.425 121.355 13.515 ;
        RECT 120.145 11.715 120.665 12.255 ;
        RECT 120.835 11.885 121.355 12.425 ;
        RECT 121.525 12.350 121.815 13.515 ;
        RECT 121.985 12.425 123.655 13.515 ;
        RECT 121.985 11.735 122.735 12.255 ;
        RECT 122.905 11.905 123.655 12.425 ;
        RECT 124.285 12.425 125.495 13.515 ;
        RECT 124.285 11.885 124.805 12.425 ;
        RECT 109.105 10.965 114.450 11.510 ;
        RECT 114.625 10.965 119.970 11.510 ;
        RECT 120.145 10.965 121.355 11.715 ;
        RECT 121.525 10.965 121.815 11.690 ;
        RECT 121.985 10.965 123.655 11.735 ;
        RECT 124.975 11.715 125.495 12.255 ;
        RECT 124.285 10.965 125.495 11.715 ;
        RECT 5.520 10.795 125.580 10.965 ;
      LAYER met1 ;
        RECT 5.520 130.320 125.580 130.800 ;
        RECT 33.205 129.780 33.495 129.825 ;
        RECT 34.570 129.780 34.890 129.840 ;
        RECT 35.950 129.825 36.270 129.840 ;
        RECT 33.205 129.640 34.890 129.780 ;
        RECT 33.205 129.595 33.495 129.640 ;
        RECT 34.570 129.580 34.890 129.640 ;
        RECT 35.485 129.780 36.270 129.825 ;
        RECT 39.085 129.780 39.375 129.825 ;
        RECT 35.485 129.640 39.375 129.780 ;
        RECT 35.485 129.595 36.270 129.640 ;
        RECT 35.950 129.580 36.270 129.595 ;
        RECT 38.785 129.595 39.375 129.640 ;
        RECT 61.245 129.780 61.895 129.825 ;
        RECT 62.630 129.780 62.950 129.840 ;
        RECT 64.845 129.780 65.135 129.825 ;
        RECT 61.245 129.640 65.135 129.780 ;
        RECT 61.245 129.595 61.895 129.640 ;
        RECT 13.885 129.440 14.175 129.485 ;
        RECT 18.470 129.440 18.790 129.500 ;
        RECT 13.885 129.300 18.790 129.440 ;
        RECT 13.885 129.255 14.175 129.300 ;
        RECT 18.470 129.240 18.790 129.300 ;
        RECT 32.290 129.440 32.580 129.485 ;
        RECT 34.125 129.440 34.415 129.485 ;
        RECT 37.705 129.440 37.995 129.485 ;
        RECT 32.290 129.300 37.995 129.440 ;
        RECT 32.290 129.255 32.580 129.300 ;
        RECT 34.125 129.255 34.415 129.300 ;
        RECT 37.705 129.255 37.995 129.300 ;
        RECT 38.785 129.280 39.075 129.595 ;
        RECT 62.630 129.580 62.950 129.640 ;
        RECT 64.545 129.595 65.135 129.640 ;
        RECT 114.145 129.780 114.795 129.825 ;
        RECT 117.745 129.780 118.035 129.825 ;
        RECT 119.670 129.780 119.990 129.840 ;
        RECT 114.145 129.640 119.990 129.780 ;
        RECT 114.145 129.595 114.795 129.640 ;
        RECT 117.445 129.595 118.035 129.640 ;
        RECT 58.050 129.440 58.340 129.485 ;
        RECT 59.885 129.440 60.175 129.485 ;
        RECT 63.465 129.440 63.755 129.485 ;
        RECT 58.050 129.300 63.755 129.440 ;
        RECT 58.050 129.255 58.340 129.300 ;
        RECT 59.885 129.255 60.175 129.300 ;
        RECT 63.465 129.255 63.755 129.300 ;
        RECT 64.545 129.280 64.835 129.595 ;
        RECT 110.950 129.440 111.240 129.485 ;
        RECT 112.785 129.440 113.075 129.485 ;
        RECT 116.365 129.440 116.655 129.485 ;
        RECT 110.950 129.300 116.655 129.440 ;
        RECT 110.950 129.255 111.240 129.300 ;
        RECT 112.785 129.255 113.075 129.300 ;
        RECT 116.365 129.255 116.655 129.300 ;
        RECT 117.445 129.280 117.735 129.595 ;
        RECT 119.670 129.580 119.990 129.640 ;
        RECT 120.130 129.780 120.450 129.840 ;
        RECT 120.605 129.780 120.895 129.825 ;
        RECT 120.130 129.640 120.895 129.780 ;
        RECT 120.130 129.580 120.450 129.640 ;
        RECT 120.605 129.595 120.895 129.640 ;
        RECT 31.810 128.900 32.130 129.160 ;
        RECT 36.410 129.100 36.730 129.160 ;
        RECT 41.945 129.100 42.235 129.145 ;
        RECT 36.410 128.960 42.235 129.100 ;
        RECT 36.410 128.900 36.730 128.960 ;
        RECT 41.945 128.915 42.235 128.960 ;
        RECT 57.570 128.900 57.890 129.160 ;
        RECT 58.950 128.900 59.270 129.160 ;
        RECT 62.170 129.100 62.490 129.160 ;
        RECT 67.705 129.100 67.995 129.145 ;
        RECT 62.170 128.960 67.995 129.100 ;
        RECT 62.170 128.900 62.490 128.960 ;
        RECT 67.705 128.915 67.995 128.960 ;
        RECT 110.010 129.100 110.330 129.160 ;
        RECT 110.485 129.100 110.775 129.145 ;
        RECT 110.010 128.960 110.775 129.100 ;
        RECT 110.010 128.900 110.330 128.960 ;
        RECT 110.485 128.915 110.775 128.960 ;
        RECT 111.850 128.900 112.170 129.160 ;
        RECT 32.695 128.760 32.985 128.805 ;
        RECT 34.585 128.760 34.875 128.805 ;
        RECT 37.705 128.760 37.995 128.805 ;
        RECT 32.695 128.620 37.995 128.760 ;
        RECT 32.695 128.575 32.985 128.620 ;
        RECT 34.585 128.575 34.875 128.620 ;
        RECT 37.705 128.575 37.995 128.620 ;
        RECT 58.455 128.760 58.745 128.805 ;
        RECT 60.345 128.760 60.635 128.805 ;
        RECT 63.465 128.760 63.755 128.805 ;
        RECT 58.455 128.620 63.755 128.760 ;
        RECT 58.455 128.575 58.745 128.620 ;
        RECT 60.345 128.575 60.635 128.620 ;
        RECT 63.465 128.575 63.755 128.620 ;
        RECT 111.355 128.760 111.645 128.805 ;
        RECT 113.245 128.760 113.535 128.805 ;
        RECT 116.365 128.760 116.655 128.805 ;
        RECT 111.355 128.620 116.655 128.760 ;
        RECT 111.355 128.575 111.645 128.620 ;
        RECT 113.245 128.575 113.535 128.620 ;
        RECT 116.365 128.575 116.655 128.620 ;
        RECT 13.410 128.220 13.730 128.480 ;
        RECT 5.520 127.600 125.580 128.080 ;
        RECT 107.250 127.400 107.570 127.460 ;
        RECT 107.250 127.260 117.140 127.400 ;
        RECT 107.250 127.200 107.570 127.260 ;
        RECT 8.775 127.060 9.065 127.105 ;
        RECT 10.665 127.060 10.955 127.105 ;
        RECT 13.785 127.060 14.075 127.105 ;
        RECT 8.775 126.920 14.075 127.060 ;
        RECT 8.775 126.875 9.065 126.920 ;
        RECT 10.665 126.875 10.955 126.920 ;
        RECT 13.785 126.875 14.075 126.920 ;
        RECT 23.955 127.060 24.245 127.105 ;
        RECT 25.845 127.060 26.135 127.105 ;
        RECT 28.965 127.060 29.255 127.105 ;
        RECT 23.955 126.920 29.255 127.060 ;
        RECT 23.955 126.875 24.245 126.920 ;
        RECT 25.845 126.875 26.135 126.920 ;
        RECT 28.965 126.875 29.255 126.920 ;
        RECT 34.535 127.060 34.825 127.105 ;
        RECT 36.425 127.060 36.715 127.105 ;
        RECT 39.545 127.060 39.835 127.105 ;
        RECT 34.535 126.920 39.835 127.060 ;
        RECT 34.535 126.875 34.825 126.920 ;
        RECT 36.425 126.875 36.715 126.920 ;
        RECT 39.545 126.875 39.835 126.920 ;
        RECT 49.715 127.060 50.005 127.105 ;
        RECT 51.605 127.060 51.895 127.105 ;
        RECT 54.725 127.060 55.015 127.105 ;
        RECT 49.715 126.920 55.015 127.060 ;
        RECT 49.715 126.875 50.005 126.920 ;
        RECT 51.605 126.875 51.895 126.920 ;
        RECT 54.725 126.875 55.015 126.920 ;
        RECT 60.295 127.060 60.585 127.105 ;
        RECT 62.185 127.060 62.475 127.105 ;
        RECT 65.305 127.060 65.595 127.105 ;
        RECT 60.295 126.920 65.595 127.060 ;
        RECT 60.295 126.875 60.585 126.920 ;
        RECT 62.185 126.875 62.475 126.920 ;
        RECT 65.305 126.875 65.595 126.920 ;
        RECT 74.555 127.060 74.845 127.105 ;
        RECT 76.445 127.060 76.735 127.105 ;
        RECT 79.565 127.060 79.855 127.105 ;
        RECT 74.555 126.920 79.855 127.060 ;
        RECT 74.555 126.875 74.845 126.920 ;
        RECT 76.445 126.875 76.735 126.920 ;
        RECT 79.565 126.875 79.855 126.920 ;
        RECT 85.135 127.060 85.425 127.105 ;
        RECT 87.025 127.060 87.315 127.105 ;
        RECT 90.145 127.060 90.435 127.105 ;
        RECT 85.135 126.920 90.435 127.060 ;
        RECT 85.135 126.875 85.425 126.920 ;
        RECT 87.025 126.875 87.315 126.920 ;
        RECT 90.145 126.875 90.435 126.920 ;
        RECT 97.095 127.060 97.385 127.105 ;
        RECT 98.985 127.060 99.275 127.105 ;
        RECT 102.105 127.060 102.395 127.105 ;
        RECT 97.095 126.920 102.395 127.060 ;
        RECT 97.095 126.875 97.385 126.920 ;
        RECT 98.985 126.875 99.275 126.920 ;
        RECT 102.105 126.875 102.395 126.920 ;
        RECT 107.675 127.060 107.965 127.105 ;
        RECT 109.565 127.060 109.855 127.105 ;
        RECT 112.685 127.060 112.975 127.105 ;
        RECT 107.675 126.920 112.975 127.060 ;
        RECT 107.675 126.875 107.965 126.920 ;
        RECT 109.565 126.875 109.855 126.920 ;
        RECT 112.685 126.875 112.975 126.920 ;
        RECT 7.905 126.720 8.195 126.765 ;
        RECT 12.030 126.720 12.350 126.780 ;
        RECT 23.085 126.720 23.375 126.765 ;
        RECT 31.810 126.720 32.130 126.780 ;
        RECT 7.905 126.580 32.130 126.720 ;
        RECT 7.905 126.535 8.195 126.580 ;
        RECT 12.030 126.520 12.350 126.580 ;
        RECT 23.085 126.535 23.375 126.580 ;
        RECT 31.810 126.520 32.130 126.580 ;
        RECT 42.850 126.720 43.170 126.780 ;
        RECT 43.785 126.720 44.075 126.765 ;
        RECT 42.850 126.580 44.075 126.720 ;
        RECT 42.850 126.520 43.170 126.580 ;
        RECT 43.785 126.535 44.075 126.580 ;
        RECT 48.370 126.720 48.690 126.780 ;
        RECT 48.845 126.720 49.135 126.765 ;
        RECT 57.570 126.720 57.890 126.780 ;
        RECT 59.425 126.720 59.715 126.765 ;
        RECT 48.370 126.580 59.715 126.720 ;
        RECT 48.370 126.520 48.690 126.580 ;
        RECT 48.845 126.535 49.135 126.580 ;
        RECT 57.570 126.520 57.890 126.580 ;
        RECT 59.425 126.535 59.715 126.580 ;
        RECT 68.610 126.720 68.930 126.780 ;
        RECT 69.545 126.720 69.835 126.765 ;
        RECT 68.610 126.580 69.835 126.720 ;
        RECT 68.610 126.520 68.930 126.580 ;
        RECT 69.545 126.535 69.835 126.580 ;
        RECT 81.490 126.720 81.810 126.780 ;
        RECT 83.805 126.720 84.095 126.765 ;
        RECT 81.490 126.580 84.095 126.720 ;
        RECT 81.490 126.520 81.810 126.580 ;
        RECT 83.805 126.535 84.095 126.580 ;
        RECT 87.930 126.720 88.250 126.780 ;
        RECT 94.385 126.720 94.675 126.765 ;
        RECT 87.930 126.580 94.675 126.720 ;
        RECT 87.930 126.520 88.250 126.580 ;
        RECT 94.385 126.535 94.675 126.580 ;
        RECT 96.225 126.720 96.515 126.765 ;
        RECT 106.805 126.720 107.095 126.765 ;
        RECT 110.010 126.720 110.330 126.780 ;
        RECT 117.000 126.765 117.140 127.260 ;
        RECT 96.225 126.580 110.330 126.720 ;
        RECT 96.225 126.535 96.515 126.580 ;
        RECT 106.805 126.535 107.095 126.580 ;
        RECT 110.010 126.520 110.330 126.580 ;
        RECT 116.925 126.535 117.215 126.765 ;
        RECT 8.370 126.380 8.660 126.425 ;
        RECT 10.205 126.380 10.495 126.425 ;
        RECT 13.785 126.380 14.075 126.425 ;
        RECT 8.370 126.240 14.075 126.380 ;
        RECT 8.370 126.195 8.660 126.240 ;
        RECT 10.205 126.195 10.495 126.240 ;
        RECT 13.785 126.195 14.075 126.240 ;
        RECT 14.865 126.085 15.155 126.400 ;
        RECT 17.090 126.380 17.410 126.440 ;
        RECT 18.025 126.380 18.315 126.425 ;
        RECT 17.090 126.240 18.315 126.380 ;
        RECT 17.090 126.180 17.410 126.240 ;
        RECT 18.025 126.195 18.315 126.240 ;
        RECT 23.550 126.380 23.840 126.425 ;
        RECT 25.385 126.380 25.675 126.425 ;
        RECT 28.965 126.380 29.255 126.425 ;
        RECT 23.550 126.240 29.255 126.380 ;
        RECT 23.550 126.195 23.840 126.240 ;
        RECT 25.385 126.195 25.675 126.240 ;
        RECT 28.965 126.195 29.255 126.240 ;
        RECT 29.970 126.400 30.290 126.440 ;
        RECT 29.970 126.180 30.335 126.400 ;
        RECT 31.350 126.380 31.670 126.440 ;
        RECT 33.205 126.380 33.495 126.425 ;
        RECT 31.350 126.240 33.495 126.380 ;
        RECT 31.350 126.180 31.670 126.240 ;
        RECT 33.205 126.195 33.495 126.240 ;
        RECT 33.650 126.180 33.970 126.440 ;
        RECT 34.130 126.380 34.420 126.425 ;
        RECT 35.965 126.380 36.255 126.425 ;
        RECT 39.545 126.380 39.835 126.425 ;
        RECT 34.130 126.240 39.835 126.380 ;
        RECT 34.130 126.195 34.420 126.240 ;
        RECT 35.965 126.195 36.255 126.240 ;
        RECT 39.545 126.195 39.835 126.240 ;
        RECT 40.550 126.400 40.870 126.440 ;
        RECT 40.550 126.180 40.915 126.400 ;
        RECT 46.530 126.180 46.850 126.440 ;
        RECT 49.310 126.380 49.600 126.425 ;
        RECT 51.145 126.380 51.435 126.425 ;
        RECT 54.725 126.380 55.015 126.425 ;
        RECT 49.310 126.240 55.015 126.380 ;
        RECT 49.310 126.195 49.600 126.240 ;
        RECT 51.145 126.195 51.435 126.240 ;
        RECT 54.725 126.195 55.015 126.240 ;
        RECT 9.285 125.855 9.575 126.085 ;
        RECT 11.565 126.040 12.215 126.085 ;
        RECT 14.865 126.040 15.455 126.085 ;
        RECT 17.550 126.040 17.870 126.100 ;
        RECT 30.045 126.085 30.335 126.180 ;
        RECT 11.565 125.900 17.870 126.040 ;
        RECT 11.565 125.855 12.215 125.900 ;
        RECT 15.165 125.855 15.455 125.900 ;
        RECT 9.360 125.700 9.500 125.855 ;
        RECT 17.550 125.840 17.870 125.900 ;
        RECT 24.465 125.855 24.755 126.085 ;
        RECT 26.745 126.040 27.395 126.085 ;
        RECT 30.045 126.040 30.635 126.085 ;
        RECT 26.745 125.900 30.635 126.040 ;
        RECT 26.745 125.855 27.395 125.900 ;
        RECT 30.345 125.855 30.635 125.900 ;
        RECT 20.310 125.700 20.630 125.760 ;
        RECT 9.360 125.560 20.630 125.700 ;
        RECT 24.540 125.700 24.680 125.855 ;
        RECT 35.030 125.840 35.350 126.100 ;
        RECT 40.625 126.085 40.915 126.180 ;
        RECT 37.325 126.040 37.975 126.085 ;
        RECT 40.625 126.040 41.215 126.085 ;
        RECT 37.325 125.900 41.215 126.040 ;
        RECT 37.325 125.855 37.975 125.900 ;
        RECT 40.925 125.855 41.215 125.900 ;
        RECT 50.210 125.840 50.530 126.100 ;
        RECT 55.805 126.085 56.095 126.400 ;
        RECT 57.110 126.380 57.430 126.440 ;
        RECT 58.965 126.380 59.255 126.425 ;
        RECT 57.110 126.240 59.255 126.380 ;
        RECT 57.110 126.180 57.430 126.240 ;
        RECT 58.965 126.195 59.255 126.240 ;
        RECT 59.890 126.380 60.180 126.425 ;
        RECT 61.725 126.380 62.015 126.425 ;
        RECT 65.305 126.380 65.595 126.425 ;
        RECT 59.890 126.240 65.595 126.380 ;
        RECT 59.890 126.195 60.180 126.240 ;
        RECT 61.725 126.195 62.015 126.240 ;
        RECT 65.305 126.195 65.595 126.240 ;
        RECT 52.505 126.040 53.155 126.085 ;
        RECT 55.805 126.040 56.395 126.085 ;
        RECT 56.650 126.040 56.970 126.100 ;
        RECT 52.505 125.900 56.970 126.040 ;
        RECT 52.505 125.855 53.155 125.900 ;
        RECT 56.105 125.855 56.395 125.900 ;
        RECT 56.650 125.840 56.970 125.900 ;
        RECT 60.805 126.040 61.095 126.085 ;
        RECT 62.170 126.040 62.490 126.100 ;
        RECT 66.385 126.085 66.675 126.400 ;
        RECT 67.690 126.380 68.010 126.440 ;
        RECT 73.685 126.380 73.975 126.425 ;
        RECT 67.690 126.240 73.975 126.380 ;
        RECT 67.690 126.180 68.010 126.240 ;
        RECT 73.685 126.195 73.975 126.240 ;
        RECT 74.150 126.380 74.440 126.425 ;
        RECT 75.985 126.380 76.275 126.425 ;
        RECT 79.565 126.380 79.855 126.425 ;
        RECT 74.150 126.240 79.855 126.380 ;
        RECT 74.150 126.195 74.440 126.240 ;
        RECT 75.985 126.195 76.275 126.240 ;
        RECT 79.565 126.195 79.855 126.240 ;
        RECT 60.805 125.900 62.490 126.040 ;
        RECT 60.805 125.855 61.095 125.900 ;
        RECT 62.170 125.840 62.490 125.900 ;
        RECT 63.085 126.040 63.735 126.085 ;
        RECT 66.385 126.040 66.975 126.085 ;
        RECT 68.610 126.040 68.930 126.100 ;
        RECT 63.085 125.900 68.930 126.040 ;
        RECT 63.085 125.855 63.735 125.900 ;
        RECT 66.685 125.855 66.975 125.900 ;
        RECT 68.610 125.840 68.930 125.900 ;
        RECT 75.065 126.040 75.355 126.085 ;
        RECT 76.430 126.040 76.750 126.100 ;
        RECT 75.065 125.900 76.750 126.040 ;
        RECT 75.065 125.855 75.355 125.900 ;
        RECT 76.430 125.840 76.750 125.900 ;
        RECT 77.345 126.040 77.995 126.085 ;
        RECT 80.110 126.040 80.430 126.100 ;
        RECT 80.645 126.085 80.935 126.400 ;
        RECT 84.265 126.195 84.555 126.425 ;
        RECT 84.730 126.380 85.020 126.425 ;
        RECT 86.565 126.380 86.855 126.425 ;
        RECT 90.145 126.380 90.435 126.425 ;
        RECT 84.730 126.240 90.435 126.380 ;
        RECT 84.730 126.195 85.020 126.240 ;
        RECT 86.565 126.195 86.855 126.240 ;
        RECT 90.145 126.195 90.435 126.240 ;
        RECT 80.645 126.040 81.235 126.085 ;
        RECT 77.345 125.900 81.235 126.040 ;
        RECT 77.345 125.855 77.995 125.900 ;
        RECT 80.110 125.840 80.430 125.900 ;
        RECT 80.945 125.855 81.235 125.900 ;
        RECT 27.670 125.700 27.990 125.760 ;
        RECT 24.540 125.560 27.990 125.700 ;
        RECT 20.310 125.500 20.630 125.560 ;
        RECT 27.670 125.500 27.990 125.560 ;
        RECT 47.005 125.700 47.295 125.745 ;
        RECT 49.290 125.700 49.610 125.760 ;
        RECT 47.005 125.560 49.610 125.700 ;
        RECT 84.340 125.700 84.480 126.195 ;
        RECT 85.645 126.040 85.935 126.085 ;
        RECT 86.090 126.040 86.410 126.100 ;
        RECT 85.645 125.900 86.410 126.040 ;
        RECT 85.645 125.855 85.935 125.900 ;
        RECT 86.090 125.840 86.410 125.900 ;
        RECT 87.925 126.040 88.575 126.085 ;
        RECT 90.690 126.040 91.010 126.100 ;
        RECT 91.225 126.085 91.515 126.400 ;
        RECT 96.690 126.380 96.980 126.425 ;
        RECT 98.525 126.380 98.815 126.425 ;
        RECT 102.105 126.380 102.395 126.425 ;
        RECT 96.690 126.240 102.395 126.380 ;
        RECT 96.690 126.195 96.980 126.240 ;
        RECT 98.525 126.195 98.815 126.240 ;
        RECT 102.105 126.195 102.395 126.240 ;
        RECT 91.225 126.040 91.815 126.085 ;
        RECT 87.925 125.900 91.815 126.040 ;
        RECT 87.925 125.855 88.575 125.900 ;
        RECT 90.690 125.840 91.010 125.900 ;
        RECT 91.525 125.855 91.815 125.900 ;
        RECT 97.590 125.840 97.910 126.100 ;
        RECT 98.050 126.040 98.370 126.100 ;
        RECT 103.185 126.085 103.475 126.400 ;
        RECT 107.270 126.380 107.560 126.425 ;
        RECT 109.105 126.380 109.395 126.425 ;
        RECT 112.685 126.380 112.975 126.425 ;
        RECT 107.270 126.240 112.975 126.380 ;
        RECT 107.270 126.195 107.560 126.240 ;
        RECT 109.105 126.195 109.395 126.240 ;
        RECT 112.685 126.195 112.975 126.240 ;
        RECT 99.885 126.040 100.535 126.085 ;
        RECT 103.185 126.040 103.775 126.085 ;
        RECT 98.050 125.900 103.775 126.040 ;
        RECT 98.050 125.840 98.370 125.900 ;
        RECT 99.885 125.855 100.535 125.900 ;
        RECT 103.485 125.855 103.775 125.900 ;
        RECT 106.345 125.855 106.635 126.085 ;
        RECT 106.790 126.040 107.110 126.100 ;
        RECT 110.470 126.085 110.790 126.100 ;
        RECT 113.765 126.085 114.055 126.400 ;
        RECT 108.185 126.040 108.475 126.085 ;
        RECT 106.790 125.900 108.475 126.040 ;
        RECT 87.010 125.700 87.330 125.760 ;
        RECT 84.340 125.560 87.330 125.700 ;
        RECT 47.005 125.515 47.295 125.560 ;
        RECT 49.290 125.500 49.610 125.560 ;
        RECT 87.010 125.500 87.330 125.560 ;
        RECT 102.650 125.700 102.970 125.760 ;
        RECT 106.420 125.700 106.560 125.855 ;
        RECT 106.790 125.840 107.110 125.900 ;
        RECT 108.185 125.855 108.475 125.900 ;
        RECT 110.465 126.040 111.115 126.085 ;
        RECT 113.765 126.040 114.355 126.085 ;
        RECT 110.465 125.900 114.355 126.040 ;
        RECT 110.465 125.855 111.115 125.900 ;
        RECT 114.065 125.855 114.355 125.900 ;
        RECT 110.470 125.840 110.790 125.855 ;
        RECT 102.650 125.560 106.560 125.700 ;
        RECT 102.650 125.500 102.970 125.560 ;
        RECT 5.520 124.880 125.580 125.360 ;
        RECT 47.910 124.680 48.230 124.740 ;
        RECT 41.560 124.540 48.230 124.680 ;
        RECT 13.410 124.385 13.730 124.400 ;
        RECT 9.845 124.340 10.135 124.385 ;
        RECT 13.085 124.340 13.735 124.385 ;
        RECT 9.845 124.200 13.735 124.340 ;
        RECT 9.845 124.155 10.435 124.200 ;
        RECT 13.085 124.155 13.735 124.200 ;
        RECT 23.065 124.340 23.715 124.385 ;
        RECT 26.665 124.340 26.955 124.385 ;
        RECT 23.065 124.200 26.955 124.340 ;
        RECT 23.065 124.155 23.715 124.200 ;
        RECT 26.365 124.155 26.955 124.200 ;
        RECT 33.650 124.340 33.970 124.400 ;
        RECT 41.560 124.340 41.700 124.540 ;
        RECT 47.910 124.480 48.230 124.540 ;
        RECT 50.210 124.680 50.530 124.740 ;
        RECT 54.825 124.680 55.115 124.725 ;
        RECT 50.210 124.540 55.115 124.680 ;
        RECT 50.210 124.480 50.530 124.540 ;
        RECT 54.825 124.495 55.115 124.540 ;
        RECT 58.950 124.480 59.270 124.740 ;
        RECT 110.470 124.680 110.790 124.740 ;
        RECT 108.720 124.540 110.790 124.680 ;
        RECT 33.650 124.200 41.700 124.340 ;
        RECT 6.985 124.000 7.275 124.045 ;
        RECT 8.810 124.000 9.130 124.060 ;
        RECT 6.985 123.860 9.130 124.000 ;
        RECT 6.985 123.815 7.275 123.860 ;
        RECT 8.810 123.800 9.130 123.860 ;
        RECT 10.145 123.840 10.435 124.155 ;
        RECT 13.410 124.140 13.730 124.155 ;
        RECT 26.365 124.060 26.655 124.155 ;
        RECT 33.650 124.140 33.970 124.200 ;
        RECT 11.225 124.000 11.515 124.045 ;
        RECT 14.805 124.000 15.095 124.045 ;
        RECT 16.640 124.000 16.930 124.045 ;
        RECT 11.225 123.860 16.930 124.000 ;
        RECT 11.225 123.815 11.515 123.860 ;
        RECT 14.805 123.815 15.095 123.860 ;
        RECT 16.640 123.815 16.930 123.860 ;
        RECT 17.550 124.000 17.870 124.060 ;
        RECT 18.025 124.000 18.315 124.045 ;
        RECT 17.550 123.860 18.315 124.000 ;
        RECT 17.550 123.800 17.870 123.860 ;
        RECT 18.025 123.815 18.315 123.860 ;
        RECT 18.470 123.800 18.790 124.060 ;
        RECT 19.870 124.000 20.160 124.045 ;
        RECT 21.705 124.000 21.995 124.045 ;
        RECT 25.285 124.000 25.575 124.045 ;
        RECT 19.870 123.860 25.575 124.000 ;
        RECT 19.870 123.815 20.160 123.860 ;
        RECT 21.705 123.815 21.995 123.860 ;
        RECT 25.285 123.815 25.575 123.860 ;
        RECT 26.290 123.840 26.655 124.060 ;
        RECT 29.970 124.000 30.290 124.060 ;
        RECT 30.445 124.000 30.735 124.045 ;
        RECT 29.970 123.860 30.735 124.000 ;
        RECT 26.290 123.800 26.610 123.840 ;
        RECT 29.970 123.800 30.290 123.860 ;
        RECT 30.445 123.815 30.735 123.860 ;
        RECT 30.890 124.000 31.210 124.060 ;
        RECT 35.505 124.000 35.795 124.045 ;
        RECT 30.890 123.860 35.795 124.000 ;
        RECT 30.890 123.800 31.210 123.860 ;
        RECT 35.505 123.815 35.795 123.860 ;
        RECT 12.490 123.660 12.810 123.720 ;
        RECT 15.725 123.660 16.015 123.705 ;
        RECT 12.490 123.520 16.015 123.660 ;
        RECT 12.490 123.460 12.810 123.520 ;
        RECT 15.725 123.475 16.015 123.520 ;
        RECT 17.090 123.660 17.410 123.720 ;
        RECT 19.405 123.660 19.695 123.705 ;
        RECT 17.090 123.520 19.695 123.660 ;
        RECT 17.090 123.460 17.410 123.520 ;
        RECT 19.405 123.475 19.695 123.520 ;
        RECT 20.785 123.660 21.075 123.705 ;
        RECT 23.530 123.660 23.850 123.720 ;
        RECT 20.785 123.520 23.850 123.660 ;
        RECT 20.785 123.475 21.075 123.520 ;
        RECT 23.530 123.460 23.850 123.520 ;
        RECT 23.990 123.660 24.310 123.720 ;
        RECT 29.525 123.660 29.815 123.705 ;
        RECT 23.990 123.520 29.815 123.660 ;
        RECT 35.580 123.660 35.720 123.815 ;
        RECT 35.950 123.800 36.270 124.060 ;
        RECT 40.550 123.800 40.870 124.060 ;
        RECT 41.560 124.045 41.700 124.200 ;
        RECT 45.145 124.340 45.795 124.385 ;
        RECT 48.745 124.340 49.035 124.385 ;
        RECT 49.290 124.340 49.610 124.400 ;
        RECT 71.365 124.340 72.015 124.385 ;
        RECT 74.965 124.340 75.255 124.385 ;
        RECT 45.145 124.200 49.610 124.340 ;
        RECT 45.145 124.155 45.795 124.200 ;
        RECT 48.445 124.155 49.035 124.200 ;
        RECT 41.025 123.815 41.315 124.045 ;
        RECT 41.485 123.815 41.775 124.045 ;
        RECT 41.950 124.000 42.240 124.045 ;
        RECT 43.785 124.000 44.075 124.045 ;
        RECT 47.365 124.000 47.655 124.045 ;
        RECT 41.950 123.860 47.655 124.000 ;
        RECT 41.950 123.815 42.240 123.860 ;
        RECT 43.785 123.815 44.075 123.860 ;
        RECT 47.365 123.815 47.655 123.860 ;
        RECT 48.445 123.840 48.735 124.155 ;
        RECT 49.290 124.140 49.610 124.200 ;
        RECT 55.360 124.200 58.720 124.340 ;
        RECT 49.750 124.000 50.070 124.060 ;
        RECT 51.605 124.000 51.895 124.045 ;
        RECT 49.750 123.860 51.895 124.000 ;
        RECT 41.100 123.660 41.240 123.815 ;
        RECT 49.750 123.800 50.070 123.860 ;
        RECT 51.605 123.815 51.895 123.860 ;
        RECT 53.430 124.000 53.750 124.060 ;
        RECT 55.360 124.000 55.500 124.200 ;
        RECT 53.430 123.860 55.500 124.000 ;
        RECT 55.745 124.000 56.035 124.045 ;
        RECT 57.570 124.000 57.890 124.060 ;
        RECT 55.745 123.860 57.890 124.000 ;
        RECT 53.430 123.800 53.750 123.860 ;
        RECT 55.745 123.815 56.035 123.860 ;
        RECT 57.570 123.800 57.890 123.860 ;
        RECT 58.045 123.815 58.335 124.045 ;
        RECT 58.580 124.000 58.720 124.200 ;
        RECT 71.365 124.200 75.255 124.340 ;
        RECT 71.365 124.155 72.015 124.200 ;
        RECT 74.665 124.155 75.255 124.200 ;
        RECT 90.685 124.340 91.335 124.385 ;
        RECT 94.285 124.340 94.575 124.385 ;
        RECT 90.685 124.200 94.575 124.340 ;
        RECT 90.685 124.155 91.335 124.200 ;
        RECT 93.985 124.155 94.575 124.200 ;
        RECT 59.425 124.000 59.715 124.045 ;
        RECT 58.580 123.860 59.715 124.000 ;
        RECT 59.425 123.815 59.715 123.860 ;
        RECT 59.885 124.000 60.175 124.045 ;
        RECT 62.630 124.000 62.950 124.060 ;
        RECT 59.885 123.860 62.950 124.000 ;
        RECT 59.885 123.815 60.175 123.860 ;
        RECT 35.580 123.520 41.240 123.660 ;
        RECT 23.990 123.460 24.310 123.520 ;
        RECT 29.525 123.475 29.815 123.520 ;
        RECT 11.225 123.320 11.515 123.365 ;
        RECT 14.345 123.320 14.635 123.365 ;
        RECT 16.235 123.320 16.525 123.365 ;
        RECT 11.225 123.180 16.525 123.320 ;
        RECT 11.225 123.135 11.515 123.180 ;
        RECT 14.345 123.135 14.635 123.180 ;
        RECT 16.235 123.135 16.525 123.180 ;
        RECT 20.275 123.320 20.565 123.365 ;
        RECT 22.165 123.320 22.455 123.365 ;
        RECT 25.285 123.320 25.575 123.365 ;
        RECT 20.275 123.180 25.575 123.320 ;
        RECT 20.275 123.135 20.565 123.180 ;
        RECT 22.165 123.135 22.455 123.180 ;
        RECT 25.285 123.135 25.575 123.180 ;
        RECT 41.100 122.980 41.240 123.520 ;
        RECT 42.865 123.660 43.155 123.705 ;
        RECT 45.610 123.660 45.930 123.720 ;
        RECT 42.865 123.520 45.930 123.660 ;
        RECT 42.865 123.475 43.155 123.520 ;
        RECT 45.610 123.460 45.930 123.520 ;
        RECT 46.530 123.660 46.850 123.720 ;
        RECT 53.520 123.660 53.660 123.800 ;
        RECT 46.530 123.520 53.660 123.660 ;
        RECT 53.905 123.660 54.195 123.705 ;
        RECT 56.650 123.660 56.970 123.720 ;
        RECT 53.905 123.520 56.970 123.660 ;
        RECT 46.530 123.460 46.850 123.520 ;
        RECT 53.905 123.475 54.195 123.520 ;
        RECT 56.650 123.460 56.970 123.520 ;
        RECT 42.355 123.320 42.645 123.365 ;
        RECT 44.245 123.320 44.535 123.365 ;
        RECT 47.365 123.320 47.655 123.365 ;
        RECT 42.355 123.180 47.655 123.320 ;
        RECT 42.355 123.135 42.645 123.180 ;
        RECT 44.245 123.135 44.535 123.180 ;
        RECT 47.365 123.135 47.655 123.180 ;
        RECT 46.530 122.980 46.850 123.040 ;
        RECT 41.100 122.840 46.850 122.980 ;
        RECT 46.530 122.780 46.850 122.840 ;
        RECT 52.970 122.980 53.290 123.040 ;
        RECT 58.120 122.980 58.260 123.815 ;
        RECT 62.630 123.800 62.950 123.860 ;
        RECT 68.170 124.000 68.460 124.045 ;
        RECT 70.005 124.000 70.295 124.045 ;
        RECT 73.585 124.000 73.875 124.045 ;
        RECT 68.170 123.860 73.875 124.000 ;
        RECT 68.170 123.815 68.460 123.860 ;
        RECT 70.005 123.815 70.295 123.860 ;
        RECT 73.585 123.815 73.875 123.860 ;
        RECT 74.665 124.000 74.955 124.155 ;
        RECT 93.985 124.060 94.275 124.155 ;
        RECT 78.745 124.000 79.035 124.045 ;
        RECT 74.665 123.860 79.035 124.000 ;
        RECT 74.665 123.840 74.955 123.860 ;
        RECT 78.745 123.815 79.035 123.860 ;
        RECT 79.205 124.000 79.495 124.045 ;
        RECT 80.585 124.000 80.875 124.045 ;
        RECT 82.870 124.000 83.190 124.060 ;
        RECT 85.185 124.000 85.475 124.045 ;
        RECT 79.205 123.860 85.475 124.000 ;
        RECT 79.205 123.815 79.495 123.860 ;
        RECT 80.585 123.815 80.875 123.860 ;
        RECT 82.870 123.800 83.190 123.860 ;
        RECT 85.185 123.815 85.475 123.860 ;
        RECT 87.490 124.000 87.780 124.045 ;
        RECT 89.325 124.000 89.615 124.045 ;
        RECT 92.905 124.000 93.195 124.045 ;
        RECT 87.490 123.860 93.195 124.000 ;
        RECT 87.490 123.815 87.780 123.860 ;
        RECT 89.325 123.815 89.615 123.860 ;
        RECT 92.905 123.815 93.195 123.860 ;
        RECT 93.910 123.840 94.275 124.060 ;
        RECT 93.910 123.800 94.230 123.840 ;
        RECT 97.605 123.815 97.895 124.045 ;
        RECT 67.690 123.460 68.010 123.720 ;
        RECT 69.070 123.460 69.390 123.720 ;
        RECT 75.050 123.660 75.370 123.720 ;
        RECT 77.825 123.660 78.115 123.705 ;
        RECT 75.050 123.520 78.115 123.660 ;
        RECT 75.050 123.460 75.370 123.520 ;
        RECT 77.825 123.475 78.115 123.520 ;
        RECT 80.110 123.460 80.430 123.720 ;
        RECT 87.010 123.460 87.330 123.720 ;
        RECT 88.390 123.460 88.710 123.720 ;
        RECT 94.370 123.660 94.690 123.720 ;
        RECT 97.145 123.660 97.435 123.705 ;
        RECT 94.370 123.520 97.435 123.660 ;
        RECT 94.370 123.460 94.690 123.520 ;
        RECT 97.145 123.475 97.435 123.520 ;
        RECT 97.680 123.660 97.820 123.815 ;
        RECT 98.050 123.800 98.370 124.060 ;
        RECT 104.965 124.000 105.255 124.045 ;
        RECT 107.250 124.000 107.570 124.060 ;
        RECT 108.720 124.000 108.860 124.540 ;
        RECT 110.470 124.480 110.790 124.540 ;
        RECT 110.010 124.340 110.330 124.400 ;
        RECT 112.770 124.385 113.090 124.400 ;
        RECT 109.180 124.200 110.330 124.340 ;
        RECT 109.180 124.045 109.320 124.200 ;
        RECT 110.010 124.140 110.330 124.200 ;
        RECT 112.765 124.340 113.415 124.385 ;
        RECT 116.365 124.340 116.655 124.385 ;
        RECT 112.765 124.200 116.655 124.340 ;
        RECT 112.765 124.155 113.415 124.200 ;
        RECT 116.065 124.155 116.655 124.200 ;
        RECT 112.770 124.140 113.090 124.155 ;
        RECT 104.965 123.860 107.570 124.000 ;
        RECT 104.965 123.815 105.255 123.860 ;
        RECT 105.040 123.660 105.180 123.815 ;
        RECT 107.250 123.800 107.570 123.860 ;
        RECT 107.800 123.860 108.860 124.000 ;
        RECT 97.680 123.520 105.180 123.660 ;
        RECT 105.425 123.660 105.715 123.705 ;
        RECT 107.800 123.660 107.940 123.860 ;
        RECT 109.105 123.815 109.395 124.045 ;
        RECT 109.570 124.000 109.860 124.045 ;
        RECT 111.405 124.000 111.695 124.045 ;
        RECT 114.985 124.000 115.275 124.045 ;
        RECT 109.570 123.860 115.275 124.000 ;
        RECT 109.570 123.815 109.860 123.860 ;
        RECT 111.405 123.815 111.695 123.860 ;
        RECT 114.985 123.815 115.275 123.860 ;
        RECT 116.065 123.840 116.355 124.155 ;
        RECT 119.670 124.000 119.990 124.060 ;
        RECT 120.145 124.000 120.435 124.045 ;
        RECT 119.670 123.860 120.435 124.000 ;
        RECT 119.670 123.800 119.990 123.860 ;
        RECT 120.145 123.815 120.435 123.860 ;
        RECT 120.590 124.000 120.910 124.060 ;
        RECT 121.065 124.000 121.355 124.045 ;
        RECT 120.590 123.860 121.355 124.000 ;
        RECT 120.590 123.800 120.910 123.860 ;
        RECT 121.065 123.815 121.355 123.860 ;
        RECT 105.425 123.520 107.940 123.660 ;
        RECT 108.170 123.660 108.490 123.720 ;
        RECT 110.485 123.660 110.775 123.705 ;
        RECT 108.170 123.520 110.775 123.660 ;
        RECT 68.575 123.320 68.865 123.365 ;
        RECT 70.465 123.320 70.755 123.365 ;
        RECT 73.585 123.320 73.875 123.365 ;
        RECT 68.575 123.180 73.875 123.320 ;
        RECT 68.575 123.135 68.865 123.180 ;
        RECT 70.465 123.135 70.755 123.180 ;
        RECT 73.585 123.135 73.875 123.180 ;
        RECT 87.895 123.320 88.185 123.365 ;
        RECT 89.785 123.320 90.075 123.365 ;
        RECT 92.905 123.320 93.195 123.365 ;
        RECT 87.895 123.180 93.195 123.320 ;
        RECT 87.895 123.135 88.185 123.180 ;
        RECT 89.785 123.135 90.075 123.180 ;
        RECT 92.905 123.135 93.195 123.180 ;
        RECT 94.830 123.320 95.150 123.380 ;
        RECT 97.680 123.320 97.820 123.520 ;
        RECT 105.425 123.475 105.715 123.520 ;
        RECT 108.170 123.460 108.490 123.520 ;
        RECT 110.485 123.475 110.775 123.520 ;
        RECT 113.690 123.660 114.010 123.720 ;
        RECT 119.225 123.660 119.515 123.705 ;
        RECT 113.690 123.520 119.515 123.660 ;
        RECT 113.690 123.460 114.010 123.520 ;
        RECT 119.225 123.475 119.515 123.520 ;
        RECT 94.830 123.180 97.820 123.320 ;
        RECT 109.975 123.320 110.265 123.365 ;
        RECT 111.865 123.320 112.155 123.365 ;
        RECT 114.985 123.320 115.275 123.365 ;
        RECT 109.975 123.180 115.275 123.320 ;
        RECT 94.830 123.120 95.150 123.180 ;
        RECT 109.975 123.135 110.265 123.180 ;
        RECT 111.865 123.135 112.155 123.180 ;
        RECT 114.985 123.135 115.275 123.180 ;
        RECT 52.970 122.840 58.260 122.980 ;
        RECT 85.645 122.980 85.935 123.025 ;
        RECT 90.690 122.980 91.010 123.040 ;
        RECT 85.645 122.840 91.010 122.980 ;
        RECT 52.970 122.780 53.290 122.840 ;
        RECT 85.645 122.795 85.935 122.840 ;
        RECT 90.690 122.780 91.010 122.840 ;
        RECT 107.725 122.980 108.015 123.025 ;
        RECT 112.770 122.980 113.090 123.040 ;
        RECT 107.725 122.840 113.090 122.980 ;
        RECT 107.725 122.795 108.015 122.840 ;
        RECT 112.770 122.780 113.090 122.840 ;
        RECT 118.750 122.980 119.070 123.040 ;
        RECT 121.525 122.980 121.815 123.025 ;
        RECT 118.750 122.840 121.815 122.980 ;
        RECT 118.750 122.780 119.070 122.840 ;
        RECT 121.525 122.795 121.815 122.840 ;
        RECT 5.520 122.160 125.580 122.640 ;
        RECT 20.310 121.960 20.630 122.020 ;
        RECT 21.245 121.960 21.535 122.005 ;
        RECT 20.310 121.820 21.535 121.960 ;
        RECT 20.310 121.760 20.630 121.820 ;
        RECT 21.245 121.775 21.535 121.820 ;
        RECT 23.530 121.760 23.850 122.020 ;
        RECT 25.385 121.960 25.675 122.005 ;
        RECT 26.290 121.960 26.610 122.020 ;
        RECT 25.385 121.820 26.610 121.960 ;
        RECT 25.385 121.775 25.675 121.820 ;
        RECT 26.290 121.760 26.610 121.820 ;
        RECT 27.670 121.760 27.990 122.020 ;
        RECT 34.570 121.760 34.890 122.020 ;
        RECT 35.030 121.960 35.350 122.020 ;
        RECT 40.565 121.960 40.855 122.005 ;
        RECT 35.030 121.820 40.855 121.960 ;
        RECT 35.030 121.760 35.350 121.820 ;
        RECT 40.565 121.775 40.855 121.820 ;
        RECT 45.610 121.760 45.930 122.020 ;
        RECT 62.170 121.960 62.490 122.020 ;
        RECT 67.705 121.960 67.995 122.005 ;
        RECT 62.170 121.820 67.995 121.960 ;
        RECT 62.170 121.760 62.490 121.820 ;
        RECT 67.705 121.775 67.995 121.820 ;
        RECT 69.070 121.960 69.390 122.020 ;
        RECT 75.525 121.960 75.815 122.005 ;
        RECT 69.070 121.820 75.815 121.960 ;
        RECT 69.070 121.760 69.390 121.820 ;
        RECT 75.525 121.775 75.815 121.820 ;
        RECT 76.430 121.960 76.750 122.020 ;
        RECT 78.745 121.960 79.035 122.005 ;
        RECT 76.430 121.820 79.035 121.960 ;
        RECT 76.430 121.760 76.750 121.820 ;
        RECT 78.745 121.775 79.035 121.820 ;
        RECT 85.185 121.960 85.475 122.005 ;
        RECT 86.550 121.960 86.870 122.020 ;
        RECT 85.185 121.820 86.870 121.960 ;
        RECT 85.185 121.775 85.475 121.820 ;
        RECT 86.550 121.760 86.870 121.820 ;
        RECT 88.390 121.960 88.710 122.020 ;
        RECT 89.325 121.960 89.615 122.005 ;
        RECT 88.390 121.820 89.615 121.960 ;
        RECT 88.390 121.760 88.710 121.820 ;
        RECT 89.325 121.775 89.615 121.820 ;
        RECT 93.910 121.760 94.230 122.020 ;
        RECT 103.125 121.960 103.415 122.005 ;
        RECT 106.790 121.960 107.110 122.020 ;
        RECT 103.125 121.820 107.110 121.960 ;
        RECT 103.125 121.775 103.415 121.820 ;
        RECT 106.790 121.760 107.110 121.820 ;
        RECT 108.170 121.760 108.490 122.020 ;
        RECT 120.590 121.960 120.910 122.020 ;
        RECT 108.720 121.820 120.910 121.960 ;
        RECT 11.225 121.620 11.515 121.665 ;
        RECT 14.345 121.620 14.635 121.665 ;
        RECT 16.235 121.620 16.525 121.665 ;
        RECT 58.950 121.620 59.270 121.680 ;
        RECT 11.225 121.480 16.525 121.620 ;
        RECT 11.225 121.435 11.515 121.480 ;
        RECT 14.345 121.435 14.635 121.480 ;
        RECT 16.235 121.435 16.525 121.480 ;
        RECT 41.560 121.480 59.270 121.620 ;
        RECT 4.210 121.280 4.530 121.340 ;
        RECT 6.985 121.280 7.275 121.325 ;
        RECT 4.210 121.140 7.275 121.280 ;
        RECT 4.210 121.080 4.530 121.140 ;
        RECT 6.985 121.095 7.275 121.140 ;
        RECT 12.030 121.280 12.350 121.340 ;
        RECT 17.090 121.280 17.410 121.340 ;
        RECT 12.030 121.140 17.410 121.280 ;
        RECT 12.030 121.080 12.350 121.140 ;
        RECT 17.090 121.080 17.410 121.140 ;
        RECT 18.470 121.280 18.790 121.340 ;
        RECT 30.890 121.280 31.210 121.340 ;
        RECT 18.470 121.140 31.210 121.280 ;
        RECT 18.470 121.080 18.790 121.140 ;
        RECT 10.145 120.645 10.435 120.960 ;
        RECT 11.225 120.940 11.515 120.985 ;
        RECT 14.805 120.940 15.095 120.985 ;
        RECT 16.640 120.940 16.930 120.985 ;
        RECT 11.225 120.800 16.930 120.940 ;
        RECT 11.225 120.755 11.515 120.800 ;
        RECT 14.805 120.755 15.095 120.800 ;
        RECT 16.640 120.755 16.930 120.800 ;
        RECT 22.150 120.740 22.470 121.000 ;
        RECT 25.920 120.985 26.060 121.140 ;
        RECT 30.890 121.080 31.210 121.140 ;
        RECT 24.465 120.755 24.755 120.985 ;
        RECT 25.845 120.755 26.135 120.985 ;
        RECT 13.410 120.645 13.730 120.660 ;
        RECT 9.845 120.600 10.435 120.645 ;
        RECT 13.085 120.600 13.735 120.645 ;
        RECT 9.845 120.460 13.735 120.600 ;
        RECT 9.845 120.415 10.135 120.460 ;
        RECT 13.085 120.415 13.735 120.460 ;
        RECT 15.725 120.415 16.015 120.645 ;
        RECT 24.540 120.600 24.680 120.755 ;
        RECT 28.590 120.740 28.910 121.000 ;
        RECT 35.490 120.740 35.810 121.000 ;
        RECT 41.560 120.985 41.700 121.480 ;
        RECT 58.950 121.420 59.270 121.480 ;
        RECT 68.610 121.620 68.930 121.680 ;
        RECT 70.925 121.620 71.215 121.665 ;
        RECT 68.610 121.480 71.215 121.620 ;
        RECT 68.610 121.420 68.930 121.480 ;
        RECT 70.925 121.435 71.215 121.480 ;
        RECT 93.005 121.620 93.295 121.665 ;
        RECT 97.590 121.620 97.910 121.680 ;
        RECT 93.005 121.480 97.910 121.620 ;
        RECT 93.005 121.435 93.295 121.480 ;
        RECT 97.590 121.420 97.910 121.480 ;
        RECT 107.250 121.620 107.570 121.680 ;
        RECT 108.720 121.620 108.860 121.820 ;
        RECT 120.590 121.760 120.910 121.820 ;
        RECT 107.250 121.480 108.860 121.620 ;
        RECT 111.815 121.620 112.105 121.665 ;
        RECT 113.705 121.620 113.995 121.665 ;
        RECT 116.825 121.620 117.115 121.665 ;
        RECT 111.815 121.480 117.115 121.620 ;
        RECT 107.250 121.420 107.570 121.480 ;
        RECT 111.815 121.435 112.105 121.480 ;
        RECT 113.705 121.435 113.995 121.480 ;
        RECT 116.825 121.435 117.115 121.480 ;
        RECT 53.430 121.080 53.750 121.340 ;
        RECT 74.145 121.280 74.435 121.325 ;
        RECT 82.870 121.280 83.190 121.340 ;
        RECT 108.170 121.280 108.490 121.340 ;
        RECT 74.145 121.140 94.600 121.280 ;
        RECT 74.145 121.095 74.435 121.140 ;
        RECT 41.485 120.755 41.775 120.985 ;
        RECT 46.530 120.740 46.850 121.000 ;
        RECT 54.825 120.755 55.115 120.985 ;
        RECT 26.750 120.600 27.070 120.660 ;
        RECT 24.540 120.460 27.070 120.600 ;
        RECT 54.900 120.600 55.040 120.755 ;
        RECT 58.490 120.740 58.810 121.000 ;
        RECT 68.150 120.940 68.470 121.000 ;
        RECT 68.625 120.940 68.915 120.985 ;
        RECT 68.150 120.800 68.915 120.940 ;
        RECT 68.150 120.740 68.470 120.800 ;
        RECT 68.625 120.755 68.915 120.800 ;
        RECT 71.385 120.940 71.675 120.985 ;
        RECT 74.220 120.940 74.360 121.095 ;
        RECT 82.870 121.080 83.190 121.140 ;
        RECT 75.050 120.940 75.370 121.000 ;
        RECT 71.385 120.800 74.360 120.940 ;
        RECT 74.680 120.800 75.370 120.940 ;
        RECT 71.385 120.755 71.675 120.800 ;
        RECT 74.680 120.600 74.820 120.800 ;
        RECT 75.050 120.740 75.370 120.800 ;
        RECT 76.430 120.740 76.750 121.000 ;
        RECT 79.665 120.940 79.955 120.985 ;
        RECT 81.490 120.940 81.810 121.000 ;
        RECT 79.665 120.800 81.810 120.940 ;
        RECT 79.665 120.755 79.955 120.800 ;
        RECT 81.490 120.740 81.810 120.800 ;
        RECT 84.265 120.940 84.555 120.985 ;
        RECT 88.390 120.940 88.710 121.000 ;
        RECT 84.265 120.800 88.710 120.940 ;
        RECT 84.265 120.755 84.555 120.800 ;
        RECT 88.390 120.740 88.710 120.800 ;
        RECT 90.230 120.740 90.550 121.000 ;
        RECT 92.070 120.740 92.390 121.000 ;
        RECT 94.460 120.985 94.600 121.140 ;
        RECT 105.960 121.140 108.490 121.280 ;
        RECT 94.385 120.940 94.675 120.985 ;
        RECT 94.830 120.940 95.150 121.000 ;
        RECT 94.385 120.800 95.150 120.940 ;
        RECT 94.385 120.755 94.675 120.800 ;
        RECT 94.830 120.740 95.150 120.800 ;
        RECT 102.205 120.940 102.495 120.985 ;
        RECT 104.490 120.940 104.810 121.000 ;
        RECT 105.960 120.985 106.100 121.140 ;
        RECT 108.170 121.080 108.490 121.140 ;
        RECT 121.065 121.280 121.355 121.325 ;
        RECT 126.570 121.280 126.890 121.340 ;
        RECT 121.065 121.140 126.890 121.280 ;
        RECT 121.065 121.095 121.355 121.140 ;
        RECT 126.570 121.080 126.890 121.140 ;
        RECT 102.205 120.800 104.810 120.940 ;
        RECT 102.205 120.755 102.495 120.800 ;
        RECT 104.490 120.740 104.810 120.800 ;
        RECT 105.885 120.755 106.175 120.985 ;
        RECT 107.265 120.940 107.555 120.985 ;
        RECT 106.420 120.800 107.555 120.940 ;
        RECT 54.900 120.460 74.820 120.600 ;
        RECT 104.030 120.600 104.350 120.660 ;
        RECT 106.420 120.600 106.560 120.800 ;
        RECT 107.265 120.755 107.555 120.800 ;
        RECT 108.630 120.940 108.950 121.000 ;
        RECT 109.565 120.940 109.855 120.985 ;
        RECT 108.630 120.800 109.855 120.940 ;
        RECT 108.630 120.740 108.950 120.800 ;
        RECT 109.565 120.755 109.855 120.800 ;
        RECT 110.010 120.940 110.330 121.000 ;
        RECT 110.945 120.940 111.235 120.985 ;
        RECT 110.010 120.800 111.235 120.940 ;
        RECT 110.010 120.740 110.330 120.800 ;
        RECT 110.945 120.755 111.235 120.800 ;
        RECT 111.410 120.940 111.700 120.985 ;
        RECT 113.245 120.940 113.535 120.985 ;
        RECT 116.825 120.940 117.115 120.985 ;
        RECT 111.410 120.800 117.115 120.940 ;
        RECT 111.410 120.755 111.700 120.800 ;
        RECT 113.245 120.755 113.535 120.800 ;
        RECT 116.825 120.755 117.115 120.800 ;
        RECT 111.850 120.600 112.170 120.660 ;
        RECT 117.905 120.645 118.195 120.960 ;
        RECT 104.030 120.460 106.560 120.600 ;
        RECT 106.880 120.460 112.170 120.600 ;
        RECT 13.410 120.400 13.730 120.415 ;
        RECT 11.110 120.260 11.430 120.320 ;
        RECT 15.800 120.260 15.940 120.415 ;
        RECT 26.750 120.400 27.070 120.460 ;
        RECT 104.030 120.400 104.350 120.460 ;
        RECT 11.110 120.120 15.940 120.260 ;
        RECT 58.965 120.260 59.255 120.305 ;
        RECT 63.090 120.260 63.410 120.320 ;
        RECT 106.880 120.305 107.020 120.460 ;
        RECT 111.850 120.400 112.170 120.460 ;
        RECT 112.325 120.415 112.615 120.645 ;
        RECT 114.605 120.600 115.255 120.645 ;
        RECT 117.905 120.600 118.495 120.645 ;
        RECT 118.750 120.600 119.070 120.660 ;
        RECT 114.605 120.460 119.070 120.600 ;
        RECT 114.605 120.415 115.255 120.460 ;
        RECT 118.205 120.415 118.495 120.460 ;
        RECT 58.965 120.120 63.410 120.260 ;
        RECT 11.110 120.060 11.430 120.120 ;
        RECT 58.965 120.075 59.255 120.120 ;
        RECT 63.090 120.060 63.410 120.120 ;
        RECT 106.805 120.075 107.095 120.305 ;
        RECT 110.485 120.260 110.775 120.305 ;
        RECT 112.400 120.260 112.540 120.415 ;
        RECT 118.750 120.400 119.070 120.460 ;
        RECT 110.485 120.120 112.540 120.260 ;
        RECT 110.485 120.075 110.775 120.120 ;
        RECT 5.520 119.440 125.580 119.920 ;
        RECT 11.110 119.040 11.430 119.300 ;
        RECT 12.490 119.040 12.810 119.300 ;
        RECT 13.410 119.040 13.730 119.300 ;
        RECT 1.910 118.560 2.230 118.620 ;
        RECT 6.985 118.560 7.275 118.605 ;
        RECT 1.910 118.420 7.275 118.560 ;
        RECT 1.910 118.360 2.230 118.420 ;
        RECT 6.985 118.375 7.275 118.420 ;
        RECT 10.205 118.375 10.495 118.605 ;
        RECT 11.585 118.560 11.875 118.605 ;
        RECT 12.030 118.560 12.350 118.620 ;
        RECT 11.585 118.420 12.350 118.560 ;
        RECT 11.585 118.375 11.875 118.420 ;
        RECT 10.280 118.220 10.420 118.375 ;
        RECT 12.030 118.360 12.350 118.420 ;
        RECT 13.885 118.560 14.175 118.605 ;
        RECT 18.470 118.560 18.790 118.620 ;
        RECT 13.885 118.420 18.790 118.560 ;
        RECT 13.885 118.375 14.175 118.420 ;
        RECT 18.470 118.360 18.790 118.420 ;
        RECT 75.050 118.560 75.370 118.620 ;
        RECT 89.325 118.560 89.615 118.605 ;
        RECT 96.210 118.560 96.530 118.620 ;
        RECT 75.050 118.420 96.530 118.560 ;
        RECT 75.050 118.360 75.370 118.420 ;
        RECT 89.325 118.375 89.615 118.420 ;
        RECT 96.210 118.360 96.530 118.420 ;
        RECT 31.350 118.220 31.670 118.280 ;
        RECT 10.280 118.080 31.670 118.220 ;
        RECT 31.350 118.020 31.670 118.080 ;
        RECT 7.905 117.880 8.195 117.925 ;
        RECT 58.490 117.880 58.810 117.940 ;
        RECT 7.905 117.740 58.810 117.880 ;
        RECT 7.905 117.695 8.195 117.740 ;
        RECT 58.490 117.680 58.810 117.740 ;
        RECT 88.850 117.340 89.170 117.600 ;
        RECT 5.520 116.720 125.580 117.200 ;
        RECT 87.440 116.180 87.730 116.225 ;
        RECT 90.220 116.180 90.510 116.225 ;
        RECT 92.080 116.180 92.370 116.225 ;
        RECT 87.440 116.040 92.370 116.180 ;
        RECT 87.440 115.995 87.730 116.040 ;
        RECT 90.220 115.995 90.510 116.040 ;
        RECT 92.080 115.995 92.370 116.040 ;
        RECT 112.330 116.180 112.620 116.225 ;
        RECT 114.190 116.180 114.480 116.225 ;
        RECT 116.970 116.180 117.260 116.225 ;
        RECT 112.330 116.040 117.260 116.180 ;
        RECT 112.330 115.995 112.620 116.040 ;
        RECT 114.190 115.995 114.480 116.040 ;
        RECT 116.970 115.995 117.260 116.040 ;
        RECT 113.705 115.840 113.995 115.885 ;
        RECT 119.210 115.840 119.530 115.900 ;
        RECT 113.705 115.700 119.530 115.840 ;
        RECT 113.705 115.655 113.995 115.700 ;
        RECT 119.210 115.640 119.530 115.700 ;
        RECT 16.170 115.300 16.490 115.560 ;
        RECT 47.925 115.500 48.215 115.545 ;
        RECT 48.370 115.500 48.690 115.560 ;
        RECT 47.925 115.360 48.690 115.500 ;
        RECT 47.925 115.315 48.215 115.360 ;
        RECT 48.370 115.300 48.690 115.360 ;
        RECT 55.745 115.500 56.035 115.545 ;
        RECT 57.570 115.500 57.890 115.560 ;
        RECT 55.745 115.360 57.890 115.500 ;
        RECT 55.745 115.315 56.035 115.360 ;
        RECT 57.570 115.300 57.890 115.360 ;
        RECT 60.805 115.500 61.095 115.545 ;
        RECT 61.710 115.500 62.030 115.560 ;
        RECT 60.805 115.360 62.030 115.500 ;
        RECT 60.805 115.315 61.095 115.360 ;
        RECT 61.710 115.300 62.030 115.360 ;
        RECT 87.440 115.500 87.730 115.545 ;
        RECT 87.440 115.360 89.975 115.500 ;
        RECT 87.440 115.315 87.730 115.360 ;
        RECT 88.850 115.205 89.170 115.220 ;
        RECT 85.580 115.160 85.870 115.205 ;
        RECT 88.840 115.160 89.170 115.205 ;
        RECT 85.580 115.020 89.170 115.160 ;
        RECT 85.580 114.975 85.870 115.020 ;
        RECT 88.840 114.975 89.170 115.020 ;
        RECT 89.760 115.205 89.975 115.360 ;
        RECT 90.690 115.300 91.010 115.560 ;
        RECT 92.545 115.500 92.835 115.545 ;
        RECT 95.290 115.500 95.610 115.560 ;
        RECT 92.545 115.360 95.610 115.500 ;
        RECT 92.545 115.315 92.835 115.360 ;
        RECT 95.290 115.300 95.610 115.360 ;
        RECT 96.210 115.300 96.530 115.560 ;
        RECT 97.605 115.500 97.895 115.545 ;
        RECT 100.365 115.500 100.655 115.545 ;
        RECT 102.190 115.500 102.510 115.560 ;
        RECT 97.605 115.360 102.510 115.500 ;
        RECT 97.605 115.315 97.895 115.360 ;
        RECT 100.365 115.315 100.655 115.360 ;
        RECT 102.190 115.300 102.510 115.360 ;
        RECT 103.570 115.300 103.890 115.560 ;
        RECT 110.010 115.500 110.330 115.560 ;
        RECT 111.865 115.500 112.155 115.545 ;
        RECT 116.970 115.500 117.260 115.545 ;
        RECT 110.010 115.360 112.155 115.500 ;
        RECT 110.010 115.300 110.330 115.360 ;
        RECT 111.865 115.315 112.155 115.360 ;
        RECT 114.725 115.360 117.260 115.500 ;
        RECT 114.725 115.205 114.940 115.360 ;
        RECT 116.970 115.315 117.260 115.360 ;
        RECT 89.760 115.160 90.050 115.205 ;
        RECT 91.620 115.160 91.910 115.205 ;
        RECT 89.760 115.020 91.910 115.160 ;
        RECT 89.760 114.975 90.050 115.020 ;
        RECT 91.620 114.975 91.910 115.020 ;
        RECT 112.790 115.160 113.080 115.205 ;
        RECT 114.650 115.160 114.940 115.205 ;
        RECT 112.790 115.020 114.940 115.160 ;
        RECT 112.790 114.975 113.080 115.020 ;
        RECT 114.650 114.975 114.940 115.020 ;
        RECT 115.570 115.160 115.860 115.205 ;
        RECT 118.830 115.160 119.120 115.205 ;
        RECT 122.430 115.160 122.750 115.220 ;
        RECT 115.570 115.020 122.750 115.160 ;
        RECT 115.570 114.975 115.860 115.020 ;
        RECT 118.830 114.975 119.120 115.020 ;
        RECT 88.850 114.960 89.170 114.975 ;
        RECT 122.430 114.960 122.750 115.020 ;
        RECT 13.410 114.820 13.730 114.880 ;
        RECT 15.265 114.820 15.555 114.865 ;
        RECT 13.410 114.680 15.555 114.820 ;
        RECT 13.410 114.620 13.730 114.680 ;
        RECT 15.265 114.635 15.555 114.680 ;
        RECT 47.910 114.820 48.230 114.880 ;
        RECT 48.385 114.820 48.675 114.865 ;
        RECT 47.910 114.680 48.675 114.820 ;
        RECT 47.910 114.620 48.230 114.680 ;
        RECT 48.385 114.635 48.675 114.680 ;
        RECT 56.650 114.620 56.970 114.880 ;
        RECT 61.250 114.620 61.570 114.880 ;
        RECT 83.330 114.865 83.650 114.880 ;
        RECT 83.330 114.635 83.865 114.865 ;
        RECT 83.330 114.620 83.650 114.635 ;
        RECT 99.890 114.620 100.210 114.880 ;
        RECT 104.505 114.820 104.795 114.865 ;
        RECT 105.870 114.820 106.190 114.880 ;
        RECT 104.505 114.680 106.190 114.820 ;
        RECT 104.505 114.635 104.795 114.680 ;
        RECT 105.870 114.620 106.190 114.680 ;
        RECT 118.290 114.820 118.610 114.880 ;
        RECT 120.835 114.820 121.125 114.865 ;
        RECT 118.290 114.680 121.125 114.820 ;
        RECT 118.290 114.620 118.610 114.680 ;
        RECT 120.835 114.635 121.125 114.680 ;
        RECT 5.520 114.000 125.580 114.480 ;
        RECT 52.510 113.800 52.830 113.860 ;
        RECT 45.240 113.660 52.830 113.800 ;
        RECT 12.510 113.460 12.800 113.505 ;
        RECT 14.370 113.460 14.660 113.505 ;
        RECT 12.510 113.320 14.660 113.460 ;
        RECT 12.510 113.275 12.800 113.320 ;
        RECT 14.370 113.275 14.660 113.320 ;
        RECT 15.290 113.460 15.580 113.505 ;
        RECT 17.090 113.460 17.410 113.520 ;
        RECT 18.550 113.460 18.840 113.505 ;
        RECT 15.290 113.320 18.840 113.460 ;
        RECT 15.290 113.275 15.580 113.320 ;
        RECT 11.570 113.120 11.890 113.180 ;
        RECT 14.445 113.120 14.660 113.275 ;
        RECT 17.090 113.260 17.410 113.320 ;
        RECT 18.550 113.275 18.840 113.320 ;
        RECT 22.630 113.460 22.920 113.505 ;
        RECT 24.490 113.460 24.780 113.505 ;
        RECT 22.630 113.320 24.780 113.460 ;
        RECT 22.630 113.275 22.920 113.320 ;
        RECT 24.490 113.275 24.780 113.320 ;
        RECT 25.410 113.460 25.700 113.505 ;
        RECT 27.210 113.460 27.530 113.520 ;
        RECT 28.670 113.460 28.960 113.505 ;
        RECT 25.410 113.320 28.960 113.460 ;
        RECT 25.410 113.275 25.700 113.320 ;
        RECT 16.690 113.120 16.980 113.165 ;
        RECT 11.570 112.980 14.100 113.120 ;
        RECT 14.445 112.980 16.980 113.120 ;
        RECT 11.570 112.920 11.890 112.980 ;
        RECT 13.410 112.580 13.730 112.840 ;
        RECT 13.960 112.780 14.100 112.980 ;
        RECT 16.690 112.935 16.980 112.980 ;
        RECT 21.705 113.120 21.995 113.165 ;
        RECT 24.565 113.120 24.780 113.275 ;
        RECT 27.210 113.260 27.530 113.320 ;
        RECT 28.670 113.275 28.960 113.320 ;
        RECT 34.125 113.460 34.415 113.505 ;
        RECT 43.555 113.460 43.845 113.505 ;
        RECT 45.240 113.460 45.380 113.660 ;
        RECT 52.510 113.600 52.830 113.660 ;
        RECT 83.330 113.800 83.650 113.860 ;
        RECT 86.105 113.800 86.395 113.845 ;
        RECT 88.850 113.800 89.170 113.860 ;
        RECT 83.330 113.660 89.170 113.800 ;
        RECT 83.330 113.600 83.650 113.660 ;
        RECT 86.105 113.615 86.395 113.660 ;
        RECT 88.850 113.600 89.170 113.660 ;
        RECT 89.785 113.800 90.075 113.845 ;
        RECT 90.690 113.800 91.010 113.860 ;
        RECT 89.785 113.660 91.010 113.800 ;
        RECT 89.785 113.615 90.075 113.660 ;
        RECT 90.690 113.600 91.010 113.660 ;
        RECT 103.570 113.600 103.890 113.860 ;
        RECT 34.125 113.320 45.380 113.460 ;
        RECT 45.560 113.460 45.850 113.505 ;
        RECT 47.910 113.460 48.230 113.520 ;
        RECT 48.820 113.460 49.110 113.505 ;
        RECT 45.560 113.320 49.110 113.460 ;
        RECT 34.125 113.275 34.415 113.320 ;
        RECT 43.555 113.275 43.845 113.320 ;
        RECT 45.560 113.275 45.850 113.320 ;
        RECT 47.910 113.260 48.230 113.320 ;
        RECT 48.820 113.275 49.110 113.320 ;
        RECT 49.740 113.460 50.030 113.505 ;
        RECT 51.600 113.460 51.890 113.505 ;
        RECT 49.740 113.320 51.890 113.460 ;
        RECT 49.740 113.275 50.030 113.320 ;
        RECT 51.600 113.275 51.890 113.320 ;
        RECT 59.820 113.460 60.110 113.505 ;
        RECT 61.250 113.460 61.570 113.520 ;
        RECT 63.080 113.460 63.370 113.505 ;
        RECT 59.820 113.320 63.370 113.460 ;
        RECT 59.820 113.275 60.110 113.320 ;
        RECT 26.810 113.120 27.100 113.165 ;
        RECT 33.665 113.120 33.955 113.165 ;
        RECT 21.705 112.980 24.220 113.120 ;
        RECT 24.565 112.980 27.100 113.120 ;
        RECT 21.705 112.935 21.995 112.980 ;
        RECT 21.780 112.780 21.920 112.935 ;
        RECT 13.960 112.640 21.920 112.780 ;
        RECT 23.530 112.580 23.850 112.840 ;
        RECT 24.080 112.780 24.220 112.980 ;
        RECT 26.810 112.935 27.100 112.980 ;
        RECT 32.360 112.980 33.955 113.120 ;
        RECT 27.670 112.780 27.990 112.840 ;
        RECT 24.080 112.640 27.990 112.780 ;
        RECT 27.670 112.580 27.990 112.640 ;
        RECT 32.360 112.500 32.500 112.980 ;
        RECT 33.665 112.935 33.955 112.980 ;
        RECT 36.870 112.920 37.190 113.180 ;
        RECT 38.725 112.935 39.015 113.165 ;
        RECT 34.570 112.580 34.890 112.840 ;
        RECT 38.800 112.780 38.940 112.935 ;
        RECT 41.010 112.920 41.330 113.180 ;
        RECT 42.405 112.935 42.695 113.165 ;
        RECT 47.420 113.120 47.710 113.165 ;
        RECT 49.740 113.120 49.955 113.275 ;
        RECT 61.250 113.260 61.570 113.320 ;
        RECT 63.080 113.275 63.370 113.320 ;
        RECT 64.000 113.460 64.290 113.505 ;
        RECT 65.860 113.460 66.150 113.505 ;
        RECT 64.000 113.320 66.150 113.460 ;
        RECT 64.000 113.275 64.290 113.320 ;
        RECT 65.860 113.275 66.150 113.320 ;
        RECT 70.930 113.460 71.220 113.505 ;
        RECT 72.790 113.460 73.080 113.505 ;
        RECT 70.930 113.320 73.080 113.460 ;
        RECT 70.930 113.275 71.220 113.320 ;
        RECT 72.790 113.275 73.080 113.320 ;
        RECT 73.710 113.460 74.000 113.505 ;
        RECT 75.510 113.460 75.830 113.520 ;
        RECT 76.970 113.460 77.260 113.505 ;
        RECT 73.710 113.320 77.260 113.460 ;
        RECT 73.710 113.275 74.000 113.320 ;
        RECT 52.525 113.120 52.815 113.165 ;
        RECT 47.420 112.980 49.955 113.120 ;
        RECT 50.300 112.980 52.815 113.120 ;
        RECT 47.420 112.935 47.710 112.980 ;
        RECT 41.930 112.780 42.250 112.840 ;
        RECT 38.800 112.640 42.250 112.780 ;
        RECT 42.480 112.780 42.620 112.935 ;
        RECT 48.830 112.780 49.150 112.840 ;
        RECT 50.300 112.780 50.440 112.980 ;
        RECT 52.525 112.935 52.815 112.980 ;
        RECT 54.825 113.120 55.115 113.165 ;
        RECT 58.950 113.120 59.270 113.180 ;
        RECT 54.825 112.980 59.270 113.120 ;
        RECT 54.825 112.935 55.115 112.980 ;
        RECT 58.950 112.920 59.270 112.980 ;
        RECT 61.680 113.120 61.970 113.165 ;
        RECT 64.000 113.120 64.215 113.275 ;
        RECT 61.680 112.980 64.215 113.120 ;
        RECT 72.865 113.120 73.080 113.275 ;
        RECT 75.510 113.260 75.830 113.320 ;
        RECT 76.970 113.275 77.260 113.320 ;
        RECT 94.850 113.460 95.140 113.505 ;
        RECT 96.710 113.460 97.000 113.505 ;
        RECT 94.850 113.320 97.000 113.460 ;
        RECT 94.850 113.275 95.140 113.320 ;
        RECT 96.710 113.275 97.000 113.320 ;
        RECT 97.630 113.460 97.920 113.505 ;
        RECT 99.890 113.460 100.210 113.520 ;
        RECT 117.830 113.505 118.150 113.520 ;
        RECT 100.890 113.460 101.180 113.505 ;
        RECT 97.630 113.320 101.180 113.460 ;
        RECT 97.630 113.275 97.920 113.320 ;
        RECT 75.110 113.120 75.400 113.165 ;
        RECT 72.865 112.980 75.400 113.120 ;
        RECT 61.680 112.935 61.970 112.980 ;
        RECT 75.110 112.935 75.400 112.980 ;
        RECT 82.870 113.120 83.190 113.180 ;
        RECT 83.345 113.120 83.635 113.165 ;
        RECT 82.870 112.980 83.635 113.120 ;
        RECT 82.870 112.920 83.190 112.980 ;
        RECT 83.345 112.935 83.635 112.980 ;
        RECT 86.565 113.120 86.855 113.165 ;
        RECT 87.470 113.120 87.790 113.180 ;
        RECT 88.865 113.120 89.155 113.165 ;
        RECT 86.565 112.980 87.790 113.120 ;
        RECT 86.565 112.935 86.855 112.980 ;
        RECT 87.470 112.920 87.790 112.980 ;
        RECT 88.480 112.980 89.155 113.120 ;
        RECT 42.480 112.640 50.440 112.780 ;
        RECT 41.930 112.580 42.250 112.640 ;
        RECT 48.830 112.580 49.150 112.640 ;
        RECT 50.670 112.580 50.990 112.840 ;
        RECT 53.445 112.595 53.735 112.825 ;
        RECT 53.890 112.780 54.210 112.840 ;
        RECT 54.365 112.780 54.655 112.825 ;
        RECT 53.890 112.640 54.655 112.780 ;
        RECT 12.050 112.440 12.340 112.485 ;
        RECT 13.910 112.440 14.200 112.485 ;
        RECT 16.690 112.440 16.980 112.485 ;
        RECT 12.050 112.300 16.980 112.440 ;
        RECT 12.050 112.255 12.340 112.300 ;
        RECT 13.910 112.255 14.200 112.300 ;
        RECT 16.690 112.255 16.980 112.300 ;
        RECT 22.170 112.440 22.460 112.485 ;
        RECT 24.030 112.440 24.320 112.485 ;
        RECT 26.810 112.440 27.100 112.485 ;
        RECT 22.170 112.300 27.100 112.440 ;
        RECT 22.170 112.255 22.460 112.300 ;
        RECT 24.030 112.255 24.320 112.300 ;
        RECT 26.810 112.255 27.100 112.300 ;
        RECT 30.675 112.440 30.965 112.485 ;
        RECT 32.270 112.440 32.590 112.500 ;
        RECT 30.675 112.300 32.590 112.440 ;
        RECT 30.675 112.255 30.965 112.300 ;
        RECT 32.270 112.240 32.590 112.300 ;
        RECT 38.710 112.440 39.030 112.500 ;
        RECT 40.565 112.440 40.855 112.485 ;
        RECT 38.710 112.300 40.855 112.440 ;
        RECT 38.710 112.240 39.030 112.300 ;
        RECT 40.565 112.255 40.855 112.300 ;
        RECT 47.420 112.440 47.710 112.485 ;
        RECT 50.200 112.440 50.490 112.485 ;
        RECT 52.060 112.440 52.350 112.485 ;
        RECT 47.420 112.300 52.350 112.440 ;
        RECT 53.520 112.440 53.660 112.595 ;
        RECT 53.890 112.580 54.210 112.640 ;
        RECT 54.365 112.595 54.655 112.640 ;
        RECT 56.650 112.780 56.970 112.840 ;
        RECT 64.945 112.780 65.235 112.825 ;
        RECT 56.650 112.640 65.235 112.780 ;
        RECT 56.650 112.580 56.970 112.640 ;
        RECT 64.945 112.595 65.235 112.640 ;
        RECT 65.390 112.780 65.710 112.840 ;
        RECT 66.785 112.780 67.075 112.825 ;
        RECT 67.690 112.780 68.010 112.840 ;
        RECT 70.005 112.780 70.295 112.825 ;
        RECT 65.390 112.640 70.295 112.780 ;
        RECT 65.390 112.580 65.710 112.640 ;
        RECT 66.785 112.595 67.075 112.640 ;
        RECT 67.690 112.580 68.010 112.640 ;
        RECT 70.005 112.595 70.295 112.640 ;
        RECT 71.830 112.580 72.150 112.840 ;
        RECT 85.645 112.595 85.935 112.825 ;
        RECT 60.790 112.440 61.110 112.500 ;
        RECT 53.520 112.300 61.110 112.440 ;
        RECT 47.420 112.255 47.710 112.300 ;
        RECT 50.200 112.255 50.490 112.300 ;
        RECT 52.060 112.255 52.350 112.300 ;
        RECT 60.790 112.240 61.110 112.300 ;
        RECT 61.680 112.440 61.970 112.485 ;
        RECT 64.460 112.440 64.750 112.485 ;
        RECT 66.320 112.440 66.610 112.485 ;
        RECT 61.680 112.300 66.610 112.440 ;
        RECT 61.680 112.255 61.970 112.300 ;
        RECT 64.460 112.255 64.750 112.300 ;
        RECT 66.320 112.255 66.610 112.300 ;
        RECT 70.470 112.440 70.760 112.485 ;
        RECT 72.330 112.440 72.620 112.485 ;
        RECT 75.110 112.440 75.400 112.485 ;
        RECT 70.470 112.300 75.400 112.440 ;
        RECT 85.720 112.440 85.860 112.595 ;
        RECT 86.550 112.440 86.870 112.500 ;
        RECT 88.480 112.485 88.620 112.980 ;
        RECT 88.865 112.935 89.155 112.980 ;
        RECT 92.530 112.920 92.850 113.180 ;
        RECT 95.765 113.120 96.055 113.165 ;
        RECT 93.540 112.980 96.055 113.120 ;
        RECT 96.785 113.120 97.000 113.275 ;
        RECT 99.890 113.260 100.210 113.320 ;
        RECT 100.890 113.275 101.180 113.320 ;
        RECT 111.870 113.460 112.160 113.505 ;
        RECT 113.730 113.460 114.020 113.505 ;
        RECT 111.870 113.320 114.020 113.460 ;
        RECT 111.870 113.275 112.160 113.320 ;
        RECT 113.730 113.275 114.020 113.320 ;
        RECT 114.650 113.460 114.940 113.505 ;
        RECT 117.830 113.460 118.200 113.505 ;
        RECT 114.650 113.320 118.200 113.460 ;
        RECT 114.650 113.275 114.940 113.320 ;
        RECT 117.830 113.275 118.200 113.320 ;
        RECT 99.030 113.120 99.320 113.165 ;
        RECT 96.785 112.980 99.320 113.120 ;
        RECT 93.540 112.485 93.680 112.980 ;
        RECT 95.765 112.935 96.055 112.980 ;
        RECT 99.030 112.935 99.320 112.980 ;
        RECT 105.410 112.920 105.730 113.180 ;
        RECT 113.805 113.120 114.020 113.275 ;
        RECT 117.830 113.260 118.150 113.275 ;
        RECT 116.050 113.120 116.340 113.165 ;
        RECT 113.805 112.980 116.340 113.120 ;
        RECT 116.050 112.935 116.340 112.980 ;
        RECT 93.925 112.780 94.215 112.825 ;
        RECT 95.290 112.780 95.610 112.840 ;
        RECT 93.925 112.640 95.610 112.780 ;
        RECT 93.925 112.595 94.215 112.640 ;
        RECT 95.290 112.580 95.610 112.640 ;
        RECT 96.670 112.780 96.990 112.840 ;
        RECT 102.895 112.780 103.185 112.825 ;
        RECT 105.885 112.780 106.175 112.825 ;
        RECT 96.670 112.640 106.175 112.780 ;
        RECT 96.670 112.580 96.990 112.640 ;
        RECT 102.895 112.595 103.185 112.640 ;
        RECT 105.885 112.595 106.175 112.640 ;
        RECT 106.345 112.595 106.635 112.825 ;
        RECT 110.010 112.780 110.330 112.840 ;
        RECT 110.945 112.780 111.235 112.825 ;
        RECT 110.010 112.640 111.235 112.780 ;
        RECT 85.720 112.300 86.870 112.440 ;
        RECT 70.470 112.255 70.760 112.300 ;
        RECT 72.330 112.255 72.620 112.300 ;
        RECT 75.110 112.255 75.400 112.300 ;
        RECT 86.550 112.240 86.870 112.300 ;
        RECT 88.405 112.255 88.695 112.485 ;
        RECT 93.465 112.255 93.755 112.485 ;
        RECT 94.390 112.440 94.680 112.485 ;
        RECT 96.250 112.440 96.540 112.485 ;
        RECT 99.030 112.440 99.320 112.485 ;
        RECT 94.390 112.300 99.320 112.440 ;
        RECT 94.390 112.255 94.680 112.300 ;
        RECT 96.250 112.255 96.540 112.300 ;
        RECT 99.030 112.255 99.320 112.300 ;
        RECT 103.570 112.440 103.890 112.500 ;
        RECT 106.420 112.440 106.560 112.595 ;
        RECT 110.010 112.580 110.330 112.640 ;
        RECT 110.945 112.595 111.235 112.640 ;
        RECT 112.770 112.580 113.090 112.840 ;
        RECT 103.570 112.300 106.560 112.440 ;
        RECT 111.410 112.440 111.700 112.485 ;
        RECT 113.270 112.440 113.560 112.485 ;
        RECT 116.050 112.440 116.340 112.485 ;
        RECT 111.410 112.300 116.340 112.440 ;
        RECT 103.570 112.240 103.890 112.300 ;
        RECT 111.410 112.255 111.700 112.300 ;
        RECT 113.270 112.255 113.560 112.300 ;
        RECT 116.050 112.255 116.340 112.300 ;
        RECT 20.555 112.100 20.845 112.145 ;
        RECT 21.690 112.100 22.010 112.160 ;
        RECT 20.555 111.960 22.010 112.100 ;
        RECT 20.555 111.915 20.845 111.960 ;
        RECT 21.690 111.900 22.010 111.960 ;
        RECT 31.810 111.900 32.130 112.160 ;
        RECT 35.950 111.900 36.270 112.160 ;
        RECT 39.170 112.100 39.490 112.160 ;
        RECT 39.645 112.100 39.935 112.145 ;
        RECT 39.170 111.960 39.935 112.100 ;
        RECT 39.170 111.900 39.490 111.960 ;
        RECT 39.645 111.915 39.935 111.960 ;
        RECT 41.010 112.100 41.330 112.160 ;
        RECT 48.370 112.100 48.690 112.160 ;
        RECT 41.010 111.960 48.690 112.100 ;
        RECT 41.010 111.900 41.330 111.960 ;
        RECT 48.370 111.900 48.690 111.960 ;
        RECT 56.650 111.900 56.970 112.160 ;
        RECT 57.815 112.100 58.105 112.145 ;
        RECT 59.410 112.100 59.730 112.160 ;
        RECT 57.815 111.960 59.730 112.100 ;
        RECT 57.815 111.915 58.105 111.960 ;
        RECT 59.410 111.900 59.730 111.960 ;
        RECT 76.890 112.100 77.210 112.160 ;
        RECT 78.975 112.100 79.265 112.145 ;
        RECT 76.890 111.960 79.265 112.100 ;
        RECT 76.890 111.900 77.210 111.960 ;
        RECT 78.975 111.915 79.265 111.960 ;
        RECT 83.790 111.900 84.110 112.160 ;
        RECT 117.370 112.100 117.690 112.160 ;
        RECT 119.915 112.100 120.205 112.145 ;
        RECT 117.370 111.960 120.205 112.100 ;
        RECT 117.370 111.900 117.690 111.960 ;
        RECT 119.915 111.915 120.205 111.960 ;
        RECT 5.520 111.280 125.580 111.760 ;
        RECT 16.170 111.080 16.490 111.140 ;
        RECT 18.945 111.080 19.235 111.125 ;
        RECT 16.170 110.940 19.235 111.080 ;
        RECT 16.170 110.880 16.490 110.940 ;
        RECT 18.945 110.895 19.235 110.940 ;
        RECT 23.530 110.880 23.850 111.140 ;
        RECT 47.005 111.080 47.295 111.125 ;
        RECT 48.830 111.080 49.150 111.140 ;
        RECT 47.005 110.940 49.150 111.080 ;
        RECT 47.005 110.895 47.295 110.940 ;
        RECT 32.270 110.740 32.590 110.800 ;
        RECT 22.240 110.600 32.590 110.740 ;
        RECT 16.645 110.400 16.935 110.445 ;
        RECT 17.090 110.400 17.410 110.460 ;
        RECT 16.645 110.260 17.410 110.400 ;
        RECT 16.645 110.215 16.935 110.260 ;
        RECT 17.090 110.200 17.410 110.260 ;
        RECT 20.770 110.400 21.090 110.460 ;
        RECT 21.705 110.400 21.995 110.445 ;
        RECT 20.770 110.260 21.995 110.400 ;
        RECT 20.770 110.200 21.090 110.260 ;
        RECT 21.705 110.215 21.995 110.260 ;
        RECT 16.170 109.860 16.490 110.120 ;
        RECT 21.245 110.060 21.535 110.105 ;
        RECT 22.240 110.060 22.380 110.600 ;
        RECT 32.270 110.540 32.590 110.600 ;
        RECT 34.590 110.740 34.880 110.785 ;
        RECT 36.450 110.740 36.740 110.785 ;
        RECT 39.230 110.740 39.520 110.785 ;
        RECT 34.590 110.600 39.520 110.740 ;
        RECT 34.590 110.555 34.880 110.600 ;
        RECT 36.450 110.555 36.740 110.600 ;
        RECT 39.230 110.555 39.520 110.600 ;
        RECT 47.080 110.460 47.220 110.895 ;
        RECT 48.830 110.880 49.150 110.940 ;
        RECT 69.545 111.080 69.835 111.125 ;
        RECT 71.830 111.080 72.150 111.140 ;
        RECT 69.545 110.940 72.150 111.080 ;
        RECT 69.545 110.895 69.835 110.940 ;
        RECT 71.830 110.880 72.150 110.940 ;
        RECT 92.530 111.080 92.850 111.140 ;
        RECT 96.225 111.080 96.515 111.125 ;
        RECT 92.530 110.940 96.515 111.080 ;
        RECT 92.530 110.880 92.850 110.940 ;
        RECT 96.225 110.895 96.515 110.940 ;
        RECT 119.210 110.880 119.530 111.140 ;
        RECT 54.830 110.740 55.120 110.785 ;
        RECT 56.690 110.740 56.980 110.785 ;
        RECT 59.470 110.740 59.760 110.785 ;
        RECT 54.830 110.600 59.760 110.740 ;
        RECT 54.830 110.555 55.120 110.600 ;
        RECT 56.690 110.555 56.980 110.600 ;
        RECT 59.470 110.555 59.760 110.600 ;
        RECT 70.930 110.740 71.220 110.785 ;
        RECT 72.790 110.740 73.080 110.785 ;
        RECT 75.570 110.740 75.860 110.785 ;
        RECT 70.930 110.600 75.860 110.740 ;
        RECT 70.930 110.555 71.220 110.600 ;
        RECT 72.790 110.555 73.080 110.600 ;
        RECT 75.570 110.555 75.860 110.600 ;
        RECT 80.590 110.740 80.880 110.785 ;
        RECT 82.450 110.740 82.740 110.785 ;
        RECT 85.230 110.740 85.520 110.785 ;
        RECT 80.590 110.600 85.520 110.740 ;
        RECT 80.590 110.555 80.880 110.600 ;
        RECT 82.450 110.555 82.740 110.600 ;
        RECT 85.230 110.555 85.520 110.600 ;
        RECT 87.470 110.740 87.790 110.800 ;
        RECT 89.095 110.740 89.385 110.785 ;
        RECT 87.470 110.600 89.385 110.740 ;
        RECT 87.470 110.540 87.790 110.600 ;
        RECT 89.095 110.555 89.385 110.600 ;
        RECT 104.510 110.740 104.800 110.785 ;
        RECT 106.370 110.740 106.660 110.785 ;
        RECT 109.150 110.740 109.440 110.785 ;
        RECT 104.510 110.600 109.440 110.740 ;
        RECT 104.510 110.555 104.800 110.600 ;
        RECT 106.370 110.555 106.660 110.600 ;
        RECT 109.150 110.555 109.440 110.600 ;
        RECT 34.125 110.400 34.415 110.445 ;
        RECT 46.990 110.400 47.310 110.460 ;
        RECT 54.365 110.400 54.655 110.445 ;
        RECT 34.125 110.260 54.655 110.400 ;
        RECT 34.125 110.215 34.415 110.260 ;
        RECT 46.990 110.200 47.310 110.260 ;
        RECT 54.365 110.215 54.655 110.260 ;
        RECT 56.205 110.400 56.495 110.445 ;
        RECT 57.110 110.400 57.430 110.460 ;
        RECT 56.205 110.260 57.430 110.400 ;
        RECT 56.205 110.215 56.495 110.260 ;
        RECT 57.110 110.200 57.430 110.260 ;
        RECT 61.710 110.400 62.030 110.460 ;
        RECT 65.390 110.400 65.710 110.460 ;
        RECT 70.465 110.400 70.755 110.445 ;
        RECT 80.125 110.400 80.415 110.445 ;
        RECT 87.010 110.400 87.330 110.460 ;
        RECT 98.510 110.400 98.830 110.460 ;
        RECT 98.985 110.400 99.275 110.445 ;
        RECT 103.110 110.400 103.430 110.460 ;
        RECT 61.710 110.260 65.160 110.400 ;
        RECT 61.710 110.200 62.030 110.260 ;
        RECT 21.245 109.920 22.380 110.060 ;
        RECT 24.465 110.060 24.755 110.105 ;
        RECT 31.810 110.060 32.130 110.120 ;
        RECT 24.465 109.920 32.130 110.060 ;
        RECT 21.245 109.875 21.535 109.920 ;
        RECT 24.465 109.875 24.755 109.920 ;
        RECT 31.810 109.860 32.130 109.920 ;
        RECT 35.950 109.860 36.270 110.120 ;
        RECT 65.020 110.105 65.160 110.260 ;
        RECT 65.390 110.260 90.000 110.400 ;
        RECT 65.390 110.200 65.710 110.260 ;
        RECT 70.465 110.215 70.755 110.260 ;
        RECT 80.125 110.215 80.415 110.260 ;
        RECT 87.010 110.200 87.330 110.260 ;
        RECT 39.230 110.060 39.520 110.105 ;
        RECT 59.470 110.060 59.760 110.105 ;
        RECT 36.985 109.920 39.520 110.060 ;
        RECT 33.650 109.520 33.970 109.780 ;
        RECT 36.985 109.765 37.200 109.920 ;
        RECT 39.230 109.875 39.520 109.920 ;
        RECT 57.225 109.920 59.760 110.060 ;
        RECT 35.050 109.720 35.340 109.765 ;
        RECT 36.910 109.720 37.200 109.765 ;
        RECT 35.050 109.580 37.200 109.720 ;
        RECT 35.050 109.535 35.340 109.580 ;
        RECT 36.910 109.535 37.200 109.580 ;
        RECT 37.830 109.720 38.120 109.765 ;
        RECT 38.710 109.720 39.030 109.780 ;
        RECT 41.090 109.720 41.380 109.765 ;
        RECT 37.830 109.580 41.380 109.720 ;
        RECT 37.830 109.535 38.120 109.580 ;
        RECT 38.710 109.520 39.030 109.580 ;
        RECT 41.090 109.535 41.380 109.580 ;
        RECT 53.430 109.520 53.750 109.780 ;
        RECT 57.225 109.765 57.440 109.920 ;
        RECT 59.470 109.875 59.760 109.920 ;
        RECT 64.945 110.060 65.235 110.105 ;
        RECT 66.310 110.060 66.630 110.120 ;
        RECT 64.945 109.920 66.630 110.060 ;
        RECT 64.945 109.875 65.235 109.920 ;
        RECT 66.310 109.860 66.630 109.920 ;
        RECT 68.610 109.860 68.930 110.120 ;
        RECT 70.910 110.060 71.230 110.120 ;
        RECT 72.305 110.060 72.595 110.105 ;
        RECT 75.570 110.060 75.860 110.105 ;
        RECT 70.910 109.920 72.595 110.060 ;
        RECT 70.910 109.860 71.230 109.920 ;
        RECT 72.305 109.875 72.595 109.920 ;
        RECT 73.325 109.920 75.860 110.060 ;
        RECT 73.325 109.765 73.540 109.920 ;
        RECT 75.570 109.875 75.860 109.920 ;
        RECT 80.570 110.060 80.890 110.120 ;
        RECT 89.860 110.105 90.000 110.260 ;
        RECT 98.510 110.260 103.430 110.400 ;
        RECT 98.510 110.200 98.830 110.260 ;
        RECT 98.985 110.215 99.275 110.260 ;
        RECT 103.110 110.200 103.430 110.260 ;
        RECT 104.045 110.400 104.335 110.445 ;
        RECT 110.010 110.400 110.330 110.460 ;
        RECT 104.045 110.260 110.330 110.400 ;
        RECT 104.045 110.215 104.335 110.260 ;
        RECT 110.010 110.200 110.330 110.260 ;
        RECT 114.150 110.400 114.470 110.460 ;
        RECT 116.465 110.400 116.755 110.445 ;
        RECT 114.150 110.260 116.755 110.400 ;
        RECT 114.150 110.200 114.470 110.260 ;
        RECT 116.465 110.215 116.755 110.260 ;
        RECT 117.830 110.400 118.150 110.460 ;
        RECT 118.305 110.400 118.595 110.445 ;
        RECT 117.830 110.260 118.595 110.400 ;
        RECT 117.830 110.200 118.150 110.260 ;
        RECT 118.305 110.215 118.595 110.260 ;
        RECT 122.430 110.200 122.750 110.460 ;
        RECT 81.965 110.060 82.255 110.105 ;
        RECT 85.230 110.060 85.520 110.105 ;
        RECT 80.570 109.920 82.255 110.060 ;
        RECT 80.570 109.860 80.890 109.920 ;
        RECT 81.965 109.875 82.255 109.920 ;
        RECT 82.985 109.920 85.520 110.060 ;
        RECT 55.290 109.720 55.580 109.765 ;
        RECT 57.150 109.720 57.440 109.765 ;
        RECT 55.290 109.580 57.440 109.720 ;
        RECT 55.290 109.535 55.580 109.580 ;
        RECT 57.150 109.535 57.440 109.580 ;
        RECT 58.070 109.720 58.360 109.765 ;
        RECT 61.330 109.720 61.620 109.765 ;
        RECT 64.485 109.720 64.775 109.765 ;
        RECT 58.070 109.580 64.775 109.720 ;
        RECT 58.070 109.535 58.360 109.580 ;
        RECT 61.330 109.535 61.620 109.580 ;
        RECT 64.485 109.535 64.775 109.580 ;
        RECT 71.390 109.720 71.680 109.765 ;
        RECT 73.250 109.720 73.540 109.765 ;
        RECT 71.390 109.580 73.540 109.720 ;
        RECT 71.390 109.535 71.680 109.580 ;
        RECT 73.250 109.535 73.540 109.580 ;
        RECT 74.130 109.765 74.450 109.780 ;
        RECT 82.985 109.765 83.200 109.920 ;
        RECT 85.230 109.875 85.520 109.920 ;
        RECT 89.785 109.875 90.075 110.105 ;
        RECT 105.870 109.860 106.190 110.120 ;
        RECT 109.150 110.060 109.440 110.105 ;
        RECT 113.015 110.060 113.305 110.105 ;
        RECT 116.005 110.060 116.295 110.105 ;
        RECT 106.905 109.920 109.440 110.060 ;
        RECT 74.130 109.720 74.460 109.765 ;
        RECT 77.430 109.720 77.720 109.765 ;
        RECT 74.130 109.580 77.720 109.720 ;
        RECT 74.130 109.535 74.460 109.580 ;
        RECT 77.430 109.535 77.720 109.580 ;
        RECT 81.050 109.720 81.340 109.765 ;
        RECT 82.910 109.720 83.200 109.765 ;
        RECT 81.050 109.580 83.200 109.720 ;
        RECT 81.050 109.535 81.340 109.580 ;
        RECT 82.910 109.535 83.200 109.580 ;
        RECT 83.790 109.765 84.110 109.780 ;
        RECT 106.905 109.765 107.120 109.920 ;
        RECT 109.150 109.875 109.440 109.920 ;
        RECT 111.480 110.030 113.305 110.060 ;
        RECT 113.780 110.030 116.295 110.060 ;
        RECT 111.480 109.920 116.295 110.030 ;
        RECT 83.790 109.720 84.120 109.765 ;
        RECT 87.090 109.720 87.380 109.765 ;
        RECT 83.790 109.580 87.380 109.720 ;
        RECT 83.790 109.535 84.120 109.580 ;
        RECT 87.090 109.535 87.380 109.580 ;
        RECT 104.970 109.720 105.260 109.765 ;
        RECT 106.830 109.720 107.120 109.765 ;
        RECT 104.970 109.580 107.120 109.720 ;
        RECT 104.970 109.535 105.260 109.580 ;
        RECT 106.830 109.535 107.120 109.580 ;
        RECT 107.750 109.720 108.040 109.765 ;
        RECT 109.550 109.720 109.870 109.780 ;
        RECT 111.010 109.720 111.300 109.765 ;
        RECT 107.750 109.580 111.300 109.720 ;
        RECT 107.750 109.535 108.040 109.580 ;
        RECT 74.130 109.520 74.450 109.535 ;
        RECT 83.790 109.520 84.110 109.535 ;
        RECT 109.550 109.520 109.870 109.580 ;
        RECT 111.010 109.535 111.300 109.580 ;
        RECT 20.785 109.380 21.075 109.425 ;
        RECT 21.690 109.380 22.010 109.440 ;
        RECT 20.785 109.240 22.010 109.380 ;
        RECT 20.785 109.195 21.075 109.240 ;
        RECT 21.690 109.180 22.010 109.240 ;
        RECT 27.225 109.380 27.515 109.425 ;
        RECT 27.670 109.380 27.990 109.440 ;
        RECT 27.225 109.240 27.990 109.380 ;
        RECT 27.225 109.195 27.515 109.240 ;
        RECT 27.670 109.180 27.990 109.240 ;
        RECT 36.410 109.380 36.730 109.440 ;
        RECT 43.095 109.380 43.385 109.425 ;
        RECT 36.410 109.240 43.385 109.380 ;
        RECT 36.410 109.180 36.730 109.240 ;
        RECT 43.095 109.195 43.385 109.240 ;
        RECT 58.950 109.380 59.270 109.440 ;
        RECT 63.335 109.380 63.625 109.425 ;
        RECT 58.950 109.240 63.625 109.380 ;
        RECT 58.950 109.180 59.270 109.240 ;
        RECT 63.335 109.195 63.625 109.240 ;
        RECT 75.970 109.380 76.290 109.440 ;
        RECT 79.435 109.380 79.725 109.425 ;
        RECT 75.970 109.240 79.725 109.380 ;
        RECT 75.970 109.180 76.290 109.240 ;
        RECT 79.435 109.195 79.725 109.240 ;
        RECT 96.670 109.380 96.990 109.440 ;
        RECT 98.065 109.380 98.355 109.425 ;
        RECT 96.670 109.240 98.355 109.380 ;
        RECT 96.670 109.180 96.990 109.240 ;
        RECT 98.065 109.195 98.355 109.240 ;
        RECT 98.525 109.380 98.815 109.425 ;
        RECT 98.970 109.380 99.290 109.440 ;
        RECT 98.525 109.240 99.290 109.380 ;
        RECT 98.525 109.195 98.815 109.240 ;
        RECT 98.970 109.180 99.290 109.240 ;
        RECT 105.410 109.380 105.730 109.440 ;
        RECT 111.480 109.380 111.620 109.920 ;
        RECT 112.860 109.890 113.920 109.920 ;
        RECT 113.015 109.875 113.305 109.890 ;
        RECT 116.005 109.875 116.295 109.920 ;
        RECT 118.750 109.860 119.070 110.120 ;
        RECT 119.210 110.060 119.530 110.120 ;
        RECT 120.145 110.060 120.435 110.105 ;
        RECT 119.210 109.920 120.435 110.060 ;
        RECT 119.210 109.860 119.530 109.920 ;
        RECT 120.145 109.875 120.435 109.920 ;
        RECT 121.985 109.875 122.275 110.105 ;
        RECT 118.840 109.720 118.980 109.860 ;
        RECT 122.060 109.720 122.200 109.875 ;
        RECT 118.840 109.580 122.200 109.720 ;
        RECT 105.410 109.240 111.620 109.380 ;
        RECT 105.410 109.180 105.730 109.240 ;
        RECT 113.690 109.180 114.010 109.440 ;
        RECT 115.545 109.380 115.835 109.425 ;
        RECT 116.910 109.380 117.230 109.440 ;
        RECT 115.545 109.240 117.230 109.380 ;
        RECT 115.545 109.195 115.835 109.240 ;
        RECT 116.910 109.180 117.230 109.240 ;
        RECT 5.520 108.560 125.580 109.040 ;
        RECT 27.210 108.360 27.530 108.420 ;
        RECT 28.605 108.360 28.895 108.405 ;
        RECT 27.210 108.220 28.895 108.360 ;
        RECT 27.210 108.160 27.530 108.220 ;
        RECT 28.605 108.175 28.895 108.220 ;
        RECT 36.870 108.360 37.190 108.420 ;
        RECT 37.345 108.360 37.635 108.405 ;
        RECT 36.870 108.220 37.635 108.360 ;
        RECT 36.870 108.160 37.190 108.220 ;
        RECT 37.345 108.175 37.635 108.220 ;
        RECT 50.225 108.360 50.515 108.405 ;
        RECT 50.670 108.360 50.990 108.420 ;
        RECT 50.225 108.220 50.990 108.360 ;
        RECT 50.225 108.175 50.515 108.220 ;
        RECT 50.670 108.160 50.990 108.220 ;
        RECT 55.285 108.360 55.575 108.405 ;
        RECT 57.110 108.360 57.430 108.420 ;
        RECT 55.285 108.220 57.430 108.360 ;
        RECT 55.285 108.175 55.575 108.220 ;
        RECT 57.110 108.160 57.430 108.220 ;
        RECT 57.570 108.160 57.890 108.420 ;
        RECT 59.410 108.160 59.730 108.420 ;
        RECT 70.465 108.360 70.755 108.405 ;
        RECT 70.910 108.360 71.230 108.420 ;
        RECT 70.465 108.220 71.230 108.360 ;
        RECT 70.465 108.175 70.755 108.220 ;
        RECT 70.910 108.160 71.230 108.220 ;
        RECT 72.305 108.360 72.595 108.405 ;
        RECT 74.130 108.360 74.450 108.420 ;
        RECT 72.305 108.220 74.450 108.360 ;
        RECT 72.305 108.175 72.595 108.220 ;
        RECT 74.130 108.160 74.450 108.220 ;
        RECT 75.510 108.360 75.830 108.420 ;
        RECT 78.745 108.360 79.035 108.405 ;
        RECT 75.510 108.220 79.035 108.360 ;
        RECT 75.510 108.160 75.830 108.220 ;
        RECT 78.745 108.175 79.035 108.220 ;
        RECT 80.570 108.160 80.890 108.420 ;
        RECT 109.550 108.160 109.870 108.420 ;
        RECT 111.865 108.360 112.155 108.405 ;
        RECT 112.770 108.360 113.090 108.420 ;
        RECT 111.865 108.220 113.090 108.360 ;
        RECT 111.865 108.175 112.155 108.220 ;
        RECT 112.770 108.160 113.090 108.220 ;
        RECT 119.210 108.160 119.530 108.420 ;
        RECT 39.190 108.020 39.480 108.065 ;
        RECT 41.050 108.020 41.340 108.065 ;
        RECT 16.260 107.880 29.280 108.020 ;
        RECT 16.260 107.740 16.400 107.880 ;
        RECT 29.140 107.740 29.280 107.880 ;
        RECT 39.190 107.880 41.340 108.020 ;
        RECT 39.190 107.835 39.480 107.880 ;
        RECT 41.050 107.835 41.340 107.880 ;
        RECT 41.970 108.020 42.260 108.065 ;
        RECT 45.230 108.020 45.520 108.065 ;
        RECT 48.385 108.020 48.675 108.065 ;
        RECT 52.985 108.020 53.275 108.065 ;
        RECT 59.500 108.020 59.640 108.160 ;
        RECT 41.970 107.880 48.675 108.020 ;
        RECT 41.970 107.835 42.260 107.880 ;
        RECT 45.230 107.835 45.520 107.880 ;
        RECT 48.385 107.835 48.675 107.880 ;
        RECT 48.920 107.880 52.280 108.020 ;
        RECT 12.950 107.480 13.270 107.740 ;
        RECT 14.345 107.495 14.635 107.725 ;
        RECT 14.420 107.340 14.560 107.495 ;
        RECT 16.170 107.480 16.490 107.740 ;
        RECT 18.470 107.480 18.790 107.740 ;
        RECT 18.945 107.680 19.235 107.725 ;
        RECT 20.770 107.680 21.090 107.740 ;
        RECT 18.945 107.540 21.090 107.680 ;
        RECT 18.945 107.495 19.235 107.540 ;
        RECT 20.770 107.480 21.090 107.540 ;
        RECT 23.530 107.480 23.850 107.740 ;
        RECT 25.385 107.680 25.675 107.725 ;
        RECT 27.670 107.680 27.990 107.740 ;
        RECT 25.385 107.540 27.990 107.680 ;
        RECT 25.385 107.495 25.675 107.540 ;
        RECT 27.670 107.480 27.990 107.540 ;
        RECT 29.050 107.680 29.370 107.740 ;
        RECT 29.525 107.680 29.815 107.725 ;
        RECT 29.050 107.540 29.815 107.680 ;
        RECT 29.050 107.480 29.370 107.540 ;
        RECT 29.525 107.495 29.815 107.540 ;
        RECT 29.970 107.680 30.290 107.740 ;
        RECT 35.045 107.680 35.335 107.725 ;
        RECT 29.970 107.540 35.335 107.680 ;
        RECT 29.970 107.480 30.290 107.540 ;
        RECT 35.045 107.495 35.335 107.540 ;
        RECT 35.505 107.680 35.795 107.725 ;
        RECT 36.410 107.680 36.730 107.740 ;
        RECT 35.505 107.540 36.730 107.680 ;
        RECT 35.505 107.495 35.795 107.540 ;
        RECT 36.410 107.480 36.730 107.540 ;
        RECT 38.265 107.680 38.555 107.725 ;
        RECT 41.125 107.680 41.340 107.835 ;
        RECT 48.920 107.740 49.060 107.880 ;
        RECT 43.370 107.680 43.660 107.725 ;
        RECT 38.265 107.540 40.780 107.680 ;
        RECT 41.125 107.540 43.660 107.680 ;
        RECT 38.265 107.495 38.555 107.540 ;
        RECT 19.865 107.340 20.155 107.385 ;
        RECT 21.230 107.340 21.550 107.400 ;
        RECT 14.420 107.200 16.860 107.340 ;
        RECT 16.720 107.045 16.860 107.200 ;
        RECT 19.865 107.200 21.550 107.340 ;
        RECT 19.865 107.155 20.155 107.200 ;
        RECT 21.230 107.140 21.550 107.200 ;
        RECT 34.570 107.140 34.890 107.400 ;
        RECT 39.170 107.340 39.490 107.400 ;
        RECT 40.105 107.340 40.395 107.385 ;
        RECT 39.170 107.200 40.395 107.340 ;
        RECT 40.640 107.340 40.780 107.540 ;
        RECT 43.370 107.495 43.660 107.540 ;
        RECT 48.830 107.480 49.150 107.740 ;
        RECT 49.305 107.680 49.595 107.725 ;
        RECT 49.305 107.540 50.900 107.680 ;
        RECT 49.305 107.495 49.595 107.540 ;
        RECT 44.690 107.340 45.010 107.400 ;
        RECT 46.990 107.340 47.310 107.400 ;
        RECT 40.640 107.200 47.310 107.340 ;
        RECT 39.170 107.140 39.490 107.200 ;
        RECT 40.105 107.155 40.395 107.200 ;
        RECT 44.690 107.140 45.010 107.200 ;
        RECT 46.990 107.140 47.310 107.200 ;
        RECT 50.760 107.045 50.900 107.540 ;
        RECT 16.645 106.815 16.935 107.045 ;
        RECT 38.730 107.000 39.020 107.045 ;
        RECT 40.590 107.000 40.880 107.045 ;
        RECT 43.370 107.000 43.660 107.045 ;
        RECT 38.730 106.860 43.660 107.000 ;
        RECT 38.730 106.815 39.020 106.860 ;
        RECT 40.590 106.815 40.880 106.860 ;
        RECT 43.370 106.815 43.660 106.860 ;
        RECT 50.685 106.815 50.975 107.045 ;
        RECT 52.140 107.000 52.280 107.880 ;
        RECT 52.985 107.880 59.640 108.020 ;
        RECT 52.985 107.835 53.275 107.880 ;
        RECT 75.970 107.820 76.290 108.080 ;
        RECT 76.445 108.020 76.735 108.065 ;
        RECT 76.890 108.020 77.210 108.080 ;
        RECT 82.870 108.020 83.190 108.080 ;
        RECT 76.445 107.880 77.210 108.020 ;
        RECT 76.445 107.835 76.735 107.880 ;
        RECT 76.890 107.820 77.210 107.880 ;
        RECT 79.280 107.880 83.190 108.020 ;
        RECT 52.510 107.480 52.830 107.740 ;
        RECT 56.205 107.680 56.495 107.725 ;
        RECT 56.650 107.680 56.970 107.740 ;
        RECT 69.070 107.680 69.390 107.740 ;
        RECT 69.545 107.680 69.835 107.725 ;
        RECT 56.205 107.540 56.970 107.680 ;
        RECT 56.205 107.495 56.495 107.540 ;
        RECT 56.650 107.480 56.970 107.540 ;
        RECT 57.200 107.540 61.020 107.680 ;
        RECT 53.905 107.340 54.195 107.385 ;
        RECT 55.270 107.340 55.590 107.400 ;
        RECT 57.200 107.340 57.340 107.540 ;
        RECT 60.880 107.400 61.020 107.540 ;
        RECT 69.070 107.540 69.835 107.680 ;
        RECT 69.070 107.480 69.390 107.540 ;
        RECT 69.545 107.495 69.835 107.540 ;
        RECT 71.830 107.680 72.150 107.740 ;
        RECT 79.280 107.725 79.420 107.880 ;
        RECT 82.870 107.820 83.190 107.880 ;
        RECT 96.690 108.020 96.980 108.065 ;
        RECT 98.550 108.020 98.840 108.065 ;
        RECT 96.690 107.880 98.840 108.020 ;
        RECT 96.690 107.835 96.980 107.880 ;
        RECT 98.550 107.835 98.840 107.880 ;
        RECT 99.470 108.020 99.760 108.065 ;
        RECT 102.730 108.020 103.020 108.065 ;
        RECT 105.885 108.020 106.175 108.065 ;
        RECT 99.470 107.880 106.175 108.020 ;
        RECT 99.470 107.835 99.760 107.880 ;
        RECT 102.730 107.835 103.020 107.880 ;
        RECT 105.885 107.835 106.175 107.880 ;
        RECT 79.205 107.680 79.495 107.725 ;
        RECT 71.830 107.540 79.495 107.680 ;
        RECT 71.830 107.480 72.150 107.540 ;
        RECT 79.205 107.495 79.495 107.540 ;
        RECT 79.650 107.480 79.970 107.740 ;
        RECT 83.330 107.480 83.650 107.740 ;
        RECT 98.625 107.680 98.840 107.835 ;
        RECT 100.870 107.680 101.160 107.725 ;
        RECT 98.625 107.540 101.160 107.680 ;
        RECT 100.870 107.495 101.160 107.540 ;
        RECT 101.730 107.680 102.050 107.740 ;
        RECT 106.345 107.680 106.635 107.725 ;
        RECT 110.025 107.680 110.315 107.725 ;
        RECT 101.730 107.540 110.315 107.680 ;
        RECT 101.730 107.480 102.050 107.540 ;
        RECT 106.345 107.495 106.635 107.540 ;
        RECT 110.025 107.495 110.315 107.540 ;
        RECT 112.785 107.680 113.075 107.725 ;
        RECT 113.690 107.680 114.010 107.740 ;
        RECT 112.785 107.540 114.010 107.680 ;
        RECT 112.785 107.495 113.075 107.540 ;
        RECT 113.690 107.480 114.010 107.540 ;
        RECT 114.150 107.680 114.470 107.740 ;
        RECT 117.385 107.680 117.675 107.725 ;
        RECT 118.290 107.680 118.610 107.740 ;
        RECT 114.150 107.540 118.610 107.680 ;
        RECT 114.150 107.480 114.470 107.540 ;
        RECT 117.385 107.495 117.675 107.540 ;
        RECT 118.290 107.480 118.610 107.540 ;
        RECT 53.905 107.200 57.340 107.340 ;
        RECT 58.950 107.340 59.270 107.400 ;
        RECT 59.870 107.340 60.190 107.400 ;
        RECT 58.950 107.200 60.190 107.340 ;
        RECT 53.905 107.155 54.195 107.200 ;
        RECT 55.270 107.140 55.590 107.200 ;
        RECT 58.950 107.140 59.270 107.200 ;
        RECT 59.870 107.140 60.190 107.200 ;
        RECT 60.790 107.140 61.110 107.400 ;
        RECT 74.590 107.340 74.910 107.400 ;
        RECT 77.365 107.340 77.655 107.385 ;
        RECT 86.550 107.340 86.870 107.400 ;
        RECT 74.590 107.200 86.870 107.340 ;
        RECT 74.590 107.140 74.910 107.200 ;
        RECT 77.365 107.155 77.655 107.200 ;
        RECT 86.550 107.140 86.870 107.200 ;
        RECT 95.750 107.140 96.070 107.400 ;
        RECT 97.130 107.340 97.450 107.400 ;
        RECT 97.605 107.340 97.895 107.385 ;
        RECT 97.130 107.200 97.895 107.340 ;
        RECT 97.130 107.140 97.450 107.200 ;
        RECT 97.605 107.155 97.895 107.200 ;
        RECT 114.610 107.340 114.930 107.400 ;
        RECT 116.005 107.340 116.295 107.385 ;
        RECT 114.610 107.200 116.295 107.340 ;
        RECT 114.610 107.140 114.930 107.200 ;
        RECT 116.005 107.155 116.295 107.200 ;
        RECT 116.910 107.140 117.230 107.400 ;
        RECT 61.710 107.000 62.030 107.060 ;
        RECT 52.140 106.860 62.030 107.000 ;
        RECT 61.710 106.800 62.030 106.860 ;
        RECT 68.610 107.000 68.930 107.060 ;
        RECT 74.145 107.000 74.435 107.045 ;
        RECT 68.610 106.860 74.435 107.000 ;
        RECT 68.610 106.800 68.930 106.860 ;
        RECT 74.145 106.815 74.435 106.860 ;
        RECT 96.230 107.000 96.520 107.045 ;
        RECT 98.090 107.000 98.380 107.045 ;
        RECT 100.870 107.000 101.160 107.045 ;
        RECT 96.230 106.860 101.160 107.000 ;
        RECT 96.230 106.815 96.520 106.860 ;
        RECT 98.090 106.815 98.380 106.860 ;
        RECT 100.870 106.815 101.160 106.860 ;
        RECT 8.810 106.660 9.130 106.720 ;
        RECT 12.045 106.660 12.335 106.705 ;
        RECT 8.810 106.520 12.335 106.660 ;
        RECT 8.810 106.460 9.130 106.520 ;
        RECT 12.045 106.475 12.335 106.520 ;
        RECT 12.490 106.660 12.810 106.720 ;
        RECT 13.425 106.660 13.715 106.705 ;
        RECT 12.490 106.520 13.715 106.660 ;
        RECT 12.490 106.460 12.810 106.520 ;
        RECT 13.425 106.475 13.715 106.520 ;
        RECT 15.710 106.460 16.030 106.720 ;
        RECT 24.465 106.660 24.755 106.705 ;
        RECT 26.750 106.660 27.070 106.720 ;
        RECT 24.465 106.520 27.070 106.660 ;
        RECT 24.465 106.475 24.755 106.520 ;
        RECT 26.750 106.460 27.070 106.520 ;
        RECT 29.510 106.660 29.830 106.720 ;
        RECT 29.985 106.660 30.275 106.705 ;
        RECT 29.510 106.520 30.275 106.660 ;
        RECT 29.510 106.460 29.830 106.520 ;
        RECT 29.985 106.475 30.275 106.520 ;
        RECT 47.235 106.660 47.525 106.705 ;
        RECT 48.370 106.660 48.690 106.720 ;
        RECT 53.890 106.660 54.210 106.720 ;
        RECT 47.235 106.520 54.210 106.660 ;
        RECT 47.235 106.475 47.525 106.520 ;
        RECT 48.370 106.460 48.690 106.520 ;
        RECT 53.890 106.460 54.210 106.520 ;
        RECT 87.010 106.660 87.330 106.720 ;
        RECT 89.785 106.660 90.075 106.705 ;
        RECT 87.010 106.520 90.075 106.660 ;
        RECT 87.010 106.460 87.330 106.520 ;
        RECT 89.785 106.475 90.075 106.520 ;
        RECT 98.970 106.660 99.290 106.720 ;
        RECT 104.735 106.660 105.025 106.705 ;
        RECT 98.970 106.520 105.025 106.660 ;
        RECT 98.970 106.460 99.290 106.520 ;
        RECT 104.735 106.475 105.025 106.520 ;
        RECT 5.520 105.840 125.580 106.320 ;
        RECT 12.950 105.640 13.270 105.700 ;
        RECT 18.945 105.640 19.235 105.685 ;
        RECT 12.950 105.500 19.235 105.640 ;
        RECT 12.950 105.440 13.270 105.500 ;
        RECT 18.945 105.455 19.235 105.500 ;
        RECT 21.230 105.640 21.550 105.700 ;
        RECT 23.990 105.640 24.310 105.700 ;
        RECT 41.930 105.640 42.250 105.700 ;
        RECT 44.705 105.640 44.995 105.685 ;
        RECT 21.230 105.500 34.800 105.640 ;
        RECT 21.230 105.440 21.550 105.500 ;
        RECT 8.830 105.300 9.120 105.345 ;
        RECT 10.690 105.300 10.980 105.345 ;
        RECT 13.470 105.300 13.760 105.345 ;
        RECT 8.830 105.160 13.760 105.300 ;
        RECT 8.830 105.115 9.120 105.160 ;
        RECT 10.690 105.115 10.980 105.160 ;
        RECT 13.470 105.115 13.760 105.160 ;
        RECT 8.365 104.960 8.655 105.005 ;
        RECT 11.570 104.960 11.890 105.020 ;
        RECT 22.240 105.005 22.380 105.500 ;
        RECT 23.990 105.440 24.310 105.500 ;
        RECT 34.660 105.360 34.800 105.500 ;
        RECT 41.930 105.500 44.995 105.640 ;
        RECT 41.930 105.440 42.250 105.500 ;
        RECT 44.705 105.455 44.995 105.500 ;
        RECT 69.070 105.640 69.390 105.700 ;
        RECT 71.385 105.640 71.675 105.685 ;
        RECT 69.070 105.500 71.675 105.640 ;
        RECT 69.070 105.440 69.390 105.500 ;
        RECT 71.385 105.455 71.675 105.500 ;
        RECT 79.650 105.640 79.970 105.700 ;
        RECT 83.345 105.640 83.635 105.685 ;
        RECT 79.650 105.500 83.635 105.640 ;
        RECT 79.650 105.440 79.970 105.500 ;
        RECT 83.345 105.455 83.635 105.500 ;
        RECT 97.130 105.440 97.450 105.700 ;
        RECT 25.390 105.300 25.680 105.345 ;
        RECT 27.250 105.300 27.540 105.345 ;
        RECT 30.030 105.300 30.320 105.345 ;
        RECT 25.390 105.160 30.320 105.300 ;
        RECT 25.390 105.115 25.680 105.160 ;
        RECT 27.250 105.115 27.540 105.160 ;
        RECT 30.030 105.115 30.320 105.160 ;
        RECT 34.570 105.300 34.890 105.360 ;
        RECT 52.510 105.300 52.830 105.360 ;
        RECT 86.550 105.300 86.870 105.360 ;
        RECT 34.570 105.160 48.140 105.300 ;
        RECT 34.570 105.100 34.890 105.160 ;
        RECT 8.365 104.820 11.890 104.960 ;
        RECT 8.365 104.775 8.655 104.820 ;
        RECT 11.570 104.760 11.890 104.820 ;
        RECT 22.165 104.775 22.455 105.005 ;
        RECT 24.925 104.960 25.215 105.005 ;
        RECT 27.670 104.960 27.990 105.020 ;
        RECT 24.925 104.820 27.990 104.960 ;
        RECT 24.925 104.775 25.215 104.820 ;
        RECT 27.670 104.760 27.990 104.820 ;
        RECT 36.410 104.960 36.730 105.020 ;
        RECT 48.000 105.005 48.140 105.160 ;
        RECT 52.510 105.160 61.020 105.300 ;
        RECT 52.510 105.100 52.830 105.160 ;
        RECT 47.005 104.960 47.295 105.005 ;
        RECT 36.410 104.820 47.295 104.960 ;
        RECT 36.410 104.760 36.730 104.820 ;
        RECT 47.005 104.775 47.295 104.820 ;
        RECT 47.925 104.960 48.215 105.005 ;
        RECT 55.270 104.960 55.590 105.020 ;
        RECT 47.925 104.820 55.590 104.960 ;
        RECT 47.925 104.775 48.215 104.820 ;
        RECT 55.270 104.760 55.590 104.820 ;
        RECT 56.665 104.960 56.955 105.005 ;
        RECT 59.410 104.960 59.730 105.020 ;
        RECT 60.880 105.005 61.020 105.160 ;
        RECT 86.180 105.160 86.870 105.300 ;
        RECT 56.665 104.820 59.730 104.960 ;
        RECT 56.665 104.775 56.955 104.820 ;
        RECT 59.410 104.760 59.730 104.820 ;
        RECT 60.805 104.775 61.095 105.005 ;
        RECT 74.590 104.760 74.910 105.020 ;
        RECT 86.180 105.005 86.320 105.160 ;
        RECT 86.550 105.100 86.870 105.160 ;
        RECT 97.605 105.115 97.895 105.345 ;
        RECT 86.105 104.775 86.395 105.005 ;
        RECT 91.165 104.960 91.455 105.005 ;
        RECT 96.670 104.960 96.990 105.020 ;
        RECT 91.165 104.820 96.990 104.960 ;
        RECT 91.165 104.775 91.455 104.820 ;
        RECT 96.670 104.760 96.990 104.820 ;
        RECT 8.810 104.620 9.130 104.680 ;
        RECT 10.205 104.620 10.495 104.665 ;
        RECT 13.470 104.620 13.760 104.665 ;
        RECT 8.810 104.480 10.495 104.620 ;
        RECT 8.810 104.420 9.130 104.480 ;
        RECT 10.205 104.435 10.495 104.480 ;
        RECT 11.225 104.480 13.760 104.620 ;
        RECT 11.225 104.325 11.440 104.480 ;
        RECT 13.470 104.435 13.760 104.480 ;
        RECT 26.750 104.420 27.070 104.680 ;
        RECT 30.030 104.620 30.320 104.665 ;
        RECT 27.785 104.480 30.320 104.620 ;
        RECT 9.290 104.280 9.580 104.325 ;
        RECT 11.150 104.280 11.440 104.325 ;
        RECT 9.290 104.140 11.440 104.280 ;
        RECT 9.290 104.095 9.580 104.140 ;
        RECT 11.150 104.095 11.440 104.140 ;
        RECT 12.070 104.280 12.360 104.325 ;
        RECT 14.790 104.280 15.110 104.340 ;
        RECT 27.785 104.325 28.000 104.480 ;
        RECT 30.030 104.435 30.320 104.480 ;
        RECT 46.545 104.620 46.835 104.665 ;
        RECT 48.370 104.620 48.690 104.680 ;
        RECT 46.545 104.480 48.690 104.620 ;
        RECT 46.545 104.435 46.835 104.480 ;
        RECT 48.370 104.420 48.690 104.480 ;
        RECT 57.585 104.620 57.875 104.665 ;
        RECT 58.950 104.620 59.270 104.680 ;
        RECT 59.885 104.620 60.175 104.665 ;
        RECT 57.585 104.480 60.175 104.620 ;
        RECT 57.585 104.435 57.875 104.480 ;
        RECT 58.950 104.420 59.270 104.480 ;
        RECT 59.885 104.435 60.175 104.480 ;
        RECT 73.685 104.620 73.975 104.665 ;
        RECT 75.970 104.620 76.290 104.680 ;
        RECT 73.685 104.480 76.290 104.620 ;
        RECT 73.685 104.435 73.975 104.480 ;
        RECT 75.970 104.420 76.290 104.480 ;
        RECT 76.890 104.620 77.210 104.680 ;
        RECT 81.950 104.620 82.270 104.680 ;
        RECT 85.185 104.620 85.475 104.665 ;
        RECT 76.890 104.480 85.475 104.620 ;
        RECT 76.890 104.420 77.210 104.480 ;
        RECT 81.950 104.420 82.270 104.480 ;
        RECT 85.185 104.435 85.475 104.480 ;
        RECT 85.645 104.620 85.935 104.665 ;
        RECT 86.550 104.620 86.870 104.680 ;
        RECT 87.470 104.620 87.790 104.680 ;
        RECT 85.645 104.480 87.790 104.620 ;
        RECT 85.645 104.435 85.935 104.480 ;
        RECT 86.550 104.420 86.870 104.480 ;
        RECT 87.470 104.420 87.790 104.480 ;
        RECT 90.245 104.620 90.535 104.665 ;
        RECT 92.530 104.620 92.850 104.680 ;
        RECT 90.245 104.480 92.850 104.620 ;
        RECT 90.245 104.435 90.535 104.480 ;
        RECT 92.530 104.420 92.850 104.480 ;
        RECT 93.465 104.435 93.755 104.665 ;
        RECT 96.225 104.620 96.515 104.665 ;
        RECT 97.680 104.620 97.820 105.115 ;
        RECT 98.510 104.960 98.830 105.020 ;
        RECT 100.350 104.960 100.670 105.020 ;
        RECT 114.150 104.960 114.470 105.020 ;
        RECT 98.510 104.820 114.470 104.960 ;
        RECT 98.510 104.760 98.830 104.820 ;
        RECT 100.350 104.760 100.670 104.820 ;
        RECT 114.150 104.760 114.470 104.820 ;
        RECT 96.225 104.480 97.820 104.620 ;
        RECT 96.225 104.435 96.515 104.480 ;
        RECT 15.330 104.280 15.620 104.325 ;
        RECT 12.070 104.140 15.620 104.280 ;
        RECT 12.070 104.095 12.360 104.140 ;
        RECT 14.790 104.080 15.110 104.140 ;
        RECT 15.330 104.095 15.620 104.140 ;
        RECT 25.850 104.280 26.140 104.325 ;
        RECT 27.710 104.280 28.000 104.325 ;
        RECT 25.850 104.140 28.000 104.280 ;
        RECT 25.850 104.095 26.140 104.140 ;
        RECT 27.710 104.095 28.000 104.140 ;
        RECT 28.630 104.280 28.920 104.325 ;
        RECT 29.510 104.280 29.830 104.340 ;
        RECT 31.890 104.280 32.180 104.325 ;
        RECT 28.630 104.140 32.180 104.280 ;
        RECT 28.630 104.095 28.920 104.140 ;
        RECT 29.510 104.080 29.830 104.140 ;
        RECT 31.890 104.095 32.180 104.140 ;
        RECT 58.505 104.280 58.795 104.325 ;
        RECT 59.410 104.280 59.730 104.340 ;
        RECT 58.505 104.140 59.730 104.280 ;
        RECT 58.505 104.095 58.795 104.140 ;
        RECT 59.410 104.080 59.730 104.140 ;
        RECT 73.225 104.280 73.515 104.325 ;
        RECT 75.050 104.280 75.370 104.340 ;
        RECT 73.225 104.140 75.370 104.280 ;
        RECT 93.540 104.280 93.680 104.435 ;
        RECT 103.110 104.420 103.430 104.680 ;
        RECT 105.410 104.280 105.730 104.340 ;
        RECT 93.540 104.140 105.730 104.280 ;
        RECT 73.225 104.095 73.515 104.140 ;
        RECT 75.050 104.080 75.370 104.140 ;
        RECT 105.410 104.080 105.730 104.140 ;
        RECT 17.335 103.940 17.625 103.985 ;
        RECT 20.770 103.940 21.090 104.000 ;
        RECT 17.335 103.800 21.090 103.940 ;
        RECT 17.335 103.755 17.625 103.800 ;
        RECT 20.770 103.740 21.090 103.800 ;
        RECT 21.245 103.940 21.535 103.985 ;
        RECT 21.690 103.940 22.010 104.000 ;
        RECT 21.245 103.800 22.010 103.940 ;
        RECT 21.245 103.755 21.535 103.800 ;
        RECT 21.690 103.740 22.010 103.800 ;
        RECT 29.970 103.940 30.290 104.000 ;
        RECT 33.895 103.940 34.185 103.985 ;
        RECT 29.970 103.800 34.185 103.940 ;
        RECT 29.970 103.740 30.290 103.800 ;
        RECT 33.895 103.755 34.185 103.800 ;
        RECT 58.965 103.940 59.255 103.985 ;
        RECT 60.330 103.940 60.650 104.000 ;
        RECT 58.965 103.800 60.650 103.940 ;
        RECT 58.965 103.755 59.255 103.800 ;
        RECT 60.330 103.740 60.650 103.800 ;
        RECT 88.850 103.940 89.170 104.000 ;
        RECT 89.325 103.940 89.615 103.985 ;
        RECT 88.850 103.800 89.615 103.940 ;
        RECT 88.850 103.740 89.170 103.800 ;
        RECT 89.325 103.755 89.615 103.800 ;
        RECT 91.610 103.740 91.930 104.000 ;
        RECT 99.430 103.740 99.750 104.000 ;
        RECT 99.905 103.940 100.195 103.985 ;
        RECT 102.650 103.940 102.970 104.000 ;
        RECT 99.905 103.800 102.970 103.940 ;
        RECT 99.905 103.755 100.195 103.800 ;
        RECT 102.650 103.740 102.970 103.800 ;
        RECT 109.565 103.940 109.855 103.985 ;
        RECT 110.010 103.940 110.330 104.000 ;
        RECT 109.565 103.800 110.330 103.940 ;
        RECT 109.565 103.755 109.855 103.800 ;
        RECT 110.010 103.740 110.330 103.800 ;
        RECT 5.520 103.120 125.580 103.600 ;
        RECT 18.470 102.920 18.790 102.980 ;
        RECT 19.175 102.920 19.465 102.965 ;
        RECT 23.530 102.920 23.850 102.980 ;
        RECT 24.925 102.920 25.215 102.965 ;
        RECT 18.470 102.780 22.380 102.920 ;
        RECT 18.470 102.720 18.790 102.780 ;
        RECT 19.175 102.735 19.465 102.780 ;
        RECT 11.130 102.580 11.420 102.625 ;
        RECT 12.990 102.580 13.280 102.625 ;
        RECT 11.130 102.440 13.280 102.580 ;
        RECT 11.130 102.395 11.420 102.440 ;
        RECT 12.990 102.395 13.280 102.440 ;
        RECT 13.910 102.580 14.200 102.625 ;
        RECT 15.710 102.580 16.030 102.640 ;
        RECT 17.170 102.580 17.460 102.625 ;
        RECT 13.910 102.440 17.460 102.580 ;
        RECT 22.240 102.580 22.380 102.780 ;
        RECT 23.530 102.780 25.215 102.920 ;
        RECT 23.530 102.720 23.850 102.780 ;
        RECT 24.925 102.735 25.215 102.780 ;
        RECT 26.765 102.920 27.055 102.965 ;
        RECT 28.130 102.920 28.450 102.980 ;
        RECT 29.970 102.920 30.290 102.980 ;
        RECT 26.765 102.780 30.290 102.920 ;
        RECT 26.765 102.735 27.055 102.780 ;
        RECT 28.130 102.720 28.450 102.780 ;
        RECT 29.970 102.720 30.290 102.780 ;
        RECT 88.390 102.720 88.710 102.980 ;
        RECT 90.230 102.920 90.550 102.980 ;
        RECT 91.165 102.920 91.455 102.965 ;
        RECT 90.230 102.780 91.455 102.920 ;
        RECT 90.230 102.720 90.550 102.780 ;
        RECT 91.165 102.735 91.455 102.780 ;
        RECT 27.225 102.580 27.515 102.625 ;
        RECT 22.240 102.440 27.515 102.580 ;
        RECT 13.910 102.395 14.200 102.440 ;
        RECT 10.205 102.240 10.495 102.285 ;
        RECT 11.570 102.240 11.890 102.300 ;
        RECT 10.205 102.100 11.890 102.240 ;
        RECT 10.205 102.055 10.495 102.100 ;
        RECT 11.570 102.040 11.890 102.100 ;
        RECT 12.045 102.240 12.335 102.285 ;
        RECT 12.490 102.240 12.810 102.300 ;
        RECT 12.045 102.100 12.810 102.240 ;
        RECT 13.065 102.240 13.280 102.395 ;
        RECT 15.710 102.380 16.030 102.440 ;
        RECT 17.170 102.395 17.460 102.440 ;
        RECT 27.225 102.395 27.515 102.440 ;
        RECT 60.790 102.580 61.110 102.640 ;
        RECT 62.185 102.580 62.475 102.625 ;
        RECT 99.430 102.580 99.750 102.640 ;
        RECT 60.790 102.440 62.475 102.580 ;
        RECT 60.790 102.380 61.110 102.440 ;
        RECT 62.185 102.395 62.475 102.440 ;
        RECT 94.000 102.440 99.750 102.580 ;
        RECT 15.310 102.240 15.600 102.285 ;
        RECT 13.065 102.100 15.600 102.240 ;
        RECT 12.045 102.055 12.335 102.100 ;
        RECT 12.490 102.040 12.810 102.100 ;
        RECT 15.310 102.055 15.600 102.100 ;
        RECT 43.310 102.240 43.630 102.300 ;
        RECT 47.925 102.240 48.215 102.285 ;
        RECT 43.310 102.100 48.215 102.240 ;
        RECT 43.310 102.040 43.630 102.100 ;
        RECT 47.925 102.055 48.215 102.100 ;
        RECT 53.890 102.240 54.210 102.300 ;
        RECT 54.825 102.240 55.115 102.285 ;
        RECT 53.890 102.100 55.115 102.240 ;
        RECT 53.890 102.040 54.210 102.100 ;
        RECT 54.825 102.055 55.115 102.100 ;
        RECT 55.745 102.240 56.035 102.285 ;
        RECT 58.505 102.240 58.795 102.285 ;
        RECT 58.950 102.240 59.270 102.300 ;
        RECT 55.745 102.100 59.270 102.240 ;
        RECT 55.745 102.055 56.035 102.100 ;
        RECT 58.505 102.055 58.795 102.100 ;
        RECT 58.950 102.040 59.270 102.100 ;
        RECT 59.425 102.240 59.715 102.285 ;
        RECT 59.870 102.240 60.190 102.300 ;
        RECT 59.425 102.100 60.190 102.240 ;
        RECT 59.425 102.055 59.715 102.100 ;
        RECT 59.870 102.040 60.190 102.100 ;
        RECT 64.025 102.240 64.315 102.285 ;
        RECT 64.930 102.240 65.250 102.300 ;
        RECT 64.025 102.100 65.250 102.240 ;
        RECT 64.025 102.055 64.315 102.100 ;
        RECT 64.930 102.040 65.250 102.100 ;
        RECT 84.250 102.240 84.570 102.300 ;
        RECT 86.105 102.240 86.395 102.285 ;
        RECT 84.250 102.100 86.395 102.240 ;
        RECT 84.250 102.040 84.570 102.100 ;
        RECT 86.105 102.055 86.395 102.100 ;
        RECT 87.470 102.040 87.790 102.300 ;
        RECT 87.930 102.240 88.250 102.300 ;
        RECT 88.865 102.240 89.155 102.285 ;
        RECT 87.930 102.100 89.155 102.240 ;
        RECT 87.930 102.040 88.250 102.100 ;
        RECT 88.865 102.055 89.155 102.100 ;
        RECT 90.230 102.040 90.550 102.300 ;
        RECT 92.530 102.240 92.850 102.300 ;
        RECT 94.000 102.285 94.140 102.440 ;
        RECT 99.430 102.380 99.750 102.440 ;
        RECT 93.005 102.240 93.295 102.285 ;
        RECT 92.530 102.100 93.295 102.240 ;
        RECT 92.530 102.040 92.850 102.100 ;
        RECT 93.005 102.055 93.295 102.100 ;
        RECT 93.925 102.055 94.215 102.285 ;
        RECT 95.305 102.055 95.595 102.285 ;
        RECT 101.730 102.240 102.050 102.300 ;
        RECT 111.405 102.240 111.695 102.285 ;
        RECT 118.750 102.240 119.070 102.300 ;
        RECT 101.730 102.100 119.070 102.240 ;
        RECT 23.990 101.900 24.310 101.960 ;
        RECT 27.685 101.900 27.975 101.945 ;
        RECT 23.990 101.760 27.975 101.900 ;
        RECT 23.990 101.700 24.310 101.760 ;
        RECT 27.685 101.715 27.975 101.760 ;
        RECT 87.025 101.900 87.315 101.945 ;
        RECT 88.390 101.900 88.710 101.960 ;
        RECT 87.025 101.760 88.710 101.900 ;
        RECT 87.025 101.715 87.315 101.760 ;
        RECT 88.390 101.700 88.710 101.760 ;
        RECT 89.770 101.700 90.090 101.960 ;
        RECT 93.080 101.900 93.220 102.055 ;
        RECT 94.830 101.900 95.150 101.960 ;
        RECT 95.380 101.900 95.520 102.055 ;
        RECT 101.730 102.040 102.050 102.100 ;
        RECT 111.405 102.055 111.695 102.100 ;
        RECT 118.750 102.040 119.070 102.100 ;
        RECT 90.320 101.760 92.760 101.900 ;
        RECT 93.080 101.760 95.520 101.900 ;
        RECT 96.225 101.900 96.515 101.945 ;
        RECT 116.910 101.900 117.230 101.960 ;
        RECT 96.225 101.760 117.230 101.900 ;
        RECT 10.670 101.560 10.960 101.605 ;
        RECT 12.530 101.560 12.820 101.605 ;
        RECT 15.310 101.560 15.600 101.605 ;
        RECT 10.670 101.420 15.600 101.560 ;
        RECT 10.670 101.375 10.960 101.420 ;
        RECT 12.530 101.375 12.820 101.420 ;
        RECT 15.310 101.375 15.600 101.420 ;
        RECT 69.070 101.560 69.390 101.620 ;
        RECT 90.320 101.560 90.460 101.760 ;
        RECT 69.070 101.420 90.460 101.560 ;
        RECT 90.690 101.560 91.010 101.620 ;
        RECT 92.085 101.560 92.375 101.605 ;
        RECT 90.690 101.420 92.375 101.560 ;
        RECT 92.620 101.560 92.760 101.760 ;
        RECT 94.830 101.700 95.150 101.760 ;
        RECT 96.225 101.715 96.515 101.760 ;
        RECT 116.910 101.700 117.230 101.760 ;
        RECT 98.970 101.560 99.290 101.620 ;
        RECT 100.350 101.560 100.670 101.620 ;
        RECT 92.620 101.420 100.670 101.560 ;
        RECT 69.070 101.360 69.390 101.420 ;
        RECT 90.690 101.360 91.010 101.420 ;
        RECT 92.085 101.375 92.375 101.420 ;
        RECT 98.970 101.360 99.290 101.420 ;
        RECT 100.350 101.360 100.670 101.420 ;
        RECT 48.370 101.020 48.690 101.280 ;
        RECT 56.650 101.020 56.970 101.280 ;
        RECT 57.570 101.020 57.890 101.280 ;
        RECT 87.485 101.220 87.775 101.265 ;
        RECT 88.850 101.220 89.170 101.280 ;
        RECT 87.485 101.080 89.170 101.220 ;
        RECT 87.485 101.035 87.775 101.080 ;
        RECT 88.850 101.020 89.170 101.080 ;
        RECT 89.325 101.220 89.615 101.265 ;
        RECT 91.610 101.220 91.930 101.280 ;
        RECT 89.325 101.080 91.930 101.220 ;
        RECT 89.325 101.035 89.615 101.080 ;
        RECT 91.610 101.020 91.930 101.080 ;
        RECT 94.370 101.020 94.690 101.280 ;
        RECT 110.930 101.020 111.250 101.280 ;
        RECT 5.520 100.400 125.580 100.880 ;
        RECT 14.790 100.000 15.110 100.260 ;
        RECT 37.420 100.060 50.440 100.200 ;
        RECT 21.690 99.860 22.010 99.920 ;
        RECT 21.690 99.720 27.900 99.860 ;
        RECT 21.690 99.660 22.010 99.720 ;
        RECT 20.770 99.520 21.090 99.580 ;
        RECT 27.760 99.565 27.900 99.720 ;
        RECT 21.245 99.520 21.535 99.565 ;
        RECT 20.770 99.380 21.535 99.520 ;
        RECT 20.770 99.320 21.090 99.380 ;
        RECT 21.245 99.335 21.535 99.380 ;
        RECT 22.240 99.380 24.680 99.520 ;
        RECT 15.265 99.180 15.555 99.225 ;
        RECT 16.170 99.180 16.490 99.240 ;
        RECT 22.240 99.225 22.380 99.380 ;
        RECT 24.540 99.225 24.680 99.380 ;
        RECT 27.685 99.335 27.975 99.565 ;
        RECT 28.130 99.320 28.450 99.580 ;
        RECT 32.270 99.320 32.590 99.580 ;
        RECT 36.410 99.320 36.730 99.580 ;
        RECT 37.420 99.225 37.560 100.060 ;
        RECT 45.170 99.860 45.460 99.905 ;
        RECT 47.030 99.860 47.320 99.905 ;
        RECT 49.810 99.860 50.100 99.905 ;
        RECT 45.170 99.720 50.100 99.860 ;
        RECT 50.300 99.860 50.440 100.060 ;
        RECT 56.650 100.000 56.970 100.260 ;
        RECT 58.045 100.200 58.335 100.245 ;
        RECT 58.490 100.200 58.810 100.260 ;
        RECT 58.045 100.060 58.810 100.200 ;
        RECT 58.045 100.015 58.335 100.060 ;
        RECT 58.490 100.000 58.810 100.060 ;
        RECT 69.070 100.000 69.390 100.260 ;
        RECT 84.250 100.000 84.570 100.260 ;
        RECT 86.180 100.060 87.240 100.200 ;
        RECT 63.550 99.860 63.870 99.920 ;
        RECT 50.300 99.720 63.870 99.860 ;
        RECT 45.170 99.675 45.460 99.720 ;
        RECT 47.030 99.675 47.320 99.720 ;
        RECT 49.810 99.675 50.100 99.720 ;
        RECT 63.550 99.660 63.870 99.720 ;
        RECT 67.690 99.860 68.010 99.920 ;
        RECT 72.305 99.860 72.595 99.905 ;
        RECT 67.690 99.720 72.595 99.860 ;
        RECT 67.690 99.660 68.010 99.720 ;
        RECT 72.305 99.675 72.595 99.720 ;
        RECT 79.190 99.860 79.510 99.920 ;
        RECT 82.410 99.860 82.730 99.920 ;
        RECT 86.180 99.860 86.320 100.060 ;
        RECT 79.190 99.720 86.320 99.860 ;
        RECT 79.190 99.660 79.510 99.720 ;
        RECT 82.410 99.660 82.730 99.720 ;
        RECT 86.550 99.660 86.870 99.920 ;
        RECT 41.470 99.520 41.790 99.580 ;
        RECT 44.690 99.520 45.010 99.580 ;
        RECT 41.470 99.380 45.010 99.520 ;
        RECT 41.470 99.320 41.790 99.380 ;
        RECT 44.690 99.320 45.010 99.380 ;
        RECT 53.890 99.520 54.210 99.580 ;
        RECT 56.205 99.520 56.495 99.565 ;
        RECT 53.890 99.380 56.495 99.520 ;
        RECT 53.890 99.320 54.210 99.380 ;
        RECT 56.205 99.335 56.495 99.380 ;
        RECT 75.970 99.520 76.290 99.580 ;
        RECT 86.640 99.520 86.780 99.660 ;
        RECT 75.970 99.380 78.500 99.520 ;
        RECT 75.970 99.320 76.290 99.380 ;
        RECT 15.265 99.040 16.490 99.180 ;
        RECT 15.265 98.995 15.555 99.040 ;
        RECT 16.170 98.980 16.490 99.040 ;
        RECT 22.165 98.995 22.455 99.225 ;
        RECT 23.545 98.995 23.835 99.225 ;
        RECT 24.465 99.180 24.755 99.225 ;
        RECT 26.765 99.180 27.055 99.225 ;
        RECT 24.465 99.040 27.055 99.180 ;
        RECT 24.465 98.995 24.755 99.040 ;
        RECT 26.765 98.995 27.055 99.040 ;
        RECT 29.065 99.180 29.355 99.225 ;
        RECT 31.365 99.180 31.655 99.225 ;
        RECT 37.345 99.180 37.635 99.225 ;
        RECT 29.065 99.040 37.635 99.180 ;
        RECT 29.065 98.995 29.355 99.040 ;
        RECT 31.365 98.995 31.655 99.040 ;
        RECT 37.345 98.995 37.635 99.040 ;
        RECT 18.470 98.840 18.790 98.900 ;
        RECT 23.620 98.840 23.760 98.995 ;
        RECT 18.470 98.700 23.760 98.840 ;
        RECT 26.840 98.840 26.980 98.995 ;
        RECT 29.140 98.840 29.280 98.995 ;
        RECT 38.710 98.980 39.030 99.240 ;
        RECT 46.545 99.180 46.835 99.225 ;
        RECT 46.990 99.180 47.310 99.240 ;
        RECT 49.810 99.180 50.100 99.225 ;
        RECT 46.545 99.040 47.310 99.180 ;
        RECT 46.545 98.995 46.835 99.040 ;
        RECT 46.990 98.980 47.310 99.040 ;
        RECT 47.565 99.040 50.100 99.180 ;
        RECT 47.565 98.885 47.780 99.040 ;
        RECT 49.810 98.995 50.100 99.040 ;
        RECT 53.430 99.180 53.750 99.240 ;
        RECT 55.745 99.180 56.035 99.225 ;
        RECT 53.430 99.040 56.035 99.180 ;
        RECT 53.430 98.980 53.750 99.040 ;
        RECT 55.745 98.995 56.035 99.040 ;
        RECT 57.110 98.980 57.430 99.240 ;
        RECT 71.830 98.980 72.150 99.240 ;
        RECT 73.210 98.980 73.530 99.240 ;
        RECT 78.360 99.225 78.500 99.380 ;
        RECT 78.820 99.380 85.400 99.520 ;
        RECT 78.820 99.240 78.960 99.380 ;
        RECT 77.365 98.995 77.655 99.225 ;
        RECT 78.285 98.995 78.575 99.225 ;
        RECT 26.840 98.700 29.280 98.840 ;
        RECT 45.630 98.840 45.920 98.885 ;
        RECT 47.490 98.840 47.780 98.885 ;
        RECT 45.630 98.700 47.780 98.840 ;
        RECT 18.470 98.640 18.790 98.700 ;
        RECT 45.630 98.655 45.920 98.700 ;
        RECT 47.490 98.655 47.780 98.700 ;
        RECT 48.370 98.885 48.690 98.900 ;
        RECT 48.370 98.840 48.700 98.885 ;
        RECT 51.670 98.840 51.960 98.885 ;
        RECT 48.370 98.700 51.960 98.840 ;
        RECT 48.370 98.655 48.700 98.700 ;
        RECT 51.670 98.655 51.960 98.700 ;
        RECT 64.930 98.840 65.250 98.900 ;
        RECT 67.705 98.840 67.995 98.885 ;
        RECT 64.930 98.700 67.995 98.840 ;
        RECT 71.920 98.840 72.060 98.980 ;
        RECT 74.130 98.840 74.450 98.900 ;
        RECT 71.920 98.700 74.450 98.840 ;
        RECT 48.370 98.640 48.690 98.655 ;
        RECT 64.930 98.640 65.250 98.700 ;
        RECT 67.705 98.655 67.995 98.700 ;
        RECT 74.130 98.640 74.450 98.700 ;
        RECT 75.970 98.840 76.290 98.900 ;
        RECT 77.440 98.840 77.580 98.995 ;
        RECT 78.730 98.980 79.050 99.240 ;
        RECT 79.190 98.980 79.510 99.240 ;
        RECT 81.045 98.995 81.335 99.225 ;
        RECT 81.120 98.840 81.260 98.995 ;
        RECT 81.950 98.980 82.270 99.240 ;
        RECT 82.500 99.225 82.640 99.380 ;
        RECT 82.425 98.995 82.715 99.225 ;
        RECT 82.870 98.980 83.190 99.240 ;
        RECT 84.725 98.995 85.015 99.225 ;
        RECT 84.800 98.840 84.940 98.995 ;
        RECT 75.970 98.700 84.940 98.840 ;
        RECT 85.260 98.840 85.400 99.380 ;
        RECT 85.720 99.380 86.780 99.520 ;
        RECT 85.720 99.225 85.860 99.380 ;
        RECT 85.645 98.995 85.935 99.225 ;
        RECT 86.105 98.995 86.395 99.225 ;
        RECT 86.565 99.180 86.855 99.225 ;
        RECT 87.100 99.180 87.240 100.060 ;
        RECT 87.930 100.000 88.250 100.260 ;
        RECT 105.890 99.860 106.180 99.905 ;
        RECT 107.750 99.860 108.040 99.905 ;
        RECT 110.530 99.860 110.820 99.905 ;
        RECT 105.890 99.720 110.820 99.860 ;
        RECT 105.890 99.675 106.180 99.720 ;
        RECT 107.750 99.675 108.040 99.720 ;
        RECT 110.530 99.675 110.820 99.720 ;
        RECT 95.750 99.520 96.070 99.580 ;
        RECT 105.425 99.520 105.715 99.565 ;
        RECT 110.010 99.520 110.330 99.580 ;
        RECT 95.750 99.380 110.330 99.520 ;
        RECT 95.750 99.320 96.070 99.380 ;
        RECT 105.425 99.335 105.715 99.380 ;
        RECT 110.010 99.320 110.330 99.380 ;
        RECT 114.150 99.520 114.470 99.580 ;
        RECT 115.545 99.520 115.835 99.565 ;
        RECT 114.150 99.380 115.835 99.520 ;
        RECT 114.150 99.320 114.470 99.380 ;
        RECT 115.545 99.335 115.835 99.380 ;
        RECT 118.750 99.520 119.070 99.580 ;
        RECT 118.750 99.380 122.200 99.520 ;
        RECT 118.750 99.320 119.070 99.380 ;
        RECT 86.565 99.040 87.240 99.180 ;
        RECT 94.385 99.180 94.675 99.225 ;
        RECT 94.830 99.180 95.150 99.240 ;
        RECT 94.385 99.040 95.150 99.180 ;
        RECT 86.565 98.995 86.855 99.040 ;
        RECT 94.385 98.995 94.675 99.040 ;
        RECT 86.180 98.840 86.320 98.995 ;
        RECT 94.830 98.980 95.150 99.040 ;
        RECT 95.305 98.995 95.595 99.225 ;
        RECT 85.260 98.700 86.320 98.840 ;
        RECT 95.380 98.840 95.520 98.995 ;
        RECT 98.050 98.980 98.370 99.240 ;
        RECT 101.730 98.980 102.050 99.240 ;
        RECT 107.250 98.980 107.570 99.240 ;
        RECT 122.060 99.225 122.200 99.380 ;
        RECT 110.530 99.180 110.820 99.225 ;
        RECT 120.145 99.180 120.435 99.225 ;
        RECT 108.285 99.040 110.820 99.180 ;
        RECT 102.650 98.840 102.970 98.900 ;
        RECT 108.285 98.885 108.500 99.040 ;
        RECT 110.530 98.995 110.820 99.040 ;
        RECT 118.840 99.040 120.435 99.180 ;
        RECT 95.380 98.700 102.970 98.840 ;
        RECT 75.970 98.640 76.290 98.700 ;
        RECT 82.500 98.560 82.640 98.700 ;
        RECT 102.650 98.640 102.970 98.700 ;
        RECT 106.350 98.840 106.640 98.885 ;
        RECT 108.210 98.840 108.500 98.885 ;
        RECT 106.350 98.700 108.500 98.840 ;
        RECT 106.350 98.655 106.640 98.700 ;
        RECT 108.210 98.655 108.500 98.700 ;
        RECT 109.130 98.840 109.420 98.885 ;
        RECT 110.930 98.840 111.250 98.900 ;
        RECT 112.390 98.840 112.680 98.885 ;
        RECT 109.130 98.700 112.680 98.840 ;
        RECT 109.130 98.655 109.420 98.700 ;
        RECT 110.930 98.640 111.250 98.700 ;
        RECT 112.390 98.655 112.680 98.700 ;
        RECT 113.690 98.840 114.010 98.900 ;
        RECT 116.465 98.840 116.755 98.885 ;
        RECT 113.690 98.700 116.755 98.840 ;
        RECT 113.690 98.640 114.010 98.700 ;
        RECT 116.465 98.655 116.755 98.700 ;
        RECT 23.085 98.500 23.375 98.545 ;
        RECT 23.530 98.500 23.850 98.560 ;
        RECT 23.085 98.360 23.850 98.500 ;
        RECT 23.085 98.315 23.375 98.360 ;
        RECT 23.530 98.300 23.850 98.360 ;
        RECT 23.990 98.500 24.310 98.560 ;
        RECT 25.385 98.500 25.675 98.545 ;
        RECT 23.990 98.360 25.675 98.500 ;
        RECT 23.990 98.300 24.310 98.360 ;
        RECT 25.385 98.315 25.675 98.360 ;
        RECT 25.845 98.500 26.135 98.545 ;
        RECT 26.750 98.500 27.070 98.560 ;
        RECT 25.845 98.360 27.070 98.500 ;
        RECT 25.845 98.315 26.135 98.360 ;
        RECT 26.750 98.300 27.070 98.360 ;
        RECT 29.970 98.300 30.290 98.560 ;
        RECT 30.445 98.500 30.735 98.545 ;
        RECT 31.350 98.500 31.670 98.560 ;
        RECT 30.445 98.360 31.670 98.500 ;
        RECT 30.445 98.315 30.735 98.360 ;
        RECT 31.350 98.300 31.670 98.360 ;
        RECT 38.250 98.300 38.570 98.560 ;
        RECT 39.170 98.500 39.490 98.560 ;
        RECT 39.645 98.500 39.935 98.545 ;
        RECT 39.170 98.360 39.935 98.500 ;
        RECT 39.170 98.300 39.490 98.360 ;
        RECT 39.645 98.315 39.935 98.360 ;
        RECT 50.670 98.500 50.990 98.560 ;
        RECT 53.675 98.500 53.965 98.545 ;
        RECT 56.650 98.500 56.970 98.560 ;
        RECT 50.670 98.360 56.970 98.500 ;
        RECT 50.670 98.300 50.990 98.360 ;
        RECT 53.675 98.315 53.965 98.360 ;
        RECT 56.650 98.300 56.970 98.360 ;
        RECT 58.490 98.500 58.810 98.560 ;
        RECT 67.230 98.500 67.550 98.560 ;
        RECT 58.490 98.360 67.550 98.500 ;
        RECT 58.490 98.300 58.810 98.360 ;
        RECT 67.230 98.300 67.550 98.360 ;
        RECT 71.370 98.300 71.690 98.560 ;
        RECT 80.570 98.300 80.890 98.560 ;
        RECT 82.410 98.300 82.730 98.560 ;
        RECT 82.870 98.500 83.190 98.560 ;
        RECT 93.465 98.500 93.755 98.545 ;
        RECT 82.870 98.360 93.755 98.500 ;
        RECT 82.870 98.300 83.190 98.360 ;
        RECT 93.465 98.315 93.755 98.360 ;
        RECT 97.145 98.500 97.435 98.545 ;
        RECT 97.590 98.500 97.910 98.560 ;
        RECT 97.145 98.360 97.910 98.500 ;
        RECT 97.145 98.315 97.435 98.360 ;
        RECT 97.590 98.300 97.910 98.360 ;
        RECT 101.270 98.300 101.590 98.560 ;
        RECT 101.730 98.500 102.050 98.560 ;
        RECT 111.390 98.500 111.710 98.560 ;
        RECT 114.395 98.500 114.685 98.545 ;
        RECT 101.730 98.360 114.685 98.500 ;
        RECT 101.730 98.300 102.050 98.360 ;
        RECT 111.390 98.300 111.710 98.360 ;
        RECT 114.395 98.315 114.685 98.360 ;
        RECT 116.910 98.300 117.230 98.560 ;
        RECT 118.840 98.545 118.980 99.040 ;
        RECT 120.145 98.995 120.435 99.040 ;
        RECT 121.985 98.995 122.275 99.225 ;
        RECT 118.765 98.315 119.055 98.545 ;
        RECT 119.210 98.300 119.530 98.560 ;
        RECT 122.430 98.300 122.750 98.560 ;
        RECT 5.520 97.680 125.580 98.160 ;
        RECT 41.470 97.480 41.790 97.540 ;
        RECT 37.880 97.340 41.790 97.480 ;
        RECT 14.345 96.800 14.635 96.845 ;
        RECT 17.090 96.800 17.410 96.860 ;
        RECT 14.345 96.660 17.410 96.800 ;
        RECT 14.345 96.615 14.635 96.660 ;
        RECT 17.090 96.600 17.410 96.660 ;
        RECT 29.050 96.800 29.370 96.860 ;
        RECT 33.665 96.800 33.955 96.845 ;
        RECT 37.345 96.800 37.635 96.845 ;
        RECT 37.880 96.800 38.020 97.340 ;
        RECT 41.470 97.280 41.790 97.340 ;
        RECT 46.990 97.280 47.310 97.540 ;
        RECT 48.385 97.295 48.675 97.525 ;
        RECT 38.270 97.140 38.560 97.185 ;
        RECT 40.130 97.140 40.420 97.185 ;
        RECT 38.270 97.000 40.420 97.140 ;
        RECT 38.270 96.955 38.560 97.000 ;
        RECT 40.130 96.955 40.420 97.000 ;
        RECT 41.050 97.140 41.340 97.185 ;
        RECT 42.850 97.140 43.170 97.200 ;
        RECT 44.310 97.140 44.600 97.185 ;
        RECT 41.050 97.000 44.600 97.140 ;
        RECT 41.050 96.955 41.340 97.000 ;
        RECT 29.050 96.660 37.100 96.800 ;
        RECT 29.050 96.600 29.370 96.660 ;
        RECT 33.665 96.615 33.955 96.660 ;
        RECT 36.960 96.460 37.100 96.660 ;
        RECT 37.345 96.660 38.020 96.800 ;
        RECT 37.345 96.615 37.635 96.660 ;
        RECT 39.170 96.600 39.490 96.860 ;
        RECT 40.205 96.800 40.420 96.955 ;
        RECT 42.850 96.940 43.170 97.000 ;
        RECT 44.310 96.955 44.600 97.000 ;
        RECT 42.450 96.800 42.740 96.845 ;
        RECT 40.205 96.660 42.740 96.800 ;
        RECT 42.450 96.615 42.740 96.660 ;
        RECT 47.925 96.800 48.215 96.845 ;
        RECT 48.460 96.800 48.600 97.295 ;
        RECT 50.670 97.280 50.990 97.540 ;
        RECT 53.430 97.280 53.750 97.540 ;
        RECT 56.650 97.480 56.970 97.540 ;
        RECT 56.650 97.340 58.720 97.480 ;
        RECT 56.650 97.280 56.970 97.340 ;
        RECT 50.300 97.000 55.960 97.140 ;
        RECT 50.300 96.845 50.440 97.000 ;
        RECT 55.820 96.845 55.960 97.000 ;
        RECT 50.225 96.800 50.515 96.845 ;
        RECT 47.925 96.660 48.600 96.800 ;
        RECT 48.920 96.660 50.515 96.800 ;
        RECT 47.925 96.615 48.215 96.660 ;
        RECT 43.310 96.460 43.630 96.520 ;
        RECT 48.920 96.460 49.060 96.660 ;
        RECT 50.225 96.615 50.515 96.660 ;
        RECT 54.825 96.615 55.115 96.845 ;
        RECT 55.285 96.615 55.575 96.845 ;
        RECT 55.745 96.615 56.035 96.845 ;
        RECT 56.190 96.800 56.510 96.860 ;
        RECT 58.580 96.845 58.720 97.340 ;
        RECT 64.930 97.280 65.250 97.540 ;
        RECT 67.230 97.480 67.550 97.540 ;
        RECT 81.490 97.480 81.810 97.540 ;
        RECT 83.345 97.480 83.635 97.525 ;
        RECT 67.230 97.340 74.360 97.480 ;
        RECT 67.230 97.280 67.550 97.340 ;
        RECT 61.250 97.140 61.570 97.200 ;
        RECT 66.790 97.140 67.080 97.185 ;
        RECT 68.650 97.140 68.940 97.185 ;
        RECT 59.040 97.000 66.540 97.140 ;
        RECT 59.040 96.845 59.180 97.000 ;
        RECT 61.250 96.940 61.570 97.000 ;
        RECT 56.665 96.800 56.955 96.845 ;
        RECT 57.585 96.800 57.875 96.845 ;
        RECT 56.190 96.660 57.875 96.800 ;
        RECT 36.960 96.320 43.630 96.460 ;
        RECT 43.310 96.260 43.630 96.320 ;
        RECT 48.000 96.320 49.060 96.460 ;
        RECT 51.605 96.460 51.895 96.505 ;
        RECT 52.050 96.460 52.370 96.520 ;
        RECT 51.605 96.320 52.370 96.460 ;
        RECT 37.810 96.120 38.100 96.165 ;
        RECT 39.670 96.120 39.960 96.165 ;
        RECT 42.450 96.120 42.740 96.165 ;
        RECT 37.810 95.980 42.740 96.120 ;
        RECT 37.810 95.935 38.100 95.980 ;
        RECT 39.670 95.935 39.960 95.980 ;
        RECT 42.450 95.935 42.740 95.980 ;
        RECT 12.030 95.780 12.350 95.840 ;
        RECT 13.425 95.780 13.715 95.825 ;
        RECT 12.030 95.640 13.715 95.780 ;
        RECT 12.030 95.580 12.350 95.640 ;
        RECT 13.425 95.595 13.715 95.640 ;
        RECT 33.190 95.580 33.510 95.840 ;
        RECT 41.930 95.780 42.250 95.840 ;
        RECT 46.315 95.780 46.605 95.825 ;
        RECT 48.000 95.780 48.140 96.320 ;
        RECT 51.605 96.275 51.895 96.320 ;
        RECT 52.050 96.260 52.370 96.320 ;
        RECT 54.900 96.120 55.040 96.615 ;
        RECT 55.360 96.460 55.500 96.615 ;
        RECT 56.190 96.600 56.510 96.660 ;
        RECT 56.665 96.615 56.955 96.660 ;
        RECT 57.585 96.615 57.875 96.660 ;
        RECT 58.505 96.615 58.795 96.845 ;
        RECT 58.965 96.615 59.255 96.845 ;
        RECT 59.425 96.800 59.715 96.845 ;
        RECT 61.710 96.800 62.030 96.860 ;
        RECT 59.425 96.660 62.030 96.800 ;
        RECT 59.425 96.615 59.715 96.660 ;
        RECT 59.040 96.460 59.180 96.615 ;
        RECT 55.360 96.320 59.180 96.460 ;
        RECT 59.500 96.120 59.640 96.615 ;
        RECT 61.710 96.600 62.030 96.660 ;
        RECT 64.025 96.800 64.315 96.845 ;
        RECT 64.470 96.800 64.790 96.860 ;
        RECT 64.025 96.660 64.790 96.800 ;
        RECT 66.400 96.800 66.540 97.000 ;
        RECT 66.790 97.000 68.940 97.140 ;
        RECT 66.790 96.955 67.080 97.000 ;
        RECT 68.650 96.955 68.940 97.000 ;
        RECT 69.570 97.140 69.860 97.185 ;
        RECT 71.370 97.140 71.690 97.200 ;
        RECT 72.830 97.140 73.120 97.185 ;
        RECT 69.570 97.000 73.120 97.140 ;
        RECT 69.570 96.955 69.860 97.000 ;
        RECT 66.400 96.660 67.460 96.800 ;
        RECT 64.025 96.615 64.315 96.660 ;
        RECT 64.470 96.600 64.790 96.660 ;
        RECT 63.090 96.260 63.410 96.520 ;
        RECT 65.390 96.460 65.710 96.520 ;
        RECT 65.865 96.460 66.155 96.505 ;
        RECT 65.390 96.320 66.155 96.460 ;
        RECT 67.320 96.460 67.460 96.660 ;
        RECT 67.690 96.600 68.010 96.860 ;
        RECT 68.725 96.800 68.940 96.955 ;
        RECT 71.370 96.940 71.690 97.000 ;
        RECT 72.830 96.955 73.120 97.000 ;
        RECT 70.970 96.800 71.260 96.845 ;
        RECT 68.725 96.660 71.260 96.800 ;
        RECT 74.220 96.800 74.360 97.340 ;
        RECT 81.490 97.340 83.635 97.480 ;
        RECT 81.490 97.280 81.810 97.340 ;
        RECT 83.345 97.295 83.635 97.340 ;
        RECT 92.070 97.480 92.390 97.540 ;
        RECT 93.005 97.480 93.295 97.525 ;
        RECT 92.070 97.340 93.295 97.480 ;
        RECT 92.070 97.280 92.390 97.340 ;
        RECT 93.005 97.295 93.295 97.340 ;
        RECT 110.945 97.480 111.235 97.525 ;
        RECT 111.390 97.480 111.710 97.540 ;
        RECT 119.210 97.480 119.530 97.540 ;
        RECT 110.945 97.340 111.710 97.480 ;
        RECT 110.945 97.295 111.235 97.340 ;
        RECT 111.390 97.280 111.710 97.340 ;
        RECT 114.240 97.340 119.530 97.480 ;
        RECT 75.050 97.185 75.370 97.200 ;
        RECT 74.835 97.140 75.370 97.185 ;
        RECT 80.570 97.140 80.890 97.200 ;
        RECT 85.645 97.140 85.935 97.185 ;
        RECT 74.615 97.000 76.660 97.140 ;
        RECT 74.835 96.955 75.370 97.000 ;
        RECT 75.050 96.940 75.370 96.955 ;
        RECT 75.525 96.800 75.815 96.845 ;
        RECT 75.970 96.800 76.290 96.860 ;
        RECT 76.520 96.845 76.660 97.000 ;
        RECT 80.570 97.000 85.935 97.140 ;
        RECT 80.570 96.940 80.890 97.000 ;
        RECT 85.645 96.955 85.935 97.000 ;
        RECT 93.450 97.140 93.770 97.200 ;
        RECT 96.690 97.140 96.980 97.185 ;
        RECT 98.550 97.140 98.840 97.185 ;
        RECT 93.450 97.000 94.600 97.140 ;
        RECT 93.450 96.940 93.770 97.000 ;
        RECT 74.220 96.660 76.290 96.800 ;
        RECT 70.970 96.615 71.260 96.660 ;
        RECT 75.525 96.615 75.815 96.660 ;
        RECT 75.970 96.600 76.290 96.660 ;
        RECT 76.445 96.615 76.735 96.845 ;
        RECT 76.905 96.615 77.195 96.845 ;
        RECT 77.365 96.800 77.655 96.845 ;
        RECT 79.190 96.800 79.510 96.860 ;
        RECT 81.030 96.800 81.350 96.860 ;
        RECT 77.365 96.660 81.350 96.800 ;
        RECT 77.365 96.615 77.655 96.660 ;
        RECT 76.980 96.460 77.120 96.615 ;
        RECT 79.190 96.600 79.510 96.660 ;
        RECT 81.030 96.600 81.350 96.660 ;
        RECT 83.790 96.800 84.110 96.860 ;
        RECT 84.265 96.800 84.555 96.845 ;
        RECT 83.790 96.660 84.555 96.800 ;
        RECT 83.790 96.600 84.110 96.660 ;
        RECT 84.265 96.615 84.555 96.660 ;
        RECT 84.725 96.800 85.015 96.845 ;
        RECT 88.850 96.800 89.170 96.860 ;
        RECT 84.725 96.660 89.170 96.800 ;
        RECT 84.725 96.615 85.015 96.660 ;
        RECT 88.850 96.600 89.170 96.660 ;
        RECT 93.910 96.600 94.230 96.860 ;
        RECT 94.460 96.845 94.600 97.000 ;
        RECT 96.690 97.000 98.840 97.140 ;
        RECT 96.690 96.955 96.980 97.000 ;
        RECT 98.550 96.955 98.840 97.000 ;
        RECT 99.470 97.140 99.760 97.185 ;
        RECT 101.270 97.140 101.590 97.200 ;
        RECT 102.730 97.140 103.020 97.185 ;
        RECT 99.470 97.000 103.020 97.140 ;
        RECT 99.470 96.955 99.760 97.000 ;
        RECT 94.385 96.615 94.675 96.845 ;
        RECT 95.290 96.600 95.610 96.860 ;
        RECT 95.750 96.600 96.070 96.860 ;
        RECT 97.590 96.600 97.910 96.860 ;
        RECT 98.625 96.800 98.840 96.955 ;
        RECT 101.270 96.940 101.590 97.000 ;
        RECT 102.730 96.955 103.020 97.000 ;
        RECT 110.010 97.140 110.330 97.200 ;
        RECT 110.010 97.000 113.920 97.140 ;
        RECT 110.010 96.940 110.330 97.000 ;
        RECT 100.870 96.800 101.160 96.845 ;
        RECT 98.625 96.660 101.160 96.800 ;
        RECT 100.870 96.615 101.160 96.660 ;
        RECT 102.190 96.800 102.510 96.860 ;
        RECT 105.425 96.800 105.715 96.845 ;
        RECT 102.190 96.660 105.715 96.800 ;
        RECT 102.190 96.600 102.510 96.660 ;
        RECT 105.425 96.615 105.715 96.660 ;
        RECT 106.345 96.615 106.635 96.845 ;
        RECT 78.730 96.460 79.050 96.520 ;
        RECT 85.630 96.460 85.950 96.520 ;
        RECT 105.870 96.460 106.190 96.520 ;
        RECT 106.420 96.460 106.560 96.615 ;
        RECT 111.390 96.600 111.710 96.860 ;
        RECT 113.780 96.845 113.920 97.000 ;
        RECT 113.705 96.615 113.995 96.845 ;
        RECT 114.240 96.800 114.380 97.340 ;
        RECT 119.210 97.280 119.530 97.340 ;
        RECT 114.630 97.140 114.920 97.185 ;
        RECT 116.490 97.140 116.780 97.185 ;
        RECT 114.630 97.000 116.780 97.140 ;
        RECT 114.630 96.955 114.920 97.000 ;
        RECT 116.490 96.955 116.780 97.000 ;
        RECT 117.410 97.140 117.700 97.185 ;
        RECT 120.670 97.140 120.960 97.185 ;
        RECT 122.430 97.140 122.750 97.200 ;
        RECT 117.410 97.000 122.750 97.140 ;
        RECT 117.410 96.955 117.700 97.000 ;
        RECT 120.670 96.955 120.960 97.000 ;
        RECT 115.545 96.800 115.835 96.845 ;
        RECT 114.240 96.660 115.835 96.800 ;
        RECT 116.565 96.800 116.780 96.955 ;
        RECT 122.430 96.940 122.750 97.000 ;
        RECT 118.810 96.800 119.100 96.845 ;
        RECT 116.565 96.660 119.100 96.800 ;
        RECT 115.545 96.615 115.835 96.660 ;
        RECT 118.810 96.615 119.100 96.660 ;
        RECT 67.320 96.320 85.950 96.460 ;
        RECT 65.390 96.260 65.710 96.320 ;
        RECT 65.865 96.275 66.155 96.320 ;
        RECT 78.730 96.260 79.050 96.320 ;
        RECT 85.630 96.260 85.950 96.320 ;
        RECT 95.840 96.320 106.560 96.460 ;
        RECT 107.265 96.460 107.555 96.505 ;
        RECT 112.325 96.460 112.615 96.505 ;
        RECT 114.610 96.460 114.930 96.520 ;
        RECT 107.265 96.320 110.470 96.460 ;
        RECT 54.900 95.980 59.640 96.120 ;
        RECT 63.180 96.120 63.320 96.260 ;
        RECT 64.010 96.120 64.330 96.180 ;
        RECT 63.180 95.980 64.330 96.120 ;
        RECT 64.010 95.920 64.330 95.980 ;
        RECT 66.330 96.120 66.620 96.165 ;
        RECT 68.190 96.120 68.480 96.165 ;
        RECT 70.970 96.120 71.260 96.165 ;
        RECT 95.840 96.120 95.980 96.320 ;
        RECT 105.870 96.260 106.190 96.320 ;
        RECT 107.265 96.275 107.555 96.320 ;
        RECT 66.330 95.980 71.260 96.120 ;
        RECT 66.330 95.935 66.620 95.980 ;
        RECT 68.190 95.935 68.480 95.980 ;
        RECT 70.970 95.935 71.260 95.980 ;
        RECT 78.360 95.980 95.980 96.120 ;
        RECT 96.230 96.120 96.520 96.165 ;
        RECT 98.090 96.120 98.380 96.165 ;
        RECT 100.870 96.120 101.160 96.165 ;
        RECT 96.230 95.980 101.160 96.120 ;
        RECT 110.330 96.120 110.470 96.320 ;
        RECT 112.325 96.320 114.930 96.460 ;
        RECT 112.325 96.275 112.615 96.320 ;
        RECT 114.610 96.260 114.930 96.320 ;
        RECT 113.690 96.120 114.010 96.180 ;
        RECT 110.330 95.980 114.010 96.120 ;
        RECT 41.930 95.640 48.140 95.780 ;
        RECT 41.930 95.580 42.250 95.640 ;
        RECT 46.315 95.595 46.605 95.640 ;
        RECT 60.790 95.580 61.110 95.840 ;
        RECT 63.550 95.780 63.870 95.840 ;
        RECT 78.360 95.780 78.500 95.980 ;
        RECT 96.230 95.935 96.520 95.980 ;
        RECT 98.090 95.935 98.380 95.980 ;
        RECT 100.870 95.935 101.160 95.980 ;
        RECT 113.690 95.920 114.010 95.980 ;
        RECT 114.170 96.120 114.460 96.165 ;
        RECT 116.030 96.120 116.320 96.165 ;
        RECT 118.810 96.120 119.100 96.165 ;
        RECT 114.170 95.980 119.100 96.120 ;
        RECT 114.170 95.935 114.460 95.980 ;
        RECT 116.030 95.935 116.320 95.980 ;
        RECT 118.810 95.935 119.100 95.980 ;
        RECT 63.550 95.640 78.500 95.780 ;
        RECT 78.745 95.780 79.035 95.825 ;
        RECT 80.570 95.780 80.890 95.840 ;
        RECT 78.745 95.640 80.890 95.780 ;
        RECT 63.550 95.580 63.870 95.640 ;
        RECT 78.745 95.595 79.035 95.640 ;
        RECT 80.570 95.580 80.890 95.640 ;
        RECT 85.645 95.780 85.935 95.825 ;
        RECT 90.690 95.780 91.010 95.840 ;
        RECT 85.645 95.640 91.010 95.780 ;
        RECT 85.645 95.595 85.935 95.640 ;
        RECT 90.690 95.580 91.010 95.640 ;
        RECT 94.370 95.580 94.690 95.840 ;
        RECT 102.650 95.780 102.970 95.840 ;
        RECT 104.735 95.780 105.025 95.825 ;
        RECT 102.650 95.640 105.025 95.780 ;
        RECT 102.650 95.580 102.970 95.640 ;
        RECT 104.735 95.595 105.025 95.640 ;
        RECT 107.710 95.780 108.030 95.840 ;
        RECT 109.105 95.780 109.395 95.825 ;
        RECT 107.710 95.640 109.395 95.780 ;
        RECT 107.710 95.580 108.030 95.640 ;
        RECT 109.105 95.595 109.395 95.640 ;
        RECT 116.910 95.780 117.230 95.840 ;
        RECT 122.675 95.780 122.965 95.825 ;
        RECT 116.910 95.640 122.965 95.780 ;
        RECT 116.910 95.580 117.230 95.640 ;
        RECT 122.675 95.595 122.965 95.640 ;
        RECT 5.520 94.960 125.580 95.440 ;
        RECT 38.265 94.760 38.555 94.805 ;
        RECT 38.710 94.760 39.030 94.820 ;
        RECT 38.265 94.620 39.030 94.760 ;
        RECT 38.265 94.575 38.555 94.620 ;
        RECT 38.710 94.560 39.030 94.620 ;
        RECT 42.850 94.560 43.170 94.820 ;
        RECT 46.530 94.760 46.850 94.820 ;
        RECT 56.665 94.760 56.955 94.805 ;
        RECT 46.530 94.620 56.955 94.760 ;
        RECT 46.530 94.560 46.850 94.620 ;
        RECT 56.665 94.575 56.955 94.620 ;
        RECT 57.570 94.560 57.890 94.820 ;
        RECT 73.210 94.760 73.530 94.820 ;
        RECT 74.145 94.760 74.435 94.805 ;
        RECT 73.210 94.620 74.435 94.760 ;
        RECT 73.210 94.560 73.530 94.620 ;
        RECT 74.145 94.575 74.435 94.620 ;
        RECT 76.430 94.760 76.750 94.820 ;
        RECT 78.285 94.760 78.575 94.805 ;
        RECT 76.430 94.620 78.575 94.760 ;
        RECT 76.430 94.560 76.750 94.620 ;
        RECT 78.285 94.575 78.575 94.620 ;
        RECT 80.585 94.760 80.875 94.805 ;
        RECT 82.870 94.760 83.190 94.820 ;
        RECT 80.585 94.620 83.190 94.760 ;
        RECT 80.585 94.575 80.875 94.620 ;
        RECT 82.870 94.560 83.190 94.620 ;
        RECT 87.485 94.760 87.775 94.805 ;
        RECT 95.290 94.760 95.610 94.820 ;
        RECT 87.485 94.620 95.610 94.760 ;
        RECT 87.485 94.575 87.775 94.620 ;
        RECT 95.290 94.560 95.610 94.620 ;
        RECT 97.605 94.760 97.895 94.805 ;
        RECT 98.050 94.760 98.370 94.820 ;
        RECT 97.605 94.620 98.370 94.760 ;
        RECT 97.605 94.575 97.895 94.620 ;
        RECT 98.050 94.560 98.370 94.620 ;
        RECT 106.805 94.760 107.095 94.805 ;
        RECT 107.250 94.760 107.570 94.820 ;
        RECT 106.805 94.620 107.570 94.760 ;
        RECT 106.805 94.575 107.095 94.620 ;
        RECT 107.250 94.560 107.570 94.620 ;
        RECT 9.290 94.420 9.580 94.465 ;
        RECT 11.150 94.420 11.440 94.465 ;
        RECT 13.930 94.420 14.220 94.465 ;
        RECT 9.290 94.280 14.220 94.420 ;
        RECT 9.290 94.235 9.580 94.280 ;
        RECT 11.150 94.235 11.440 94.280 ;
        RECT 13.930 94.235 14.220 94.280 ;
        RECT 27.225 94.235 27.515 94.465 ;
        RECT 28.150 94.420 28.440 94.465 ;
        RECT 30.010 94.420 30.300 94.465 ;
        RECT 32.790 94.420 33.080 94.465 ;
        RECT 28.150 94.280 33.080 94.420 ;
        RECT 28.150 94.235 28.440 94.280 ;
        RECT 30.010 94.235 30.300 94.280 ;
        RECT 32.790 94.235 33.080 94.280 ;
        RECT 58.950 94.420 59.270 94.480 ;
        RECT 65.405 94.420 65.695 94.465 ;
        RECT 74.590 94.420 74.910 94.480 ;
        RECT 58.950 94.280 65.695 94.420 ;
        RECT 7.430 94.080 7.750 94.140 ;
        RECT 8.825 94.080 9.115 94.125 ;
        RECT 11.570 94.080 11.890 94.140 ;
        RECT 7.430 93.940 11.890 94.080 ;
        RECT 27.300 94.080 27.440 94.235 ;
        RECT 58.950 94.220 59.270 94.280 ;
        RECT 65.405 94.235 65.695 94.280 ;
        RECT 71.460 94.280 74.910 94.420 ;
        RECT 29.525 94.080 29.815 94.125 ;
        RECT 27.300 93.940 29.815 94.080 ;
        RECT 7.430 93.880 7.750 93.940 ;
        RECT 8.825 93.895 9.115 93.940 ;
        RECT 11.570 93.880 11.890 93.940 ;
        RECT 29.525 93.895 29.815 93.940 ;
        RECT 39.170 94.080 39.490 94.140 ;
        RECT 41.025 94.080 41.315 94.125 ;
        RECT 39.170 93.940 41.315 94.080 ;
        RECT 39.170 93.880 39.490 93.940 ;
        RECT 41.025 93.895 41.315 93.940 ;
        RECT 58.505 94.080 58.795 94.125 ;
        RECT 60.330 94.080 60.650 94.140 ;
        RECT 58.505 93.940 60.650 94.080 ;
        RECT 58.505 93.895 58.795 93.940 ;
        RECT 60.330 93.880 60.650 93.940 ;
        RECT 10.665 93.740 10.955 93.785 ;
        RECT 11.110 93.740 11.430 93.800 ;
        RECT 13.930 93.740 14.220 93.785 ;
        RECT 10.665 93.600 11.430 93.740 ;
        RECT 10.665 93.555 10.955 93.600 ;
        RECT 11.110 93.540 11.430 93.600 ;
        RECT 11.685 93.600 14.220 93.740 ;
        RECT 11.685 93.445 11.900 93.600 ;
        RECT 13.930 93.555 14.220 93.600 ;
        RECT 26.305 93.555 26.595 93.785 ;
        RECT 9.750 93.400 10.040 93.445 ;
        RECT 11.610 93.400 11.900 93.445 ;
        RECT 9.750 93.260 11.900 93.400 ;
        RECT 9.750 93.215 10.040 93.260 ;
        RECT 11.610 93.215 11.900 93.260 ;
        RECT 12.530 93.400 12.820 93.445 ;
        RECT 15.790 93.400 16.080 93.445 ;
        RECT 21.690 93.400 22.010 93.460 ;
        RECT 12.530 93.260 22.010 93.400 ;
        RECT 12.530 93.215 12.820 93.260 ;
        RECT 15.790 93.215 16.080 93.260 ;
        RECT 21.690 93.200 22.010 93.260 ;
        RECT 17.795 93.060 18.085 93.105 ;
        RECT 20.770 93.060 21.090 93.120 ;
        RECT 17.795 92.920 21.090 93.060 ;
        RECT 26.380 93.060 26.520 93.555 ;
        RECT 27.670 93.540 27.990 93.800 ;
        RECT 32.790 93.740 33.080 93.785 ;
        RECT 30.545 93.600 33.080 93.740 ;
        RECT 30.545 93.445 30.760 93.600 ;
        RECT 32.790 93.555 33.080 93.600 ;
        RECT 40.565 93.740 40.855 93.785 ;
        RECT 41.930 93.740 42.250 93.800 ;
        RECT 40.565 93.600 42.250 93.740 ;
        RECT 40.565 93.555 40.855 93.600 ;
        RECT 41.930 93.540 42.250 93.600 ;
        RECT 43.310 93.540 43.630 93.800 ;
        RECT 57.570 93.540 57.890 93.800 ;
        RECT 58.965 93.740 59.255 93.785 ;
        RECT 60.790 93.740 61.110 93.800 ;
        RECT 58.965 93.600 61.110 93.740 ;
        RECT 58.965 93.555 59.255 93.600 ;
        RECT 60.790 93.540 61.110 93.600 ;
        RECT 28.610 93.400 28.900 93.445 ;
        RECT 30.470 93.400 30.760 93.445 ;
        RECT 28.610 93.260 30.760 93.400 ;
        RECT 28.610 93.215 28.900 93.260 ;
        RECT 30.470 93.215 30.760 93.260 ;
        RECT 31.390 93.400 31.680 93.445 ;
        RECT 33.190 93.400 33.510 93.460 ;
        RECT 34.650 93.400 34.940 93.445 ;
        RECT 31.390 93.260 34.940 93.400 ;
        RECT 31.390 93.215 31.680 93.260 ;
        RECT 33.190 93.200 33.510 93.260 ;
        RECT 34.650 93.215 34.940 93.260 ;
        RECT 64.470 93.200 64.790 93.460 ;
        RECT 65.480 93.400 65.620 94.235 ;
        RECT 71.460 94.125 71.600 94.280 ;
        RECT 74.590 94.220 74.910 94.280 ;
        RECT 71.385 93.895 71.675 94.125 ;
        RECT 71.845 94.080 72.135 94.125 ;
        RECT 75.050 94.080 75.370 94.140 ;
        RECT 71.845 93.940 75.370 94.080 ;
        RECT 71.845 93.895 72.135 93.940 ;
        RECT 75.050 93.880 75.370 93.940 ;
        RECT 80.110 93.880 80.430 94.140 ;
        RECT 81.030 94.080 81.350 94.140 ;
        RECT 98.970 94.080 99.290 94.140 ;
        RECT 100.365 94.080 100.655 94.125 ;
        RECT 81.030 93.940 86.320 94.080 ;
        RECT 81.030 93.880 81.350 93.940 ;
        RECT 79.190 93.540 79.510 93.800 ;
        RECT 80.570 93.540 80.890 93.800 ;
        RECT 82.410 93.740 82.730 93.800 ;
        RECT 84.265 93.740 84.555 93.785 ;
        RECT 82.410 93.600 84.555 93.740 ;
        RECT 82.410 93.540 82.730 93.600 ;
        RECT 84.265 93.555 84.555 93.600 ;
        RECT 85.185 93.555 85.475 93.785 ;
        RECT 85.260 93.400 85.400 93.555 ;
        RECT 85.630 93.540 85.950 93.800 ;
        RECT 86.180 93.785 86.320 93.940 ;
        RECT 98.970 93.940 100.655 94.080 ;
        RECT 98.970 93.880 99.290 93.940 ;
        RECT 100.365 93.895 100.655 93.940 ;
        RECT 86.105 93.555 86.395 93.785 ;
        RECT 94.385 93.740 94.675 93.785 ;
        RECT 94.830 93.740 95.150 93.800 ;
        RECT 87.560 93.600 95.150 93.740 ;
        RECT 86.550 93.400 86.870 93.460 ;
        RECT 65.480 93.260 84.940 93.400 ;
        RECT 85.260 93.260 86.870 93.400 ;
        RECT 31.810 93.060 32.130 93.120 ;
        RECT 26.380 92.920 32.130 93.060 ;
        RECT 17.795 92.875 18.085 92.920 ;
        RECT 20.770 92.860 21.090 92.920 ;
        RECT 31.810 92.860 32.130 92.920 ;
        RECT 35.490 93.060 35.810 93.120 ;
        RECT 36.655 93.060 36.945 93.105 ;
        RECT 40.105 93.060 40.395 93.105 ;
        RECT 35.490 92.920 40.395 93.060 ;
        RECT 35.490 92.860 35.810 92.920 ;
        RECT 36.655 92.875 36.945 92.920 ;
        RECT 40.105 92.875 40.395 92.920 ;
        RECT 56.190 93.060 56.510 93.120 ;
        RECT 58.950 93.060 59.270 93.120 ;
        RECT 60.790 93.060 61.110 93.120 ;
        RECT 56.190 92.920 61.110 93.060 ;
        RECT 56.190 92.860 56.510 92.920 ;
        RECT 58.950 92.860 59.270 92.920 ;
        RECT 60.790 92.860 61.110 92.920 ;
        RECT 72.305 93.060 72.595 93.105 ;
        RECT 74.590 93.060 74.910 93.120 ;
        RECT 72.305 92.920 74.910 93.060 ;
        RECT 84.800 93.060 84.940 93.260 ;
        RECT 86.550 93.200 86.870 93.260 ;
        RECT 87.560 93.060 87.700 93.600 ;
        RECT 94.385 93.555 94.675 93.600 ;
        RECT 94.830 93.540 95.150 93.600 ;
        RECT 95.305 93.740 95.595 93.785 ;
        RECT 99.905 93.740 100.195 93.785 ;
        RECT 101.730 93.740 102.050 93.800 ;
        RECT 95.305 93.600 102.050 93.740 ;
        RECT 95.305 93.555 95.595 93.600 ;
        RECT 99.905 93.555 100.195 93.600 ;
        RECT 101.730 93.540 102.050 93.600 ;
        RECT 107.710 93.540 108.030 93.800 ;
        RECT 118.750 93.540 119.070 93.800 ;
        RECT 99.445 93.400 99.735 93.445 ;
        RECT 102.650 93.400 102.970 93.460 ;
        RECT 99.445 93.260 102.970 93.400 ;
        RECT 99.445 93.215 99.735 93.260 ;
        RECT 102.650 93.200 102.970 93.260 ;
        RECT 84.800 92.920 87.700 93.060 ;
        RECT 87.930 93.060 88.250 93.120 ;
        RECT 93.465 93.060 93.755 93.105 ;
        RECT 87.930 92.920 93.755 93.060 ;
        RECT 72.305 92.875 72.595 92.920 ;
        RECT 74.590 92.860 74.910 92.920 ;
        RECT 87.930 92.860 88.250 92.920 ;
        RECT 93.465 92.875 93.755 92.920 ;
        RECT 118.290 92.860 118.610 93.120 ;
        RECT 5.520 92.240 125.580 92.720 ;
        RECT 17.090 91.840 17.410 92.100 ;
        RECT 19.405 92.040 19.695 92.085 ;
        RECT 20.770 92.040 21.090 92.100 ;
        RECT 19.405 91.900 21.090 92.040 ;
        RECT 19.405 91.855 19.695 91.900 ;
        RECT 20.770 91.840 21.090 91.900 ;
        RECT 21.690 91.840 22.010 92.100 ;
        RECT 23.990 92.040 24.310 92.100 ;
        RECT 25.370 92.040 25.690 92.100 ;
        RECT 23.990 91.900 25.690 92.040 ;
        RECT 23.990 91.840 24.310 91.900 ;
        RECT 25.370 91.840 25.690 91.900 ;
        RECT 26.765 92.040 27.055 92.085 ;
        RECT 27.210 92.040 27.530 92.100 ;
        RECT 26.765 91.900 27.530 92.040 ;
        RECT 26.765 91.855 27.055 91.900 ;
        RECT 27.210 91.840 27.530 91.900 ;
        RECT 28.590 91.840 28.910 92.100 ;
        RECT 31.810 91.840 32.130 92.100 ;
        RECT 34.125 92.040 34.415 92.085 ;
        RECT 34.570 92.040 34.890 92.100 ;
        RECT 35.490 92.040 35.810 92.100 ;
        RECT 34.125 91.900 35.810 92.040 ;
        RECT 34.125 91.855 34.415 91.900 ;
        RECT 34.570 91.840 34.890 91.900 ;
        RECT 35.490 91.840 35.810 91.900 ;
        RECT 58.490 92.040 58.810 92.100 ;
        RECT 59.885 92.040 60.175 92.085 ;
        RECT 58.490 91.900 60.175 92.040 ;
        RECT 58.490 91.840 58.810 91.900 ;
        RECT 59.885 91.855 60.175 91.900 ;
        RECT 74.590 91.840 74.910 92.100 ;
        RECT 86.550 92.040 86.870 92.100 ;
        RECT 89.310 92.040 89.630 92.100 ;
        RECT 86.550 91.900 89.630 92.040 ;
        RECT 86.550 91.840 86.870 91.900 ;
        RECT 89.310 91.840 89.630 91.900 ;
        RECT 8.370 91.700 8.660 91.745 ;
        RECT 10.230 91.700 10.520 91.745 ;
        RECT 8.370 91.560 10.520 91.700 ;
        RECT 8.370 91.515 8.660 91.560 ;
        RECT 10.230 91.515 10.520 91.560 ;
        RECT 11.150 91.700 11.440 91.745 ;
        RECT 12.950 91.700 13.270 91.760 ;
        RECT 14.410 91.700 14.700 91.745 ;
        RECT 11.150 91.560 14.700 91.700 ;
        RECT 20.860 91.700 21.000 91.840 ;
        RECT 33.665 91.700 33.955 91.745 ;
        RECT 20.860 91.560 33.955 91.700 ;
        RECT 11.150 91.515 11.440 91.560 ;
        RECT 7.430 91.160 7.750 91.420 ;
        RECT 10.305 91.360 10.520 91.515 ;
        RECT 12.950 91.500 13.270 91.560 ;
        RECT 14.410 91.515 14.700 91.560 ;
        RECT 33.665 91.515 33.955 91.560 ;
        RECT 63.550 91.500 63.870 91.760 ;
        RECT 64.470 91.700 64.790 91.760 ;
        RECT 68.150 91.700 68.470 91.760 ;
        RECT 64.470 91.560 68.470 91.700 ;
        RECT 64.470 91.500 64.790 91.560 ;
        RECT 68.150 91.500 68.470 91.560 ;
        RECT 69.065 91.700 69.715 91.745 ;
        RECT 72.665 91.700 72.955 91.745 ;
        RECT 75.050 91.700 75.370 91.760 ;
        RECT 69.065 91.560 75.370 91.700 ;
        RECT 69.065 91.515 69.715 91.560 ;
        RECT 72.365 91.515 72.955 91.560 ;
        RECT 12.550 91.360 12.840 91.405 ;
        RECT 10.305 91.220 12.840 91.360 ;
        RECT 12.550 91.175 12.840 91.220 ;
        RECT 16.415 91.360 16.705 91.405 ;
        RECT 18.930 91.360 19.250 91.420 ;
        RECT 16.415 91.220 19.250 91.360 ;
        RECT 16.415 91.175 16.705 91.220 ;
        RECT 18.930 91.160 19.250 91.220 ;
        RECT 20.310 91.360 20.630 91.420 ;
        RECT 22.165 91.360 22.455 91.405 ;
        RECT 20.310 91.220 22.455 91.360 ;
        RECT 20.310 91.160 20.630 91.220 ;
        RECT 22.165 91.175 22.455 91.220 ;
        RECT 24.450 91.160 24.770 91.420 ;
        RECT 25.845 91.360 26.135 91.405 ;
        RECT 27.210 91.360 27.530 91.420 ;
        RECT 25.845 91.220 27.530 91.360 ;
        RECT 25.845 91.175 26.135 91.220 ;
        RECT 27.210 91.160 27.530 91.220 ;
        RECT 29.510 91.160 29.830 91.420 ;
        RECT 30.890 91.160 31.210 91.420 ;
        RECT 57.570 91.160 57.890 91.420 ;
        RECT 58.950 91.160 59.270 91.420 ;
        RECT 65.390 91.160 65.710 91.420 ;
        RECT 65.870 91.360 66.160 91.405 ;
        RECT 67.705 91.360 67.995 91.405 ;
        RECT 71.285 91.360 71.575 91.405 ;
        RECT 65.870 91.220 71.575 91.360 ;
        RECT 65.870 91.175 66.160 91.220 ;
        RECT 67.705 91.175 67.995 91.220 ;
        RECT 71.285 91.175 71.575 91.220 ;
        RECT 72.365 91.200 72.655 91.515 ;
        RECT 75.050 91.500 75.370 91.560 ;
        RECT 78.730 91.700 79.050 91.760 ;
        RECT 81.505 91.700 81.795 91.745 ;
        RECT 85.645 91.700 85.935 91.745 ;
        RECT 78.730 91.560 79.880 91.700 ;
        RECT 78.730 91.500 79.050 91.560 ;
        RECT 75.970 91.360 76.290 91.420 ;
        RECT 79.740 91.405 79.880 91.560 ;
        RECT 81.505 91.560 85.935 91.700 ;
        RECT 81.505 91.515 81.795 91.560 ;
        RECT 85.645 91.515 85.935 91.560 ;
        RECT 78.285 91.360 78.575 91.405 ;
        RECT 75.970 91.220 78.575 91.360 ;
        RECT 75.970 91.160 76.290 91.220 ;
        RECT 78.285 91.175 78.575 91.220 ;
        RECT 79.205 91.175 79.495 91.405 ;
        RECT 79.665 91.175 79.955 91.405 ;
        RECT 80.125 91.360 80.415 91.405 ;
        RECT 80.570 91.360 80.890 91.420 ;
        RECT 80.125 91.220 80.890 91.360 ;
        RECT 80.125 91.175 80.415 91.220 ;
        RECT 8.810 91.020 9.130 91.080 ;
        RECT 9.285 91.020 9.575 91.065 ;
        RECT 8.810 90.880 9.575 91.020 ;
        RECT 8.810 90.820 9.130 90.880 ;
        RECT 9.285 90.835 9.575 90.880 ;
        RECT 17.090 91.020 17.410 91.080 ;
        RECT 19.865 91.020 20.155 91.065 ;
        RECT 17.090 90.880 20.155 91.020 ;
        RECT 17.090 90.820 17.410 90.880 ;
        RECT 19.865 90.835 20.155 90.880 ;
        RECT 7.910 90.680 8.200 90.725 ;
        RECT 9.770 90.680 10.060 90.725 ;
        RECT 12.550 90.680 12.840 90.725 ;
        RECT 7.910 90.540 12.840 90.680 ;
        RECT 7.910 90.495 8.200 90.540 ;
        RECT 9.770 90.495 10.060 90.540 ;
        RECT 12.550 90.495 12.840 90.540 ;
        RECT 19.940 90.340 20.080 90.835 ;
        RECT 24.910 90.820 25.230 91.080 ;
        RECT 30.430 90.820 30.750 91.080 ;
        RECT 34.585 90.835 34.875 91.065 ;
        RECT 25.370 90.680 25.690 90.740 ;
        RECT 26.290 90.680 26.610 90.740 ;
        RECT 34.660 90.680 34.800 90.835 ;
        RECT 58.490 90.820 58.810 91.080 ;
        RECT 66.770 90.820 67.090 91.080 ;
        RECT 74.145 91.020 74.435 91.065 ;
        RECT 77.365 91.020 77.655 91.065 ;
        RECT 79.280 91.020 79.420 91.175 ;
        RECT 80.570 91.160 80.890 91.220 ;
        RECT 83.330 91.360 83.650 91.420 ;
        RECT 84.265 91.360 84.555 91.405 ;
        RECT 92.545 91.360 92.835 91.405 ;
        RECT 83.330 91.220 84.555 91.360 ;
        RECT 83.330 91.160 83.650 91.220 ;
        RECT 84.265 91.175 84.555 91.220 ;
        RECT 91.240 91.220 92.835 91.360 ;
        RECT 74.145 90.880 79.420 91.020 ;
        RECT 85.185 91.020 85.475 91.065 ;
        RECT 86.550 91.020 86.870 91.080 ;
        RECT 85.185 90.880 86.870 91.020 ;
        RECT 74.145 90.835 74.435 90.880 ;
        RECT 77.365 90.835 77.655 90.880 ;
        RECT 85.185 90.835 85.475 90.880 ;
        RECT 86.550 90.820 86.870 90.880 ;
        RECT 87.945 90.835 88.235 91.065 ;
        RECT 88.865 91.020 89.155 91.065 ;
        RECT 90.690 91.020 91.010 91.080 ;
        RECT 88.865 90.880 91.010 91.020 ;
        RECT 88.865 90.835 89.155 90.880 ;
        RECT 39.170 90.680 39.490 90.740 ;
        RECT 52.050 90.680 52.370 90.740 ;
        RECT 25.370 90.540 26.060 90.680 ;
        RECT 25.370 90.480 25.690 90.540 ;
        RECT 24.910 90.340 25.230 90.400 ;
        RECT 25.920 90.385 26.060 90.540 ;
        RECT 26.290 90.540 52.370 90.680 ;
        RECT 26.290 90.480 26.610 90.540 ;
        RECT 39.170 90.480 39.490 90.540 ;
        RECT 52.050 90.480 52.370 90.540 ;
        RECT 66.275 90.680 66.565 90.725 ;
        RECT 68.165 90.680 68.455 90.725 ;
        RECT 71.285 90.680 71.575 90.725 ;
        RECT 66.275 90.540 71.575 90.680 ;
        RECT 66.275 90.495 66.565 90.540 ;
        RECT 68.165 90.495 68.455 90.540 ;
        RECT 71.285 90.495 71.575 90.540 ;
        RECT 75.510 90.680 75.830 90.740 ;
        RECT 88.020 90.680 88.160 90.835 ;
        RECT 90.690 90.820 91.010 90.880 ;
        RECT 91.240 90.725 91.380 91.220 ;
        RECT 92.545 91.175 92.835 91.220 ;
        RECT 93.925 91.360 94.215 91.405 ;
        RECT 94.370 91.360 94.690 91.420 ;
        RECT 96.210 91.360 96.530 91.420 ;
        RECT 93.925 91.220 96.530 91.360 ;
        RECT 93.925 91.175 94.215 91.220 ;
        RECT 94.370 91.160 94.690 91.220 ;
        RECT 96.210 91.160 96.530 91.220 ;
        RECT 116.005 91.360 116.295 91.405 ;
        RECT 117.370 91.360 117.690 91.420 ;
        RECT 119.685 91.360 119.975 91.405 ;
        RECT 116.005 91.220 119.975 91.360 ;
        RECT 116.005 91.175 116.295 91.220 ;
        RECT 117.370 91.160 117.690 91.220 ;
        RECT 119.685 91.175 119.975 91.220 ;
        RECT 120.145 91.360 120.435 91.405 ;
        RECT 120.590 91.360 120.910 91.420 ;
        RECT 120.145 91.220 120.910 91.360 ;
        RECT 120.145 91.175 120.435 91.220 ;
        RECT 120.590 91.160 120.910 91.220 ;
        RECT 110.930 91.020 111.250 91.080 ;
        RECT 116.450 91.020 116.770 91.080 ;
        RECT 110.930 90.880 116.770 91.020 ;
        RECT 110.930 90.820 111.250 90.880 ;
        RECT 116.450 90.820 116.770 90.880 ;
        RECT 116.925 91.020 117.215 91.065 ;
        RECT 118.765 91.020 119.055 91.065 ;
        RECT 116.925 90.880 119.055 91.020 ;
        RECT 116.925 90.835 117.215 90.880 ;
        RECT 118.765 90.835 119.055 90.880 ;
        RECT 75.510 90.540 88.160 90.680 ;
        RECT 75.510 90.480 75.830 90.540 ;
        RECT 91.165 90.495 91.455 90.725 ;
        RECT 114.610 90.680 114.930 90.740 ;
        RECT 117.000 90.680 117.140 90.835 ;
        RECT 114.610 90.540 117.140 90.680 ;
        RECT 114.610 90.480 114.930 90.540 ;
        RECT 19.940 90.200 25.230 90.340 ;
        RECT 24.910 90.140 25.230 90.200 ;
        RECT 25.845 90.155 26.135 90.385 ;
        RECT 29.970 90.140 30.290 90.400 ;
        RECT 58.965 90.340 59.255 90.385 ;
        RECT 59.410 90.340 59.730 90.400 ;
        RECT 58.965 90.200 59.730 90.340 ;
        RECT 58.965 90.155 59.255 90.200 ;
        RECT 59.410 90.140 59.730 90.200 ;
        RECT 68.610 90.340 68.930 90.400 ;
        RECT 83.345 90.340 83.635 90.385 ;
        RECT 68.610 90.200 83.635 90.340 ;
        RECT 68.610 90.140 68.930 90.200 ;
        RECT 83.345 90.155 83.635 90.200 ;
        RECT 85.645 90.340 85.935 90.385 ;
        RECT 87.930 90.340 88.250 90.400 ;
        RECT 85.645 90.200 88.250 90.340 ;
        RECT 85.645 90.155 85.935 90.200 ;
        RECT 87.930 90.140 88.250 90.200 ;
        RECT 91.610 90.140 91.930 90.400 ;
        RECT 92.990 90.340 93.310 90.400 ;
        RECT 93.465 90.340 93.755 90.385 ;
        RECT 92.990 90.200 93.755 90.340 ;
        RECT 92.990 90.140 93.310 90.200 ;
        RECT 93.465 90.155 93.755 90.200 ;
        RECT 110.470 90.340 110.790 90.400 ;
        RECT 114.165 90.340 114.455 90.385 ;
        RECT 110.470 90.200 114.455 90.340 ;
        RECT 110.470 90.140 110.790 90.200 ;
        RECT 114.165 90.155 114.455 90.200 ;
        RECT 121.985 90.340 122.275 90.385 ;
        RECT 122.890 90.340 123.210 90.400 ;
        RECT 121.985 90.200 123.210 90.340 ;
        RECT 121.985 90.155 122.275 90.200 ;
        RECT 122.890 90.140 123.210 90.200 ;
        RECT 5.520 89.520 125.580 90.000 ;
        RECT 8.810 89.320 9.130 89.380 ;
        RECT 10.665 89.320 10.955 89.365 ;
        RECT 8.810 89.180 10.955 89.320 ;
        RECT 8.810 89.120 9.130 89.180 ;
        RECT 10.665 89.135 10.955 89.180 ;
        RECT 12.950 89.120 13.270 89.380 ;
        RECT 24.450 89.120 24.770 89.380 ;
        RECT 29.065 89.320 29.355 89.365 ;
        RECT 30.890 89.320 31.210 89.380 ;
        RECT 29.065 89.180 31.210 89.320 ;
        RECT 29.065 89.135 29.355 89.180 ;
        RECT 30.890 89.120 31.210 89.180 ;
        RECT 38.250 89.120 38.570 89.380 ;
        RECT 57.570 89.120 57.890 89.380 ;
        RECT 66.770 89.320 67.090 89.380 ;
        RECT 67.705 89.320 67.995 89.365 ;
        RECT 66.770 89.180 67.995 89.320 ;
        RECT 66.770 89.120 67.090 89.180 ;
        RECT 67.705 89.135 67.995 89.180 ;
        RECT 75.050 89.120 75.370 89.380 ;
        RECT 90.690 89.320 91.010 89.380 ;
        RECT 92.530 89.320 92.850 89.380 ;
        RECT 95.075 89.320 95.365 89.365 ;
        RECT 111.390 89.320 111.710 89.380 ;
        RECT 90.690 89.180 95.365 89.320 ;
        RECT 90.690 89.120 91.010 89.180 ;
        RECT 92.530 89.120 92.850 89.180 ;
        RECT 95.075 89.135 95.365 89.180 ;
        RECT 109.180 89.180 117.600 89.320 ;
        RECT 35.950 88.980 36.270 89.040 ;
        RECT 39.645 88.980 39.935 89.025 ;
        RECT 53.445 88.980 53.735 89.025 ;
        RECT 61.710 88.980 62.030 89.040 ;
        RECT 35.950 88.840 39.935 88.980 ;
        RECT 35.950 88.780 36.270 88.840 ;
        RECT 39.645 88.795 39.935 88.840 ;
        RECT 46.160 88.840 53.735 88.980 ;
        RECT 17.090 88.440 17.410 88.700 ;
        RECT 20.770 88.640 21.090 88.700 ;
        RECT 36.410 88.640 36.730 88.700 ;
        RECT 37.805 88.640 38.095 88.685 ;
        RECT 20.770 88.500 26.980 88.640 ;
        RECT 20.770 88.440 21.090 88.500 ;
        RECT 11.585 88.115 11.875 88.345 ;
        RECT 13.425 88.300 13.715 88.345 ;
        RECT 18.010 88.300 18.330 88.360 ;
        RECT 20.310 88.300 20.630 88.360 ;
        RECT 13.425 88.160 20.630 88.300 ;
        RECT 13.425 88.115 13.715 88.160 ;
        RECT 11.660 87.960 11.800 88.115 ;
        RECT 18.010 88.100 18.330 88.160 ;
        RECT 20.310 88.100 20.630 88.160 ;
        RECT 21.245 88.300 21.535 88.345 ;
        RECT 21.690 88.300 22.010 88.360 ;
        RECT 21.245 88.160 22.010 88.300 ;
        RECT 21.245 88.115 21.535 88.160 ;
        RECT 21.690 88.100 22.010 88.160 ;
        RECT 22.165 88.115 22.455 88.345 ;
        RECT 22.625 88.115 22.915 88.345 ;
        RECT 23.085 88.300 23.375 88.345 ;
        RECT 23.990 88.300 24.310 88.360 ;
        RECT 23.085 88.160 24.310 88.300 ;
        RECT 23.085 88.115 23.375 88.160 ;
        RECT 16.185 87.960 16.475 88.005 ;
        RECT 18.930 87.960 19.250 88.020 ;
        RECT 22.240 87.960 22.380 88.115 ;
        RECT 11.660 87.820 14.100 87.960 ;
        RECT 13.960 87.665 14.100 87.820 ;
        RECT 16.185 87.820 22.380 87.960 ;
        RECT 22.700 87.960 22.840 88.115 ;
        RECT 23.990 88.100 24.310 88.160 ;
        RECT 25.830 88.100 26.150 88.360 ;
        RECT 26.840 88.345 26.980 88.500 ;
        RECT 36.410 88.500 38.095 88.640 ;
        RECT 36.410 88.440 36.730 88.500 ;
        RECT 37.805 88.455 38.095 88.500 ;
        RECT 26.765 88.115 27.055 88.345 ;
        RECT 27.240 88.115 27.530 88.345 ;
        RECT 27.685 88.300 27.975 88.345 ;
        RECT 28.590 88.300 28.910 88.360 ;
        RECT 27.685 88.160 28.910 88.300 ;
        RECT 27.685 88.115 27.975 88.160 ;
        RECT 27.300 87.960 27.440 88.115 ;
        RECT 28.590 88.100 28.910 88.160 ;
        RECT 33.650 88.100 33.970 88.360 ;
        RECT 34.570 88.100 34.890 88.360 ;
        RECT 35.045 88.115 35.335 88.345 ;
        RECT 29.050 87.960 29.370 88.020 ;
        RECT 35.120 87.960 35.260 88.115 ;
        RECT 35.490 88.100 35.810 88.360 ;
        RECT 38.710 88.100 39.030 88.360 ;
        RECT 46.160 88.345 46.300 88.840 ;
        RECT 53.445 88.795 53.735 88.840 ;
        RECT 59.040 88.840 62.030 88.980 ;
        RECT 47.910 88.640 48.230 88.700 ;
        RECT 51.605 88.640 51.895 88.685 ;
        RECT 47.910 88.500 51.895 88.640 ;
        RECT 47.910 88.440 48.230 88.500 ;
        RECT 51.605 88.455 51.895 88.500 ;
        RECT 52.050 88.640 52.370 88.700 ;
        RECT 56.205 88.640 56.495 88.685 ;
        RECT 52.050 88.500 56.495 88.640 ;
        RECT 52.050 88.440 52.370 88.500 ;
        RECT 56.205 88.455 56.495 88.500 ;
        RECT 46.085 88.115 46.375 88.345 ;
        RECT 48.385 88.300 48.675 88.345 ;
        RECT 55.285 88.300 55.575 88.345 ;
        RECT 56.650 88.300 56.970 88.360 ;
        RECT 48.385 88.160 49.520 88.300 ;
        RECT 48.385 88.115 48.675 88.160 ;
        RECT 22.700 87.820 35.260 87.960 ;
        RECT 16.185 87.775 16.475 87.820 ;
        RECT 18.930 87.760 19.250 87.820 ;
        RECT 29.050 87.760 29.370 87.820 ;
        RECT 13.885 87.435 14.175 87.665 ;
        RECT 15.710 87.420 16.030 87.680 ;
        RECT 21.690 87.620 22.010 87.680 ;
        RECT 23.070 87.620 23.390 87.680 ;
        RECT 25.830 87.620 26.150 87.680 ;
        RECT 33.650 87.620 33.970 87.680 ;
        RECT 21.690 87.480 33.970 87.620 ;
        RECT 35.120 87.620 35.260 87.820 ;
        RECT 36.885 87.960 37.175 88.005 ;
        RECT 37.345 87.960 37.635 88.005 ;
        RECT 36.885 87.820 37.635 87.960 ;
        RECT 36.885 87.775 37.175 87.820 ;
        RECT 37.345 87.775 37.635 87.820 ;
        RECT 41.930 87.620 42.250 87.680 ;
        RECT 35.120 87.480 42.250 87.620 ;
        RECT 21.690 87.420 22.010 87.480 ;
        RECT 23.070 87.420 23.390 87.480 ;
        RECT 25.830 87.420 26.150 87.480 ;
        RECT 33.650 87.420 33.970 87.480 ;
        RECT 41.930 87.420 42.250 87.480 ;
        RECT 46.990 87.420 47.310 87.680 ;
        RECT 47.450 87.420 47.770 87.680 ;
        RECT 49.380 87.665 49.520 88.160 ;
        RECT 55.285 88.160 56.970 88.300 ;
        RECT 55.285 88.115 55.575 88.160 ;
        RECT 56.650 88.100 56.970 88.160 ;
        RECT 58.490 88.300 58.810 88.360 ;
        RECT 59.040 88.345 59.180 88.840 ;
        RECT 61.710 88.780 62.030 88.840 ;
        RECT 75.510 88.780 75.830 89.040 ;
        RECT 86.570 88.980 86.860 89.025 ;
        RECT 88.430 88.980 88.720 89.025 ;
        RECT 91.210 88.980 91.500 89.025 ;
        RECT 86.570 88.840 91.500 88.980 ;
        RECT 86.570 88.795 86.860 88.840 ;
        RECT 88.430 88.795 88.720 88.840 ;
        RECT 91.210 88.795 91.500 88.840 ;
        RECT 61.250 88.640 61.570 88.700 ;
        RECT 59.500 88.500 61.570 88.640 ;
        RECT 59.500 88.345 59.640 88.500 ;
        RECT 61.250 88.440 61.570 88.500 ;
        RECT 72.290 88.640 72.610 88.700 ;
        RECT 73.685 88.640 73.975 88.685 ;
        RECT 75.600 88.640 75.740 88.780 ;
        RECT 72.290 88.500 75.740 88.640 ;
        RECT 86.105 88.640 86.395 88.685 ;
        RECT 87.010 88.640 87.330 88.700 ;
        RECT 86.105 88.500 87.330 88.640 ;
        RECT 72.290 88.440 72.610 88.500 ;
        RECT 73.685 88.455 73.975 88.500 ;
        RECT 86.105 88.455 86.395 88.500 ;
        RECT 87.010 88.440 87.330 88.500 ;
        RECT 87.945 88.640 88.235 88.685 ;
        RECT 91.610 88.640 91.930 88.700 ;
        RECT 109.180 88.685 109.320 89.180 ;
        RECT 111.390 89.120 111.710 89.180 ;
        RECT 112.330 88.980 112.620 89.025 ;
        RECT 114.190 88.980 114.480 89.025 ;
        RECT 116.970 88.980 117.260 89.025 ;
        RECT 112.330 88.840 117.260 88.980 ;
        RECT 117.460 88.980 117.600 89.180 ;
        RECT 117.460 88.840 120.820 88.980 ;
        RECT 112.330 88.795 112.620 88.840 ;
        RECT 114.190 88.795 114.480 88.840 ;
        RECT 116.970 88.795 117.260 88.840 ;
        RECT 120.680 88.700 120.820 88.840 ;
        RECT 87.945 88.500 91.930 88.640 ;
        RECT 87.945 88.455 88.235 88.500 ;
        RECT 91.610 88.440 91.930 88.500 ;
        RECT 105.960 88.500 108.400 88.640 ;
        RECT 105.960 88.360 106.100 88.500 ;
        RECT 58.965 88.300 59.255 88.345 ;
        RECT 58.490 88.160 59.255 88.300 ;
        RECT 58.490 88.100 58.810 88.160 ;
        RECT 58.965 88.115 59.255 88.160 ;
        RECT 59.425 88.115 59.715 88.345 ;
        RECT 59.885 88.115 60.175 88.345 ;
        RECT 51.145 87.960 51.435 88.005 ;
        RECT 53.890 87.960 54.210 88.020 ;
        RECT 55.745 87.960 56.035 88.005 ;
        RECT 59.960 87.960 60.100 88.115 ;
        RECT 60.790 88.100 61.110 88.360 ;
        RECT 68.625 88.300 68.915 88.345 ;
        RECT 72.765 88.300 73.055 88.345 ;
        RECT 74.590 88.300 74.910 88.360 ;
        RECT 68.625 88.160 70.680 88.300 ;
        RECT 68.625 88.115 68.915 88.160 ;
        RECT 51.145 87.820 60.100 87.960 ;
        RECT 51.145 87.775 51.435 87.820 ;
        RECT 53.890 87.760 54.210 87.820 ;
        RECT 55.745 87.775 56.035 87.820 ;
        RECT 70.540 87.665 70.680 88.160 ;
        RECT 72.765 88.160 74.910 88.300 ;
        RECT 72.765 88.115 73.055 88.160 ;
        RECT 74.590 88.100 74.910 88.160 ;
        RECT 75.050 88.300 75.370 88.360 ;
        RECT 75.525 88.300 75.815 88.345 ;
        RECT 91.210 88.300 91.500 88.345 ;
        RECT 75.050 88.160 75.815 88.300 ;
        RECT 75.050 88.100 75.370 88.160 ;
        RECT 75.525 88.115 75.815 88.160 ;
        RECT 88.965 88.160 91.500 88.300 ;
        RECT 88.965 88.005 89.180 88.160 ;
        RECT 91.210 88.115 91.500 88.160 ;
        RECT 105.870 88.100 106.190 88.360 ;
        RECT 108.260 88.345 108.400 88.500 ;
        RECT 109.105 88.455 109.395 88.685 ;
        RECT 110.010 88.640 110.330 88.700 ;
        RECT 111.865 88.640 112.155 88.685 ;
        RECT 110.010 88.500 112.155 88.640 ;
        RECT 110.010 88.440 110.330 88.500 ;
        RECT 111.865 88.455 112.155 88.500 ;
        RECT 120.590 88.440 120.910 88.700 ;
        RECT 106.805 88.115 107.095 88.345 ;
        RECT 108.185 88.115 108.475 88.345 ;
        RECT 92.990 88.005 93.310 88.020 ;
        RECT 87.030 87.960 87.320 88.005 ;
        RECT 88.890 87.960 89.180 88.005 ;
        RECT 87.030 87.820 89.180 87.960 ;
        RECT 87.030 87.775 87.320 87.820 ;
        RECT 88.890 87.775 89.180 87.820 ;
        RECT 89.810 87.960 90.100 88.005 ;
        RECT 92.990 87.960 93.360 88.005 ;
        RECT 89.810 87.820 93.360 87.960 ;
        RECT 106.880 87.960 107.020 88.115 ;
        RECT 110.470 88.100 110.790 88.360 ;
        RECT 113.705 88.300 113.995 88.345 ;
        RECT 116.970 88.300 117.260 88.345 ;
        RECT 111.480 88.160 113.995 88.300 ;
        RECT 110.930 87.960 111.250 88.020 ;
        RECT 106.880 87.820 111.250 87.960 ;
        RECT 89.810 87.775 90.100 87.820 ;
        RECT 92.990 87.775 93.360 87.820 ;
        RECT 92.990 87.760 93.310 87.775 ;
        RECT 110.930 87.760 111.250 87.820 ;
        RECT 49.305 87.435 49.595 87.665 ;
        RECT 70.465 87.435 70.755 87.665 ;
        RECT 72.305 87.620 72.595 87.665 ;
        RECT 77.810 87.620 78.130 87.680 ;
        RECT 72.305 87.480 78.130 87.620 ;
        RECT 72.305 87.435 72.595 87.480 ;
        RECT 77.810 87.420 78.130 87.480 ;
        RECT 104.950 87.420 105.270 87.680 ;
        RECT 106.330 87.620 106.650 87.680 ;
        RECT 111.480 87.665 111.620 88.160 ;
        RECT 113.705 88.115 113.995 88.160 ;
        RECT 114.725 88.160 117.260 88.300 ;
        RECT 114.725 88.005 114.940 88.160 ;
        RECT 116.970 88.115 117.260 88.160 ;
        RECT 122.890 88.100 123.210 88.360 ;
        RECT 112.790 87.960 113.080 88.005 ;
        RECT 114.650 87.960 114.940 88.005 ;
        RECT 112.790 87.820 114.940 87.960 ;
        RECT 112.790 87.775 113.080 87.820 ;
        RECT 114.650 87.775 114.940 87.820 ;
        RECT 115.570 87.960 115.860 88.005 ;
        RECT 117.830 87.960 118.150 88.020 ;
        RECT 118.830 87.960 119.120 88.005 ;
        RECT 115.570 87.820 119.120 87.960 ;
        RECT 115.570 87.775 115.860 87.820 ;
        RECT 117.830 87.760 118.150 87.820 ;
        RECT 118.830 87.775 119.120 87.820 ;
        RECT 107.265 87.620 107.555 87.665 ;
        RECT 106.330 87.480 107.555 87.620 ;
        RECT 106.330 87.420 106.650 87.480 ;
        RECT 107.265 87.435 107.555 87.480 ;
        RECT 111.405 87.435 111.695 87.665 ;
        RECT 117.370 87.620 117.690 87.680 ;
        RECT 120.835 87.620 121.125 87.665 ;
        RECT 117.370 87.480 121.125 87.620 ;
        RECT 117.370 87.420 117.690 87.480 ;
        RECT 120.835 87.435 121.125 87.480 ;
        RECT 121.970 87.420 122.290 87.680 ;
        RECT 5.520 86.800 125.580 87.280 ;
        RECT 22.150 86.600 22.470 86.660 ;
        RECT 23.085 86.600 23.375 86.645 ;
        RECT 22.150 86.460 23.375 86.600 ;
        RECT 22.150 86.400 22.470 86.460 ;
        RECT 23.085 86.415 23.375 86.460 ;
        RECT 27.670 86.600 27.990 86.660 ;
        RECT 32.730 86.600 33.050 86.660 ;
        RECT 27.670 86.460 33.050 86.600 ;
        RECT 27.670 86.400 27.990 86.460 ;
        RECT 32.730 86.400 33.050 86.460 ;
        RECT 44.705 86.600 44.995 86.645 ;
        RECT 53.890 86.600 54.210 86.660 ;
        RECT 54.595 86.600 54.885 86.645 ;
        RECT 44.705 86.460 49.060 86.600 ;
        RECT 44.705 86.415 44.995 86.460 ;
        RECT 46.550 86.260 46.840 86.305 ;
        RECT 48.410 86.260 48.700 86.305 ;
        RECT 46.550 86.120 48.700 86.260 ;
        RECT 48.920 86.260 49.060 86.460 ;
        RECT 53.890 86.460 54.885 86.600 ;
        RECT 53.890 86.400 54.210 86.460 ;
        RECT 54.595 86.415 54.885 86.460 ;
        RECT 61.250 86.600 61.570 86.660 ;
        RECT 64.025 86.600 64.315 86.645 ;
        RECT 61.250 86.460 64.315 86.600 ;
        RECT 61.250 86.400 61.570 86.460 ;
        RECT 64.025 86.415 64.315 86.460 ;
        RECT 104.490 86.400 104.810 86.660 ;
        RECT 117.370 86.600 117.690 86.660 ;
        RECT 106.880 86.460 117.690 86.600 ;
        RECT 49.330 86.260 49.620 86.305 ;
        RECT 52.590 86.260 52.880 86.305 ;
        RECT 48.920 86.120 52.880 86.260 ;
        RECT 46.550 86.075 46.840 86.120 ;
        RECT 48.410 86.075 48.700 86.120 ;
        RECT 49.330 86.075 49.620 86.120 ;
        RECT 52.590 86.075 52.880 86.120 ;
        RECT 58.490 86.260 58.810 86.320 ;
        RECT 61.340 86.260 61.480 86.400 ;
        RECT 58.490 86.120 59.180 86.260 ;
        RECT 23.990 85.720 24.310 85.980 ;
        RECT 25.370 85.720 25.690 85.980 ;
        RECT 43.310 85.920 43.630 85.980 ;
        RECT 44.245 85.920 44.535 85.965 ;
        RECT 43.310 85.780 44.535 85.920 ;
        RECT 43.310 85.720 43.630 85.780 ;
        RECT 44.245 85.735 44.535 85.780 ;
        RECT 44.690 85.920 45.010 85.980 ;
        RECT 45.625 85.920 45.915 85.965 ;
        RECT 44.690 85.780 45.915 85.920 ;
        RECT 44.690 85.720 45.010 85.780 ;
        RECT 45.625 85.735 45.915 85.780 ;
        RECT 46.990 85.920 47.310 85.980 ;
        RECT 47.465 85.920 47.755 85.965 ;
        RECT 46.990 85.780 47.755 85.920 ;
        RECT 48.485 85.920 48.700 86.075 ;
        RECT 58.490 86.060 58.810 86.120 ;
        RECT 50.730 85.920 51.020 85.965 ;
        RECT 48.485 85.780 51.020 85.920 ;
        RECT 46.990 85.720 47.310 85.780 ;
        RECT 47.465 85.735 47.755 85.780 ;
        RECT 50.730 85.735 51.020 85.780 ;
        RECT 55.730 85.920 56.050 85.980 ;
        RECT 59.040 85.965 59.180 86.120 ;
        RECT 59.500 86.120 61.480 86.260 ;
        RECT 61.710 86.260 62.030 86.320 ;
        RECT 69.070 86.260 69.390 86.320 ;
        RECT 80.570 86.260 80.890 86.320 ;
        RECT 94.370 86.260 94.690 86.320 ;
        RECT 61.710 86.120 80.890 86.260 ;
        RECT 59.500 85.965 59.640 86.120 ;
        RECT 61.710 86.060 62.030 86.120 ;
        RECT 69.070 86.060 69.390 86.120 ;
        RECT 80.570 86.060 80.890 86.120 ;
        RECT 84.800 86.120 94.690 86.260 ;
        RECT 55.730 85.780 58.720 85.920 ;
        RECT 55.730 85.720 56.050 85.780 ;
        RECT 22.150 85.580 22.470 85.640 ;
        RECT 24.465 85.580 24.755 85.625 ;
        RECT 22.150 85.440 24.755 85.580 ;
        RECT 22.150 85.380 22.470 85.440 ;
        RECT 24.465 85.395 24.755 85.440 ;
        RECT 33.650 85.580 33.970 85.640 ;
        RECT 58.580 85.580 58.720 85.780 ;
        RECT 58.965 85.735 59.255 85.965 ;
        RECT 59.425 85.735 59.715 85.965 ;
        RECT 59.885 85.735 60.175 85.965 ;
        RECT 59.960 85.580 60.100 85.735 ;
        RECT 60.790 85.720 61.110 85.980 ;
        RECT 64.945 85.920 65.235 85.965 ;
        RECT 65.850 85.920 66.170 85.980 ;
        RECT 64.945 85.780 66.170 85.920 ;
        RECT 64.945 85.735 65.235 85.780 ;
        RECT 65.850 85.720 66.170 85.780 ;
        RECT 77.365 85.735 77.655 85.965 ;
        RECT 78.730 85.920 79.050 85.980 ;
        RECT 84.800 85.920 84.940 86.120 ;
        RECT 94.370 86.060 94.690 86.120 ;
        RECT 95.305 86.260 95.595 86.305 ;
        RECT 102.205 86.260 102.495 86.305 ;
        RECT 95.305 86.120 102.495 86.260 ;
        RECT 95.305 86.075 95.595 86.120 ;
        RECT 102.205 86.075 102.495 86.120 ;
        RECT 78.730 85.780 84.940 85.920 ;
        RECT 33.650 85.440 51.360 85.580 ;
        RECT 58.580 85.440 60.100 85.580 ;
        RECT 33.650 85.380 33.970 85.440 ;
        RECT 46.090 85.240 46.380 85.285 ;
        RECT 47.950 85.240 48.240 85.285 ;
        RECT 50.730 85.240 51.020 85.285 ;
        RECT 46.090 85.100 51.020 85.240 ;
        RECT 51.220 85.240 51.360 85.440 ;
        RECT 76.430 85.380 76.750 85.640 ;
        RECT 77.440 85.580 77.580 85.735 ;
        RECT 78.730 85.720 79.050 85.780 ;
        RECT 88.850 85.720 89.170 85.980 ;
        RECT 92.085 85.920 92.375 85.965 ;
        RECT 89.400 85.780 92.375 85.920 ;
        RECT 82.870 85.580 83.190 85.640 ;
        RECT 77.440 85.440 83.190 85.580 ;
        RECT 82.870 85.380 83.190 85.440 ;
        RECT 76.520 85.240 76.660 85.380 ;
        RECT 79.650 85.240 79.970 85.300 ;
        RECT 89.400 85.240 89.540 85.780 ;
        RECT 92.085 85.735 92.375 85.780 ;
        RECT 92.530 85.920 92.850 85.980 ;
        RECT 93.005 85.920 93.295 85.965 ;
        RECT 92.530 85.780 93.295 85.920 ;
        RECT 92.530 85.720 92.850 85.780 ;
        RECT 93.005 85.735 93.295 85.780 ;
        RECT 93.465 85.735 93.755 85.965 ;
        RECT 93.925 85.735 94.215 85.965 ;
        RECT 91.610 85.580 91.930 85.640 ;
        RECT 93.540 85.580 93.680 85.735 ;
        RECT 91.610 85.440 93.680 85.580 ;
        RECT 91.610 85.380 91.930 85.440 ;
        RECT 51.220 85.100 89.540 85.240 ;
        RECT 46.090 85.055 46.380 85.100 ;
        RECT 47.950 85.055 48.240 85.100 ;
        RECT 50.730 85.055 51.020 85.100 ;
        RECT 79.650 85.040 79.970 85.100 ;
        RECT 23.530 84.900 23.850 84.960 ;
        RECT 24.005 84.900 24.295 84.945 ;
        RECT 23.530 84.760 24.295 84.900 ;
        RECT 23.530 84.700 23.850 84.760 ;
        RECT 24.005 84.715 24.295 84.760 ;
        RECT 57.570 84.700 57.890 84.960 ;
        RECT 75.970 84.900 76.290 84.960 ;
        RECT 76.445 84.900 76.735 84.945 ;
        RECT 75.970 84.760 76.735 84.900 ;
        RECT 75.970 84.700 76.290 84.760 ;
        RECT 76.445 84.715 76.735 84.760 ;
        RECT 78.270 84.700 78.590 84.960 ;
        RECT 87.930 84.700 88.250 84.960 ;
        RECT 89.400 84.900 89.540 85.100 ;
        RECT 90.690 85.240 91.010 85.300 ;
        RECT 94.000 85.240 94.140 85.735 ;
        RECT 103.570 85.720 103.890 85.980 ;
        RECT 105.870 85.720 106.190 85.980 ;
        RECT 106.880 85.965 107.020 86.460 ;
        RECT 117.370 86.400 117.690 86.460 ;
        RECT 120.590 86.600 120.910 86.660 ;
        RECT 121.755 86.600 122.045 86.645 ;
        RECT 120.590 86.460 122.045 86.600 ;
        RECT 120.590 86.400 120.910 86.460 ;
        RECT 121.755 86.415 122.045 86.460 ;
        RECT 113.710 86.260 114.000 86.305 ;
        RECT 115.570 86.260 115.860 86.305 ;
        RECT 113.710 86.120 115.860 86.260 ;
        RECT 113.710 86.075 114.000 86.120 ;
        RECT 115.570 86.075 115.860 86.120 ;
        RECT 116.490 86.260 116.780 86.305 ;
        RECT 118.290 86.260 118.610 86.320 ;
        RECT 119.750 86.260 120.040 86.305 ;
        RECT 116.490 86.120 120.040 86.260 ;
        RECT 116.490 86.075 116.780 86.120 ;
        RECT 106.805 85.735 107.095 85.965 ;
        RECT 110.010 85.920 110.330 85.980 ;
        RECT 112.785 85.920 113.075 85.965 ;
        RECT 110.010 85.780 113.075 85.920 ;
        RECT 115.645 85.920 115.860 86.075 ;
        RECT 118.290 86.060 118.610 86.120 ;
        RECT 119.750 86.075 120.040 86.120 ;
        RECT 117.890 85.920 118.180 85.965 ;
        RECT 115.645 85.780 118.180 85.920 ;
        RECT 110.010 85.720 110.330 85.780 ;
        RECT 112.785 85.735 113.075 85.780 ;
        RECT 117.890 85.735 118.180 85.780 ;
        RECT 102.650 85.380 102.970 85.640 ;
        RECT 114.625 85.580 114.915 85.625 ;
        RECT 121.970 85.580 122.290 85.640 ;
        RECT 114.625 85.440 122.290 85.580 ;
        RECT 114.625 85.395 114.915 85.440 ;
        RECT 121.970 85.380 122.290 85.440 ;
        RECT 94.830 85.240 95.150 85.300 ;
        RECT 90.690 85.100 95.150 85.240 ;
        RECT 90.690 85.040 91.010 85.100 ;
        RECT 94.830 85.040 95.150 85.100 ;
        RECT 113.250 85.240 113.540 85.285 ;
        RECT 115.110 85.240 115.400 85.285 ;
        RECT 117.890 85.240 118.180 85.285 ;
        RECT 113.250 85.100 118.180 85.240 ;
        RECT 113.250 85.055 113.540 85.100 ;
        RECT 115.110 85.055 115.400 85.100 ;
        RECT 117.890 85.055 118.180 85.100 ;
        RECT 95.750 84.900 96.070 84.960 ;
        RECT 89.400 84.760 96.070 84.900 ;
        RECT 95.750 84.700 96.070 84.760 ;
        RECT 102.190 84.700 102.510 84.960 ;
        RECT 104.965 84.900 105.255 84.945 ;
        RECT 105.410 84.900 105.730 84.960 ;
        RECT 104.965 84.760 105.730 84.900 ;
        RECT 104.965 84.715 105.255 84.760 ;
        RECT 105.410 84.700 105.730 84.760 ;
        RECT 5.520 84.080 125.580 84.560 ;
        RECT 24.005 83.880 24.295 83.925 ;
        RECT 25.370 83.880 25.690 83.940 ;
        RECT 24.005 83.740 25.690 83.880 ;
        RECT 24.005 83.695 24.295 83.740 ;
        RECT 25.370 83.680 25.690 83.740 ;
        RECT 28.590 83.880 28.910 83.940 ;
        RECT 35.030 83.880 35.350 83.940 ;
        RECT 28.590 83.740 35.350 83.880 ;
        RECT 28.590 83.680 28.910 83.740 ;
        RECT 35.030 83.680 35.350 83.740 ;
        RECT 56.665 83.880 56.955 83.925 ;
        RECT 59.870 83.880 60.190 83.940 ;
        RECT 56.665 83.740 60.190 83.880 ;
        RECT 56.665 83.695 56.955 83.740 ;
        RECT 59.870 83.680 60.190 83.740 ;
        RECT 69.070 83.680 69.390 83.940 ;
        RECT 103.585 83.880 103.875 83.925 ;
        RECT 104.950 83.880 105.270 83.940 ;
        RECT 103.585 83.740 105.270 83.880 ;
        RECT 103.585 83.695 103.875 83.740 ;
        RECT 104.950 83.680 105.270 83.740 ;
        RECT 106.330 83.680 106.650 83.940 ;
        RECT 23.070 83.540 23.390 83.600 ;
        RECT 21.320 83.400 23.390 83.540 ;
        RECT 20.770 82.860 21.090 82.920 ;
        RECT 21.320 82.860 21.460 83.400 ;
        RECT 23.070 83.340 23.390 83.400 ;
        RECT 24.450 83.540 24.770 83.600 ;
        RECT 28.680 83.540 28.820 83.680 ;
        RECT 24.450 83.400 28.820 83.540 ;
        RECT 24.450 83.340 24.770 83.400 ;
        RECT 28.130 83.200 28.450 83.260 ;
        RECT 22.240 83.060 28.450 83.200 ;
        RECT 22.240 82.905 22.380 83.060 ;
        RECT 20.770 82.720 21.460 82.860 ;
        RECT 20.770 82.660 21.090 82.720 ;
        RECT 21.705 82.675 21.995 82.905 ;
        RECT 22.165 82.675 22.455 82.905 ;
        RECT 22.625 82.675 22.915 82.905 ;
        RECT 23.070 82.860 23.390 82.920 ;
        RECT 26.840 82.905 26.980 83.060 ;
        RECT 28.130 83.000 28.450 83.060 ;
        RECT 25.385 82.860 25.675 82.905 ;
        RECT 23.070 82.720 25.675 82.860 ;
        RECT 15.710 82.520 16.030 82.580 ;
        RECT 21.780 82.520 21.920 82.675 ;
        RECT 15.710 82.380 21.920 82.520 ;
        RECT 15.710 82.320 16.030 82.380 ;
        RECT 20.770 82.180 21.090 82.240 ;
        RECT 22.240 82.180 22.380 82.675 ;
        RECT 22.700 82.520 22.840 82.675 ;
        RECT 23.070 82.660 23.390 82.720 ;
        RECT 25.385 82.675 25.675 82.720 ;
        RECT 26.305 82.675 26.595 82.905 ;
        RECT 26.765 82.675 27.055 82.905 ;
        RECT 27.225 82.860 27.515 82.905 ;
        RECT 28.680 82.860 28.820 83.400 ;
        RECT 33.615 83.540 33.905 83.585 ;
        RECT 35.505 83.540 35.795 83.585 ;
        RECT 38.625 83.540 38.915 83.585 ;
        RECT 33.615 83.400 38.915 83.540 ;
        RECT 33.615 83.355 33.905 83.400 ;
        RECT 35.505 83.355 35.795 83.400 ;
        RECT 38.625 83.355 38.915 83.400 ;
        RECT 45.170 83.540 45.460 83.585 ;
        RECT 47.030 83.540 47.320 83.585 ;
        RECT 49.810 83.540 50.100 83.585 ;
        RECT 45.170 83.400 50.100 83.540 ;
        RECT 45.170 83.355 45.460 83.400 ;
        RECT 47.030 83.355 47.320 83.400 ;
        RECT 49.810 83.355 50.100 83.400 ;
        RECT 52.050 83.540 52.370 83.600 ;
        RECT 60.345 83.540 60.635 83.585 ;
        RECT 78.730 83.540 79.050 83.600 ;
        RECT 52.050 83.400 60.635 83.540 ;
        RECT 52.050 83.340 52.370 83.400 ;
        RECT 60.345 83.355 60.635 83.400 ;
        RECT 75.140 83.400 79.050 83.540 ;
        RECT 32.730 83.000 33.050 83.260 ;
        RECT 34.125 83.200 34.415 83.245 ;
        RECT 34.570 83.200 34.890 83.260 ;
        RECT 43.770 83.200 44.090 83.260 ;
        RECT 34.125 83.060 34.890 83.200 ;
        RECT 34.125 83.015 34.415 83.060 ;
        RECT 34.570 83.000 34.890 83.060 ;
        RECT 43.400 83.060 44.090 83.200 ;
        RECT 27.225 82.720 28.820 82.860 ;
        RECT 32.285 82.860 32.575 82.905 ;
        RECT 33.210 82.860 33.500 82.905 ;
        RECT 35.045 82.860 35.335 82.905 ;
        RECT 38.625 82.860 38.915 82.905 ;
        RECT 32.285 82.720 32.960 82.860 ;
        RECT 27.225 82.675 27.515 82.720 ;
        RECT 32.285 82.675 32.575 82.720 ;
        RECT 24.450 82.520 24.770 82.580 ;
        RECT 22.700 82.380 24.770 82.520 ;
        RECT 26.380 82.520 26.520 82.675 ;
        RECT 32.820 82.520 32.960 82.720 ;
        RECT 33.210 82.720 38.915 82.860 ;
        RECT 33.210 82.675 33.500 82.720 ;
        RECT 35.045 82.675 35.335 82.720 ;
        RECT 38.625 82.675 38.915 82.720 ;
        RECT 39.705 82.565 39.995 82.880 ;
        RECT 42.905 82.860 43.195 82.905 ;
        RECT 43.400 82.860 43.540 83.060 ;
        RECT 43.770 83.000 44.090 83.060 ;
        RECT 44.690 83.000 45.010 83.260 ;
        RECT 46.545 83.200 46.835 83.245 ;
        RECT 47.450 83.200 47.770 83.260 ;
        RECT 46.545 83.060 47.770 83.200 ;
        RECT 46.545 83.015 46.835 83.060 ;
        RECT 47.450 83.000 47.770 83.060 ;
        RECT 47.910 83.200 48.230 83.260 ;
        RECT 53.675 83.200 53.965 83.245 ;
        RECT 55.730 83.200 56.050 83.260 ;
        RECT 47.910 83.060 56.050 83.200 ;
        RECT 47.910 83.000 48.230 83.060 ;
        RECT 53.675 83.015 53.965 83.060 ;
        RECT 55.730 83.000 56.050 83.060 ;
        RECT 56.190 83.000 56.510 83.260 ;
        RECT 67.245 83.200 67.535 83.245 ;
        RECT 72.750 83.200 73.070 83.260 ;
        RECT 75.140 83.200 75.280 83.400 ;
        RECT 78.730 83.340 79.050 83.400 ;
        RECT 86.570 83.540 86.860 83.585 ;
        RECT 88.430 83.540 88.720 83.585 ;
        RECT 91.210 83.540 91.500 83.585 ;
        RECT 86.570 83.400 91.500 83.540 ;
        RECT 86.570 83.355 86.860 83.400 ;
        RECT 88.430 83.355 88.720 83.400 ;
        RECT 91.210 83.355 91.500 83.400 ;
        RECT 94.830 83.540 95.150 83.600 ;
        RECT 112.770 83.540 113.090 83.600 ;
        RECT 94.830 83.400 98.280 83.540 ;
        RECT 94.830 83.340 95.150 83.400 ;
        RECT 67.245 83.060 72.520 83.200 ;
        RECT 67.245 83.015 67.535 83.060 ;
        RECT 72.380 82.920 72.520 83.060 ;
        RECT 72.750 83.060 75.280 83.200 ;
        RECT 77.810 83.200 78.130 83.260 ;
        RECT 78.285 83.200 78.575 83.245 ;
        RECT 77.810 83.060 81.260 83.200 ;
        RECT 72.750 83.000 73.070 83.060 ;
        RECT 49.810 82.860 50.100 82.905 ;
        RECT 42.905 82.720 43.540 82.860 ;
        RECT 47.565 82.720 50.100 82.860 ;
        RECT 42.905 82.675 43.195 82.720 ;
        RECT 47.565 82.565 47.780 82.720 ;
        RECT 49.810 82.675 50.100 82.720 ;
        RECT 55.285 82.675 55.575 82.905 ;
        RECT 56.665 82.860 56.955 82.905 ;
        RECT 57.570 82.860 57.890 82.920 ;
        RECT 56.665 82.720 57.890 82.860 ;
        RECT 56.665 82.675 56.955 82.720 ;
        RECT 26.380 82.380 32.960 82.520 ;
        RECT 23.160 82.240 23.300 82.380 ;
        RECT 24.450 82.320 24.770 82.380 ;
        RECT 20.770 82.040 22.380 82.180 ;
        RECT 20.770 81.980 21.090 82.040 ;
        RECT 23.070 81.980 23.390 82.240 ;
        RECT 28.590 81.980 28.910 82.240 ;
        RECT 29.065 82.180 29.355 82.225 ;
        RECT 30.890 82.180 31.210 82.240 ;
        RECT 29.065 82.040 31.210 82.180 ;
        RECT 32.820 82.180 32.960 82.380 ;
        RECT 36.405 82.520 37.055 82.565 ;
        RECT 39.705 82.520 40.295 82.565 ;
        RECT 42.405 82.520 42.695 82.565 ;
        RECT 36.405 82.380 42.695 82.520 ;
        RECT 36.405 82.335 37.055 82.380 ;
        RECT 40.005 82.335 40.295 82.380 ;
        RECT 42.405 82.335 42.695 82.380 ;
        RECT 45.630 82.520 45.920 82.565 ;
        RECT 47.490 82.520 47.780 82.565 ;
        RECT 45.630 82.380 47.780 82.520 ;
        RECT 45.630 82.335 45.920 82.380 ;
        RECT 47.490 82.335 47.780 82.380 ;
        RECT 48.370 82.565 48.690 82.580 ;
        RECT 48.370 82.520 48.700 82.565 ;
        RECT 51.670 82.520 51.960 82.565 ;
        RECT 48.370 82.380 51.960 82.520 ;
        RECT 48.370 82.335 48.700 82.380 ;
        RECT 51.670 82.335 51.960 82.380 ;
        RECT 52.970 82.520 53.290 82.580 ;
        RECT 55.360 82.520 55.500 82.675 ;
        RECT 57.570 82.660 57.890 82.720 ;
        RECT 63.090 82.860 63.410 82.920 ;
        RECT 64.485 82.860 64.775 82.905 ;
        RECT 63.090 82.720 64.775 82.860 ;
        RECT 63.090 82.660 63.410 82.720 ;
        RECT 64.485 82.675 64.775 82.720 ;
        RECT 65.390 82.860 65.710 82.920 ;
        RECT 68.165 82.860 68.455 82.905 ;
        RECT 65.390 82.720 68.455 82.860 ;
        RECT 65.390 82.660 65.710 82.720 ;
        RECT 68.165 82.675 68.455 82.720 ;
        RECT 71.370 82.660 71.690 82.920 ;
        RECT 72.290 82.660 72.610 82.920 ;
        RECT 74.680 82.905 74.820 83.060 ;
        RECT 77.810 83.000 78.130 83.060 ;
        RECT 78.285 83.015 78.575 83.060 ;
        RECT 73.225 82.675 73.515 82.905 ;
        RECT 74.605 82.675 74.895 82.905 ;
        RECT 79.650 82.860 79.970 82.920 ;
        RECT 81.120 82.905 81.260 83.060 ;
        RECT 87.930 83.000 88.250 83.260 ;
        RECT 90.690 83.200 91.010 83.260 ;
        RECT 88.480 83.060 91.010 83.200 ;
        RECT 80.125 82.860 80.415 82.905 ;
        RECT 79.650 82.720 80.415 82.860 ;
        RECT 59.410 82.520 59.730 82.580 ;
        RECT 52.970 82.380 54.580 82.520 ;
        RECT 55.360 82.380 59.730 82.520 ;
        RECT 48.370 82.320 48.690 82.335 ;
        RECT 52.970 82.320 53.290 82.380 ;
        RECT 54.440 82.225 54.580 82.380 ;
        RECT 59.410 82.320 59.730 82.380 ;
        RECT 61.250 82.520 61.570 82.580 ;
        RECT 65.865 82.520 66.155 82.565 ;
        RECT 71.845 82.520 72.135 82.565 ;
        RECT 61.250 82.380 66.155 82.520 ;
        RECT 61.250 82.320 61.570 82.380 ;
        RECT 65.865 82.335 66.155 82.380 ;
        RECT 66.400 82.380 72.135 82.520 ;
        RECT 73.300 82.520 73.440 82.675 ;
        RECT 79.650 82.660 79.970 82.720 ;
        RECT 80.125 82.675 80.415 82.720 ;
        RECT 81.045 82.675 81.335 82.905 ;
        RECT 81.490 82.660 81.810 82.920 ;
        RECT 81.965 82.675 82.255 82.905 ;
        RECT 82.870 82.860 83.190 82.920 ;
        RECT 86.105 82.860 86.395 82.905 ;
        RECT 88.480 82.860 88.620 83.060 ;
        RECT 90.690 83.000 91.010 83.060 ;
        RECT 91.610 83.200 91.930 83.260 ;
        RECT 91.610 83.060 97.820 83.200 ;
        RECT 91.610 83.000 91.930 83.060 ;
        RECT 91.210 82.860 91.500 82.905 ;
        RECT 82.870 82.720 86.395 82.860 ;
        RECT 75.525 82.520 75.815 82.565 ;
        RECT 73.300 82.380 75.815 82.520 ;
        RECT 41.485 82.180 41.775 82.225 ;
        RECT 32.820 82.040 41.775 82.180 ;
        RECT 29.065 81.995 29.355 82.040 ;
        RECT 30.890 81.980 31.210 82.040 ;
        RECT 41.485 81.995 41.775 82.040 ;
        RECT 54.365 81.995 54.655 82.225 ;
        RECT 60.790 82.180 61.110 82.240 ;
        RECT 63.565 82.180 63.855 82.225 ;
        RECT 60.790 82.040 63.855 82.180 ;
        RECT 60.790 81.980 61.110 82.040 ;
        RECT 63.565 81.995 63.855 82.040 ;
        RECT 64.470 82.180 64.790 82.240 ;
        RECT 66.400 82.180 66.540 82.380 ;
        RECT 71.845 82.335 72.135 82.380 ;
        RECT 75.525 82.335 75.815 82.380 ;
        RECT 80.570 82.520 80.890 82.580 ;
        RECT 82.040 82.520 82.180 82.675 ;
        RECT 82.870 82.660 83.190 82.720 ;
        RECT 86.105 82.675 86.395 82.720 ;
        RECT 86.640 82.720 88.620 82.860 ;
        RECT 88.965 82.720 91.500 82.860 ;
        RECT 86.640 82.520 86.780 82.720 ;
        RECT 88.965 82.565 89.180 82.720 ;
        RECT 91.210 82.675 91.500 82.720 ;
        RECT 95.750 82.860 96.070 82.920 ;
        RECT 96.225 82.860 96.515 82.905 ;
        RECT 95.750 82.720 96.515 82.860 ;
        RECT 95.750 82.660 96.070 82.720 ;
        RECT 96.225 82.675 96.515 82.720 ;
        RECT 96.670 82.860 96.990 82.920 ;
        RECT 97.680 82.905 97.820 83.060 ;
        RECT 98.140 82.905 98.280 83.400 ;
        RECT 103.200 83.400 113.090 83.540 ;
        RECT 103.200 83.245 103.340 83.400 ;
        RECT 112.770 83.340 113.090 83.400 ;
        RECT 103.125 83.015 103.415 83.245 ;
        RECT 105.870 83.000 106.190 83.260 ;
        RECT 118.750 83.200 119.070 83.260 ;
        RECT 118.380 83.060 119.070 83.200 ;
        RECT 97.145 82.860 97.435 82.905 ;
        RECT 96.670 82.720 97.435 82.860 ;
        RECT 96.670 82.660 96.990 82.720 ;
        RECT 97.145 82.675 97.435 82.720 ;
        RECT 97.605 82.675 97.895 82.905 ;
        RECT 98.065 82.675 98.355 82.905 ;
        RECT 103.585 82.860 103.875 82.905 ;
        RECT 104.030 82.860 104.350 82.920 ;
        RECT 103.585 82.720 104.350 82.860 ;
        RECT 103.585 82.675 103.875 82.720 ;
        RECT 104.030 82.660 104.350 82.720 ;
        RECT 106.330 82.660 106.650 82.920 ;
        RECT 117.830 82.660 118.150 82.920 ;
        RECT 118.380 82.905 118.520 83.060 ;
        RECT 118.750 83.000 119.070 83.060 ;
        RECT 118.305 82.675 118.595 82.905 ;
        RECT 80.570 82.380 86.780 82.520 ;
        RECT 87.030 82.520 87.320 82.565 ;
        RECT 88.890 82.520 89.180 82.565 ;
        RECT 87.030 82.380 89.180 82.520 ;
        RECT 80.570 82.320 80.890 82.380 ;
        RECT 87.030 82.335 87.320 82.380 ;
        RECT 88.890 82.335 89.180 82.380 ;
        RECT 89.810 82.520 90.100 82.565 ;
        RECT 92.530 82.520 92.850 82.580 ;
        RECT 93.070 82.520 93.360 82.565 ;
        RECT 99.445 82.520 99.735 82.565 ;
        RECT 102.205 82.520 102.495 82.565 ;
        RECT 104.965 82.520 105.255 82.565 ;
        RECT 89.810 82.380 93.360 82.520 ;
        RECT 89.810 82.335 90.100 82.380 ;
        RECT 92.530 82.320 92.850 82.380 ;
        RECT 93.070 82.335 93.360 82.380 ;
        RECT 94.460 82.380 99.200 82.520 ;
        RECT 64.470 82.040 66.540 82.180 ;
        RECT 64.470 81.980 64.790 82.040 ;
        RECT 70.450 81.980 70.770 82.240 ;
        RECT 74.130 81.980 74.450 82.240 ;
        RECT 83.345 82.180 83.635 82.225 ;
        RECT 94.460 82.180 94.600 82.380 ;
        RECT 83.345 82.040 94.600 82.180 ;
        RECT 95.075 82.180 95.365 82.225 ;
        RECT 96.210 82.180 96.530 82.240 ;
        RECT 95.075 82.040 96.530 82.180 ;
        RECT 99.060 82.180 99.200 82.380 ;
        RECT 99.445 82.380 102.495 82.520 ;
        RECT 99.445 82.335 99.735 82.380 ;
        RECT 102.205 82.335 102.495 82.380 ;
        RECT 102.740 82.380 105.255 82.520 ;
        RECT 102.740 82.180 102.880 82.380 ;
        RECT 104.965 82.335 105.255 82.380 ;
        RECT 99.060 82.040 102.880 82.180 ;
        RECT 83.345 81.995 83.635 82.040 ;
        RECT 95.075 81.995 95.365 82.040 ;
        RECT 96.210 81.980 96.530 82.040 ;
        RECT 104.490 81.980 104.810 82.240 ;
        RECT 107.265 82.180 107.555 82.225 ;
        RECT 108.630 82.180 108.950 82.240 ;
        RECT 107.265 82.040 108.950 82.180 ;
        RECT 107.265 81.995 107.555 82.040 ;
        RECT 108.630 81.980 108.950 82.040 ;
        RECT 5.520 81.360 125.580 81.840 ;
        RECT 11.585 80.975 11.875 81.205 ;
        RECT 13.885 81.160 14.175 81.205 ;
        RECT 15.710 81.160 16.030 81.220 ;
        RECT 13.885 81.020 16.030 81.160 ;
        RECT 13.885 80.975 14.175 81.020 ;
        RECT 11.660 80.820 11.800 80.975 ;
        RECT 15.710 80.960 16.030 81.020 ;
        RECT 17.565 81.160 17.855 81.205 ;
        RECT 28.590 81.160 28.910 81.220 ;
        RECT 34.570 81.160 34.890 81.220 ;
        RECT 35.505 81.160 35.795 81.205 ;
        RECT 17.565 81.020 28.360 81.160 ;
        RECT 17.565 80.975 17.855 81.020 ;
        RECT 9.820 80.680 11.800 80.820 ;
        RECT 13.425 80.820 13.715 80.865 ;
        RECT 18.025 80.820 18.315 80.865 ;
        RECT 18.930 80.820 19.250 80.880 ;
        RECT 13.425 80.680 19.250 80.820 ;
        RECT 9.820 80.525 9.960 80.680 ;
        RECT 13.425 80.635 13.715 80.680 ;
        RECT 18.025 80.635 18.315 80.680 ;
        RECT 18.930 80.620 19.250 80.680 ;
        RECT 20.770 80.820 21.090 80.880 ;
        RECT 24.465 80.820 24.755 80.865 ;
        RECT 24.925 80.820 25.215 80.865 ;
        RECT 20.770 80.680 22.840 80.820 ;
        RECT 20.770 80.620 21.090 80.680 ;
        RECT 9.745 80.295 10.035 80.525 ;
        RECT 11.125 80.295 11.415 80.525 ;
        RECT 20.310 80.480 20.630 80.540 ;
        RECT 21.245 80.480 21.535 80.525 ;
        RECT 20.310 80.340 21.535 80.480 ;
        RECT 8.350 79.800 8.670 79.860 ;
        RECT 10.205 79.800 10.495 79.845 ;
        RECT 8.350 79.660 10.495 79.800 ;
        RECT 11.200 79.800 11.340 80.295 ;
        RECT 20.310 80.280 20.630 80.340 ;
        RECT 21.245 80.295 21.535 80.340 ;
        RECT 21.690 80.480 22.010 80.540 ;
        RECT 22.700 80.525 22.840 80.680 ;
        RECT 24.465 80.680 25.215 80.820 ;
        RECT 28.220 80.820 28.360 81.020 ;
        RECT 28.590 81.020 30.200 81.160 ;
        RECT 28.590 80.960 28.910 81.020 ;
        RECT 30.060 80.865 30.200 81.020 ;
        RECT 34.570 81.020 35.795 81.160 ;
        RECT 34.570 80.960 34.890 81.020 ;
        RECT 35.505 80.975 35.795 81.020 ;
        RECT 39.185 81.160 39.475 81.205 ;
        RECT 47.910 81.160 48.230 81.220 ;
        RECT 39.185 81.020 48.230 81.160 ;
        RECT 39.185 80.975 39.475 81.020 ;
        RECT 47.910 80.960 48.230 81.020 ;
        RECT 48.370 80.960 48.690 81.220 ;
        RECT 61.250 80.960 61.570 81.220 ;
        RECT 77.810 81.205 78.130 81.220 ;
        RECT 66.785 81.160 67.075 81.205 ;
        RECT 66.785 81.020 77.120 81.160 ;
        RECT 66.785 80.975 67.075 81.020 ;
        RECT 28.220 80.680 29.280 80.820 ;
        RECT 24.465 80.635 24.755 80.680 ;
        RECT 24.925 80.635 25.215 80.680 ;
        RECT 22.165 80.480 22.455 80.525 ;
        RECT 21.690 80.340 22.455 80.480 ;
        RECT 21.690 80.280 22.010 80.340 ;
        RECT 22.165 80.295 22.455 80.340 ;
        RECT 22.625 80.295 22.915 80.525 ;
        RECT 23.070 80.280 23.390 80.540 ;
        RECT 23.530 80.480 23.850 80.540 ;
        RECT 26.305 80.480 26.595 80.525 ;
        RECT 23.530 80.340 26.595 80.480 ;
        RECT 23.530 80.280 23.850 80.340 ;
        RECT 26.305 80.295 26.595 80.340 ;
        RECT 27.210 80.280 27.530 80.540 ;
        RECT 28.590 80.280 28.910 80.540 ;
        RECT 29.140 80.480 29.280 80.680 ;
        RECT 29.985 80.635 30.275 80.865 ;
        RECT 30.890 80.820 31.210 80.880 ;
        RECT 39.645 80.820 39.935 80.865 ;
        RECT 30.890 80.680 39.935 80.820 ;
        RECT 30.890 80.620 31.210 80.680 ;
        RECT 39.645 80.635 39.935 80.680 ;
        RECT 41.930 80.820 42.250 80.880 ;
        RECT 66.860 80.820 67.000 80.975 ;
        RECT 41.930 80.680 67.000 80.820 ;
        RECT 69.550 80.820 69.840 80.865 ;
        RECT 71.410 80.820 71.700 80.865 ;
        RECT 69.550 80.680 71.700 80.820 ;
        RECT 41.930 80.620 42.250 80.680 ;
        RECT 69.550 80.635 69.840 80.680 ;
        RECT 71.410 80.635 71.700 80.680 ;
        RECT 72.330 80.820 72.620 80.865 ;
        RECT 74.130 80.820 74.450 80.880 ;
        RECT 75.590 80.820 75.880 80.865 ;
        RECT 72.330 80.680 75.880 80.820 ;
        RECT 76.980 80.820 77.120 81.020 ;
        RECT 77.595 80.975 78.130 81.205 ;
        RECT 81.490 81.160 81.810 81.220 ;
        RECT 77.810 80.960 78.130 80.975 ;
        RECT 81.120 81.020 81.810 81.160 ;
        RECT 81.120 80.820 81.260 81.020 ;
        RECT 81.490 80.960 81.810 81.020 ;
        RECT 82.410 81.160 82.730 81.220 ;
        RECT 83.345 81.160 83.635 81.205 ;
        RECT 82.410 81.020 83.635 81.160 ;
        RECT 82.410 80.960 82.730 81.020 ;
        RECT 83.345 80.975 83.635 81.020 ;
        RECT 87.945 81.160 88.235 81.205 ;
        RECT 88.850 81.160 89.170 81.220 ;
        RECT 87.945 81.020 89.170 81.160 ;
        RECT 87.945 80.975 88.235 81.020 ;
        RECT 88.850 80.960 89.170 81.020 ;
        RECT 89.785 81.160 90.075 81.205 ;
        RECT 92.070 81.160 92.390 81.220 ;
        RECT 89.785 81.020 92.390 81.160 ;
        RECT 89.785 80.975 90.075 81.020 ;
        RECT 92.070 80.960 92.390 81.020 ;
        RECT 92.530 80.960 92.850 81.220 ;
        RECT 98.985 81.160 99.275 81.205 ;
        RECT 108.170 81.160 108.490 81.220 ;
        RECT 98.985 81.020 108.490 81.160 ;
        RECT 98.985 80.975 99.275 81.020 ;
        RECT 108.170 80.960 108.490 81.020 ;
        RECT 85.185 80.820 85.475 80.865 ;
        RECT 90.245 80.820 90.535 80.865 ;
        RECT 96.210 80.820 96.530 80.880 ;
        RECT 76.980 80.680 84.940 80.820 ;
        RECT 72.330 80.635 72.620 80.680 ;
        RECT 30.980 80.480 31.120 80.620 ;
        RECT 29.140 80.340 31.120 80.480 ;
        RECT 36.425 80.480 36.715 80.525 ;
        RECT 43.310 80.480 43.630 80.540 ;
        RECT 47.925 80.480 48.215 80.525 ;
        RECT 36.425 80.340 37.560 80.480 ;
        RECT 36.425 80.295 36.715 80.340 ;
        RECT 14.805 80.140 15.095 80.185 ;
        RECT 17.090 80.140 17.410 80.200 ;
        RECT 18.485 80.140 18.775 80.185 ;
        RECT 14.805 80.000 18.775 80.140 ;
        RECT 14.805 79.955 15.095 80.000 ;
        RECT 17.090 79.940 17.410 80.000 ;
        RECT 18.485 79.955 18.775 80.000 ;
        RECT 25.845 80.140 26.135 80.185 ;
        RECT 27.300 80.140 27.440 80.280 ;
        RECT 25.845 80.000 27.440 80.140 ;
        RECT 25.845 79.955 26.135 80.000 ;
        RECT 29.050 79.940 29.370 80.200 ;
        RECT 15.725 79.800 16.015 79.845 ;
        RECT 27.225 79.800 27.515 79.845 ;
        RECT 11.200 79.660 16.015 79.800 ;
        RECT 8.350 79.600 8.670 79.660 ;
        RECT 10.205 79.615 10.495 79.660 ;
        RECT 15.725 79.615 16.015 79.660 ;
        RECT 20.400 79.660 27.515 79.800 ;
        RECT 8.810 79.260 9.130 79.520 ;
        RECT 12.490 79.460 12.810 79.520 ;
        RECT 20.400 79.460 20.540 79.660 ;
        RECT 27.225 79.615 27.515 79.660 ;
        RECT 27.685 79.800 27.975 79.845 ;
        RECT 32.270 79.800 32.590 79.860 ;
        RECT 37.420 79.845 37.560 80.340 ;
        RECT 43.310 80.340 48.215 80.480 ;
        RECT 43.310 80.280 43.630 80.340 ;
        RECT 47.925 80.295 48.215 80.340 ;
        RECT 61.725 80.480 62.015 80.525 ;
        RECT 62.630 80.480 62.950 80.540 ;
        RECT 61.725 80.340 62.950 80.480 ;
        RECT 61.725 80.295 62.015 80.340 ;
        RECT 62.630 80.280 62.950 80.340 ;
        RECT 63.565 80.480 63.855 80.525 ;
        RECT 65.390 80.480 65.710 80.540 ;
        RECT 63.565 80.340 65.710 80.480 ;
        RECT 63.565 80.295 63.855 80.340 ;
        RECT 65.390 80.280 65.710 80.340 ;
        RECT 65.850 80.280 66.170 80.540 ;
        RECT 70.450 80.280 70.770 80.540 ;
        RECT 71.485 80.480 71.700 80.635 ;
        RECT 74.130 80.620 74.450 80.680 ;
        RECT 75.590 80.635 75.880 80.680 ;
        RECT 73.730 80.480 74.020 80.525 ;
        RECT 71.485 80.340 74.020 80.480 ;
        RECT 73.730 80.295 74.020 80.340 ;
        RECT 80.570 80.280 80.890 80.540 ;
        RECT 81.120 80.525 81.260 80.680 ;
        RECT 81.045 80.295 81.335 80.525 ;
        RECT 81.505 80.295 81.795 80.525 ;
        RECT 39.170 80.140 39.490 80.200 ;
        RECT 40.105 80.140 40.395 80.185 ;
        RECT 39.170 80.000 40.395 80.140 ;
        RECT 39.170 79.940 39.490 80.000 ;
        RECT 40.105 79.955 40.395 80.000 ;
        RECT 62.185 79.955 62.475 80.185 ;
        RECT 63.105 80.140 63.395 80.185 ;
        RECT 65.940 80.140 66.080 80.280 ;
        RECT 63.105 80.000 66.080 80.140 ;
        RECT 63.105 79.955 63.395 80.000 ;
        RECT 27.685 79.660 32.590 79.800 ;
        RECT 27.685 79.615 27.975 79.660 ;
        RECT 32.270 79.600 32.590 79.660 ;
        RECT 37.345 79.615 37.635 79.845 ;
        RECT 62.260 79.800 62.400 79.955 ;
        RECT 68.610 79.940 68.930 80.200 ;
        RECT 71.370 80.140 71.690 80.200 ;
        RECT 79.205 80.140 79.495 80.185 ;
        RECT 81.580 80.140 81.720 80.295 ;
        RECT 82.410 80.280 82.730 80.540 ;
        RECT 84.800 80.480 84.940 80.680 ;
        RECT 85.185 80.680 96.530 80.820 ;
        RECT 85.185 80.635 85.475 80.680 ;
        RECT 90.245 80.635 90.535 80.680 ;
        RECT 96.210 80.620 96.530 80.680 ;
        RECT 91.610 80.480 91.930 80.540 ;
        RECT 84.800 80.340 91.930 80.480 ;
        RECT 91.610 80.280 91.930 80.340 ;
        RECT 93.005 80.480 93.295 80.525 ;
        RECT 94.370 80.480 94.690 80.540 ;
        RECT 93.005 80.340 94.690 80.480 ;
        RECT 93.005 80.295 93.295 80.340 ;
        RECT 94.370 80.280 94.690 80.340 ;
        RECT 96.670 80.280 96.990 80.540 ;
        RECT 98.065 80.295 98.355 80.525 ;
        RECT 81.950 80.140 82.270 80.200 ;
        RECT 85.645 80.140 85.935 80.185 ;
        RECT 71.370 80.000 81.260 80.140 ;
        RECT 81.580 80.000 85.935 80.140 ;
        RECT 71.370 79.940 71.690 80.000 ;
        RECT 79.205 79.955 79.495 80.000 ;
        RECT 64.010 79.800 64.330 79.860 ;
        RECT 62.260 79.660 64.330 79.800 ;
        RECT 64.010 79.600 64.330 79.660 ;
        RECT 69.090 79.800 69.380 79.845 ;
        RECT 70.950 79.800 71.240 79.845 ;
        RECT 73.730 79.800 74.020 79.845 ;
        RECT 69.090 79.660 74.020 79.800 ;
        RECT 81.120 79.800 81.260 80.000 ;
        RECT 81.950 79.940 82.270 80.000 ;
        RECT 85.645 79.955 85.935 80.000 ;
        RECT 86.090 80.140 86.410 80.200 ;
        RECT 90.705 80.140 90.995 80.185 ;
        RECT 86.090 80.000 90.995 80.140 ;
        RECT 86.090 79.940 86.410 80.000 ;
        RECT 90.705 79.955 90.995 80.000 ;
        RECT 97.130 79.940 97.450 80.200 ;
        RECT 98.140 80.140 98.280 80.295 ;
        RECT 97.680 80.000 98.280 80.140 ;
        RECT 97.680 79.800 97.820 80.000 ;
        RECT 105.410 79.800 105.730 79.860 ;
        RECT 81.120 79.660 97.820 79.800 ;
        RECT 98.140 79.660 105.730 79.800 ;
        RECT 69.090 79.615 69.380 79.660 ;
        RECT 70.950 79.615 71.240 79.660 ;
        RECT 73.730 79.615 74.020 79.660 ;
        RECT 12.490 79.320 20.540 79.460 ;
        RECT 26.305 79.460 26.595 79.505 ;
        RECT 26.750 79.460 27.070 79.520 ;
        RECT 26.305 79.320 27.070 79.460 ;
        RECT 12.490 79.260 12.810 79.320 ;
        RECT 26.305 79.275 26.595 79.320 ;
        RECT 26.750 79.260 27.070 79.320 ;
        RECT 29.985 79.460 30.275 79.505 ;
        RECT 31.350 79.460 31.670 79.520 ;
        RECT 29.985 79.320 31.670 79.460 ;
        RECT 29.985 79.275 30.275 79.320 ;
        RECT 31.350 79.260 31.670 79.320 ;
        RECT 35.490 79.460 35.810 79.520 ;
        RECT 64.485 79.460 64.775 79.505 ;
        RECT 80.570 79.460 80.890 79.520 ;
        RECT 35.490 79.320 80.890 79.460 ;
        RECT 35.490 79.260 35.810 79.320 ;
        RECT 64.485 79.275 64.775 79.320 ;
        RECT 80.570 79.260 80.890 79.320 ;
        RECT 87.930 79.460 88.250 79.520 ;
        RECT 89.310 79.460 89.630 79.520 ;
        RECT 98.140 79.505 98.280 79.660 ;
        RECT 105.410 79.600 105.730 79.660 ;
        RECT 87.930 79.320 89.630 79.460 ;
        RECT 87.930 79.260 88.250 79.320 ;
        RECT 89.310 79.260 89.630 79.320 ;
        RECT 98.065 79.275 98.355 79.505 ;
        RECT 5.520 78.640 125.580 79.120 ;
        RECT 15.710 78.440 16.030 78.500 ;
        RECT 16.415 78.440 16.705 78.485 ;
        RECT 15.710 78.300 16.705 78.440 ;
        RECT 15.710 78.240 16.030 78.300 ;
        RECT 16.415 78.255 16.705 78.300 ;
        RECT 18.930 78.240 19.250 78.500 ;
        RECT 72.290 78.440 72.610 78.500 ;
        RECT 81.950 78.485 82.270 78.500 ;
        RECT 72.290 78.300 81.260 78.440 ;
        RECT 72.290 78.240 72.610 78.300 ;
        RECT 7.910 78.100 8.200 78.145 ;
        RECT 9.770 78.100 10.060 78.145 ;
        RECT 12.550 78.100 12.840 78.145 ;
        RECT 7.910 77.960 12.840 78.100 ;
        RECT 7.910 77.915 8.200 77.960 ;
        RECT 9.770 77.915 10.060 77.960 ;
        RECT 12.550 77.915 12.840 77.960 ;
        RECT 73.230 78.100 73.520 78.145 ;
        RECT 75.090 78.100 75.380 78.145 ;
        RECT 77.870 78.100 78.160 78.145 ;
        RECT 73.230 77.960 78.160 78.100 ;
        RECT 81.120 78.100 81.260 78.300 ;
        RECT 81.735 78.255 82.270 78.485 ;
        RECT 81.950 78.240 82.270 78.255 ;
        RECT 103.570 78.440 103.890 78.500 ;
        RECT 104.505 78.440 104.795 78.485 ;
        RECT 103.570 78.300 104.795 78.440 ;
        RECT 103.570 78.240 103.890 78.300 ;
        RECT 104.505 78.255 104.795 78.300 ;
        RECT 86.090 78.100 86.410 78.160 ;
        RECT 81.120 77.960 86.410 78.100 ;
        RECT 73.230 77.915 73.520 77.960 ;
        RECT 75.090 77.915 75.380 77.960 ;
        RECT 77.870 77.915 78.160 77.960 ;
        RECT 86.090 77.900 86.410 77.960 ;
        RECT 104.030 78.100 104.350 78.160 ;
        RECT 104.965 78.100 105.255 78.145 ;
        RECT 104.030 77.960 105.255 78.100 ;
        RECT 104.030 77.900 104.350 77.960 ;
        RECT 104.965 77.915 105.255 77.960 ;
        RECT 111.405 77.915 111.695 78.145 ;
        RECT 112.330 78.100 112.620 78.145 ;
        RECT 114.190 78.100 114.480 78.145 ;
        RECT 116.970 78.100 117.260 78.145 ;
        RECT 112.330 77.960 117.260 78.100 ;
        RECT 112.330 77.915 112.620 77.960 ;
        RECT 114.190 77.915 114.480 77.960 ;
        RECT 116.970 77.915 117.260 77.960 ;
        RECT 8.810 77.760 9.130 77.820 ;
        RECT 9.285 77.760 9.575 77.805 ;
        RECT 68.610 77.760 68.930 77.820 ;
        RECT 72.765 77.760 73.055 77.805 ;
        RECT 82.870 77.760 83.190 77.820 ;
        RECT 111.480 77.760 111.620 77.915 ;
        RECT 113.705 77.760 113.995 77.805 ;
        RECT 8.810 77.620 9.575 77.760 ;
        RECT 8.810 77.560 9.130 77.620 ;
        RECT 9.285 77.575 9.575 77.620 ;
        RECT 18.100 77.620 23.760 77.760 ;
        RECT 18.100 77.480 18.240 77.620 ;
        RECT 7.430 77.220 7.750 77.480 ;
        RECT 12.550 77.420 12.840 77.465 ;
        RECT 10.305 77.280 12.840 77.420 ;
        RECT 10.305 77.125 10.520 77.280 ;
        RECT 12.550 77.235 12.840 77.280 ;
        RECT 18.010 77.220 18.330 77.480 ;
        RECT 21.690 77.220 22.010 77.480 ;
        RECT 23.620 77.465 23.760 77.620 ;
        RECT 68.610 77.620 83.190 77.760 ;
        RECT 68.610 77.560 68.930 77.620 ;
        RECT 72.765 77.575 73.055 77.620 ;
        RECT 82.870 77.560 83.190 77.620 ;
        RECT 101.360 77.620 108.400 77.760 ;
        RECT 111.480 77.620 113.995 77.760 ;
        RECT 101.360 77.480 101.500 77.620 ;
        RECT 23.545 77.235 23.835 77.465 ;
        RECT 63.090 77.220 63.410 77.480 ;
        RECT 74.605 77.420 74.895 77.465 ;
        RECT 75.050 77.420 75.370 77.480 ;
        RECT 77.870 77.420 78.160 77.465 ;
        RECT 74.605 77.280 75.370 77.420 ;
        RECT 74.605 77.235 74.895 77.280 ;
        RECT 75.050 77.220 75.370 77.280 ;
        RECT 75.625 77.280 78.160 77.420 ;
        RECT 75.625 77.125 75.840 77.280 ;
        RECT 77.870 77.235 78.160 77.280 ;
        RECT 82.410 77.420 82.730 77.480 ;
        RECT 101.270 77.420 101.590 77.480 ;
        RECT 82.410 77.280 101.590 77.420 ;
        RECT 82.410 77.220 82.730 77.280 ;
        RECT 101.270 77.220 101.590 77.280 ;
        RECT 102.190 77.220 102.510 77.480 ;
        RECT 102.665 77.235 102.955 77.465 ;
        RECT 103.110 77.420 103.430 77.480 ;
        RECT 104.490 77.420 104.810 77.480 ;
        RECT 108.260 77.465 108.400 77.620 ;
        RECT 113.705 77.575 113.995 77.620 ;
        RECT 106.345 77.420 106.635 77.465 ;
        RECT 103.110 77.280 106.635 77.420 ;
        RECT 8.370 77.080 8.660 77.125 ;
        RECT 10.230 77.080 10.520 77.125 ;
        RECT 8.370 76.940 10.520 77.080 ;
        RECT 8.370 76.895 8.660 76.940 ;
        RECT 10.230 76.895 10.520 76.940 ;
        RECT 11.150 77.080 11.440 77.125 ;
        RECT 14.410 77.080 14.700 77.125 ;
        RECT 17.565 77.080 17.855 77.125 ;
        RECT 11.150 76.940 17.855 77.080 ;
        RECT 11.150 76.895 11.440 76.940 ;
        RECT 14.410 76.895 14.700 76.940 ;
        RECT 17.565 76.895 17.855 76.940 ;
        RECT 73.690 77.080 73.980 77.125 ;
        RECT 75.550 77.080 75.840 77.125 ;
        RECT 73.690 76.940 75.840 77.080 ;
        RECT 73.690 76.895 73.980 76.940 ;
        RECT 75.550 76.895 75.840 76.940 ;
        RECT 76.470 77.080 76.760 77.125 ;
        RECT 78.270 77.080 78.590 77.140 ;
        RECT 79.730 77.080 80.020 77.125 ;
        RECT 76.470 76.940 80.020 77.080 ;
        RECT 76.470 76.895 76.760 76.940 ;
        RECT 78.270 76.880 78.590 76.940 ;
        RECT 79.730 76.895 80.020 76.940 ;
        RECT 100.810 77.080 101.130 77.140 ;
        RECT 102.740 77.080 102.880 77.235 ;
        RECT 103.110 77.220 103.430 77.280 ;
        RECT 104.490 77.220 104.810 77.280 ;
        RECT 106.345 77.235 106.635 77.280 ;
        RECT 106.805 77.235 107.095 77.465 ;
        RECT 107.265 77.235 107.555 77.465 ;
        RECT 108.185 77.235 108.475 77.465 ;
        RECT 104.030 77.080 104.350 77.140 ;
        RECT 106.880 77.080 107.020 77.235 ;
        RECT 100.810 76.940 107.020 77.080 ;
        RECT 107.340 77.080 107.480 77.235 ;
        RECT 110.470 77.220 110.790 77.480 ;
        RECT 111.865 77.420 112.155 77.465 ;
        RECT 112.310 77.420 112.630 77.480 ;
        RECT 116.970 77.420 117.260 77.465 ;
        RECT 111.865 77.280 112.630 77.420 ;
        RECT 111.865 77.235 112.155 77.280 ;
        RECT 112.310 77.220 112.630 77.280 ;
        RECT 114.725 77.280 117.260 77.420 ;
        RECT 114.725 77.125 114.940 77.280 ;
        RECT 116.970 77.235 117.260 77.280 ;
        RECT 112.790 77.080 113.080 77.125 ;
        RECT 114.650 77.080 114.940 77.125 ;
        RECT 107.340 76.940 110.470 77.080 ;
        RECT 100.810 76.880 101.130 76.940 ;
        RECT 104.030 76.880 104.350 76.940 ;
        RECT 23.070 76.540 23.390 76.800 ;
        RECT 34.570 76.740 34.890 76.800 ;
        RECT 64.025 76.740 64.315 76.785 ;
        RECT 82.410 76.740 82.730 76.800 ;
        RECT 34.570 76.600 82.730 76.740 ;
        RECT 110.330 76.740 110.470 76.940 ;
        RECT 112.790 76.940 114.940 77.080 ;
        RECT 112.790 76.895 113.080 76.940 ;
        RECT 114.650 76.895 114.940 76.940 ;
        RECT 115.570 77.080 115.860 77.125 ;
        RECT 117.370 77.080 117.690 77.140 ;
        RECT 118.830 77.080 119.120 77.125 ;
        RECT 115.570 76.940 119.120 77.080 ;
        RECT 115.570 76.895 115.860 76.940 ;
        RECT 117.370 76.880 117.690 76.940 ;
        RECT 118.830 76.895 119.120 76.940 ;
        RECT 114.150 76.740 114.470 76.800 ;
        RECT 120.835 76.740 121.125 76.785 ;
        RECT 110.330 76.600 121.125 76.740 ;
        RECT 34.570 76.540 34.890 76.600 ;
        RECT 64.025 76.555 64.315 76.600 ;
        RECT 82.410 76.540 82.730 76.600 ;
        RECT 114.150 76.540 114.470 76.600 ;
        RECT 120.835 76.555 121.125 76.600 ;
        RECT 5.520 75.920 125.580 76.400 ;
        RECT 8.350 75.720 8.670 75.780 ;
        RECT 17.105 75.720 17.395 75.765 ;
        RECT 21.690 75.720 22.010 75.780 ;
        RECT 8.350 75.580 9.960 75.720 ;
        RECT 8.350 75.520 8.670 75.580 ;
        RECT 9.820 75.425 9.960 75.580 ;
        RECT 17.105 75.580 22.010 75.720 ;
        RECT 17.105 75.535 17.395 75.580 ;
        RECT 21.690 75.520 22.010 75.580 ;
        RECT 23.530 75.520 23.850 75.780 ;
        RECT 25.370 75.720 25.690 75.780 ;
        RECT 27.225 75.720 27.515 75.765 ;
        RECT 28.590 75.720 28.910 75.780 ;
        RECT 25.370 75.580 26.060 75.720 ;
        RECT 25.370 75.520 25.690 75.580 ;
        RECT 9.745 75.195 10.035 75.425 ;
        RECT 12.025 75.380 12.675 75.425 ;
        RECT 15.625 75.380 15.915 75.425 ;
        RECT 23.070 75.380 23.390 75.440 ;
        RECT 24.450 75.380 24.770 75.440 ;
        RECT 12.025 75.240 23.390 75.380 ;
        RECT 12.025 75.195 12.675 75.240 ;
        RECT 15.325 75.195 15.915 75.240 ;
        RECT 7.430 75.040 7.750 75.100 ;
        RECT 8.365 75.040 8.655 75.085 ;
        RECT 7.430 74.900 8.655 75.040 ;
        RECT 7.430 74.840 7.750 74.900 ;
        RECT 8.365 74.855 8.655 74.900 ;
        RECT 8.830 75.040 9.120 75.085 ;
        RECT 10.665 75.040 10.955 75.085 ;
        RECT 14.245 75.040 14.535 75.085 ;
        RECT 8.830 74.900 14.535 75.040 ;
        RECT 8.830 74.855 9.120 74.900 ;
        RECT 10.665 74.855 10.955 74.900 ;
        RECT 14.245 74.855 14.535 74.900 ;
        RECT 15.325 74.880 15.615 75.195 ;
        RECT 23.070 75.180 23.390 75.240 ;
        RECT 23.620 75.240 24.770 75.380 ;
        RECT 25.920 75.380 26.060 75.580 ;
        RECT 27.225 75.580 28.910 75.720 ;
        RECT 27.225 75.535 27.515 75.580 ;
        RECT 28.590 75.520 28.910 75.580 ;
        RECT 29.510 75.720 29.830 75.780 ;
        RECT 30.905 75.720 31.195 75.765 ;
        RECT 35.950 75.720 36.270 75.780 ;
        RECT 29.510 75.580 31.195 75.720 ;
        RECT 29.510 75.520 29.830 75.580 ;
        RECT 30.905 75.535 31.195 75.580 ;
        RECT 31.440 75.580 36.270 75.720 ;
        RECT 31.440 75.380 31.580 75.580 ;
        RECT 35.950 75.520 36.270 75.580 ;
        RECT 37.805 75.720 38.095 75.765 ;
        RECT 38.710 75.720 39.030 75.780 ;
        RECT 37.805 75.580 39.030 75.720 ;
        RECT 37.805 75.535 38.095 75.580 ;
        RECT 38.710 75.520 39.030 75.580 ;
        RECT 56.665 75.720 56.955 75.765 ;
        RECT 57.110 75.720 57.430 75.780 ;
        RECT 56.665 75.580 57.430 75.720 ;
        RECT 56.665 75.535 56.955 75.580 ;
        RECT 57.110 75.520 57.430 75.580 ;
        RECT 57.585 75.720 57.875 75.765 ;
        RECT 58.030 75.720 58.350 75.780 ;
        RECT 59.870 75.720 60.190 75.780 ;
        RECT 57.585 75.580 58.350 75.720 ;
        RECT 57.585 75.535 57.875 75.580 ;
        RECT 58.030 75.520 58.350 75.580 ;
        RECT 59.040 75.580 60.190 75.720 ;
        RECT 40.105 75.380 40.395 75.425 ;
        RECT 25.920 75.240 31.580 75.380 ;
        RECT 35.580 75.240 40.395 75.380 ;
        RECT 16.170 75.040 16.490 75.100 ;
        RECT 18.485 75.040 18.775 75.085 ;
        RECT 16.170 74.900 18.775 75.040 ;
        RECT 16.170 74.840 16.490 74.900 ;
        RECT 18.485 74.855 18.775 74.900 ;
        RECT 19.850 74.840 20.170 75.100 ;
        RECT 20.310 74.840 20.630 75.100 ;
        RECT 21.245 74.855 21.535 75.085 ;
        RECT 21.705 74.855 21.995 75.085 ;
        RECT 22.165 75.040 22.455 75.085 ;
        RECT 23.620 75.040 23.760 75.240 ;
        RECT 24.450 75.180 24.770 75.240 ;
        RECT 22.165 74.900 23.760 75.040 ;
        RECT 22.165 74.855 22.455 74.900 ;
        RECT 24.005 74.855 24.295 75.085 ;
        RECT 9.235 74.360 9.525 74.405 ;
        RECT 11.125 74.360 11.415 74.405 ;
        RECT 14.245 74.360 14.535 74.405 ;
        RECT 9.235 74.220 14.535 74.360 ;
        RECT 9.235 74.175 9.525 74.220 ;
        RECT 11.125 74.175 11.415 74.220 ;
        RECT 14.245 74.175 14.535 74.220 ;
        RECT 16.170 74.360 16.490 74.420 ;
        RECT 21.320 74.360 21.460 74.855 ;
        RECT 21.780 74.700 21.920 74.855 ;
        RECT 23.070 74.700 23.390 74.760 ;
        RECT 21.780 74.560 23.390 74.700 ;
        RECT 23.070 74.500 23.390 74.560 ;
        RECT 16.170 74.220 21.460 74.360 ;
        RECT 23.530 74.360 23.850 74.420 ;
        RECT 24.080 74.360 24.220 74.855 ;
        RECT 24.910 74.840 25.230 75.100 ;
        RECT 25.370 74.840 25.690 75.100 ;
        RECT 25.845 74.855 26.135 75.085 ;
        RECT 27.715 75.070 28.005 75.085 ;
        RECT 27.715 74.930 28.360 75.070 ;
        RECT 27.715 74.855 28.005 74.930 ;
        RECT 24.450 74.700 24.770 74.760 ;
        RECT 25.920 74.700 26.060 74.855 ;
        RECT 24.450 74.560 26.060 74.700 ;
        RECT 24.450 74.500 24.770 74.560 ;
        RECT 28.220 74.360 28.360 74.930 ;
        RECT 28.590 74.840 28.910 75.100 ;
        RECT 29.140 75.085 29.280 75.240 ;
        RECT 29.065 74.855 29.355 75.085 ;
        RECT 29.525 75.055 29.815 75.085 ;
        RECT 29.525 75.040 30.660 75.055 ;
        RECT 29.525 74.915 31.120 75.040 ;
        RECT 29.525 74.855 29.815 74.915 ;
        RECT 30.520 74.900 31.120 74.915 ;
        RECT 30.980 74.760 31.120 74.900 ;
        RECT 34.570 74.840 34.890 75.100 ;
        RECT 35.030 75.040 35.350 75.100 ;
        RECT 35.580 75.085 35.720 75.240 ;
        RECT 40.105 75.195 40.395 75.240 ;
        RECT 40.565 75.380 40.855 75.425 ;
        RECT 52.050 75.380 52.370 75.440 ;
        RECT 59.040 75.380 59.180 75.580 ;
        RECT 59.870 75.520 60.190 75.580 ;
        RECT 64.010 75.720 64.330 75.780 ;
        RECT 93.910 75.720 94.230 75.780 ;
        RECT 94.385 75.720 94.675 75.765 ;
        RECT 64.010 75.580 93.680 75.720 ;
        RECT 64.010 75.520 64.330 75.580 ;
        RECT 61.250 75.380 61.570 75.440 ;
        RECT 40.565 75.240 54.580 75.380 ;
        RECT 40.565 75.195 40.855 75.240 ;
        RECT 52.050 75.180 52.370 75.240 ;
        RECT 35.505 75.040 35.795 75.085 ;
        RECT 35.030 74.900 35.795 75.040 ;
        RECT 35.030 74.840 35.350 74.900 ;
        RECT 35.505 74.855 35.795 74.900 ;
        RECT 35.950 74.840 36.270 75.100 ;
        RECT 36.425 74.855 36.715 75.085 ;
        RECT 43.770 75.040 44.090 75.100 ;
        RECT 47.450 75.040 47.770 75.100 ;
        RECT 49.305 75.040 49.595 75.085 ;
        RECT 43.770 74.900 49.595 75.040 ;
        RECT 30.890 74.700 31.210 74.760 ;
        RECT 36.500 74.700 36.640 74.855 ;
        RECT 43.770 74.840 44.090 74.900 ;
        RECT 47.450 74.840 47.770 74.900 ;
        RECT 49.305 74.855 49.595 74.900 ;
        RECT 53.445 75.040 53.735 75.085 ;
        RECT 53.890 75.040 54.210 75.100 ;
        RECT 54.440 75.085 54.580 75.240 ;
        RECT 54.900 75.240 59.640 75.380 ;
        RECT 54.900 75.085 55.040 75.240 ;
        RECT 53.445 74.900 54.210 75.040 ;
        RECT 53.445 74.855 53.735 74.900 ;
        RECT 53.890 74.840 54.210 74.900 ;
        RECT 54.365 74.855 54.655 75.085 ;
        RECT 54.825 74.855 55.115 75.085 ;
        RECT 55.285 75.040 55.575 75.085 ;
        RECT 58.490 75.040 58.810 75.100 ;
        RECT 59.500 75.085 59.640 75.240 ;
        RECT 59.960 75.240 61.570 75.380 ;
        RECT 59.960 75.085 60.100 75.240 ;
        RECT 61.250 75.180 61.570 75.240 ;
        RECT 64.930 75.180 65.250 75.440 ;
        RECT 73.670 75.180 73.990 75.440 ;
        RECT 93.540 75.380 93.680 75.580 ;
        RECT 93.910 75.580 94.675 75.720 ;
        RECT 93.910 75.520 94.230 75.580 ;
        RECT 94.385 75.535 94.675 75.580 ;
        RECT 96.210 75.720 96.530 75.780 ;
        RECT 96.685 75.720 96.975 75.765 ;
        RECT 96.210 75.580 96.975 75.720 ;
        RECT 96.210 75.520 96.530 75.580 ;
        RECT 96.685 75.535 96.975 75.580 ;
        RECT 103.110 75.520 103.430 75.780 ;
        RECT 105.885 75.720 106.175 75.765 ;
        RECT 106.330 75.720 106.650 75.780 ;
        RECT 105.885 75.580 106.650 75.720 ;
        RECT 105.885 75.535 106.175 75.580 ;
        RECT 106.330 75.520 106.650 75.580 ;
        RECT 110.470 75.720 110.790 75.780 ;
        RECT 113.245 75.720 113.535 75.765 ;
        RECT 110.470 75.580 113.535 75.720 ;
        RECT 110.470 75.520 110.790 75.580 ;
        RECT 113.245 75.535 113.535 75.580 ;
        RECT 116.925 75.720 117.215 75.765 ;
        RECT 117.370 75.720 117.690 75.780 ;
        RECT 116.925 75.580 117.690 75.720 ;
        RECT 116.925 75.535 117.215 75.580 ;
        RECT 117.370 75.520 117.690 75.580 ;
        RECT 103.200 75.380 103.340 75.520 ;
        RECT 93.180 75.240 103.340 75.380 ;
        RECT 58.965 75.040 59.255 75.085 ;
        RECT 55.285 74.900 59.255 75.040 ;
        RECT 55.285 74.855 55.575 74.900 ;
        RECT 58.490 74.840 58.810 74.900 ;
        RECT 58.965 74.855 59.255 74.900 ;
        RECT 59.425 74.855 59.715 75.085 ;
        RECT 59.885 74.855 60.175 75.085 ;
        RECT 60.790 75.040 61.110 75.100 ;
        RECT 62.170 75.040 62.490 75.100 ;
        RECT 60.790 74.900 62.490 75.040 ;
        RECT 60.790 74.840 61.110 74.900 ;
        RECT 62.170 74.840 62.490 74.900 ;
        RECT 91.150 74.840 91.470 75.100 ;
        RECT 92.070 74.840 92.390 75.100 ;
        RECT 93.180 75.085 93.320 75.240 ;
        RECT 92.545 74.855 92.835 75.085 ;
        RECT 93.005 74.915 93.320 75.085 ;
        RECT 100.810 75.040 101.130 75.100 ;
        RECT 93.005 74.855 93.295 74.915 ;
        RECT 93.540 74.900 101.130 75.040 ;
        RECT 30.890 74.560 36.640 74.700 ;
        RECT 30.890 74.500 31.210 74.560 ;
        RECT 34.570 74.360 34.890 74.420 ;
        RECT 23.530 74.220 34.890 74.360 ;
        RECT 36.500 74.360 36.640 74.560 ;
        RECT 39.170 74.700 39.490 74.760 ;
        RECT 41.025 74.700 41.315 74.745 ;
        RECT 39.170 74.560 41.315 74.700 ;
        RECT 39.170 74.500 39.490 74.560 ;
        RECT 41.025 74.515 41.315 74.560 ;
        RECT 67.690 74.700 68.010 74.760 ;
        RECT 92.620 74.700 92.760 74.855 ;
        RECT 93.540 74.700 93.680 74.900 ;
        RECT 100.810 74.840 101.130 74.900 ;
        RECT 101.270 75.040 101.590 75.100 ;
        RECT 102.665 75.040 102.955 75.085 ;
        RECT 103.480 75.055 103.770 75.100 ;
        RECT 101.270 74.900 102.955 75.040 ;
        RECT 101.270 74.840 101.590 74.900 ;
        RECT 102.665 74.855 102.955 74.900 ;
        RECT 103.200 74.915 103.770 75.055 ;
        RECT 67.690 74.560 93.680 74.700 ;
        RECT 93.910 74.700 94.230 74.760 ;
        RECT 97.590 74.700 97.910 74.760 ;
        RECT 99.445 74.700 99.735 74.745 ;
        RECT 93.910 74.560 99.735 74.700 ;
        RECT 103.200 74.700 103.340 74.915 ;
        RECT 103.480 74.870 103.770 74.915 ;
        RECT 104.030 74.840 104.350 75.100 ;
        RECT 104.490 75.085 104.810 75.100 ;
        RECT 104.490 74.855 104.895 75.085 ;
        RECT 104.490 74.840 104.810 74.855 ;
        RECT 111.390 74.840 111.710 75.100 ;
        RECT 116.465 75.040 116.755 75.085 ;
        RECT 117.370 75.040 117.690 75.100 ;
        RECT 116.465 74.900 117.690 75.040 ;
        RECT 116.465 74.855 116.755 74.900 ;
        RECT 117.370 74.840 117.690 74.900 ;
        RECT 118.750 74.840 119.070 75.100 ;
        RECT 110.010 74.700 110.330 74.760 ;
        RECT 103.200 74.560 110.330 74.700 ;
        RECT 67.690 74.500 68.010 74.560 ;
        RECT 93.910 74.500 94.230 74.560 ;
        RECT 97.590 74.500 97.910 74.560 ;
        RECT 99.445 74.515 99.735 74.560 ;
        RECT 110.010 74.500 110.330 74.560 ;
        RECT 110.470 74.500 110.790 74.760 ;
        RECT 110.945 74.700 111.235 74.745 ;
        RECT 114.150 74.700 114.470 74.760 ;
        RECT 110.945 74.560 114.470 74.700 ;
        RECT 110.945 74.515 111.235 74.560 ;
        RECT 114.150 74.500 114.470 74.560 ;
        RECT 81.030 74.360 81.350 74.420 ;
        RECT 98.970 74.360 99.290 74.420 ;
        RECT 36.500 74.220 54.580 74.360 ;
        RECT 16.170 74.160 16.490 74.220 ;
        RECT 23.530 74.160 23.850 74.220 ;
        RECT 34.570 74.160 34.890 74.220 ;
        RECT 20.310 74.020 20.630 74.080 ;
        RECT 23.620 74.020 23.760 74.160 ;
        RECT 20.310 73.880 23.760 74.020 ;
        RECT 33.190 74.020 33.510 74.080 ;
        RECT 38.265 74.020 38.555 74.065 ;
        RECT 33.190 73.880 38.555 74.020 ;
        RECT 20.310 73.820 20.630 73.880 ;
        RECT 33.190 73.820 33.510 73.880 ;
        RECT 38.265 73.835 38.555 73.880 ;
        RECT 49.750 73.820 50.070 74.080 ;
        RECT 54.440 74.020 54.580 74.220 ;
        RECT 81.030 74.220 99.290 74.360 ;
        RECT 81.030 74.160 81.350 74.220 ;
        RECT 98.970 74.160 99.290 74.220 ;
        RECT 102.190 74.360 102.510 74.420 ;
        RECT 103.570 74.360 103.890 74.420 ;
        RECT 102.190 74.220 103.890 74.360 ;
        RECT 102.190 74.160 102.510 74.220 ;
        RECT 103.570 74.160 103.890 74.220 ;
        RECT 64.010 74.020 64.330 74.080 ;
        RECT 54.440 73.880 64.330 74.020 ;
        RECT 64.010 73.820 64.330 73.880 ;
        RECT 71.830 74.020 72.150 74.080 ;
        RECT 74.590 74.020 74.910 74.080 ;
        RECT 103.110 74.020 103.430 74.080 ;
        RECT 71.830 73.880 103.430 74.020 ;
        RECT 71.830 73.820 72.150 73.880 ;
        RECT 74.590 73.820 74.910 73.880 ;
        RECT 103.110 73.820 103.430 73.880 ;
        RECT 113.690 74.020 114.010 74.080 ;
        RECT 117.845 74.020 118.135 74.065 ;
        RECT 113.690 73.880 118.135 74.020 ;
        RECT 113.690 73.820 114.010 73.880 ;
        RECT 117.845 73.835 118.135 73.880 ;
        RECT 5.520 73.200 125.580 73.680 ;
        RECT 23.545 73.000 23.835 73.045 ;
        RECT 23.990 73.000 24.310 73.060 ;
        RECT 23.545 72.860 24.310 73.000 ;
        RECT 23.545 72.815 23.835 72.860 ;
        RECT 23.990 72.800 24.310 72.860 ;
        RECT 27.225 73.000 27.515 73.045 ;
        RECT 27.670 73.000 27.990 73.060 ;
        RECT 27.225 72.860 27.990 73.000 ;
        RECT 27.225 72.815 27.515 72.860 ;
        RECT 27.670 72.800 27.990 72.860 ;
        RECT 43.555 73.000 43.845 73.045 ;
        RECT 52.050 73.000 52.370 73.060 ;
        RECT 43.555 72.860 52.370 73.000 ;
        RECT 43.555 72.815 43.845 72.860 ;
        RECT 52.050 72.800 52.370 72.860 ;
        RECT 58.950 72.800 59.270 73.060 ;
        RECT 59.410 72.800 59.730 73.060 ;
        RECT 68.610 73.000 68.930 73.060 ;
        RECT 61.800 72.860 68.930 73.000 ;
        RECT 24.450 72.660 24.770 72.720 ;
        RECT 35.050 72.660 35.340 72.705 ;
        RECT 36.910 72.660 37.200 72.705 ;
        RECT 39.690 72.660 39.980 72.705 ;
        RECT 24.450 72.520 26.060 72.660 ;
        RECT 24.450 72.460 24.770 72.520 ;
        RECT 23.070 72.320 23.390 72.380 ;
        RECT 21.780 72.180 25.600 72.320 ;
        RECT 20.310 71.780 20.630 72.040 ;
        RECT 21.780 72.025 21.920 72.180 ;
        RECT 23.070 72.120 23.390 72.180 ;
        RECT 25.460 72.040 25.600 72.180 ;
        RECT 21.245 71.795 21.535 72.025 ;
        RECT 21.705 71.795 21.995 72.025 ;
        RECT 22.165 71.795 22.455 72.025 ;
        RECT 23.530 71.980 23.850 72.040 ;
        RECT 24.005 71.980 24.295 72.025 ;
        RECT 23.530 71.840 24.295 71.980 ;
        RECT 18.010 71.640 18.330 71.700 ;
        RECT 21.320 71.640 21.460 71.795 ;
        RECT 18.010 71.500 21.460 71.640 ;
        RECT 22.240 71.640 22.380 71.795 ;
        RECT 23.530 71.780 23.850 71.840 ;
        RECT 24.005 71.795 24.295 71.840 ;
        RECT 24.450 71.980 24.770 72.040 ;
        RECT 24.925 71.980 25.215 72.025 ;
        RECT 24.450 71.840 25.215 71.980 ;
        RECT 24.450 71.780 24.770 71.840 ;
        RECT 24.925 71.795 25.215 71.840 ;
        RECT 25.370 71.780 25.690 72.040 ;
        RECT 25.920 72.025 26.060 72.520 ;
        RECT 35.050 72.520 39.980 72.660 ;
        RECT 35.050 72.475 35.340 72.520 ;
        RECT 36.910 72.475 37.200 72.520 ;
        RECT 39.690 72.475 39.980 72.520 ;
        RECT 46.550 72.660 46.840 72.705 ;
        RECT 48.410 72.660 48.700 72.705 ;
        RECT 51.190 72.660 51.480 72.705 ;
        RECT 46.550 72.520 51.480 72.660 ;
        RECT 46.550 72.475 46.840 72.520 ;
        RECT 48.410 72.475 48.700 72.520 ;
        RECT 51.190 72.475 51.480 72.520 ;
        RECT 52.510 72.660 52.830 72.720 ;
        RECT 55.055 72.660 55.345 72.705 ;
        RECT 61.250 72.660 61.570 72.720 ;
        RECT 52.510 72.520 61.570 72.660 ;
        RECT 52.510 72.460 52.830 72.520 ;
        RECT 55.055 72.475 55.345 72.520 ;
        RECT 61.250 72.460 61.570 72.520 ;
        RECT 34.585 72.320 34.875 72.365 ;
        RECT 44.690 72.320 45.010 72.380 ;
        RECT 46.030 72.320 46.320 72.365 ;
        RECT 34.585 72.180 46.320 72.320 ;
        RECT 34.585 72.135 34.875 72.180 ;
        RECT 44.690 72.120 45.010 72.180 ;
        RECT 46.030 72.135 46.320 72.180 ;
        RECT 46.990 72.320 47.310 72.380 ;
        RECT 59.410 72.320 59.730 72.380 ;
        RECT 61.800 72.320 61.940 72.860 ;
        RECT 68.610 72.800 68.930 72.860 ;
        RECT 79.190 73.000 79.510 73.060 ;
        RECT 79.665 73.000 79.955 73.045 ;
        RECT 79.190 72.860 79.955 73.000 ;
        RECT 79.190 72.800 79.510 72.860 ;
        RECT 79.665 72.815 79.955 72.860 ;
        RECT 83.330 72.800 83.650 73.060 ;
        RECT 83.790 72.800 84.110 73.060 ;
        RECT 87.010 73.000 87.330 73.060 ;
        RECT 84.340 72.860 87.330 73.000 ;
        RECT 64.025 72.660 64.315 72.705 ;
        RECT 84.340 72.660 84.480 72.860 ;
        RECT 87.010 72.800 87.330 72.860 ;
        RECT 87.470 72.800 87.790 73.060 ;
        RECT 90.230 73.000 90.550 73.060 ;
        RECT 91.165 73.000 91.455 73.045 ;
        RECT 90.230 72.860 91.455 73.000 ;
        RECT 90.230 72.800 90.550 72.860 ;
        RECT 91.165 72.815 91.455 72.860 ;
        RECT 96.225 73.000 96.515 73.045 ;
        RECT 97.130 73.000 97.450 73.060 ;
        RECT 96.225 72.860 97.450 73.000 ;
        RECT 96.225 72.815 96.515 72.860 ;
        RECT 97.130 72.800 97.450 72.860 ;
        RECT 46.990 72.180 59.730 72.320 ;
        RECT 46.990 72.120 47.310 72.180 ;
        RECT 59.410 72.120 59.730 72.180 ;
        RECT 60.880 72.180 61.940 72.320 ;
        RECT 62.720 72.520 64.315 72.660 ;
        RECT 25.845 71.980 26.135 72.025 ;
        RECT 30.890 71.980 31.210 72.040 ;
        RECT 25.845 71.840 31.210 71.980 ;
        RECT 25.845 71.795 26.135 71.840 ;
        RECT 25.920 71.640 26.060 71.795 ;
        RECT 30.890 71.780 31.210 71.840 ;
        RECT 33.190 71.780 33.510 72.040 ;
        RECT 36.425 71.980 36.715 72.025 ;
        RECT 39.690 71.980 39.980 72.025 ;
        RECT 34.200 71.840 36.715 71.980 ;
        RECT 22.240 71.500 26.060 71.640 ;
        RECT 18.010 71.440 18.330 71.500 ;
        RECT 20.770 71.300 21.090 71.360 ;
        RECT 24.910 71.300 25.230 71.360 ;
        RECT 34.200 71.345 34.340 71.840 ;
        RECT 36.425 71.795 36.715 71.840 ;
        RECT 37.445 71.840 39.980 71.980 ;
        RECT 37.445 71.685 37.660 71.840 ;
        RECT 39.690 71.795 39.980 71.840 ;
        RECT 45.625 71.990 45.915 72.025 ;
        RECT 45.625 71.980 46.300 71.990 ;
        RECT 47.450 71.980 47.770 72.040 ;
        RECT 45.625 71.850 47.770 71.980 ;
        RECT 45.625 71.795 45.915 71.850 ;
        RECT 46.160 71.840 47.770 71.850 ;
        RECT 47.450 71.780 47.770 71.840 ;
        RECT 47.910 71.780 48.230 72.040 ;
        RECT 51.190 71.980 51.480 72.025 ;
        RECT 48.945 71.840 51.480 71.980 ;
        RECT 48.945 71.685 49.160 71.840 ;
        RECT 51.190 71.795 51.480 71.840 ;
        RECT 53.890 71.980 54.210 72.040 ;
        RECT 55.745 71.980 56.035 72.025 ;
        RECT 53.890 71.840 56.035 71.980 ;
        RECT 53.890 71.780 54.210 71.840 ;
        RECT 55.745 71.795 56.035 71.840 ;
        RECT 56.665 71.795 56.955 72.025 ;
        RECT 57.125 71.795 57.415 72.025 ;
        RECT 57.585 71.980 57.875 72.025 ;
        RECT 58.490 71.980 58.810 72.040 ;
        RECT 60.880 72.025 61.020 72.180 ;
        RECT 60.805 71.980 61.095 72.025 ;
        RECT 57.585 71.840 61.095 71.980 ;
        RECT 57.585 71.795 57.875 71.840 ;
        RECT 35.510 71.640 35.800 71.685 ;
        RECT 37.370 71.640 37.660 71.685 ;
        RECT 35.510 71.500 37.660 71.640 ;
        RECT 35.510 71.455 35.800 71.500 ;
        RECT 37.370 71.455 37.660 71.500 ;
        RECT 38.290 71.640 38.580 71.685 ;
        RECT 41.550 71.640 41.840 71.685 ;
        RECT 45.165 71.640 45.455 71.685 ;
        RECT 38.290 71.500 45.455 71.640 ;
        RECT 38.290 71.455 38.580 71.500 ;
        RECT 41.550 71.455 41.840 71.500 ;
        RECT 45.165 71.455 45.455 71.500 ;
        RECT 47.010 71.640 47.300 71.685 ;
        RECT 48.870 71.640 49.160 71.685 ;
        RECT 47.010 71.500 49.160 71.640 ;
        RECT 47.010 71.455 47.300 71.500 ;
        RECT 48.870 71.455 49.160 71.500 ;
        RECT 49.750 71.685 50.070 71.700 ;
        RECT 49.750 71.640 50.080 71.685 ;
        RECT 53.050 71.640 53.340 71.685 ;
        RECT 49.750 71.500 53.340 71.640 ;
        RECT 49.750 71.455 50.080 71.500 ;
        RECT 53.050 71.455 53.340 71.500 ;
        RECT 49.750 71.440 50.070 71.455 ;
        RECT 20.770 71.160 25.230 71.300 ;
        RECT 20.770 71.100 21.090 71.160 ;
        RECT 24.910 71.100 25.230 71.160 ;
        RECT 34.125 71.115 34.415 71.345 ;
        RECT 56.740 71.300 56.880 71.795 ;
        RECT 57.200 71.640 57.340 71.795 ;
        RECT 58.490 71.780 58.810 71.840 ;
        RECT 60.805 71.795 61.095 71.840 ;
        RECT 61.265 71.795 61.555 72.025 ;
        RECT 59.870 71.640 60.190 71.700 ;
        RECT 61.340 71.640 61.480 71.795 ;
        RECT 61.710 71.780 62.030 72.040 ;
        RECT 62.170 71.980 62.490 72.040 ;
        RECT 62.720 72.025 62.860 72.520 ;
        RECT 64.025 72.475 64.315 72.520 ;
        RECT 79.740 72.520 84.480 72.660 ;
        RECT 85.170 72.660 85.490 72.720 ;
        RECT 88.850 72.660 89.170 72.720 ;
        RECT 101.750 72.660 102.040 72.705 ;
        RECT 103.610 72.660 103.900 72.705 ;
        RECT 106.390 72.660 106.680 72.705 ;
        RECT 85.170 72.520 92.760 72.660 ;
        RECT 64.100 72.320 64.240 72.475 ;
        RECT 79.740 72.320 79.880 72.520 ;
        RECT 85.170 72.460 85.490 72.520 ;
        RECT 88.850 72.460 89.170 72.520 ;
        RECT 92.620 72.320 92.760 72.520 ;
        RECT 101.750 72.520 106.680 72.660 ;
        RECT 101.750 72.475 102.040 72.520 ;
        RECT 103.610 72.475 103.900 72.520 ;
        RECT 106.390 72.475 106.680 72.520 ;
        RECT 112.330 72.660 112.620 72.705 ;
        RECT 114.190 72.660 114.480 72.705 ;
        RECT 116.970 72.660 117.260 72.705 ;
        RECT 112.330 72.520 117.260 72.660 ;
        RECT 112.330 72.475 112.620 72.520 ;
        RECT 114.190 72.475 114.480 72.520 ;
        RECT 116.970 72.475 117.260 72.520 ;
        RECT 97.130 72.320 97.450 72.380 ;
        RECT 101.285 72.320 101.575 72.365 ;
        RECT 64.100 72.180 79.880 72.320 ;
        RECT 62.645 71.980 62.935 72.025 ;
        RECT 62.170 71.840 62.935 71.980 ;
        RECT 62.170 71.780 62.490 71.840 ;
        RECT 62.645 71.795 62.935 71.840 ;
        RECT 63.090 71.780 63.410 72.040 ;
        RECT 69.070 71.980 69.390 72.040 ;
        RECT 70.465 71.980 70.755 72.025 ;
        RECT 69.070 71.840 70.755 71.980 ;
        RECT 69.070 71.780 69.390 71.840 ;
        RECT 70.465 71.795 70.755 71.840 ;
        RECT 71.830 71.780 72.150 72.040 ;
        RECT 76.520 72.025 76.660 72.180 ;
        RECT 76.445 71.795 76.735 72.025 ;
        RECT 77.365 71.795 77.655 72.025 ;
        RECT 77.440 71.640 77.580 71.795 ;
        RECT 77.810 71.780 78.130 72.040 ;
        RECT 78.270 71.980 78.590 72.040 ;
        RECT 79.740 71.980 79.880 72.180 ;
        RECT 81.580 72.180 91.840 72.320 ;
        RECT 81.580 72.040 81.720 72.180 ;
        RECT 80.125 71.980 80.415 72.025 ;
        RECT 78.270 71.840 79.420 71.980 ;
        RECT 79.740 71.840 80.415 71.980 ;
        RECT 78.270 71.780 78.590 71.840 ;
        RECT 78.730 71.640 79.050 71.700 ;
        RECT 57.200 71.500 63.320 71.640 ;
        RECT 77.440 71.500 79.050 71.640 ;
        RECT 79.280 71.640 79.420 71.840 ;
        RECT 80.125 71.795 80.415 71.840 ;
        RECT 81.030 71.780 81.350 72.040 ;
        RECT 81.490 71.780 81.810 72.040 ;
        RECT 81.965 71.980 82.255 72.025 ;
        RECT 85.170 71.980 85.490 72.040 ;
        RECT 85.720 72.025 85.860 72.180 ;
        RECT 81.965 71.840 85.490 71.980 ;
        RECT 81.965 71.795 82.255 71.840 ;
        RECT 82.040 71.640 82.180 71.795 ;
        RECT 85.170 71.780 85.490 71.840 ;
        RECT 85.645 71.795 85.935 72.025 ;
        RECT 86.105 71.795 86.395 72.025 ;
        RECT 79.280 71.500 82.180 71.640 ;
        RECT 83.790 71.640 84.110 71.700 ;
        RECT 86.180 71.640 86.320 71.795 ;
        RECT 87.010 71.780 87.330 72.040 ;
        RECT 88.850 71.780 89.170 72.040 ;
        RECT 89.400 72.025 89.540 72.180 ;
        RECT 89.325 71.795 89.615 72.025 ;
        RECT 89.785 71.795 90.075 72.025 ;
        RECT 90.705 71.980 90.995 72.025 ;
        RECT 91.150 71.980 91.470 72.040 ;
        RECT 90.320 71.840 91.470 71.980 ;
        RECT 83.790 71.500 86.320 71.640 ;
        RECT 59.870 71.440 60.190 71.500 ;
        RECT 63.180 71.360 63.320 71.500 ;
        RECT 78.730 71.440 79.050 71.500 ;
        RECT 83.790 71.440 84.110 71.500 ;
        RECT 57.110 71.300 57.430 71.360 ;
        RECT 56.740 71.160 57.430 71.300 ;
        RECT 57.110 71.100 57.430 71.160 ;
        RECT 63.090 71.300 63.410 71.360 ;
        RECT 77.810 71.300 78.130 71.360 ;
        RECT 81.490 71.300 81.810 71.360 ;
        RECT 63.090 71.160 81.810 71.300 ;
        RECT 87.100 71.300 87.240 71.780 ;
        RECT 87.470 71.640 87.790 71.700 ;
        RECT 89.860 71.640 90.000 71.795 ;
        RECT 87.470 71.500 90.000 71.640 ;
        RECT 87.470 71.440 87.790 71.500 ;
        RECT 90.320 71.300 90.460 71.840 ;
        RECT 90.705 71.795 90.995 71.840 ;
        RECT 91.150 71.780 91.470 71.840 ;
        RECT 91.700 71.640 91.840 72.180 ;
        RECT 92.620 72.180 96.670 72.320 ;
        RECT 92.620 72.025 92.760 72.180 ;
        RECT 92.545 71.795 92.835 72.025 ;
        RECT 93.005 71.795 93.295 72.025 ;
        RECT 93.465 71.980 93.755 72.025 ;
        RECT 93.910 71.980 94.230 72.040 ;
        RECT 93.465 71.840 94.230 71.980 ;
        RECT 93.465 71.795 93.755 71.840 ;
        RECT 93.080 71.640 93.220 71.795 ;
        RECT 93.910 71.780 94.230 71.840 ;
        RECT 94.370 71.780 94.690 72.040 ;
        RECT 96.530 71.980 96.670 72.180 ;
        RECT 97.130 72.180 110.470 72.320 ;
        RECT 97.130 72.120 97.450 72.180 ;
        RECT 101.285 72.135 101.575 72.180 ;
        RECT 97.605 71.980 97.895 72.025 ;
        RECT 96.530 71.840 97.895 71.980 ;
        RECT 97.605 71.795 97.895 71.840 ;
        RECT 98.065 71.795 98.355 72.025 ;
        RECT 98.525 71.795 98.815 72.025 ;
        RECT 99.445 71.795 99.735 72.025 ;
        RECT 98.140 71.640 98.280 71.795 ;
        RECT 91.700 71.500 98.280 71.640 ;
        RECT 94.370 71.300 94.690 71.360 ;
        RECT 87.100 71.160 94.690 71.300 ;
        RECT 98.600 71.300 98.740 71.795 ;
        RECT 99.520 71.640 99.660 71.795 ;
        RECT 99.890 71.780 100.210 72.040 ;
        RECT 103.125 71.980 103.415 72.025 ;
        RECT 106.390 71.980 106.680 72.025 ;
        RECT 100.900 71.840 103.415 71.980 ;
        RECT 100.350 71.640 100.670 71.700 ;
        RECT 99.520 71.500 100.670 71.640 ;
        RECT 100.350 71.440 100.670 71.500 ;
        RECT 99.430 71.300 99.750 71.360 ;
        RECT 100.900 71.345 101.040 71.840 ;
        RECT 103.125 71.795 103.415 71.840 ;
        RECT 104.145 71.840 106.680 71.980 ;
        RECT 110.330 71.980 110.470 72.180 ;
        RECT 113.690 72.120 114.010 72.380 ;
        RECT 117.370 72.120 117.690 72.380 ;
        RECT 111.865 71.980 112.155 72.025 ;
        RECT 112.310 71.980 112.630 72.040 ;
        RECT 116.970 71.980 117.260 72.025 ;
        RECT 110.330 71.840 112.630 71.980 ;
        RECT 104.145 71.685 104.360 71.840 ;
        RECT 106.390 71.795 106.680 71.840 ;
        RECT 111.865 71.795 112.155 71.840 ;
        RECT 112.310 71.780 112.630 71.840 ;
        RECT 114.725 71.840 117.260 71.980 ;
        RECT 117.460 71.980 117.600 72.120 ;
        RECT 121.050 71.980 121.370 72.040 ;
        RECT 121.985 71.980 122.275 72.025 ;
        RECT 117.460 71.840 122.275 71.980 ;
        RECT 102.210 71.640 102.500 71.685 ;
        RECT 104.070 71.640 104.360 71.685 ;
        RECT 102.210 71.500 104.360 71.640 ;
        RECT 102.210 71.455 102.500 71.500 ;
        RECT 104.070 71.455 104.360 71.500 ;
        RECT 104.990 71.640 105.280 71.685 ;
        RECT 106.790 71.640 107.110 71.700 ;
        RECT 114.725 71.685 114.940 71.840 ;
        RECT 116.970 71.795 117.260 71.840 ;
        RECT 121.050 71.780 121.370 71.840 ;
        RECT 121.985 71.795 122.275 71.840 ;
        RECT 108.250 71.640 108.540 71.685 ;
        RECT 104.990 71.500 108.540 71.640 ;
        RECT 104.990 71.455 105.280 71.500 ;
        RECT 106.790 71.440 107.110 71.500 ;
        RECT 108.250 71.455 108.540 71.500 ;
        RECT 112.790 71.640 113.080 71.685 ;
        RECT 114.650 71.640 114.940 71.685 ;
        RECT 112.790 71.500 114.940 71.640 ;
        RECT 112.790 71.455 113.080 71.500 ;
        RECT 114.650 71.455 114.940 71.500 ;
        RECT 115.570 71.640 115.860 71.685 ;
        RECT 118.830 71.640 119.120 71.685 ;
        RECT 122.445 71.640 122.735 71.685 ;
        RECT 115.570 71.500 122.735 71.640 ;
        RECT 115.570 71.455 115.860 71.500 ;
        RECT 118.830 71.455 119.120 71.500 ;
        RECT 122.445 71.455 122.735 71.500 ;
        RECT 98.600 71.160 99.750 71.300 ;
        RECT 63.090 71.100 63.410 71.160 ;
        RECT 77.810 71.100 78.130 71.160 ;
        RECT 81.490 71.100 81.810 71.160 ;
        RECT 94.370 71.100 94.690 71.160 ;
        RECT 99.430 71.100 99.750 71.160 ;
        RECT 100.825 71.115 101.115 71.345 ;
        RECT 103.570 71.300 103.890 71.360 ;
        RECT 110.255 71.300 110.545 71.345 ;
        RECT 111.390 71.300 111.710 71.360 ;
        RECT 103.570 71.160 111.710 71.300 ;
        RECT 103.570 71.100 103.890 71.160 ;
        RECT 110.255 71.115 110.545 71.160 ;
        RECT 111.390 71.100 111.710 71.160 ;
        RECT 116.910 71.300 117.230 71.360 ;
        RECT 120.835 71.300 121.125 71.345 ;
        RECT 116.910 71.160 121.125 71.300 ;
        RECT 116.910 71.100 117.230 71.160 ;
        RECT 120.835 71.115 121.125 71.160 ;
        RECT 5.520 70.480 125.580 70.960 ;
        RECT 35.950 70.280 36.270 70.340 ;
        RECT 17.640 70.140 36.270 70.280 ;
        RECT 17.640 70.000 17.780 70.140 ;
        RECT 35.950 70.080 36.270 70.140 ;
        RECT 47.910 70.280 48.230 70.340 ;
        RECT 48.845 70.280 49.135 70.325 ;
        RECT 47.910 70.140 49.135 70.280 ;
        RECT 47.910 70.080 48.230 70.140 ;
        RECT 48.845 70.095 49.135 70.140 ;
        RECT 50.225 70.095 50.515 70.325 ;
        RECT 15.265 69.940 15.555 69.985 ;
        RECT 17.550 69.940 17.870 70.000 ;
        RECT 35.490 69.985 35.810 70.000 ;
        RECT 15.265 69.800 17.870 69.940 ;
        RECT 15.265 69.755 15.555 69.800 ;
        RECT 17.550 69.740 17.870 69.800 ;
        RECT 32.750 69.940 33.040 69.985 ;
        RECT 34.610 69.940 34.900 69.985 ;
        RECT 32.750 69.800 34.900 69.940 ;
        RECT 32.750 69.755 33.040 69.800 ;
        RECT 34.610 69.755 34.900 69.800 ;
        RECT 13.870 69.600 14.190 69.660 ;
        RECT 19.850 69.600 20.170 69.660 ;
        RECT 13.870 69.460 20.170 69.600 ;
        RECT 13.870 69.400 14.190 69.460 ;
        RECT 19.850 69.400 20.170 69.460 ;
        RECT 29.970 69.400 30.290 69.660 ;
        RECT 31.825 69.600 32.115 69.645 ;
        RECT 30.520 69.460 32.115 69.600 ;
        RECT 22.610 69.260 22.930 69.320 ;
        RECT 30.520 69.260 30.660 69.460 ;
        RECT 31.825 69.415 32.115 69.460 ;
        RECT 33.665 69.415 33.955 69.645 ;
        RECT 34.685 69.600 34.900 69.755 ;
        RECT 35.490 69.940 35.820 69.985 ;
        RECT 38.790 69.940 39.080 69.985 ;
        RECT 35.490 69.800 39.080 69.940 ;
        RECT 35.490 69.755 35.820 69.800 ;
        RECT 38.790 69.755 39.080 69.800 ;
        RECT 35.490 69.740 35.810 69.755 ;
        RECT 36.930 69.600 37.220 69.645 ;
        RECT 34.685 69.460 37.220 69.600 ;
        RECT 36.930 69.415 37.220 69.460 ;
        RECT 49.765 69.600 50.055 69.645 ;
        RECT 50.300 69.600 50.440 70.095 ;
        RECT 52.050 70.080 52.370 70.340 ;
        RECT 52.510 70.080 52.830 70.340 ;
        RECT 62.645 70.280 62.935 70.325 ;
        RECT 63.090 70.280 63.410 70.340 ;
        RECT 62.645 70.140 63.410 70.280 ;
        RECT 62.645 70.095 62.935 70.140 ;
        RECT 63.090 70.080 63.410 70.140 ;
        RECT 64.010 70.280 64.330 70.340 ;
        RECT 64.485 70.280 64.775 70.325 ;
        RECT 64.010 70.140 64.775 70.280 ;
        RECT 64.010 70.080 64.330 70.140 ;
        RECT 64.485 70.095 64.775 70.140 ;
        RECT 68.610 70.280 68.930 70.340 ;
        RECT 78.270 70.280 78.590 70.340 ;
        RECT 68.610 70.140 78.590 70.280 ;
        RECT 68.610 70.080 68.930 70.140 ;
        RECT 78.270 70.080 78.590 70.140 ;
        RECT 92.070 70.280 92.390 70.340 ;
        RECT 95.765 70.280 96.055 70.325 ;
        RECT 92.070 70.140 96.055 70.280 ;
        RECT 92.070 70.080 92.390 70.140 ;
        RECT 95.765 70.095 96.055 70.140 ;
        RECT 75.525 69.940 75.815 69.985 ;
        RECT 88.850 69.940 89.170 70.000 ;
        RECT 63.640 69.800 66.080 69.940 ;
        RECT 49.765 69.460 50.440 69.600 ;
        RECT 63.090 69.600 63.410 69.660 ;
        RECT 63.640 69.645 63.780 69.800 ;
        RECT 63.565 69.600 63.855 69.645 ;
        RECT 63.090 69.460 63.855 69.600 ;
        RECT 49.765 69.415 50.055 69.460 ;
        RECT 33.740 69.260 33.880 69.415 ;
        RECT 63.090 69.400 63.410 69.460 ;
        RECT 63.565 69.415 63.855 69.460 ;
        RECT 64.010 69.600 64.330 69.660 ;
        RECT 65.940 69.645 66.080 69.800 ;
        RECT 75.525 69.800 89.170 69.940 ;
        RECT 75.525 69.755 75.815 69.800 ;
        RECT 88.850 69.740 89.170 69.800 ;
        RECT 65.405 69.600 65.695 69.645 ;
        RECT 64.010 69.460 65.695 69.600 ;
        RECT 64.010 69.400 64.330 69.460 ;
        RECT 65.405 69.415 65.695 69.460 ;
        RECT 65.865 69.415 66.155 69.645 ;
        RECT 67.705 69.415 67.995 69.645 ;
        RECT 75.985 69.600 76.275 69.645 ;
        RECT 81.490 69.600 81.810 69.660 ;
        RECT 75.985 69.460 81.810 69.600 ;
        RECT 75.985 69.415 76.275 69.460 ;
        RECT 22.610 69.120 30.660 69.260 ;
        RECT 31.900 69.120 33.880 69.260 ;
        RECT 35.030 69.260 35.350 69.320 ;
        RECT 40.795 69.260 41.085 69.305 ;
        RECT 35.030 69.120 41.085 69.260 ;
        RECT 22.610 69.060 22.930 69.120 ;
        RECT 30.905 68.920 31.195 68.965 ;
        RECT 31.900 68.920 32.040 69.120 ;
        RECT 35.030 69.060 35.350 69.120 ;
        RECT 40.795 69.075 41.085 69.120 ;
        RECT 53.445 69.075 53.735 69.305 ;
        RECT 65.480 69.260 65.620 69.415 ;
        RECT 67.780 69.260 67.920 69.415 ;
        RECT 81.490 69.400 81.810 69.460 ;
        RECT 84.250 69.600 84.570 69.660 ;
        RECT 89.785 69.600 90.075 69.645 ;
        RECT 84.250 69.460 90.075 69.600 ;
        RECT 84.250 69.400 84.570 69.460 ;
        RECT 89.785 69.415 90.075 69.460 ;
        RECT 65.480 69.120 67.920 69.260 ;
        RECT 75.510 69.260 75.830 69.320 ;
        RECT 76.445 69.260 76.735 69.305 ;
        RECT 81.030 69.260 81.350 69.320 ;
        RECT 75.510 69.120 81.350 69.260 ;
        RECT 30.905 68.780 32.040 68.920 ;
        RECT 32.290 68.920 32.580 68.965 ;
        RECT 34.150 68.920 34.440 68.965 ;
        RECT 36.930 68.920 37.220 68.965 ;
        RECT 32.290 68.780 37.220 68.920 ;
        RECT 30.905 68.735 31.195 68.780 ;
        RECT 32.290 68.735 32.580 68.780 ;
        RECT 34.150 68.735 34.440 68.780 ;
        RECT 36.930 68.735 37.220 68.780 ;
        RECT 39.170 68.920 39.490 68.980 ;
        RECT 53.520 68.920 53.660 69.075 ;
        RECT 75.510 69.060 75.830 69.120 ;
        RECT 76.445 69.075 76.735 69.120 ;
        RECT 81.030 69.060 81.350 69.120 ;
        RECT 83.790 69.260 84.110 69.320 ;
        RECT 86.105 69.260 86.395 69.305 ;
        RECT 83.790 69.120 86.395 69.260 ;
        RECT 83.790 69.060 84.110 69.120 ;
        RECT 86.105 69.075 86.395 69.120 ;
        RECT 90.690 69.260 91.010 69.320 ;
        RECT 94.845 69.260 95.135 69.305 ;
        RECT 90.690 69.120 95.135 69.260 ;
        RECT 95.840 69.260 95.980 70.095 ;
        RECT 96.210 70.080 96.530 70.340 ;
        RECT 98.065 70.095 98.355 70.325 ;
        RECT 99.890 70.280 100.210 70.340 ;
        RECT 101.285 70.280 101.575 70.325 ;
        RECT 99.890 70.140 101.575 70.280 ;
        RECT 98.140 69.600 98.280 70.095 ;
        RECT 99.890 70.080 100.210 70.140 ;
        RECT 101.285 70.095 101.575 70.140 ;
        RECT 103.125 70.095 103.415 70.325 ;
        RECT 99.445 69.600 99.735 69.645 ;
        RECT 103.200 69.630 103.340 70.095 ;
        RECT 103.570 70.080 103.890 70.340 ;
        RECT 106.790 70.080 107.110 70.340 ;
        RECT 118.750 70.080 119.070 70.340 ;
        RECT 117.370 69.940 117.690 70.000 ;
        RECT 113.780 69.800 117.690 69.940 ;
        RECT 102.740 69.600 103.340 69.630 ;
        RECT 98.140 69.460 99.735 69.600 ;
        RECT 99.445 69.415 99.735 69.460 ;
        RECT 102.280 69.490 103.340 69.600 ;
        RECT 103.570 69.600 103.890 69.660 ;
        RECT 107.265 69.600 107.555 69.645 ;
        RECT 113.780 69.600 113.920 69.800 ;
        RECT 117.370 69.740 117.690 69.800 ;
        RECT 102.280 69.460 102.880 69.490 ;
        RECT 103.570 69.460 113.920 69.600 ;
        RECT 114.150 69.600 114.470 69.660 ;
        RECT 116.925 69.600 117.215 69.645 ;
        RECT 114.150 69.460 117.215 69.600 ;
        RECT 102.280 69.320 102.420 69.460 ;
        RECT 103.570 69.400 103.890 69.460 ;
        RECT 107.265 69.415 107.555 69.460 ;
        RECT 114.150 69.400 114.470 69.460 ;
        RECT 116.925 69.415 117.215 69.460 ;
        RECT 102.190 69.260 102.510 69.320 ;
        RECT 95.840 69.120 102.510 69.260 ;
        RECT 90.690 69.060 91.010 69.120 ;
        RECT 94.845 69.075 95.135 69.120 ;
        RECT 55.270 68.920 55.590 68.980 ;
        RECT 39.170 68.780 55.590 68.920 ;
        RECT 39.170 68.720 39.490 68.780 ;
        RECT 55.270 68.720 55.590 68.780 ;
        RECT 78.730 68.920 79.050 68.980 ;
        RECT 85.630 68.920 85.950 68.980 ;
        RECT 78.730 68.780 85.950 68.920 ;
        RECT 94.920 68.920 95.060 69.075 ;
        RECT 102.190 69.060 102.510 69.120 ;
        RECT 104.505 69.075 104.795 69.305 ;
        RECT 115.545 69.075 115.835 69.305 ;
        RECT 116.465 69.260 116.755 69.305 ;
        RECT 116.080 69.120 116.755 69.260 ;
        RECT 104.580 68.920 104.720 69.075 ;
        RECT 110.470 68.920 110.790 68.980 ;
        RECT 115.070 68.920 115.390 68.980 ;
        RECT 115.620 68.920 115.760 69.075 ;
        RECT 94.920 68.780 115.760 68.920 ;
        RECT 78.730 68.720 79.050 68.780 ;
        RECT 85.630 68.720 85.950 68.780 ;
        RECT 110.470 68.720 110.790 68.780 ;
        RECT 115.070 68.720 115.390 68.780 ;
        RECT 59.410 68.580 59.730 68.640 ;
        RECT 66.785 68.580 67.075 68.625 ;
        RECT 67.690 68.580 68.010 68.640 ;
        RECT 59.410 68.440 68.010 68.580 ;
        RECT 59.410 68.380 59.730 68.440 ;
        RECT 66.785 68.395 67.075 68.440 ;
        RECT 67.690 68.380 68.010 68.440 ;
        RECT 69.070 68.580 69.390 68.640 ;
        RECT 73.685 68.580 73.975 68.625 ;
        RECT 69.070 68.440 73.975 68.580 ;
        RECT 69.070 68.380 69.390 68.440 ;
        RECT 73.685 68.395 73.975 68.440 ;
        RECT 83.330 68.380 83.650 68.640 ;
        RECT 87.010 68.380 87.330 68.640 ;
        RECT 88.850 68.580 89.170 68.640 ;
        RECT 98.050 68.580 98.370 68.640 ;
        RECT 88.850 68.440 98.370 68.580 ;
        RECT 88.850 68.380 89.170 68.440 ;
        RECT 98.050 68.380 98.370 68.440 ;
        RECT 98.510 68.380 98.830 68.640 ;
        RECT 99.430 68.580 99.750 68.640 ;
        RECT 116.080 68.580 116.220 69.120 ;
        RECT 116.465 69.075 116.755 69.120 ;
        RECT 116.450 68.580 116.770 68.640 ;
        RECT 99.430 68.440 116.770 68.580 ;
        RECT 99.430 68.380 99.750 68.440 ;
        RECT 116.450 68.380 116.770 68.440 ;
        RECT 5.520 67.760 125.580 68.240 ;
        RECT 29.970 67.560 30.290 67.620 ;
        RECT 31.365 67.560 31.655 67.605 ;
        RECT 29.970 67.420 31.655 67.560 ;
        RECT 29.970 67.360 30.290 67.420 ;
        RECT 31.365 67.375 31.655 67.420 ;
        RECT 35.490 67.560 35.810 67.620 ;
        RECT 35.965 67.560 36.255 67.605 ;
        RECT 35.490 67.420 36.255 67.560 ;
        RECT 35.490 67.360 35.810 67.420 ;
        RECT 35.965 67.375 36.255 67.420 ;
        RECT 67.705 67.560 67.995 67.605 ;
        RECT 75.510 67.560 75.830 67.620 ;
        RECT 67.705 67.420 75.830 67.560 ;
        RECT 67.705 67.375 67.995 67.420 ;
        RECT 75.510 67.360 75.830 67.420 ;
        RECT 76.890 67.560 77.210 67.620 ;
        RECT 79.665 67.560 79.955 67.605 ;
        RECT 76.890 67.420 79.955 67.560 ;
        RECT 76.890 67.360 77.210 67.420 ;
        RECT 79.665 67.375 79.955 67.420 ;
        RECT 80.570 67.560 80.890 67.620 ;
        RECT 101.730 67.560 102.050 67.620 ;
        RECT 80.570 67.420 102.050 67.560 ;
        RECT 80.570 67.360 80.890 67.420 ;
        RECT 101.730 67.360 102.050 67.420 ;
        RECT 102.190 67.560 102.510 67.620 ;
        RECT 105.195 67.560 105.485 67.605 ;
        RECT 102.190 67.420 105.485 67.560 ;
        RECT 102.190 67.360 102.510 67.420 ;
        RECT 105.195 67.375 105.485 67.420 ;
        RECT 14.345 67.220 14.635 67.265 ;
        RECT 13.960 67.080 14.635 67.220 ;
        RECT 13.960 66.925 14.100 67.080 ;
        RECT 14.345 67.035 14.635 67.080 ;
        RECT 22.240 67.080 34.340 67.220 ;
        RECT 13.885 66.695 14.175 66.925 ;
        RECT 17.105 66.880 17.395 66.925 ;
        RECT 20.310 66.880 20.630 66.940 ;
        RECT 22.240 66.925 22.380 67.080 ;
        RECT 22.165 66.880 22.455 66.925 ;
        RECT 17.105 66.740 22.455 66.880 ;
        RECT 17.105 66.695 17.395 66.740 ;
        RECT 20.310 66.680 20.630 66.740 ;
        RECT 22.165 66.695 22.455 66.740 ;
        RECT 23.990 66.680 24.310 66.940 ;
        RECT 34.200 66.925 34.340 67.080 ;
        RECT 51.145 67.035 51.435 67.265 ;
        RECT 34.125 66.880 34.415 66.925 ;
        RECT 39.170 66.880 39.490 66.940 ;
        RECT 34.125 66.740 39.490 66.880 ;
        RECT 34.125 66.695 34.415 66.740 ;
        RECT 39.170 66.680 39.490 66.740 ;
        RECT 16.170 66.340 16.490 66.600 ;
        RECT 17.550 66.540 17.870 66.600 ;
        RECT 20.785 66.540 21.075 66.585 ;
        RECT 17.550 66.400 21.075 66.540 ;
        RECT 17.550 66.340 17.870 66.400 ;
        RECT 20.785 66.355 21.075 66.400 ;
        RECT 28.130 66.340 28.450 66.600 ;
        RECT 33.665 66.540 33.955 66.585 ;
        RECT 35.030 66.540 35.350 66.600 ;
        RECT 33.665 66.400 35.350 66.540 ;
        RECT 33.665 66.355 33.955 66.400 ;
        RECT 35.030 66.340 35.350 66.400 ;
        RECT 35.505 66.540 35.795 66.585 ;
        RECT 35.950 66.540 36.270 66.600 ;
        RECT 44.705 66.540 44.995 66.585 ;
        RECT 47.450 66.540 47.770 66.600 ;
        RECT 35.505 66.400 47.770 66.540 ;
        RECT 35.505 66.355 35.795 66.400 ;
        RECT 35.950 66.340 36.270 66.400 ;
        RECT 44.705 66.355 44.995 66.400 ;
        RECT 47.450 66.340 47.770 66.400 ;
        RECT 49.765 66.540 50.055 66.585 ;
        RECT 51.220 66.540 51.360 67.035 ;
        RECT 62.170 67.020 62.490 67.280 ;
        RECT 68.610 67.020 68.930 67.280 ;
        RECT 71.335 67.220 71.625 67.265 ;
        RECT 73.225 67.220 73.515 67.265 ;
        RECT 76.345 67.220 76.635 67.265 ;
        RECT 81.950 67.220 82.270 67.280 ;
        RECT 90.690 67.220 91.010 67.280 ;
        RECT 71.335 67.080 76.635 67.220 ;
        RECT 71.335 67.035 71.625 67.080 ;
        RECT 73.225 67.035 73.515 67.080 ;
        RECT 76.345 67.035 76.635 67.080 ;
        RECT 76.980 67.080 82.270 67.220 ;
        RECT 54.365 66.880 54.655 66.925 ;
        RECT 55.270 66.880 55.590 66.940 ;
        RECT 60.790 66.880 61.110 66.940 ;
        RECT 64.930 66.880 65.250 66.940 ;
        RECT 68.700 66.880 68.840 67.020 ;
        RECT 54.365 66.740 61.110 66.880 ;
        RECT 54.365 66.695 54.655 66.740 ;
        RECT 55.270 66.680 55.590 66.740 ;
        RECT 60.790 66.680 61.110 66.740 ;
        RECT 63.180 66.740 68.840 66.880 ;
        RECT 70.465 66.880 70.755 66.925 ;
        RECT 72.290 66.880 72.610 66.940 ;
        RECT 76.980 66.880 77.120 67.080 ;
        RECT 81.950 67.020 82.270 67.080 ;
        RECT 82.500 67.080 91.010 67.220 ;
        RECT 70.465 66.740 77.120 66.880 ;
        RECT 78.730 66.880 79.050 66.940 ;
        RECT 79.205 66.880 79.495 66.925 ;
        RECT 78.730 66.740 79.495 66.880 ;
        RECT 49.765 66.400 51.360 66.540 ;
        RECT 52.510 66.540 52.830 66.600 ;
        RECT 52.985 66.540 53.275 66.585 ;
        RECT 52.510 66.400 53.275 66.540 ;
        RECT 49.765 66.355 50.055 66.400 ;
        RECT 52.510 66.340 52.830 66.400 ;
        RECT 52.985 66.355 53.275 66.400 ;
        RECT 53.445 66.540 53.735 66.585 ;
        RECT 57.110 66.540 57.430 66.600 ;
        RECT 53.445 66.400 57.430 66.540 ;
        RECT 53.445 66.355 53.735 66.400 ;
        RECT 57.110 66.340 57.430 66.400 ;
        RECT 61.250 66.540 61.570 66.600 ;
        RECT 62.630 66.540 62.950 66.600 ;
        RECT 63.180 66.585 63.320 66.740 ;
        RECT 64.930 66.680 65.250 66.740 ;
        RECT 70.465 66.695 70.755 66.740 ;
        RECT 72.290 66.680 72.610 66.740 ;
        RECT 78.730 66.680 79.050 66.740 ;
        RECT 79.205 66.695 79.495 66.740 ;
        RECT 81.030 66.880 81.350 66.940 ;
        RECT 82.500 66.925 82.640 67.080 ;
        RECT 82.425 66.880 82.715 66.925 ;
        RECT 81.030 66.740 82.715 66.880 ;
        RECT 81.030 66.680 81.350 66.740 ;
        RECT 82.425 66.695 82.715 66.740 ;
        RECT 85.630 66.880 85.950 66.940 ;
        RECT 88.020 66.925 88.160 67.080 ;
        RECT 90.690 67.020 91.010 67.080 ;
        RECT 91.165 67.220 91.455 67.265 ;
        RECT 96.690 67.220 96.980 67.265 ;
        RECT 98.550 67.220 98.840 67.265 ;
        RECT 101.330 67.220 101.620 67.265 ;
        RECT 91.165 67.080 91.840 67.220 ;
        RECT 91.165 67.035 91.455 67.080 ;
        RECT 91.700 66.925 91.840 67.080 ;
        RECT 96.690 67.080 101.620 67.220 ;
        RECT 96.690 67.035 96.980 67.080 ;
        RECT 98.550 67.035 98.840 67.080 ;
        RECT 101.330 67.035 101.620 67.080 ;
        RECT 118.305 67.035 118.595 67.265 ;
        RECT 86.565 66.880 86.855 66.925 ;
        RECT 85.630 66.740 86.855 66.880 ;
        RECT 85.630 66.680 85.950 66.740 ;
        RECT 86.565 66.695 86.855 66.740 ;
        RECT 87.945 66.695 88.235 66.925 ;
        RECT 91.625 66.695 91.915 66.925 ;
        RECT 96.225 66.880 96.515 66.925 ;
        RECT 97.130 66.880 97.450 66.940 ;
        RECT 96.225 66.740 97.450 66.880 ;
        RECT 96.225 66.695 96.515 66.740 ;
        RECT 97.130 66.680 97.450 66.740 ;
        RECT 115.070 66.680 115.390 66.940 ;
        RECT 61.250 66.400 62.950 66.540 ;
        RECT 61.250 66.340 61.570 66.400 ;
        RECT 62.630 66.340 62.950 66.400 ;
        RECT 63.105 66.355 63.395 66.585 ;
        RECT 64.485 66.540 64.775 66.585 ;
        RECT 66.770 66.540 67.090 66.600 ;
        RECT 64.485 66.400 67.090 66.540 ;
        RECT 64.485 66.355 64.775 66.400 ;
        RECT 66.770 66.340 67.090 66.400 ;
        RECT 68.625 66.540 68.915 66.585 ;
        RECT 69.070 66.540 69.390 66.600 ;
        RECT 68.625 66.400 69.390 66.540 ;
        RECT 68.625 66.355 68.915 66.400 ;
        RECT 69.070 66.340 69.390 66.400 ;
        RECT 70.930 66.540 71.220 66.585 ;
        RECT 72.765 66.540 73.055 66.585 ;
        RECT 76.345 66.540 76.635 66.585 ;
        RECT 70.930 66.400 76.635 66.540 ;
        RECT 70.930 66.355 71.220 66.400 ;
        RECT 72.765 66.355 73.055 66.400 ;
        RECT 76.345 66.355 76.635 66.400 ;
        RECT 11.110 66.200 11.430 66.260 ;
        RECT 47.925 66.200 48.215 66.245 ;
        RECT 49.290 66.200 49.610 66.260 ;
        RECT 11.110 66.060 19.160 66.200 ;
        RECT 11.110 66.000 11.430 66.060 ;
        RECT 10.650 65.660 10.970 65.920 ;
        RECT 16.645 65.860 16.935 65.905 ;
        RECT 17.090 65.860 17.410 65.920 ;
        RECT 19.020 65.905 19.160 66.060 ;
        RECT 47.925 66.060 49.610 66.200 ;
        RECT 47.925 66.015 48.215 66.060 ;
        RECT 49.290 66.000 49.610 66.060 ;
        RECT 66.310 66.000 66.630 66.260 ;
        RECT 74.130 66.245 74.450 66.260 ;
        RECT 77.425 66.245 77.715 66.560 ;
        RECT 81.490 66.540 81.810 66.600 ;
        RECT 83.805 66.540 84.095 66.585 ;
        RECT 81.490 66.400 84.095 66.540 ;
        RECT 81.490 66.340 81.810 66.400 ;
        RECT 83.805 66.355 84.095 66.400 ;
        RECT 88.865 66.540 89.155 66.585 ;
        RECT 97.590 66.540 97.910 66.600 ;
        RECT 88.865 66.400 97.910 66.540 ;
        RECT 88.865 66.355 89.155 66.400 ;
        RECT 97.590 66.340 97.910 66.400 ;
        RECT 98.065 66.540 98.355 66.585 ;
        RECT 98.510 66.540 98.830 66.600 ;
        RECT 101.330 66.540 101.620 66.585 ;
        RECT 98.065 66.400 98.830 66.540 ;
        RECT 98.065 66.355 98.355 66.400 ;
        RECT 98.510 66.340 98.830 66.400 ;
        RECT 99.085 66.400 101.620 66.540 ;
        RECT 71.845 66.015 72.135 66.245 ;
        RECT 74.125 66.200 74.775 66.245 ;
        RECT 77.425 66.200 78.015 66.245 ;
        RECT 74.125 66.060 78.015 66.200 ;
        RECT 74.125 66.015 74.775 66.060 ;
        RECT 77.725 66.015 78.015 66.060 ;
        RECT 81.965 66.200 82.255 66.245 ;
        RECT 87.010 66.200 87.330 66.260 ;
        RECT 99.085 66.245 99.300 66.400 ;
        RECT 101.330 66.355 101.620 66.400 ;
        RECT 110.010 66.540 110.330 66.600 ;
        RECT 116.005 66.540 116.295 66.585 ;
        RECT 110.010 66.400 116.295 66.540 ;
        RECT 110.010 66.340 110.330 66.400 ;
        RECT 116.005 66.355 116.295 66.400 ;
        RECT 116.450 66.340 116.770 66.600 ;
        RECT 118.380 66.540 118.520 67.035 ;
        RECT 119.685 66.540 119.975 66.585 ;
        RECT 118.380 66.400 119.975 66.540 ;
        RECT 119.685 66.355 119.975 66.400 ;
        RECT 121.050 66.340 121.370 66.600 ;
        RECT 81.965 66.060 87.330 66.200 ;
        RECT 81.965 66.015 82.255 66.060 ;
        RECT 16.645 65.720 17.410 65.860 ;
        RECT 16.645 65.675 16.935 65.720 ;
        RECT 17.090 65.660 17.410 65.720 ;
        RECT 18.945 65.675 19.235 65.905 ;
        RECT 21.245 65.860 21.535 65.905 ;
        RECT 26.750 65.860 27.070 65.920 ;
        RECT 27.225 65.860 27.515 65.905 ;
        RECT 21.245 65.720 27.515 65.860 ;
        RECT 21.245 65.675 21.535 65.720 ;
        RECT 26.750 65.660 27.070 65.720 ;
        RECT 27.225 65.675 27.515 65.720 ;
        RECT 29.510 65.860 29.830 65.920 ;
        RECT 30.905 65.860 31.195 65.905 ;
        RECT 29.510 65.720 31.195 65.860 ;
        RECT 29.510 65.660 29.830 65.720 ;
        RECT 30.905 65.675 31.195 65.720 ;
        RECT 33.190 65.660 33.510 65.920 ;
        RECT 45.150 65.660 45.470 65.920 ;
        RECT 48.370 65.860 48.690 65.920 ;
        RECT 48.845 65.860 49.135 65.905 ;
        RECT 48.370 65.720 49.135 65.860 ;
        RECT 48.370 65.660 48.690 65.720 ;
        RECT 48.845 65.675 49.135 65.720 ;
        RECT 69.545 65.860 69.835 65.905 ;
        RECT 71.920 65.860 72.060 66.015 ;
        RECT 74.130 66.000 74.450 66.015 ;
        RECT 87.010 66.000 87.330 66.060 ;
        RECT 97.150 66.200 97.440 66.245 ;
        RECT 99.010 66.200 99.300 66.245 ;
        RECT 97.150 66.060 99.300 66.200 ;
        RECT 97.150 66.015 97.440 66.060 ;
        RECT 99.010 66.015 99.300 66.060 ;
        RECT 99.930 66.200 100.220 66.245 ;
        RECT 100.810 66.200 101.130 66.260 ;
        RECT 103.190 66.200 103.480 66.245 ;
        RECT 99.930 66.060 103.480 66.200 ;
        RECT 99.930 66.015 100.220 66.060 ;
        RECT 100.810 66.000 101.130 66.060 ;
        RECT 103.190 66.015 103.480 66.060 ;
        RECT 69.545 65.720 72.060 65.860 ;
        RECT 81.030 65.860 81.350 65.920 ;
        RECT 84.250 65.860 84.570 65.920 ;
        RECT 81.030 65.720 84.570 65.860 ;
        RECT 69.545 65.675 69.835 65.720 ;
        RECT 81.030 65.660 81.350 65.720 ;
        RECT 84.250 65.660 84.570 65.720 ;
        RECT 89.310 65.660 89.630 65.920 ;
        RECT 94.370 65.860 94.690 65.920 ;
        RECT 94.845 65.860 95.135 65.905 ;
        RECT 94.370 65.720 95.135 65.860 ;
        RECT 94.370 65.660 94.690 65.720 ;
        RECT 94.845 65.675 95.135 65.720 ;
        RECT 118.750 65.660 119.070 65.920 ;
        RECT 120.130 65.860 120.450 65.920 ;
        RECT 120.605 65.860 120.895 65.905 ;
        RECT 120.130 65.720 120.895 65.860 ;
        RECT 120.130 65.660 120.450 65.720 ;
        RECT 120.605 65.675 120.895 65.720 ;
        RECT 5.520 65.040 125.580 65.520 ;
        RECT 12.045 64.840 12.335 64.885 ;
        RECT 26.305 64.840 26.595 64.885 ;
        RECT 26.750 64.840 27.070 64.900 ;
        RECT 12.045 64.700 14.100 64.840 ;
        RECT 12.045 64.655 12.335 64.700 ;
        RECT 13.960 64.545 14.100 64.700 ;
        RECT 26.305 64.700 27.070 64.840 ;
        RECT 26.305 64.655 26.595 64.700 ;
        RECT 26.750 64.640 27.070 64.700 ;
        RECT 28.130 64.640 28.450 64.900 ;
        RECT 33.190 64.640 33.510 64.900 ;
        RECT 45.150 64.840 45.470 64.900 ;
        RECT 55.055 64.840 55.345 64.885 ;
        RECT 57.110 64.840 57.430 64.900 ;
        RECT 45.150 64.700 49.520 64.840 ;
        RECT 45.150 64.640 45.470 64.700 ;
        RECT 13.885 64.315 14.175 64.545 ;
        RECT 16.165 64.500 16.815 64.545 ;
        RECT 19.765 64.500 20.055 64.545 ;
        RECT 21.230 64.500 21.550 64.560 ;
        RECT 16.165 64.360 21.550 64.500 ;
        RECT 16.165 64.315 16.815 64.360 ;
        RECT 19.465 64.315 20.055 64.360 ;
        RECT 10.650 63.960 10.970 64.220 ;
        RECT 11.110 63.960 11.430 64.220 ;
        RECT 12.970 64.160 13.260 64.205 ;
        RECT 14.805 64.160 15.095 64.205 ;
        RECT 18.385 64.160 18.675 64.205 ;
        RECT 12.970 64.020 18.675 64.160 ;
        RECT 12.970 63.975 13.260 64.020 ;
        RECT 14.805 63.975 15.095 64.020 ;
        RECT 18.385 63.975 18.675 64.020 ;
        RECT 19.465 64.000 19.755 64.315 ;
        RECT 21.230 64.300 21.550 64.360 ;
        RECT 25.845 64.500 26.135 64.545 ;
        RECT 28.590 64.500 28.910 64.560 ;
        RECT 32.730 64.500 33.050 64.560 ;
        RECT 47.010 64.500 47.300 64.545 ;
        RECT 48.870 64.500 49.160 64.545 ;
        RECT 25.845 64.360 36.180 64.500 ;
        RECT 25.845 64.315 26.135 64.360 ;
        RECT 28.590 64.300 28.910 64.360 ;
        RECT 32.730 64.300 33.050 64.360 ;
        RECT 22.610 64.160 22.930 64.220 ;
        RECT 23.990 64.160 24.310 64.220 ;
        RECT 22.610 64.020 24.310 64.160 ;
        RECT 22.610 63.960 22.930 64.020 ;
        RECT 23.990 63.960 24.310 64.020 ;
        RECT 29.510 63.960 29.830 64.220 ;
        RECT 36.040 64.205 36.180 64.360 ;
        RECT 47.010 64.360 49.160 64.500 ;
        RECT 49.380 64.500 49.520 64.700 ;
        RECT 55.055 64.700 57.430 64.840 ;
        RECT 55.055 64.655 55.345 64.700 ;
        RECT 57.110 64.640 57.430 64.700 ;
        RECT 59.410 64.840 59.730 64.900 ;
        RECT 59.885 64.840 60.175 64.885 ;
        RECT 61.710 64.840 62.030 64.900 ;
        RECT 59.410 64.700 62.030 64.840 ;
        RECT 59.410 64.640 59.730 64.700 ;
        RECT 59.885 64.655 60.175 64.700 ;
        RECT 61.710 64.640 62.030 64.700 ;
        RECT 62.170 64.840 62.490 64.900 ;
        RECT 66.310 64.840 66.630 64.900 ;
        RECT 62.170 64.700 66.630 64.840 ;
        RECT 62.170 64.640 62.490 64.700 ;
        RECT 66.310 64.640 66.630 64.700 ;
        RECT 71.385 64.840 71.675 64.885 ;
        RECT 74.130 64.840 74.450 64.900 ;
        RECT 71.385 64.700 74.450 64.840 ;
        RECT 71.385 64.655 71.675 64.700 ;
        RECT 74.130 64.640 74.450 64.700 ;
        RECT 81.030 64.640 81.350 64.900 ;
        RECT 83.345 64.840 83.635 64.885 ;
        RECT 83.790 64.840 84.110 64.900 ;
        RECT 83.345 64.700 84.110 64.840 ;
        RECT 83.345 64.655 83.635 64.700 ;
        RECT 83.790 64.640 84.110 64.700 ;
        RECT 85.185 64.840 85.475 64.885 ;
        RECT 87.010 64.840 87.330 64.900 ;
        RECT 85.185 64.700 87.330 64.840 ;
        RECT 85.185 64.655 85.475 64.700 ;
        RECT 87.010 64.640 87.330 64.700 ;
        RECT 87.470 64.840 87.790 64.900 ;
        RECT 88.850 64.840 89.170 64.900 ;
        RECT 87.470 64.700 89.170 64.840 ;
        RECT 87.470 64.640 87.790 64.700 ;
        RECT 88.850 64.640 89.170 64.700 ;
        RECT 98.050 64.840 98.370 64.900 ;
        RECT 100.365 64.840 100.655 64.885 ;
        RECT 98.050 64.700 100.655 64.840 ;
        RECT 98.050 64.640 98.370 64.700 ;
        RECT 100.365 64.655 100.655 64.700 ;
        RECT 100.810 64.840 101.130 64.900 ;
        RECT 101.285 64.840 101.575 64.885 ;
        RECT 100.810 64.700 101.575 64.840 ;
        RECT 49.790 64.500 50.080 64.545 ;
        RECT 53.050 64.500 53.340 64.545 ;
        RECT 49.380 64.360 53.340 64.500 ;
        RECT 47.010 64.315 47.300 64.360 ;
        RECT 48.870 64.315 49.160 64.360 ;
        RECT 49.790 64.315 50.080 64.360 ;
        RECT 53.050 64.315 53.340 64.360 ;
        RECT 35.965 63.975 36.255 64.205 ;
        RECT 44.690 64.160 45.010 64.220 ;
        RECT 46.085 64.160 46.375 64.205 ;
        RECT 44.690 64.020 46.375 64.160 ;
        RECT 44.690 63.960 45.010 64.020 ;
        RECT 46.085 63.975 46.375 64.020 ;
        RECT 47.925 64.160 48.215 64.205 ;
        RECT 48.370 64.160 48.690 64.220 ;
        RECT 47.925 64.020 48.690 64.160 ;
        RECT 48.945 64.160 49.160 64.315 ;
        RECT 51.190 64.160 51.480 64.205 ;
        RECT 48.945 64.020 51.480 64.160 ;
        RECT 57.200 64.160 57.340 64.640 ;
        RECT 75.965 64.500 76.615 64.545 ;
        RECT 77.350 64.500 77.670 64.560 ;
        RECT 79.565 64.500 79.855 64.545 ;
        RECT 75.965 64.360 79.855 64.500 ;
        RECT 75.965 64.315 76.615 64.360 ;
        RECT 77.350 64.300 77.670 64.360 ;
        RECT 79.265 64.315 79.855 64.360 ;
        RECT 82.870 64.500 83.190 64.560 ;
        RECT 91.605 64.500 92.255 64.545 ;
        RECT 95.205 64.500 95.495 64.545 ;
        RECT 96.670 64.500 96.990 64.560 ;
        RECT 82.870 64.360 88.160 64.500 ;
        RECT 59.425 64.160 59.715 64.205 ;
        RECT 57.200 64.020 59.715 64.160 ;
        RECT 47.925 63.975 48.215 64.020 ;
        RECT 48.370 63.960 48.690 64.020 ;
        RECT 51.190 63.975 51.480 64.020 ;
        RECT 59.425 63.975 59.715 64.020 ;
        RECT 64.010 63.960 64.330 64.220 ;
        RECT 71.830 63.960 72.150 64.220 ;
        RECT 72.290 63.960 72.610 64.220 ;
        RECT 72.770 64.160 73.060 64.205 ;
        RECT 74.605 64.160 74.895 64.205 ;
        RECT 78.185 64.160 78.475 64.205 ;
        RECT 72.770 64.020 78.475 64.160 ;
        RECT 72.770 63.975 73.060 64.020 ;
        RECT 74.605 63.975 74.895 64.020 ;
        RECT 78.185 63.975 78.475 64.020 ;
        RECT 79.265 64.000 79.555 64.315 ;
        RECT 82.870 64.300 83.190 64.360 ;
        RECT 82.425 64.160 82.715 64.205 ;
        RECT 83.330 64.160 83.650 64.220 ;
        RECT 82.425 64.020 83.650 64.160 ;
        RECT 82.425 63.975 82.715 64.020 ;
        RECT 83.330 63.960 83.650 64.020 ;
        RECT 85.645 64.160 85.935 64.205 ;
        RECT 87.470 64.160 87.790 64.220 ;
        RECT 88.020 64.205 88.160 64.360 ;
        RECT 91.605 64.360 96.990 64.500 ;
        RECT 100.440 64.500 100.580 64.655 ;
        RECT 100.810 64.640 101.130 64.700 ;
        RECT 101.285 64.655 101.575 64.700 ;
        RECT 110.010 64.840 110.330 64.900 ;
        RECT 110.945 64.840 111.235 64.885 ;
        RECT 122.215 64.840 122.505 64.885 ;
        RECT 110.010 64.700 122.505 64.840 ;
        RECT 110.010 64.640 110.330 64.700 ;
        RECT 110.945 64.655 111.235 64.700 ;
        RECT 122.215 64.655 122.505 64.700 ;
        RECT 120.130 64.545 120.450 64.560 ;
        RECT 111.405 64.500 111.695 64.545 ;
        RECT 100.440 64.360 111.695 64.500 ;
        RECT 91.605 64.315 92.255 64.360 ;
        RECT 94.905 64.315 95.495 64.360 ;
        RECT 85.645 64.020 87.790 64.160 ;
        RECT 85.645 63.975 85.935 64.020 ;
        RECT 87.470 63.960 87.790 64.020 ;
        RECT 87.945 63.975 88.235 64.205 ;
        RECT 88.410 64.160 88.700 64.205 ;
        RECT 90.245 64.160 90.535 64.205 ;
        RECT 93.825 64.160 94.115 64.205 ;
        RECT 88.410 64.020 94.115 64.160 ;
        RECT 88.410 63.975 88.700 64.020 ;
        RECT 90.245 63.975 90.535 64.020 ;
        RECT 93.825 63.975 94.115 64.020 ;
        RECT 94.905 64.000 95.195 64.315 ;
        RECT 96.670 64.300 96.990 64.360 ;
        RECT 111.405 64.315 111.695 64.360 ;
        RECT 114.170 64.500 114.460 64.545 ;
        RECT 116.030 64.500 116.320 64.545 ;
        RECT 114.170 64.360 116.320 64.500 ;
        RECT 114.170 64.315 114.460 64.360 ;
        RECT 116.030 64.315 116.320 64.360 ;
        RECT 116.950 64.500 117.240 64.545 ;
        RECT 120.130 64.500 120.500 64.545 ;
        RECT 116.950 64.360 120.500 64.500 ;
        RECT 116.950 64.315 117.240 64.360 ;
        RECT 120.130 64.315 120.500 64.360 ;
        RECT 97.605 64.160 97.895 64.205 ;
        RECT 98.970 64.160 99.290 64.220 ;
        RECT 97.605 64.020 99.290 64.160 ;
        RECT 97.605 63.975 97.895 64.020 ;
        RECT 98.970 63.960 99.290 64.020 ;
        RECT 100.825 64.160 101.115 64.205 ;
        RECT 103.110 64.160 103.430 64.220 ;
        RECT 100.825 64.020 103.430 64.160 ;
        RECT 100.825 63.975 101.115 64.020 ;
        RECT 103.110 63.960 103.430 64.020 ;
        RECT 107.265 63.975 107.555 64.205 ;
        RECT 116.105 64.160 116.320 64.315 ;
        RECT 120.130 64.300 120.450 64.315 ;
        RECT 118.350 64.160 118.640 64.205 ;
        RECT 116.105 64.020 118.640 64.160 ;
        RECT 118.350 63.975 118.640 64.020 ;
        RECT 7.430 63.820 7.750 63.880 ;
        RECT 12.505 63.820 12.795 63.865 ;
        RECT 22.700 63.820 22.840 63.960 ;
        RECT 7.430 63.680 22.840 63.820 ;
        RECT 25.385 63.820 25.675 63.865 ;
        RECT 39.170 63.820 39.490 63.880 ;
        RECT 25.385 63.680 39.490 63.820 ;
        RECT 7.430 63.620 7.750 63.680 ;
        RECT 12.505 63.635 12.795 63.680 ;
        RECT 25.385 63.635 25.675 63.680 ;
        RECT 39.170 63.620 39.490 63.680 ;
        RECT 44.230 63.620 44.550 63.880 ;
        RECT 60.790 63.620 61.110 63.880 ;
        RECT 61.710 63.820 62.030 63.880 ;
        RECT 62.185 63.820 62.475 63.865 ;
        RECT 61.710 63.680 62.475 63.820 ;
        RECT 61.710 63.620 62.030 63.680 ;
        RECT 62.185 63.635 62.475 63.680 ;
        RECT 62.645 63.820 62.935 63.865 ;
        RECT 64.470 63.820 64.790 63.880 ;
        RECT 62.645 63.680 64.790 63.820 ;
        RECT 62.645 63.635 62.935 63.680 ;
        RECT 64.470 63.620 64.790 63.680 ;
        RECT 73.670 63.620 73.990 63.880 ;
        RECT 80.570 63.820 80.890 63.880 ;
        RECT 86.105 63.820 86.395 63.865 ;
        RECT 80.570 63.680 86.395 63.820 ;
        RECT 80.570 63.620 80.890 63.680 ;
        RECT 86.105 63.635 86.395 63.680 ;
        RECT 89.325 63.820 89.615 63.865 ;
        RECT 92.990 63.820 93.310 63.880 ;
        RECT 89.325 63.680 93.310 63.820 ;
        RECT 99.060 63.820 99.200 63.960 ;
        RECT 106.330 63.820 106.650 63.880 ;
        RECT 99.060 63.680 106.650 63.820 ;
        RECT 89.325 63.635 89.615 63.680 ;
        RECT 92.990 63.620 93.310 63.680 ;
        RECT 106.330 63.620 106.650 63.680 ;
        RECT 13.375 63.480 13.665 63.525 ;
        RECT 15.265 63.480 15.555 63.525 ;
        RECT 18.385 63.480 18.675 63.525 ;
        RECT 13.375 63.340 18.675 63.480 ;
        RECT 13.375 63.295 13.665 63.340 ;
        RECT 15.265 63.295 15.555 63.340 ;
        RECT 18.385 63.295 18.675 63.340 ;
        RECT 21.245 63.480 21.535 63.525 ;
        RECT 23.530 63.480 23.850 63.540 ;
        RECT 21.245 63.340 23.850 63.480 ;
        RECT 21.245 63.295 21.535 63.340 ;
        RECT 23.530 63.280 23.850 63.340 ;
        RECT 46.550 63.480 46.840 63.525 ;
        RECT 48.410 63.480 48.700 63.525 ;
        RECT 51.190 63.480 51.480 63.525 ;
        RECT 46.550 63.340 51.480 63.480 ;
        RECT 46.550 63.295 46.840 63.340 ;
        RECT 48.410 63.295 48.700 63.340 ;
        RECT 51.190 63.295 51.480 63.340 ;
        RECT 52.050 63.480 52.370 63.540 ;
        RECT 57.585 63.480 57.875 63.525 ;
        RECT 52.050 63.340 57.875 63.480 ;
        RECT 52.050 63.280 52.370 63.340 ;
        RECT 57.585 63.295 57.875 63.340 ;
        RECT 73.175 63.480 73.465 63.525 ;
        RECT 75.065 63.480 75.355 63.525 ;
        RECT 78.185 63.480 78.475 63.525 ;
        RECT 73.175 63.340 78.475 63.480 ;
        RECT 73.175 63.295 73.465 63.340 ;
        RECT 75.065 63.295 75.355 63.340 ;
        RECT 78.185 63.295 78.475 63.340 ;
        RECT 79.190 63.480 79.510 63.540 ;
        RECT 82.870 63.480 83.190 63.540 ;
        RECT 79.190 63.340 83.190 63.480 ;
        RECT 79.190 63.280 79.510 63.340 ;
        RECT 82.870 63.280 83.190 63.340 ;
        RECT 88.815 63.480 89.105 63.525 ;
        RECT 90.705 63.480 90.995 63.525 ;
        RECT 93.825 63.480 94.115 63.525 ;
        RECT 88.815 63.340 94.115 63.480 ;
        RECT 88.815 63.295 89.105 63.340 ;
        RECT 90.705 63.295 90.995 63.340 ;
        RECT 93.825 63.295 94.115 63.340 ;
        RECT 96.685 63.480 96.975 63.525 ;
        RECT 97.590 63.480 97.910 63.540 ;
        RECT 96.685 63.340 97.910 63.480 ;
        RECT 96.685 63.295 96.975 63.340 ;
        RECT 97.590 63.280 97.910 63.340 ;
        RECT 8.810 63.140 9.130 63.200 ;
        RECT 9.745 63.140 10.035 63.185 ;
        RECT 8.810 63.000 10.035 63.140 ;
        RECT 8.810 62.940 9.130 63.000 ;
        RECT 9.745 62.955 10.035 63.000 ;
        RECT 28.590 62.940 28.910 63.200 ;
        RECT 41.485 63.140 41.775 63.185 ;
        RECT 41.930 63.140 42.250 63.200 ;
        RECT 41.485 63.000 42.250 63.140 ;
        RECT 41.485 62.955 41.775 63.000 ;
        RECT 41.930 62.940 42.250 63.000 ;
        RECT 63.090 63.140 63.410 63.200 ;
        RECT 63.565 63.140 63.855 63.185 ;
        RECT 63.090 63.000 63.855 63.140 ;
        RECT 63.090 62.940 63.410 63.000 ;
        RECT 63.565 62.955 63.855 63.000 ;
        RECT 66.770 63.140 67.090 63.200 ;
        RECT 75.970 63.140 76.290 63.200 ;
        RECT 66.770 63.000 76.290 63.140 ;
        RECT 66.770 62.940 67.090 63.000 ;
        RECT 75.970 62.940 76.290 63.000 ;
        RECT 81.490 62.940 81.810 63.200 ;
        RECT 107.340 63.140 107.480 63.975 ;
        RECT 110.470 63.820 110.790 63.880 ;
        RECT 111.865 63.820 112.155 63.865 ;
        RECT 110.470 63.680 112.155 63.820 ;
        RECT 110.470 63.620 110.790 63.680 ;
        RECT 111.865 63.635 112.155 63.680 ;
        RECT 112.310 63.820 112.630 63.880 ;
        RECT 113.245 63.820 113.535 63.865 ;
        RECT 112.310 63.680 113.535 63.820 ;
        RECT 112.310 63.620 112.630 63.680 ;
        RECT 113.245 63.635 113.535 63.680 ;
        RECT 115.085 63.820 115.375 63.865 ;
        RECT 118.750 63.820 119.070 63.880 ;
        RECT 115.085 63.680 119.070 63.820 ;
        RECT 115.085 63.635 115.375 63.680 ;
        RECT 118.750 63.620 119.070 63.680 ;
        RECT 108.185 63.480 108.475 63.525 ;
        RECT 113.710 63.480 114.000 63.525 ;
        RECT 115.570 63.480 115.860 63.525 ;
        RECT 118.350 63.480 118.640 63.525 ;
        RECT 108.185 63.340 110.470 63.480 ;
        RECT 108.185 63.295 108.475 63.340 ;
        RECT 109.105 63.140 109.395 63.185 ;
        RECT 107.340 63.000 109.395 63.140 ;
        RECT 110.330 63.140 110.470 63.340 ;
        RECT 113.710 63.340 118.640 63.480 ;
        RECT 113.710 63.295 114.000 63.340 ;
        RECT 115.570 63.295 115.860 63.340 ;
        RECT 118.350 63.295 118.640 63.340 ;
        RECT 113.230 63.140 113.550 63.200 ;
        RECT 110.330 63.000 113.550 63.140 ;
        RECT 109.105 62.955 109.395 63.000 ;
        RECT 113.230 62.940 113.550 63.000 ;
        RECT 5.520 62.320 125.580 62.800 ;
        RECT 8.810 61.920 9.130 62.180 ;
        RECT 19.850 62.120 20.170 62.180 ;
        RECT 19.850 61.980 30.660 62.120 ;
        RECT 19.850 61.920 20.170 61.980 ;
        RECT 7.430 61.440 7.750 61.500 ;
        RECT 8.365 61.440 8.655 61.485 ;
        RECT 7.430 61.300 8.655 61.440 ;
        RECT 8.900 61.440 9.040 61.920 ;
        RECT 9.235 61.780 9.525 61.825 ;
        RECT 11.125 61.780 11.415 61.825 ;
        RECT 14.245 61.780 14.535 61.825 ;
        RECT 9.235 61.640 14.535 61.780 ;
        RECT 9.235 61.595 9.525 61.640 ;
        RECT 11.125 61.595 11.415 61.640 ;
        RECT 14.245 61.595 14.535 61.640 ;
        RECT 24.875 61.780 25.165 61.825 ;
        RECT 26.765 61.780 27.055 61.825 ;
        RECT 29.885 61.780 30.175 61.825 ;
        RECT 24.875 61.640 30.175 61.780 ;
        RECT 30.520 61.780 30.660 61.980 ;
        RECT 32.730 61.920 33.050 62.180 ;
        RECT 60.790 61.920 61.110 62.180 ;
        RECT 73.670 62.120 73.990 62.180 ;
        RECT 74.145 62.120 74.435 62.165 ;
        RECT 73.670 61.980 74.435 62.120 ;
        RECT 73.670 61.920 73.990 61.980 ;
        RECT 74.145 61.935 74.435 61.980 ;
        RECT 77.350 62.120 77.670 62.180 ;
        RECT 77.825 62.120 78.115 62.165 ;
        RECT 77.350 61.980 78.115 62.120 ;
        RECT 77.350 61.920 77.670 61.980 ;
        RECT 77.825 61.935 78.115 61.980 ;
        RECT 88.865 62.120 89.155 62.165 ;
        RECT 89.310 62.120 89.630 62.180 ;
        RECT 88.865 61.980 89.630 62.120 ;
        RECT 88.865 61.935 89.155 61.980 ;
        RECT 89.310 61.920 89.630 61.980 ;
        RECT 92.990 62.120 93.310 62.180 ;
        RECT 93.925 62.120 94.215 62.165 ;
        RECT 92.990 61.980 94.215 62.120 ;
        RECT 92.990 61.920 93.310 61.980 ;
        RECT 93.925 61.935 94.215 61.980 ;
        RECT 96.670 61.920 96.990 62.180 ;
        RECT 106.330 61.920 106.650 62.180 ;
        RECT 45.170 61.780 45.460 61.825 ;
        RECT 47.030 61.780 47.320 61.825 ;
        RECT 49.810 61.780 50.100 61.825 ;
        RECT 30.520 61.640 41.700 61.780 ;
        RECT 24.875 61.595 25.165 61.640 ;
        RECT 26.765 61.595 27.055 61.640 ;
        RECT 29.885 61.595 30.175 61.640 ;
        RECT 9.745 61.440 10.035 61.485 ;
        RECT 8.900 61.300 10.035 61.440 ;
        RECT 7.430 61.240 7.750 61.300 ;
        RECT 8.365 61.255 8.655 61.300 ;
        RECT 9.745 61.255 10.035 61.300 ;
        RECT 20.310 61.440 20.630 61.500 ;
        RECT 21.705 61.440 21.995 61.485 ;
        RECT 20.310 61.300 21.995 61.440 ;
        RECT 20.310 61.240 20.630 61.300 ;
        RECT 21.705 61.255 21.995 61.300 ;
        RECT 25.385 61.440 25.675 61.485 ;
        RECT 28.590 61.440 28.910 61.500 ;
        RECT 25.385 61.300 28.910 61.440 ;
        RECT 25.385 61.255 25.675 61.300 ;
        RECT 28.590 61.240 28.910 61.300 ;
        RECT 39.170 61.440 39.490 61.500 ;
        RECT 41.025 61.440 41.315 61.485 ;
        RECT 39.170 61.300 41.315 61.440 ;
        RECT 41.560 61.440 41.700 61.640 ;
        RECT 45.170 61.640 50.100 61.780 ;
        RECT 45.170 61.595 45.460 61.640 ;
        RECT 47.030 61.595 47.320 61.640 ;
        RECT 49.810 61.595 50.100 61.640 ;
        RECT 50.670 61.780 50.990 61.840 ;
        RECT 80.075 61.780 80.365 61.825 ;
        RECT 81.965 61.780 82.255 61.825 ;
        RECT 85.085 61.780 85.375 61.825 ;
        RECT 50.670 61.640 67.460 61.780 ;
        RECT 50.670 61.580 50.990 61.640 ;
        RECT 67.320 61.485 67.460 61.640 ;
        RECT 80.075 61.640 85.375 61.780 ;
        RECT 80.075 61.595 80.365 61.640 ;
        RECT 81.965 61.595 82.255 61.640 ;
        RECT 85.085 61.595 85.375 61.640 ;
        RECT 109.205 61.780 109.495 61.825 ;
        RECT 112.325 61.780 112.615 61.825 ;
        RECT 114.215 61.780 114.505 61.825 ;
        RECT 109.205 61.640 114.505 61.780 ;
        RECT 109.205 61.595 109.495 61.640 ;
        RECT 112.325 61.595 112.615 61.640 ;
        RECT 114.215 61.595 114.505 61.640 ;
        RECT 67.245 61.440 67.535 61.485 ;
        RECT 72.750 61.440 73.070 61.500 ;
        RECT 41.560 61.300 65.160 61.440 ;
        RECT 39.170 61.240 39.490 61.300 ;
        RECT 41.025 61.255 41.315 61.300 ;
        RECT 65.020 61.160 65.160 61.300 ;
        RECT 67.245 61.300 73.070 61.440 ;
        RECT 67.245 61.255 67.535 61.300 ;
        RECT 72.750 61.240 73.070 61.300 ;
        RECT 79.190 61.440 79.510 61.500 ;
        RECT 83.330 61.440 83.650 61.500 ;
        RECT 79.190 61.300 83.650 61.440 ;
        RECT 79.190 61.240 79.510 61.300 ;
        RECT 83.330 61.240 83.650 61.300 ;
        RECT 87.945 61.440 88.235 61.485 ;
        RECT 88.850 61.440 89.170 61.500 ;
        RECT 91.625 61.440 91.915 61.485 ;
        RECT 111.850 61.440 112.170 61.500 ;
        RECT 115.085 61.440 115.375 61.485 ;
        RECT 87.945 61.300 91.915 61.440 ;
        RECT 87.945 61.255 88.235 61.300 ;
        RECT 88.850 61.240 89.170 61.300 ;
        RECT 91.625 61.255 91.915 61.300 ;
        RECT 93.540 61.300 97.360 61.440 ;
        RECT 8.830 61.100 9.120 61.145 ;
        RECT 10.665 61.100 10.955 61.145 ;
        RECT 14.245 61.100 14.535 61.145 ;
        RECT 8.830 60.960 14.535 61.100 ;
        RECT 8.830 60.915 9.120 60.960 ;
        RECT 10.665 60.915 10.955 60.960 ;
        RECT 14.245 60.915 14.535 60.960 ;
        RECT 12.490 60.805 12.810 60.820 ;
        RECT 12.025 60.760 12.810 60.805 ;
        RECT 15.325 60.805 15.615 61.120 ;
        RECT 23.990 60.900 24.310 61.160 ;
        RECT 24.470 61.100 24.760 61.145 ;
        RECT 26.305 61.100 26.595 61.145 ;
        RECT 29.885 61.100 30.175 61.145 ;
        RECT 24.470 60.960 30.175 61.100 ;
        RECT 24.470 60.915 24.760 60.960 ;
        RECT 26.305 60.915 26.595 60.960 ;
        RECT 29.885 60.915 30.175 60.960 ;
        RECT 15.325 60.760 15.915 60.805 ;
        RECT 12.025 60.620 15.915 60.760 ;
        RECT 12.025 60.575 12.810 60.620 ;
        RECT 15.625 60.575 15.915 60.620 ;
        RECT 20.770 60.760 21.090 60.820 ;
        RECT 26.750 60.760 27.070 60.820 ;
        RECT 30.965 60.805 31.255 61.120 ;
        RECT 34.125 61.100 34.415 61.145 ;
        RECT 34.570 61.100 34.890 61.160 ;
        RECT 34.125 60.960 34.890 61.100 ;
        RECT 34.125 60.915 34.415 60.960 ;
        RECT 34.570 60.900 34.890 60.960 ;
        RECT 40.565 61.100 40.855 61.145 ;
        RECT 41.930 61.100 42.250 61.160 ;
        RECT 40.565 60.960 42.250 61.100 ;
        RECT 40.565 60.915 40.855 60.960 ;
        RECT 41.930 60.900 42.250 60.960 ;
        RECT 44.690 60.900 45.010 61.160 ;
        RECT 46.545 61.100 46.835 61.145 ;
        RECT 46.990 61.100 47.310 61.160 ;
        RECT 49.810 61.100 50.100 61.145 ;
        RECT 46.545 60.960 47.310 61.100 ;
        RECT 46.545 60.915 46.835 60.960 ;
        RECT 46.990 60.900 47.310 60.960 ;
        RECT 47.565 60.960 50.100 61.100 ;
        RECT 47.565 60.805 47.780 60.960 ;
        RECT 49.810 60.915 50.100 60.960 ;
        RECT 61.265 61.100 61.555 61.145 ;
        RECT 62.170 61.100 62.490 61.160 ;
        RECT 61.265 60.960 62.490 61.100 ;
        RECT 61.265 60.915 61.555 60.960 ;
        RECT 62.170 60.900 62.490 60.960 ;
        RECT 64.930 61.100 65.250 61.160 ;
        RECT 65.865 61.100 66.155 61.145 ;
        RECT 66.310 61.100 66.630 61.160 ;
        RECT 64.930 60.960 66.630 61.100 ;
        RECT 64.930 60.900 65.250 60.960 ;
        RECT 65.865 60.915 66.155 60.960 ;
        RECT 66.310 60.900 66.630 60.960 ;
        RECT 75.065 61.100 75.355 61.145 ;
        RECT 76.890 61.100 77.210 61.160 ;
        RECT 93.540 61.145 93.680 61.300 ;
        RECT 75.065 60.960 77.210 61.100 ;
        RECT 75.065 60.915 75.355 60.960 ;
        RECT 76.890 60.900 77.210 60.960 ;
        RECT 77.365 60.915 77.655 61.145 ;
        RECT 79.670 61.100 79.960 61.145 ;
        RECT 81.505 61.100 81.795 61.145 ;
        RECT 85.085 61.100 85.375 61.145 ;
        RECT 79.670 60.960 85.375 61.100 ;
        RECT 79.670 60.915 79.960 60.960 ;
        RECT 81.505 60.915 81.795 60.960 ;
        RECT 85.085 60.915 85.375 60.960 ;
        RECT 20.770 60.620 27.070 60.760 ;
        RECT 12.490 60.560 12.810 60.575 ;
        RECT 20.770 60.560 21.090 60.620 ;
        RECT 26.750 60.560 27.070 60.620 ;
        RECT 27.665 60.760 28.315 60.805 ;
        RECT 30.965 60.760 31.555 60.805 ;
        RECT 33.665 60.760 33.955 60.805 ;
        RECT 27.665 60.620 33.955 60.760 ;
        RECT 27.665 60.575 28.315 60.620 ;
        RECT 31.265 60.575 31.555 60.620 ;
        RECT 33.665 60.575 33.955 60.620 ;
        RECT 45.630 60.760 45.920 60.805 ;
        RECT 47.490 60.760 47.780 60.805 ;
        RECT 45.630 60.620 47.780 60.760 ;
        RECT 45.630 60.575 45.920 60.620 ;
        RECT 47.490 60.575 47.780 60.620 ;
        RECT 48.410 60.760 48.700 60.805 ;
        RECT 49.290 60.760 49.610 60.820 ;
        RECT 51.670 60.760 51.960 60.805 ;
        RECT 48.410 60.620 51.960 60.760 ;
        RECT 48.410 60.575 48.700 60.620 ;
        RECT 49.290 60.560 49.610 60.620 ;
        RECT 51.670 60.575 51.960 60.620 ;
        RECT 17.105 60.420 17.395 60.465 ;
        RECT 17.550 60.420 17.870 60.480 ;
        RECT 17.105 60.280 17.870 60.420 ;
        RECT 17.105 60.235 17.395 60.280 ;
        RECT 17.550 60.220 17.870 60.280 ;
        RECT 18.930 60.220 19.250 60.480 ;
        RECT 21.245 60.420 21.535 60.465 ;
        RECT 22.610 60.420 22.930 60.480 ;
        RECT 21.245 60.280 22.930 60.420 ;
        RECT 21.245 60.235 21.535 60.280 ;
        RECT 22.610 60.220 22.930 60.280 ;
        RECT 36.870 60.420 37.190 60.480 ;
        RECT 38.265 60.420 38.555 60.465 ;
        RECT 36.870 60.280 38.555 60.420 ;
        RECT 36.870 60.220 37.190 60.280 ;
        RECT 38.265 60.235 38.555 60.280 ;
        RECT 40.105 60.420 40.395 60.465 ;
        RECT 53.675 60.420 53.965 60.465 ;
        RECT 59.410 60.420 59.730 60.480 ;
        RECT 40.105 60.280 59.730 60.420 ;
        RECT 40.105 60.235 40.395 60.280 ;
        RECT 53.675 60.235 53.965 60.280 ;
        RECT 59.410 60.220 59.730 60.280 ;
        RECT 72.290 60.420 72.610 60.480 ;
        RECT 77.440 60.420 77.580 60.915 ;
        RECT 80.585 60.760 80.875 60.805 ;
        RECT 81.030 60.760 81.350 60.820 ;
        RECT 86.165 60.805 86.455 61.120 ;
        RECT 93.465 60.915 93.755 61.145 ;
        RECT 94.370 61.100 94.690 61.160 ;
        RECT 97.220 61.145 97.360 61.300 ;
        RECT 111.850 61.300 115.375 61.440 ;
        RECT 111.850 61.240 112.170 61.300 ;
        RECT 115.085 61.255 115.375 61.300 ;
        RECT 94.845 61.100 95.135 61.145 ;
        RECT 94.370 60.960 95.135 61.100 ;
        RECT 80.585 60.620 81.350 60.760 ;
        RECT 80.585 60.575 80.875 60.620 ;
        RECT 81.030 60.560 81.350 60.620 ;
        RECT 82.865 60.760 83.515 60.805 ;
        RECT 86.165 60.760 86.755 60.805 ;
        RECT 93.005 60.760 93.295 60.805 ;
        RECT 82.865 60.620 93.295 60.760 ;
        RECT 82.865 60.575 83.515 60.620 ;
        RECT 86.465 60.575 86.755 60.620 ;
        RECT 93.005 60.575 93.295 60.620 ;
        RECT 93.540 60.420 93.680 60.915 ;
        RECT 94.370 60.900 94.690 60.960 ;
        RECT 94.845 60.915 95.135 60.960 ;
        RECT 97.145 61.100 97.435 61.145 ;
        RECT 97.590 61.100 97.910 61.160 ;
        RECT 104.490 61.100 104.810 61.160 ;
        RECT 97.145 60.960 104.810 61.100 ;
        RECT 97.145 60.915 97.435 60.960 ;
        RECT 97.590 60.900 97.910 60.960 ;
        RECT 104.490 60.900 104.810 60.960 ;
        RECT 108.125 60.805 108.415 61.120 ;
        RECT 109.205 61.100 109.495 61.145 ;
        RECT 112.785 61.100 113.075 61.145 ;
        RECT 114.620 61.100 114.910 61.145 ;
        RECT 109.205 60.960 114.910 61.100 ;
        RECT 109.205 60.915 109.495 60.960 ;
        RECT 112.785 60.915 113.075 60.960 ;
        RECT 114.620 60.915 114.910 60.960 ;
        RECT 107.825 60.760 108.415 60.805 ;
        RECT 110.930 60.805 111.250 60.820 ;
        RECT 110.930 60.760 111.715 60.805 ;
        RECT 107.825 60.620 111.715 60.760 ;
        RECT 107.825 60.575 108.115 60.620 ;
        RECT 110.930 60.575 111.715 60.620 ;
        RECT 113.230 60.760 113.550 60.820 ;
        RECT 113.705 60.760 113.995 60.805 ;
        RECT 113.230 60.620 113.995 60.760 ;
        RECT 110.930 60.560 111.250 60.575 ;
        RECT 113.230 60.560 113.550 60.620 ;
        RECT 113.705 60.575 113.995 60.620 ;
        RECT 72.290 60.280 93.680 60.420 ;
        RECT 72.290 60.220 72.610 60.280 ;
        RECT 5.520 59.600 125.580 60.080 ;
        RECT 12.490 59.200 12.810 59.460 ;
        RECT 17.090 59.200 17.410 59.460 ;
        RECT 21.230 59.200 21.550 59.460 ;
        RECT 23.545 59.400 23.835 59.445 ;
        RECT 23.990 59.400 24.310 59.460 ;
        RECT 23.545 59.260 24.310 59.400 ;
        RECT 23.545 59.215 23.835 59.260 ;
        RECT 23.990 59.200 24.310 59.260 ;
        RECT 26.750 59.400 27.070 59.460 ;
        RECT 41.945 59.400 42.235 59.445 ;
        RECT 44.230 59.400 44.550 59.460 ;
        RECT 26.750 59.260 44.550 59.400 ;
        RECT 26.750 59.200 27.070 59.260 ;
        RECT 41.945 59.215 42.235 59.260 ;
        RECT 44.230 59.200 44.550 59.260 ;
        RECT 46.990 59.200 47.310 59.460 ;
        RECT 105.870 59.400 106.190 59.460 ;
        RECT 107.265 59.400 107.555 59.445 ;
        RECT 105.870 59.260 107.555 59.400 ;
        RECT 105.870 59.200 106.190 59.260 ;
        RECT 107.265 59.215 107.555 59.260 ;
        RECT 110.930 59.200 111.250 59.460 ;
        RECT 13.425 59.060 13.715 59.105 ;
        RECT 34.570 59.060 34.890 59.120 ;
        RECT 11.660 58.920 13.715 59.060 ;
        RECT 11.660 58.765 11.800 58.920 ;
        RECT 13.425 58.875 13.715 58.920 ;
        RECT 15.340 58.920 34.890 59.060 ;
        RECT 15.340 58.780 15.480 58.920 ;
        RECT 11.585 58.535 11.875 58.765 ;
        RECT 12.965 58.720 13.255 58.765 ;
        RECT 15.250 58.720 15.570 58.780 ;
        RECT 12.965 58.580 15.570 58.720 ;
        RECT 12.965 58.535 13.255 58.580 ;
        RECT 15.250 58.520 15.570 58.580 ;
        RECT 16.645 58.720 16.935 58.765 ;
        RECT 18.930 58.720 19.250 58.780 ;
        RECT 21.780 58.765 21.920 58.920 ;
        RECT 34.570 58.860 34.890 58.920 ;
        RECT 36.865 59.060 37.515 59.105 ;
        RECT 38.250 59.060 38.570 59.120 ;
        RECT 40.465 59.060 40.755 59.105 ;
        RECT 36.865 58.920 40.755 59.060 ;
        RECT 36.865 58.875 37.515 58.920 ;
        RECT 38.250 58.860 38.570 58.920 ;
        RECT 40.165 58.875 40.755 58.920 ;
        RECT 16.645 58.580 19.250 58.720 ;
        RECT 16.645 58.535 16.935 58.580 ;
        RECT 18.930 58.520 19.250 58.580 ;
        RECT 21.705 58.535 21.995 58.765 ;
        RECT 30.890 58.520 31.210 58.780 ;
        RECT 33.670 58.720 33.960 58.765 ;
        RECT 35.505 58.720 35.795 58.765 ;
        RECT 39.085 58.720 39.375 58.765 ;
        RECT 33.670 58.580 39.375 58.720 ;
        RECT 33.670 58.535 33.960 58.580 ;
        RECT 35.505 58.535 35.795 58.580 ;
        RECT 39.085 58.535 39.375 58.580 ;
        RECT 40.165 58.560 40.455 58.875 ;
        RECT 72.290 58.860 72.610 59.120 ;
        RECT 92.070 58.860 92.390 59.120 ;
        RECT 101.285 59.060 101.575 59.105 ;
        RECT 107.710 59.060 108.030 59.120 ;
        RECT 101.285 58.920 108.030 59.060 ;
        RECT 101.285 58.875 101.575 58.920 ;
        RECT 107.710 58.860 108.030 58.920 ;
        RECT 47.925 58.720 48.215 58.765 ;
        RECT 52.050 58.720 52.370 58.780 ;
        RECT 47.925 58.580 52.370 58.720 ;
        RECT 47.925 58.535 48.215 58.580 ;
        RECT 52.050 58.520 52.370 58.580 ;
        RECT 62.170 58.720 62.490 58.780 ;
        RECT 63.105 58.720 63.395 58.765 ;
        RECT 62.170 58.580 63.395 58.720 ;
        RECT 62.170 58.520 62.490 58.580 ;
        RECT 63.105 58.535 63.395 58.580 ;
        RECT 66.310 58.720 66.630 58.780 ;
        RECT 70.925 58.720 71.215 58.765 ;
        RECT 66.310 58.580 71.215 58.720 ;
        RECT 66.310 58.520 66.630 58.580 ;
        RECT 70.925 58.535 71.215 58.580 ;
        RECT 81.965 58.535 82.255 58.765 ;
        RECT 17.550 58.380 17.870 58.440 ;
        RECT 19.865 58.380 20.155 58.425 ;
        RECT 17.550 58.240 20.155 58.380 ;
        RECT 17.550 58.180 17.870 58.240 ;
        RECT 19.865 58.195 20.155 58.240 ;
        RECT 33.205 58.380 33.495 58.425 ;
        RECT 33.205 58.240 33.880 58.380 ;
        RECT 33.205 58.195 33.495 58.240 ;
        RECT 10.665 57.700 10.955 57.745 ;
        RECT 11.570 57.700 11.890 57.760 ;
        RECT 10.665 57.560 11.890 57.700 ;
        RECT 33.740 57.700 33.880 58.240 ;
        RECT 34.570 58.180 34.890 58.440 ;
        RECT 82.040 58.380 82.180 58.535 ;
        RECT 83.330 58.380 83.650 58.440 ;
        RECT 82.040 58.240 83.650 58.380 ;
        RECT 92.160 58.380 92.300 58.860 ;
        RECT 98.510 58.720 98.830 58.780 ;
        RECT 101.730 58.720 102.050 58.780 ;
        RECT 104.045 58.720 104.335 58.765 ;
        RECT 98.510 58.580 104.335 58.720 ;
        RECT 98.510 58.520 98.830 58.580 ;
        RECT 101.730 58.520 102.050 58.580 ;
        RECT 104.045 58.535 104.335 58.580 ;
        RECT 102.190 58.380 102.510 58.440 ;
        RECT 92.160 58.240 102.510 58.380 ;
        RECT 83.330 58.180 83.650 58.240 ;
        RECT 102.190 58.180 102.510 58.240 ;
        RECT 34.075 58.040 34.365 58.085 ;
        RECT 35.965 58.040 36.255 58.085 ;
        RECT 39.085 58.040 39.375 58.085 ;
        RECT 34.075 57.900 39.375 58.040 ;
        RECT 34.075 57.855 34.365 57.900 ;
        RECT 35.965 57.855 36.255 57.900 ;
        RECT 39.085 57.855 39.375 57.900 ;
        RECT 41.930 57.700 42.250 57.760 ;
        RECT 44.690 57.700 45.010 57.760 ;
        RECT 33.740 57.560 45.010 57.700 ;
        RECT 10.665 57.515 10.955 57.560 ;
        RECT 11.570 57.500 11.890 57.560 ;
        RECT 41.930 57.500 42.250 57.560 ;
        RECT 44.690 57.500 45.010 57.560 ;
        RECT 64.485 57.700 64.775 57.745 ;
        RECT 76.430 57.700 76.750 57.760 ;
        RECT 91.150 57.700 91.470 57.760 ;
        RECT 64.485 57.560 91.470 57.700 ;
        RECT 104.120 57.700 104.260 58.535 ;
        RECT 104.950 58.520 105.270 58.780 ;
        RECT 105.410 58.520 105.730 58.780 ;
        RECT 105.870 58.720 106.190 58.780 ;
        RECT 105.870 58.580 110.470 58.720 ;
        RECT 105.870 58.520 106.190 58.580 ;
        RECT 110.330 58.380 110.470 58.580 ;
        RECT 111.390 58.520 111.710 58.780 ;
        RECT 114.150 58.380 114.470 58.440 ;
        RECT 110.330 58.240 114.470 58.380 ;
        RECT 114.150 58.180 114.470 58.240 ;
        RECT 104.490 58.040 104.810 58.100 ;
        RECT 111.390 58.040 111.710 58.100 ;
        RECT 104.490 57.900 111.710 58.040 ;
        RECT 104.490 57.840 104.810 57.900 ;
        RECT 111.390 57.840 111.710 57.900 ;
        RECT 113.690 57.700 114.010 57.760 ;
        RECT 104.120 57.560 114.010 57.700 ;
        RECT 64.485 57.515 64.775 57.560 ;
        RECT 76.430 57.500 76.750 57.560 ;
        RECT 91.150 57.500 91.470 57.560 ;
        RECT 113.690 57.500 114.010 57.560 ;
        RECT 5.520 56.880 125.580 57.360 ;
        RECT 16.170 56.680 16.490 56.740 ;
        RECT 17.105 56.680 17.395 56.725 ;
        RECT 16.170 56.540 17.395 56.680 ;
        RECT 16.170 56.480 16.490 56.540 ;
        RECT 17.105 56.495 17.395 56.540 ;
        RECT 9.235 56.340 9.525 56.385 ;
        RECT 11.125 56.340 11.415 56.385 ;
        RECT 14.245 56.340 14.535 56.385 ;
        RECT 9.235 56.200 14.535 56.340 ;
        RECT 9.235 56.155 9.525 56.200 ;
        RECT 11.125 56.155 11.415 56.200 ;
        RECT 14.245 56.155 14.535 56.200 ;
        RECT 7.430 56.000 7.750 56.060 ;
        RECT 8.365 56.000 8.655 56.045 ;
        RECT 7.430 55.860 8.655 56.000 ;
        RECT 7.430 55.800 7.750 55.860 ;
        RECT 8.365 55.815 8.655 55.860 ;
        RECT 9.745 56.000 10.035 56.045 ;
        RECT 11.570 56.000 11.890 56.060 ;
        RECT 9.745 55.860 11.890 56.000 ;
        RECT 17.180 56.000 17.320 56.495 ;
        RECT 22.610 56.480 22.930 56.740 ;
        RECT 34.570 56.680 34.890 56.740 ;
        RECT 35.965 56.680 36.255 56.725 ;
        RECT 34.570 56.540 36.255 56.680 ;
        RECT 34.570 56.480 34.890 56.540 ;
        RECT 35.965 56.495 36.255 56.540 ;
        RECT 38.250 56.680 38.570 56.740 ;
        RECT 38.725 56.680 39.015 56.725 ;
        RECT 38.250 56.540 39.015 56.680 ;
        RECT 38.250 56.480 38.570 56.540 ;
        RECT 38.725 56.495 39.015 56.540 ;
        RECT 48.370 56.680 48.690 56.740 ;
        RECT 65.865 56.680 66.155 56.725 ;
        RECT 93.005 56.680 93.295 56.725 ;
        RECT 93.450 56.680 93.770 56.740 ;
        RECT 48.370 56.540 92.300 56.680 ;
        RECT 48.370 56.480 48.690 56.540 ;
        RECT 65.865 56.495 66.155 56.540 ;
        RECT 22.150 56.340 22.470 56.400 ;
        RECT 26.305 56.340 26.595 56.385 ;
        RECT 22.150 56.200 26.595 56.340 ;
        RECT 22.150 56.140 22.470 56.200 ;
        RECT 26.305 56.155 26.595 56.200 ;
        RECT 63.550 56.340 63.870 56.400 ;
        RECT 64.025 56.340 64.315 56.385 ;
        RECT 63.550 56.200 64.315 56.340 ;
        RECT 63.550 56.140 63.870 56.200 ;
        RECT 64.025 56.155 64.315 56.200 ;
        RECT 64.470 56.140 64.790 56.400 ;
        RECT 91.610 56.140 91.930 56.400 ;
        RECT 19.405 56.000 19.695 56.045 ;
        RECT 17.180 55.860 19.695 56.000 ;
        RECT 9.745 55.815 10.035 55.860 ;
        RECT 11.570 55.800 11.890 55.860 ;
        RECT 19.405 55.815 19.695 55.860 ;
        RECT 35.030 56.000 35.350 56.060 ;
        RECT 47.910 56.000 48.230 56.060 ;
        RECT 50.225 56.000 50.515 56.045 ;
        RECT 35.030 55.860 38.480 56.000 ;
        RECT 35.030 55.800 35.350 55.860 ;
        RECT 38.340 55.720 38.480 55.860 ;
        RECT 47.910 55.860 50.515 56.000 ;
        RECT 47.910 55.800 48.230 55.860 ;
        RECT 50.225 55.815 50.515 55.860 ;
        RECT 59.870 56.000 60.190 56.060 ;
        RECT 62.170 56.000 62.490 56.060 ;
        RECT 62.645 56.000 62.935 56.045 ;
        RECT 59.870 55.860 62.935 56.000 ;
        RECT 59.870 55.800 60.190 55.860 ;
        RECT 62.170 55.800 62.490 55.860 ;
        RECT 62.645 55.815 62.935 55.860 ;
        RECT 63.105 56.000 63.395 56.045 ;
        RECT 64.560 56.000 64.700 56.140 ;
        RECT 91.700 56.000 91.840 56.140 ;
        RECT 63.105 55.860 64.700 56.000 ;
        RECT 90.320 55.860 91.840 56.000 ;
        RECT 92.160 56.000 92.300 56.540 ;
        RECT 93.005 56.540 93.770 56.680 ;
        RECT 93.005 56.495 93.295 56.540 ;
        RECT 93.450 56.480 93.770 56.540 ;
        RECT 101.745 56.680 102.035 56.725 ;
        RECT 102.650 56.680 102.970 56.740 ;
        RECT 101.745 56.540 102.970 56.680 ;
        RECT 101.745 56.495 102.035 56.540 ;
        RECT 102.650 56.480 102.970 56.540 ;
        RECT 105.870 56.000 106.190 56.060 ;
        RECT 92.160 55.860 106.190 56.000 ;
        RECT 63.105 55.815 63.395 55.860 ;
        RECT 8.830 55.660 9.120 55.705 ;
        RECT 10.665 55.660 10.955 55.705 ;
        RECT 14.245 55.660 14.535 55.705 ;
        RECT 8.830 55.520 14.535 55.660 ;
        RECT 8.830 55.475 9.120 55.520 ;
        RECT 10.665 55.475 10.955 55.520 ;
        RECT 14.245 55.475 14.535 55.520 ;
        RECT 12.025 55.320 12.675 55.365 ;
        RECT 14.790 55.320 15.110 55.380 ;
        RECT 15.325 55.365 15.615 55.680 ;
        RECT 23.070 55.460 23.390 55.720 ;
        RECT 23.990 55.460 24.310 55.720 ;
        RECT 24.465 55.475 24.755 55.705 ;
        RECT 24.925 55.660 25.215 55.705 ;
        RECT 28.590 55.660 28.910 55.720 ;
        RECT 24.925 55.520 28.910 55.660 ;
        RECT 24.925 55.475 25.215 55.520 ;
        RECT 15.325 55.320 15.915 55.365 ;
        RECT 12.025 55.180 15.915 55.320 ;
        RECT 12.025 55.135 12.675 55.180 ;
        RECT 14.790 55.120 15.110 55.180 ;
        RECT 15.625 55.135 15.915 55.180 ;
        RECT 23.530 55.320 23.850 55.380 ;
        RECT 24.540 55.320 24.680 55.475 ;
        RECT 28.590 55.460 28.910 55.520 ;
        RECT 36.870 55.460 37.190 55.720 ;
        RECT 38.250 55.460 38.570 55.720 ;
        RECT 41.025 55.660 41.315 55.705 ;
        RECT 41.930 55.660 42.250 55.720 ;
        RECT 41.025 55.520 42.250 55.660 ;
        RECT 41.025 55.475 41.315 55.520 ;
        RECT 41.930 55.460 42.250 55.520 ;
        RECT 42.850 55.660 43.170 55.720 ;
        RECT 48.370 55.660 48.690 55.720 ;
        RECT 42.850 55.520 48.690 55.660 ;
        RECT 42.850 55.460 43.170 55.520 ;
        RECT 48.370 55.460 48.690 55.520 ;
        RECT 49.305 55.660 49.595 55.705 ;
        RECT 50.670 55.660 50.990 55.720 ;
        RECT 49.305 55.520 50.990 55.660 ;
        RECT 49.305 55.475 49.595 55.520 ;
        RECT 50.670 55.460 50.990 55.520 ;
        RECT 51.590 55.460 51.910 55.720 ;
        RECT 64.470 55.660 64.790 55.720 ;
        RECT 66.785 55.660 67.075 55.705 ;
        RECT 67.245 55.660 67.535 55.705 ;
        RECT 64.470 55.520 67.535 55.660 ;
        RECT 64.470 55.460 64.790 55.520 ;
        RECT 66.785 55.475 67.075 55.520 ;
        RECT 67.245 55.475 67.535 55.520 ;
        RECT 89.785 55.660 90.075 55.705 ;
        RECT 90.320 55.660 90.460 55.860 ;
        RECT 89.785 55.520 90.460 55.660 ;
        RECT 89.785 55.475 90.075 55.520 ;
        RECT 90.690 55.460 91.010 55.720 ;
        RECT 91.165 55.475 91.455 55.705 ;
        RECT 91.625 55.660 91.915 55.705 ;
        RECT 92.160 55.660 92.300 55.860 ;
        RECT 91.625 55.520 92.300 55.660 ;
        RECT 91.625 55.475 91.915 55.520 ;
        RECT 23.530 55.180 24.680 55.320 ;
        RECT 46.990 55.320 47.310 55.380 ;
        RECT 47.925 55.320 48.215 55.365 ;
        RECT 62.185 55.320 62.475 55.365 ;
        RECT 74.590 55.320 74.910 55.380 ;
        RECT 46.990 55.180 48.215 55.320 ;
        RECT 23.530 55.120 23.850 55.180 ;
        RECT 46.990 55.120 47.310 55.180 ;
        RECT 47.925 55.135 48.215 55.180 ;
        RECT 52.600 55.180 74.910 55.320 ;
        RECT 51.590 54.980 51.910 55.040 ;
        RECT 52.600 54.980 52.740 55.180 ;
        RECT 62.185 55.135 62.475 55.180 ;
        RECT 74.590 55.120 74.910 55.180 ;
        RECT 90.230 55.320 90.550 55.380 ;
        RECT 91.240 55.320 91.380 55.475 ;
        RECT 98.510 55.460 98.830 55.720 ;
        RECT 98.970 55.660 99.290 55.720 ;
        RECT 100.440 55.705 100.580 55.860 ;
        RECT 105.870 55.800 106.190 55.860 ;
        RECT 107.710 56.000 108.030 56.060 ;
        RECT 110.945 56.000 111.235 56.045 ;
        RECT 111.850 56.000 112.170 56.060 ;
        RECT 107.710 55.860 112.170 56.000 ;
        RECT 107.710 55.800 108.030 55.860 ;
        RECT 110.945 55.815 111.235 55.860 ;
        RECT 111.850 55.800 112.170 55.860 ;
        RECT 99.445 55.660 99.735 55.705 ;
        RECT 98.970 55.520 99.735 55.660 ;
        RECT 98.970 55.460 99.290 55.520 ;
        RECT 99.445 55.475 99.735 55.520 ;
        RECT 99.905 55.475 100.195 55.705 ;
        RECT 100.365 55.475 100.655 55.705 ;
        RECT 111.390 55.660 111.710 55.720 ;
        RECT 112.325 55.660 112.615 55.705 ;
        RECT 111.390 55.520 112.615 55.660 ;
        RECT 90.230 55.180 91.380 55.320 ;
        RECT 90.230 55.120 90.550 55.180 ;
        RECT 51.590 54.840 52.740 54.980 ;
        RECT 57.570 54.980 57.890 55.040 ;
        RECT 68.165 54.980 68.455 55.025 ;
        RECT 70.450 54.980 70.770 55.040 ;
        RECT 57.570 54.840 70.770 54.980 ;
        RECT 91.240 54.980 91.380 55.180 ;
        RECT 99.980 54.980 100.120 55.475 ;
        RECT 111.390 55.460 111.710 55.520 ;
        RECT 112.325 55.475 112.615 55.520 ;
        RECT 102.190 55.120 102.510 55.380 ;
        RECT 111.850 55.120 112.170 55.380 ;
        RECT 105.410 54.980 105.730 55.040 ;
        RECT 91.240 54.840 105.730 54.980 ;
        RECT 51.590 54.780 51.910 54.840 ;
        RECT 57.570 54.780 57.890 54.840 ;
        RECT 68.165 54.795 68.455 54.840 ;
        RECT 70.450 54.780 70.770 54.840 ;
        RECT 105.410 54.780 105.730 54.840 ;
        RECT 5.520 54.160 125.580 54.640 ;
        RECT 14.790 53.760 15.110 54.020 ;
        RECT 22.610 53.760 22.930 54.020 ;
        RECT 26.305 53.960 26.595 54.005 ;
        RECT 27.210 53.960 27.530 54.020 ;
        RECT 26.305 53.820 27.530 53.960 ;
        RECT 26.305 53.775 26.595 53.820 ;
        RECT 27.210 53.760 27.530 53.820 ;
        RECT 29.050 53.960 29.370 54.020 ;
        RECT 29.985 53.960 30.275 54.005 ;
        RECT 35.030 53.960 35.350 54.020 ;
        RECT 29.050 53.820 30.275 53.960 ;
        RECT 29.050 53.760 29.370 53.820 ;
        RECT 29.985 53.775 30.275 53.820 ;
        RECT 31.900 53.820 35.350 53.960 ;
        RECT 11.585 53.620 11.875 53.665 ;
        RECT 13.870 53.620 14.190 53.680 ;
        RECT 23.530 53.620 23.850 53.680 ;
        RECT 31.350 53.620 31.670 53.680 ;
        RECT 11.585 53.480 14.190 53.620 ;
        RECT 11.585 53.435 11.875 53.480 ;
        RECT 13.870 53.420 14.190 53.480 ;
        RECT 20.860 53.480 31.670 53.620 ;
        RECT 5.590 53.280 5.910 53.340 ;
        RECT 10.665 53.280 10.955 53.325 ;
        RECT 5.590 53.140 10.955 53.280 ;
        RECT 5.590 53.080 5.910 53.140 ;
        RECT 10.665 53.095 10.955 53.140 ;
        RECT 15.250 53.080 15.570 53.340 ;
        RECT 19.405 53.280 19.695 53.325 ;
        RECT 19.405 53.140 20.080 53.280 ;
        RECT 19.405 53.095 19.695 53.140 ;
        RECT 19.940 52.260 20.080 53.140 ;
        RECT 20.310 53.080 20.630 53.340 ;
        RECT 20.860 53.325 21.000 53.480 ;
        RECT 23.530 53.420 23.850 53.480 ;
        RECT 20.785 53.095 21.075 53.325 ;
        RECT 21.245 53.280 21.535 53.325 ;
        RECT 21.245 53.140 22.840 53.280 ;
        RECT 21.245 53.095 21.535 53.140 ;
        RECT 22.700 52.600 22.840 53.140 ;
        RECT 23.070 53.080 23.390 53.340 ;
        RECT 24.540 53.325 24.680 53.480 ;
        RECT 27.300 53.340 27.440 53.480 ;
        RECT 24.005 53.095 24.295 53.325 ;
        RECT 24.465 53.095 24.755 53.325 ;
        RECT 24.925 53.095 25.215 53.325 ;
        RECT 26.765 53.095 27.055 53.325 ;
        RECT 23.530 52.940 23.850 53.000 ;
        RECT 24.080 52.940 24.220 53.095 ;
        RECT 23.530 52.800 24.220 52.940 ;
        RECT 23.530 52.740 23.850 52.800 ;
        RECT 25.000 52.600 25.140 53.095 ;
        RECT 25.830 52.940 26.150 53.000 ;
        RECT 26.840 52.940 26.980 53.095 ;
        RECT 27.210 53.080 27.530 53.340 ;
        RECT 27.670 53.080 27.990 53.340 ;
        RECT 28.220 53.325 28.360 53.480 ;
        RECT 31.350 53.420 31.670 53.480 ;
        RECT 28.145 53.095 28.435 53.325 ;
        RECT 28.590 53.280 28.910 53.340 ;
        RECT 31.900 53.280 32.040 53.820 ;
        RECT 35.030 53.760 35.350 53.820 ;
        RECT 36.410 53.760 36.730 54.020 ;
        RECT 53.430 53.960 53.750 54.020 ;
        RECT 54.825 53.960 55.115 54.005 ;
        RECT 36.960 53.820 53.200 53.960 ;
        RECT 32.270 53.620 32.590 53.680 ;
        RECT 36.960 53.620 37.100 53.820 ;
        RECT 32.270 53.480 37.100 53.620 ;
        RECT 41.025 53.620 41.315 53.665 ;
        RECT 41.930 53.620 42.250 53.680 ;
        RECT 41.025 53.480 42.250 53.620 ;
        RECT 32.270 53.420 32.590 53.480 ;
        RECT 28.590 53.140 32.040 53.280 ;
        RECT 28.590 53.080 28.910 53.140 ;
        RECT 33.205 53.095 33.495 53.325 ;
        RECT 33.650 53.280 33.970 53.340 ;
        RECT 34.660 53.325 34.800 53.480 ;
        RECT 41.025 53.435 41.315 53.480 ;
        RECT 41.930 53.420 42.250 53.480 ;
        RECT 48.830 53.420 49.150 53.680 ;
        RECT 53.060 53.620 53.200 53.820 ;
        RECT 53.430 53.820 55.115 53.960 ;
        RECT 53.430 53.760 53.750 53.820 ;
        RECT 54.825 53.775 55.115 53.820 ;
        RECT 60.805 53.960 61.095 54.005 ;
        RECT 87.945 53.960 88.235 54.005 ;
        RECT 88.390 53.960 88.710 54.020 ;
        RECT 60.805 53.820 87.700 53.960 ;
        RECT 60.805 53.775 61.095 53.820 ;
        RECT 60.880 53.620 61.020 53.775 ;
        RECT 62.645 53.620 62.935 53.665 ;
        RECT 49.380 53.480 52.740 53.620 ;
        RECT 53.060 53.480 61.020 53.620 ;
        RECT 61.340 53.480 62.935 53.620 ;
        RECT 34.125 53.280 34.415 53.325 ;
        RECT 33.650 53.140 34.415 53.280 ;
        RECT 33.280 52.940 33.420 53.095 ;
        RECT 33.650 53.080 33.970 53.140 ;
        RECT 34.125 53.095 34.415 53.140 ;
        RECT 34.585 53.095 34.875 53.325 ;
        RECT 35.030 53.280 35.350 53.340 ;
        RECT 42.850 53.280 43.170 53.340 ;
        RECT 35.030 53.140 43.170 53.280 ;
        RECT 35.030 53.080 35.350 53.140 ;
        RECT 42.850 53.080 43.170 53.140 ;
        RECT 47.450 53.280 47.770 53.340 ;
        RECT 49.380 53.280 49.520 53.480 ;
        RECT 52.600 53.325 52.740 53.480 ;
        RECT 47.450 53.140 49.520 53.280 ;
        RECT 47.450 53.080 47.770 53.140 ;
        RECT 51.605 53.095 51.895 53.325 ;
        RECT 52.525 53.095 52.815 53.325 ;
        RECT 52.985 53.095 53.275 53.325 ;
        RECT 53.445 53.280 53.735 53.325 ;
        RECT 57.570 53.280 57.890 53.340 ;
        RECT 53.445 53.140 57.890 53.280 ;
        RECT 53.445 53.095 53.735 53.140 ;
        RECT 51.130 52.940 51.450 53.000 ;
        RECT 25.830 52.800 51.450 52.940 ;
        RECT 51.680 52.940 51.820 53.095 ;
        RECT 53.060 52.940 53.200 53.095 ;
        RECT 57.570 53.080 57.890 53.140 ;
        RECT 59.870 53.080 60.190 53.340 ;
        RECT 53.890 52.940 54.210 53.000 ;
        RECT 51.680 52.800 52.740 52.940 ;
        RECT 53.060 52.800 54.210 52.940 ;
        RECT 61.340 52.940 61.480 53.480 ;
        RECT 62.645 53.435 62.935 53.480 ;
        RECT 64.945 53.620 65.235 53.665 ;
        RECT 66.770 53.620 67.090 53.680 ;
        RECT 64.945 53.480 67.090 53.620 ;
        RECT 64.945 53.435 65.235 53.480 ;
        RECT 66.770 53.420 67.090 53.480 ;
        RECT 67.690 53.420 68.010 53.680 ;
        RECT 68.150 53.620 68.470 53.680 ;
        RECT 69.545 53.620 69.835 53.665 ;
        RECT 68.150 53.480 69.835 53.620 ;
        RECT 68.150 53.420 68.470 53.480 ;
        RECT 69.545 53.435 69.835 53.480 ;
        RECT 70.450 53.620 70.770 53.680 ;
        RECT 78.730 53.620 79.050 53.680 ;
        RECT 87.560 53.620 87.700 53.820 ;
        RECT 87.945 53.820 88.710 53.960 ;
        RECT 87.945 53.775 88.235 53.820 ;
        RECT 88.390 53.760 88.710 53.820 ;
        RECT 90.230 53.760 90.550 54.020 ;
        RECT 95.305 53.960 95.595 54.005 ;
        RECT 97.130 53.960 97.450 54.020 ;
        RECT 95.305 53.820 97.450 53.960 ;
        RECT 95.305 53.775 95.595 53.820 ;
        RECT 97.130 53.760 97.450 53.820 ;
        RECT 98.970 53.960 99.290 54.020 ;
        RECT 108.185 53.960 108.475 54.005 ;
        RECT 98.970 53.820 112.540 53.960 ;
        RECT 98.970 53.760 99.290 53.820 ;
        RECT 108.185 53.775 108.475 53.820 ;
        RECT 90.320 53.620 90.460 53.760 ;
        RECT 70.450 53.480 86.780 53.620 ;
        RECT 87.560 53.480 90.460 53.620 ;
        RECT 91.150 53.620 91.470 53.680 ;
        RECT 102.190 53.620 102.510 53.680 ;
        RECT 91.150 53.480 92.300 53.620 ;
        RECT 70.450 53.420 70.770 53.480 ;
        RECT 78.730 53.420 79.050 53.480 ;
        RECT 61.725 53.280 62.015 53.325 ;
        RECT 63.550 53.280 63.870 53.340 ;
        RECT 67.780 53.280 67.920 53.420 ;
        RECT 70.005 53.280 70.295 53.325 ;
        RECT 61.725 53.140 70.295 53.280 ;
        RECT 61.725 53.095 62.015 53.140 ;
        RECT 63.550 53.080 63.870 53.140 ;
        RECT 70.005 53.095 70.295 53.140 ;
        RECT 76.890 53.280 77.210 53.340 ;
        RECT 84.725 53.280 85.015 53.325 ;
        RECT 76.890 53.140 85.015 53.280 ;
        RECT 76.890 53.080 77.210 53.140 ;
        RECT 84.725 53.095 85.015 53.140 ;
        RECT 85.645 53.095 85.935 53.325 ;
        RECT 64.930 52.940 65.250 53.000 ;
        RECT 61.340 52.800 65.250 52.940 ;
        RECT 25.830 52.740 26.150 52.800 ;
        RECT 51.130 52.740 51.450 52.800 ;
        RECT 52.600 52.660 52.740 52.800 ;
        RECT 53.890 52.740 54.210 52.800 ;
        RECT 64.930 52.740 65.250 52.800 ;
        RECT 65.405 52.940 65.695 52.985 ;
        RECT 65.850 52.940 66.170 53.000 ;
        RECT 65.405 52.800 66.170 52.940 ;
        RECT 65.405 52.755 65.695 52.800 ;
        RECT 65.850 52.740 66.170 52.800 ;
        RECT 66.310 52.740 66.630 53.000 ;
        RECT 66.770 52.940 67.090 53.000 ;
        RECT 67.245 52.940 67.535 52.985 ;
        RECT 66.770 52.800 67.535 52.940 ;
        RECT 66.770 52.740 67.090 52.800 ;
        RECT 67.245 52.755 67.535 52.800 ;
        RECT 67.705 52.755 67.995 52.985 ;
        RECT 52.510 52.600 52.830 52.660 ;
        RECT 58.965 52.600 59.255 52.645 ;
        RECT 61.250 52.600 61.570 52.660 ;
        RECT 22.700 52.460 26.520 52.600 ;
        RECT 23.070 52.260 23.390 52.320 ;
        RECT 25.830 52.260 26.150 52.320 ;
        RECT 19.940 52.120 26.150 52.260 ;
        RECT 26.380 52.260 26.520 52.460 ;
        RECT 52.510 52.460 61.570 52.600 ;
        RECT 52.510 52.400 52.830 52.460 ;
        RECT 58.965 52.415 59.255 52.460 ;
        RECT 61.250 52.400 61.570 52.460 ;
        RECT 62.630 52.400 62.950 52.660 ;
        RECT 65.940 52.600 66.080 52.740 ;
        RECT 67.780 52.600 67.920 52.755 ;
        RECT 68.150 52.740 68.470 53.000 ;
        RECT 68.625 52.940 68.915 52.985 ;
        RECT 69.070 52.940 69.390 53.000 ;
        RECT 68.625 52.800 69.390 52.940 ;
        RECT 68.625 52.755 68.915 52.800 ;
        RECT 69.070 52.740 69.390 52.800 ;
        RECT 65.940 52.460 67.920 52.600 ;
        RECT 28.590 52.260 28.910 52.320 ;
        RECT 26.380 52.120 28.910 52.260 ;
        RECT 62.720 52.260 62.860 52.400 ;
        RECT 66.310 52.260 66.630 52.320 ;
        RECT 62.720 52.120 66.630 52.260 ;
        RECT 23.070 52.060 23.390 52.120 ;
        RECT 25.830 52.060 26.150 52.120 ;
        RECT 28.590 52.060 28.910 52.120 ;
        RECT 66.310 52.060 66.630 52.120 ;
        RECT 67.230 52.260 67.550 52.320 ;
        RECT 70.925 52.260 71.215 52.305 ;
        RECT 78.270 52.260 78.590 52.320 ;
        RECT 83.790 52.260 84.110 52.320 ;
        RECT 67.230 52.120 84.110 52.260 ;
        RECT 84.800 52.260 84.940 53.095 ;
        RECT 85.720 52.940 85.860 53.095 ;
        RECT 86.090 53.080 86.410 53.340 ;
        RECT 86.640 53.325 86.780 53.480 ;
        RECT 91.150 53.420 91.470 53.480 ;
        RECT 86.565 53.280 86.855 53.325 ;
        RECT 89.310 53.280 89.630 53.340 ;
        RECT 89.785 53.280 90.075 53.325 ;
        RECT 86.565 53.140 90.075 53.280 ;
        RECT 86.565 53.095 86.855 53.140 ;
        RECT 89.310 53.080 89.630 53.140 ;
        RECT 89.785 53.095 90.075 53.140 ;
        RECT 90.245 53.095 90.535 53.325 ;
        RECT 90.705 53.095 90.995 53.325 ;
        RECT 87.010 52.940 87.330 53.000 ;
        RECT 90.320 52.940 90.460 53.095 ;
        RECT 85.720 52.800 87.330 52.940 ;
        RECT 87.010 52.740 87.330 52.800 ;
        RECT 87.560 52.800 90.460 52.940 ;
        RECT 90.780 52.940 90.920 53.095 ;
        RECT 91.610 53.080 91.930 53.340 ;
        RECT 92.160 53.325 92.300 53.480 ;
        RECT 93.080 53.480 102.510 53.620 ;
        RECT 93.080 53.325 93.220 53.480 ;
        RECT 102.190 53.420 102.510 53.480 ;
        RECT 103.105 53.620 103.755 53.665 ;
        RECT 106.705 53.620 106.995 53.665 ;
        RECT 111.850 53.620 112.170 53.680 ;
        RECT 103.105 53.480 112.170 53.620 ;
        RECT 103.105 53.435 103.755 53.480 ;
        RECT 106.405 53.435 106.995 53.480 ;
        RECT 92.085 53.095 92.375 53.325 ;
        RECT 93.005 53.095 93.295 53.325 ;
        RECT 93.465 53.095 93.755 53.325 ;
        RECT 93.925 53.095 94.215 53.325 ;
        RECT 99.910 53.280 100.200 53.325 ;
        RECT 101.745 53.280 102.035 53.325 ;
        RECT 105.325 53.280 105.615 53.325 ;
        RECT 99.910 53.140 105.615 53.280 ;
        RECT 99.910 53.095 100.200 53.140 ;
        RECT 101.745 53.095 102.035 53.140 ;
        RECT 105.325 53.095 105.615 53.140 ;
        RECT 92.530 52.940 92.850 53.000 ;
        RECT 90.780 52.800 92.850 52.940 ;
        RECT 86.090 52.600 86.410 52.660 ;
        RECT 87.560 52.600 87.700 52.800 ;
        RECT 86.090 52.460 87.700 52.600 ;
        RECT 88.405 52.600 88.695 52.645 ;
        RECT 89.770 52.600 90.090 52.660 ;
        RECT 88.405 52.460 90.090 52.600 ;
        RECT 90.320 52.600 90.460 52.800 ;
        RECT 92.530 52.740 92.850 52.800 ;
        RECT 93.540 52.600 93.680 53.095 ;
        RECT 90.320 52.460 93.680 52.600 ;
        RECT 86.090 52.400 86.410 52.460 ;
        RECT 88.405 52.415 88.695 52.460 ;
        RECT 89.770 52.400 90.090 52.460 ;
        RECT 87.470 52.260 87.790 52.320 ;
        RECT 84.800 52.120 87.790 52.260 ;
        RECT 67.230 52.060 67.550 52.120 ;
        RECT 70.925 52.075 71.215 52.120 ;
        RECT 78.270 52.060 78.590 52.120 ;
        RECT 83.790 52.060 84.110 52.120 ;
        RECT 87.470 52.060 87.790 52.120 ;
        RECT 89.310 52.260 89.630 52.320 ;
        RECT 94.000 52.260 94.140 53.095 ;
        RECT 105.870 53.080 106.190 53.340 ;
        RECT 106.405 53.120 106.695 53.435 ;
        RECT 111.850 53.420 112.170 53.480 ;
        RECT 112.400 53.325 112.540 53.820 ;
        RECT 112.770 53.760 113.090 54.020 ;
        RECT 113.690 53.620 114.010 53.680 ;
        RECT 113.690 53.480 116.220 53.620 ;
        RECT 113.690 53.420 114.010 53.480 ;
        RECT 112.325 53.095 112.615 53.325 ;
        RECT 114.150 53.080 114.470 53.340 ;
        RECT 114.625 53.095 114.915 53.325 ;
        RECT 96.225 52.940 96.515 52.985 ;
        RECT 98.050 52.940 98.370 53.000 ;
        RECT 96.225 52.800 98.370 52.940 ;
        RECT 96.225 52.755 96.515 52.800 ;
        RECT 98.050 52.740 98.370 52.800 ;
        RECT 99.445 52.755 99.735 52.985 ;
        RECT 100.825 52.940 101.115 52.985 ;
        RECT 102.650 52.940 102.970 53.000 ;
        RECT 100.825 52.800 102.970 52.940 ;
        RECT 105.960 52.940 106.100 53.080 ;
        RECT 114.700 52.940 114.840 53.095 ;
        RECT 115.070 53.080 115.390 53.340 ;
        RECT 116.080 53.325 116.220 53.480 ;
        RECT 116.005 53.095 116.295 53.325 ;
        RECT 105.960 52.800 114.840 52.940 ;
        RECT 100.825 52.755 101.115 52.800 ;
        RECT 89.310 52.120 94.140 52.260 ;
        RECT 89.310 52.060 89.630 52.120 ;
        RECT 98.970 52.060 99.290 52.320 ;
        RECT 99.520 52.260 99.660 52.755 ;
        RECT 102.650 52.740 102.970 52.800 ;
        RECT 100.315 52.600 100.605 52.645 ;
        RECT 102.205 52.600 102.495 52.645 ;
        RECT 105.325 52.600 105.615 52.645 ;
        RECT 100.315 52.460 105.615 52.600 ;
        RECT 100.315 52.415 100.605 52.460 ;
        RECT 102.205 52.415 102.495 52.460 ;
        RECT 105.325 52.415 105.615 52.460 ;
        RECT 105.870 52.600 106.190 52.660 ;
        RECT 109.105 52.600 109.395 52.645 ;
        RECT 105.870 52.460 109.395 52.600 ;
        RECT 105.870 52.400 106.190 52.460 ;
        RECT 109.105 52.415 109.395 52.460 ;
        RECT 107.710 52.260 108.030 52.320 ;
        RECT 99.520 52.120 108.030 52.260 ;
        RECT 107.710 52.060 108.030 52.120 ;
        RECT 5.520 51.440 125.580 51.920 ;
        RECT 29.065 51.240 29.355 51.285 ;
        RECT 30.430 51.240 30.750 51.300 ;
        RECT 47.910 51.240 48.230 51.300 ;
        RECT 29.065 51.100 30.750 51.240 ;
        RECT 29.065 51.055 29.355 51.100 ;
        RECT 30.430 51.040 30.750 51.100 ;
        RECT 36.040 51.100 48.230 51.240 ;
        RECT 35.505 50.560 35.795 50.605 ;
        RECT 36.040 50.560 36.180 51.100 ;
        RECT 47.910 51.040 48.230 51.100 ;
        RECT 56.205 51.240 56.495 51.285 ;
        RECT 56.650 51.240 56.970 51.300 ;
        RECT 67.230 51.240 67.550 51.300 ;
        RECT 56.205 51.100 56.970 51.240 ;
        RECT 56.205 51.055 56.495 51.100 ;
        RECT 56.650 51.040 56.970 51.100 ;
        RECT 60.880 51.100 67.550 51.240 ;
        RECT 38.265 50.900 38.555 50.945 ;
        RECT 55.745 50.900 56.035 50.945 ;
        RECT 60.330 50.900 60.650 50.960 ;
        RECT 38.265 50.760 41.700 50.900 ;
        RECT 38.265 50.715 38.555 50.760 ;
        RECT 41.560 50.605 41.700 50.760 ;
        RECT 55.745 50.760 60.650 50.900 ;
        RECT 55.745 50.715 56.035 50.760 ;
        RECT 60.330 50.700 60.650 50.760 ;
        RECT 35.505 50.420 36.180 50.560 ;
        RECT 35.505 50.375 35.795 50.420 ;
        RECT 41.485 50.375 41.775 50.605 ;
        RECT 60.880 50.560 61.020 51.100 ;
        RECT 67.230 51.040 67.550 51.100 ;
        RECT 80.110 51.040 80.430 51.300 ;
        RECT 83.790 51.240 84.110 51.300 ;
        RECT 86.090 51.240 86.410 51.300 ;
        RECT 83.790 51.100 86.410 51.240 ;
        RECT 83.790 51.040 84.110 51.100 ;
        RECT 86.090 51.040 86.410 51.100 ;
        RECT 90.690 51.240 91.010 51.300 ;
        RECT 95.290 51.240 95.610 51.300 ;
        RECT 90.690 51.100 95.610 51.240 ;
        RECT 90.690 51.040 91.010 51.100 ;
        RECT 95.290 51.040 95.610 51.100 ;
        RECT 98.050 51.040 98.370 51.300 ;
        RECT 102.205 51.240 102.495 51.285 ;
        RECT 102.650 51.240 102.970 51.300 ;
        RECT 114.150 51.240 114.470 51.300 ;
        RECT 115.070 51.240 115.390 51.300 ;
        RECT 116.465 51.240 116.755 51.285 ;
        RECT 102.205 51.100 102.970 51.240 ;
        RECT 102.205 51.055 102.495 51.100 ;
        RECT 102.650 51.040 102.970 51.100 ;
        RECT 105.040 51.100 116.755 51.240 ;
        RECT 64.010 50.900 64.330 50.960 ;
        RECT 64.485 50.900 64.775 50.945 ;
        RECT 64.010 50.760 64.775 50.900 ;
        RECT 64.010 50.700 64.330 50.760 ;
        RECT 64.485 50.715 64.775 50.760 ;
        RECT 65.480 50.760 67.000 50.900 ;
        RECT 65.480 50.620 65.620 50.760 ;
        RECT 53.980 50.420 61.020 50.560 ;
        RECT 61.710 50.560 62.030 50.620 ;
        RECT 62.185 50.560 62.475 50.605 ;
        RECT 61.710 50.420 62.475 50.560 ;
        RECT 53.980 50.280 54.120 50.420 ;
        RECT 13.870 50.020 14.190 50.280 ;
        RECT 15.265 50.220 15.555 50.265 ;
        RECT 20.770 50.220 21.090 50.280 ;
        RECT 15.265 50.080 21.090 50.220 ;
        RECT 15.265 50.035 15.555 50.080 ;
        RECT 20.770 50.020 21.090 50.080 ;
        RECT 22.150 50.020 22.470 50.280 ;
        RECT 25.830 50.020 26.150 50.280 ;
        RECT 26.765 50.035 27.055 50.265 ;
        RECT 22.240 49.880 22.380 50.020 ;
        RECT 26.840 49.880 26.980 50.035 ;
        RECT 27.210 50.020 27.530 50.280 ;
        RECT 27.685 50.220 27.975 50.265 ;
        RECT 28.590 50.220 28.910 50.280 ;
        RECT 27.685 50.080 28.910 50.220 ;
        RECT 27.685 50.035 27.975 50.080 ;
        RECT 28.590 50.020 28.910 50.080 ;
        RECT 32.270 50.020 32.590 50.280 ;
        RECT 42.865 50.220 43.155 50.265 ;
        RECT 45.625 50.220 45.915 50.265 ;
        RECT 42.865 50.080 45.915 50.220 ;
        RECT 42.865 50.035 43.155 50.080 ;
        RECT 45.625 50.035 45.915 50.080 ;
        RECT 48.370 50.020 48.690 50.280 ;
        RECT 50.670 50.220 50.990 50.280 ;
        RECT 51.605 50.220 51.895 50.265 ;
        RECT 50.670 50.080 51.895 50.220 ;
        RECT 50.670 50.020 50.990 50.080 ;
        RECT 51.605 50.035 51.895 50.080 ;
        RECT 52.510 50.020 52.830 50.280 ;
        RECT 53.430 50.020 53.750 50.280 ;
        RECT 53.890 50.020 54.210 50.280 ;
        RECT 54.365 50.220 54.655 50.265 ;
        RECT 57.570 50.220 57.890 50.280 ;
        RECT 58.120 50.265 58.260 50.420 ;
        RECT 61.710 50.360 62.030 50.420 ;
        RECT 62.185 50.375 62.475 50.420 ;
        RECT 62.630 50.360 62.950 50.620 ;
        RECT 65.390 50.560 65.710 50.620 ;
        RECT 64.100 50.420 65.710 50.560 ;
        RECT 54.365 50.080 57.890 50.220 ;
        RECT 54.365 50.035 54.655 50.080 ;
        RECT 57.570 50.020 57.890 50.080 ;
        RECT 58.045 50.035 58.335 50.265 ;
        RECT 58.490 50.020 58.810 50.280 ;
        RECT 59.425 50.220 59.715 50.265 ;
        RECT 61.250 50.220 61.570 50.280 ;
        RECT 59.425 50.080 61.570 50.220 ;
        RECT 59.425 50.035 59.715 50.080 ;
        RECT 61.250 50.020 61.570 50.080 ;
        RECT 63.105 50.035 63.395 50.265 ;
        RECT 63.580 50.230 63.870 50.265 ;
        RECT 64.100 50.230 64.240 50.420 ;
        RECT 65.390 50.360 65.710 50.420 ;
        RECT 66.310 50.360 66.630 50.620 ;
        RECT 66.860 50.560 67.000 50.760 ;
        RECT 67.690 50.700 68.010 50.960 ;
        RECT 78.270 50.700 78.590 50.960 ;
        RECT 87.435 50.900 87.725 50.945 ;
        RECT 89.325 50.900 89.615 50.945 ;
        RECT 92.445 50.900 92.735 50.945 ;
        RECT 87.435 50.760 92.735 50.900 ;
        RECT 87.435 50.715 87.725 50.760 ;
        RECT 89.325 50.715 89.615 50.760 ;
        RECT 92.445 50.715 92.735 50.760 ;
        RECT 68.150 50.560 68.470 50.620 ;
        RECT 66.860 50.420 68.470 50.560 ;
        RECT 68.150 50.360 68.470 50.420 ;
        RECT 63.580 50.090 64.240 50.230 ;
        RECT 63.580 50.035 63.870 50.090 ;
        RECT 22.240 49.740 26.980 49.880 ;
        RECT 35.965 49.880 36.255 49.925 ;
        RECT 41.470 49.880 41.790 49.940 ;
        RECT 35.965 49.740 41.790 49.880 ;
        RECT 35.965 49.695 36.255 49.740 ;
        RECT 41.470 49.680 41.790 49.740 ;
        RECT 50.210 49.680 50.530 49.940 ;
        RECT 63.180 49.880 63.320 50.035 ;
        RECT 65.850 50.020 66.170 50.280 ;
        RECT 66.770 50.020 67.090 50.280 ;
        RECT 69.070 50.020 69.390 50.280 ;
        RECT 74.590 50.020 74.910 50.280 ;
        RECT 76.890 50.020 77.210 50.280 ;
        RECT 78.360 50.265 78.500 50.700 ;
        RECT 89.770 50.560 90.090 50.620 ;
        RECT 85.260 50.420 90.090 50.560 ;
        RECT 78.730 50.265 79.050 50.290 ;
        RECT 77.720 50.220 78.010 50.265 ;
        RECT 77.670 50.035 78.010 50.220 ;
        RECT 78.300 50.035 78.590 50.265 ;
        RECT 78.730 50.035 79.265 50.265 ;
        RECT 82.870 50.220 83.190 50.280 ;
        RECT 85.260 50.265 85.400 50.420 ;
        RECT 89.770 50.360 90.090 50.420 ;
        RECT 98.510 50.560 98.830 50.620 ;
        RECT 100.365 50.560 100.655 50.605 ;
        RECT 98.510 50.420 100.655 50.560 ;
        RECT 98.510 50.360 98.830 50.420 ;
        RECT 100.365 50.375 100.655 50.420 ;
        RECT 101.285 50.560 101.575 50.605 ;
        RECT 103.570 50.560 103.890 50.620 ;
        RECT 105.040 50.605 105.180 51.100 ;
        RECT 114.150 51.040 114.470 51.100 ;
        RECT 115.070 51.040 115.390 51.100 ;
        RECT 116.465 51.055 116.755 51.100 ;
        RECT 108.595 50.900 108.885 50.945 ;
        RECT 110.485 50.900 110.775 50.945 ;
        RECT 113.605 50.900 113.895 50.945 ;
        RECT 108.595 50.760 113.895 50.900 ;
        RECT 108.595 50.715 108.885 50.760 ;
        RECT 110.485 50.715 110.775 50.760 ;
        RECT 113.605 50.715 113.895 50.760 ;
        RECT 104.045 50.560 104.335 50.605 ;
        RECT 101.285 50.420 104.335 50.560 ;
        RECT 101.285 50.375 101.575 50.420 ;
        RECT 103.570 50.360 103.890 50.420 ;
        RECT 104.045 50.375 104.335 50.420 ;
        RECT 104.965 50.375 105.255 50.605 ;
        RECT 107.710 50.360 108.030 50.620 ;
        RECT 83.345 50.220 83.635 50.265 ;
        RECT 82.870 50.080 83.635 50.220 ;
        RECT 61.800 49.740 63.320 49.880 ;
        RECT 64.010 49.880 64.330 49.940 ;
        RECT 65.940 49.880 66.080 50.020 ;
        RECT 64.010 49.740 66.080 49.880 ;
        RECT 66.310 49.880 66.630 49.940 ;
        RECT 76.980 49.880 77.120 50.020 ;
        RECT 66.310 49.740 77.120 49.880 ;
        RECT 77.670 49.880 77.810 50.035 ;
        RECT 78.730 50.030 79.050 50.035 ;
        RECT 82.870 50.020 83.190 50.080 ;
        RECT 83.345 50.035 83.635 50.080 ;
        RECT 85.185 50.035 85.475 50.265 ;
        RECT 86.565 50.035 86.855 50.265 ;
        RECT 87.030 50.220 87.320 50.265 ;
        RECT 88.865 50.220 89.155 50.265 ;
        RECT 92.445 50.220 92.735 50.265 ;
        RECT 87.030 50.080 92.735 50.220 ;
        RECT 87.030 50.035 87.320 50.080 ;
        RECT 88.865 50.035 89.155 50.080 ;
        RECT 92.445 50.035 92.735 50.080 ;
        RECT 79.650 49.880 79.970 49.940 ;
        RECT 86.640 49.880 86.780 50.035 ;
        RECT 93.525 49.925 93.815 50.240 ;
        RECT 97.145 50.220 97.435 50.265 ;
        RECT 97.590 50.220 97.910 50.280 ;
        RECT 97.145 50.080 97.910 50.220 ;
        RECT 97.145 50.035 97.435 50.080 ;
        RECT 97.590 50.020 97.910 50.080 ;
        RECT 98.970 50.220 99.290 50.280 ;
        RECT 103.125 50.220 103.415 50.265 ;
        RECT 98.970 50.080 103.415 50.220 ;
        RECT 98.970 50.020 99.290 50.080 ;
        RECT 103.125 50.035 103.415 50.080 ;
        RECT 105.425 50.220 105.715 50.265 ;
        RECT 105.870 50.220 106.190 50.280 ;
        RECT 105.425 50.080 106.190 50.220 ;
        RECT 105.425 50.035 105.715 50.080 ;
        RECT 105.870 50.020 106.190 50.080 ;
        RECT 108.190 50.220 108.480 50.265 ;
        RECT 110.025 50.220 110.315 50.265 ;
        RECT 113.605 50.220 113.895 50.265 ;
        RECT 108.190 50.080 113.895 50.220 ;
        RECT 108.190 50.035 108.480 50.080 ;
        RECT 110.025 50.035 110.315 50.080 ;
        RECT 113.605 50.035 113.895 50.080 ;
        RECT 77.670 49.740 79.970 49.880 ;
        RECT 61.800 49.600 61.940 49.740 ;
        RECT 64.010 49.680 64.330 49.740 ;
        RECT 66.310 49.680 66.630 49.740 ;
        RECT 79.650 49.680 79.970 49.740 ;
        RECT 83.420 49.740 86.780 49.880 ;
        RECT 83.420 49.600 83.560 49.740 ;
        RECT 87.945 49.695 88.235 49.925 ;
        RECT 90.225 49.880 90.875 49.925 ;
        RECT 93.525 49.880 94.115 49.925 ;
        RECT 96.685 49.880 96.975 49.925 ;
        RECT 90.225 49.740 96.975 49.880 ;
        RECT 90.225 49.695 90.875 49.740 ;
        RECT 93.825 49.695 94.115 49.740 ;
        RECT 96.685 49.695 96.975 49.740 ;
        RECT 12.030 49.540 12.350 49.600 ;
        RECT 12.965 49.540 13.255 49.585 ;
        RECT 12.030 49.400 13.255 49.540 ;
        RECT 12.030 49.340 12.350 49.400 ;
        RECT 12.965 49.355 13.255 49.400 ;
        RECT 14.330 49.340 14.650 49.600 ;
        RECT 23.070 49.540 23.390 49.600 ;
        RECT 25.385 49.540 25.675 49.585 ;
        RECT 23.070 49.400 25.675 49.540 ;
        RECT 23.070 49.340 23.390 49.400 ;
        RECT 25.385 49.355 25.675 49.400 ;
        RECT 29.510 49.340 29.830 49.600 ;
        RECT 36.410 49.340 36.730 49.600 ;
        RECT 38.710 49.340 39.030 49.600 ;
        RECT 43.770 49.340 44.090 49.600 ;
        RECT 61.710 49.340 62.030 49.600 ;
        RECT 62.170 49.540 62.490 49.600 ;
        RECT 68.625 49.540 68.915 49.585 ;
        RECT 62.170 49.400 68.915 49.540 ;
        RECT 62.170 49.340 62.490 49.400 ;
        RECT 68.625 49.355 68.915 49.400 ;
        RECT 75.970 49.340 76.290 49.600 ;
        RECT 76.430 49.540 76.750 49.600 ;
        RECT 80.585 49.540 80.875 49.585 ;
        RECT 76.430 49.400 80.875 49.540 ;
        RECT 76.430 49.340 76.750 49.400 ;
        RECT 80.585 49.355 80.875 49.400 ;
        RECT 83.330 49.340 83.650 49.600 ;
        RECT 86.105 49.540 86.395 49.585 ;
        RECT 88.020 49.540 88.160 49.695 ;
        RECT 109.090 49.680 109.410 49.940 ;
        RECT 111.850 49.925 112.170 49.940 ;
        RECT 111.385 49.880 112.170 49.925 ;
        RECT 114.685 49.925 114.975 50.240 ;
        RECT 114.685 49.880 115.275 49.925 ;
        RECT 111.385 49.740 115.275 49.880 ;
        RECT 111.385 49.695 112.170 49.740 ;
        RECT 114.985 49.695 115.275 49.740 ;
        RECT 111.850 49.680 112.170 49.695 ;
        RECT 86.105 49.400 88.160 49.540 ;
        RECT 86.105 49.355 86.395 49.400 ;
        RECT 99.890 49.340 100.210 49.600 ;
        RECT 107.265 49.540 107.555 49.585 ;
        RECT 110.930 49.540 111.250 49.600 ;
        RECT 107.265 49.400 111.250 49.540 ;
        RECT 107.265 49.355 107.555 49.400 ;
        RECT 110.930 49.340 111.250 49.400 ;
        RECT 5.520 48.720 125.580 49.200 ;
        RECT 20.770 48.320 21.090 48.580 ;
        RECT 23.070 48.320 23.390 48.580 ;
        RECT 30.445 48.520 30.735 48.565 ;
        RECT 32.270 48.520 32.590 48.580 ;
        RECT 30.445 48.380 32.590 48.520 ;
        RECT 30.445 48.335 30.735 48.380 ;
        RECT 32.270 48.320 32.590 48.380 ;
        RECT 41.470 48.520 41.790 48.580 ;
        RECT 47.450 48.520 47.770 48.580 ;
        RECT 41.470 48.380 47.770 48.520 ;
        RECT 41.470 48.320 41.790 48.380 ;
        RECT 47.450 48.320 47.770 48.380 ;
        RECT 53.890 48.320 54.210 48.580 ;
        RECT 54.810 48.520 55.130 48.580 ;
        RECT 57.570 48.520 57.890 48.580 ;
        RECT 54.810 48.380 57.890 48.520 ;
        RECT 54.810 48.320 55.130 48.380 ;
        RECT 57.570 48.320 57.890 48.380 ;
        RECT 61.710 48.520 62.030 48.580 ;
        RECT 63.550 48.520 63.870 48.580 ;
        RECT 89.310 48.520 89.630 48.580 ;
        RECT 61.710 48.380 63.870 48.520 ;
        RECT 61.710 48.320 62.030 48.380 ;
        RECT 63.550 48.320 63.870 48.380 ;
        RECT 82.960 48.380 89.630 48.520 ;
        RECT 12.965 48.180 13.255 48.225 ;
        RECT 14.330 48.180 14.650 48.240 ;
        RECT 12.965 48.040 14.650 48.180 ;
        RECT 12.965 47.995 13.255 48.040 ;
        RECT 14.330 47.980 14.650 48.040 ;
        RECT 15.245 48.180 15.895 48.225 ;
        RECT 18.010 48.180 18.330 48.240 ;
        RECT 18.845 48.180 19.135 48.225 ;
        RECT 15.245 48.040 19.135 48.180 ;
        RECT 23.160 48.180 23.300 48.320 ;
        RECT 28.605 48.180 28.895 48.225 ;
        RECT 33.650 48.180 33.970 48.240 ;
        RECT 23.160 48.040 28.895 48.180 ;
        RECT 15.245 47.995 15.895 48.040 ;
        RECT 18.010 47.980 18.330 48.040 ;
        RECT 18.545 47.995 19.135 48.040 ;
        RECT 28.605 47.995 28.895 48.040 ;
        RECT 32.820 48.040 33.970 48.180 ;
        RECT 7.430 47.840 7.750 47.900 ;
        RECT 11.585 47.840 11.875 47.885 ;
        RECT 7.430 47.700 11.875 47.840 ;
        RECT 7.430 47.640 7.750 47.700 ;
        RECT 11.585 47.655 11.875 47.700 ;
        RECT 12.050 47.840 12.340 47.885 ;
        RECT 13.885 47.840 14.175 47.885 ;
        RECT 17.465 47.840 17.755 47.885 ;
        RECT 12.050 47.700 17.755 47.840 ;
        RECT 12.050 47.655 12.340 47.700 ;
        RECT 13.885 47.655 14.175 47.700 ;
        RECT 17.465 47.655 17.755 47.700 ;
        RECT 18.545 47.680 18.835 47.995 ;
        RECT 21.230 47.840 21.550 47.900 ;
        RECT 22.625 47.840 22.915 47.885 ;
        RECT 21.230 47.700 22.915 47.840 ;
        RECT 21.230 47.640 21.550 47.700 ;
        RECT 22.625 47.655 22.915 47.700 ;
        RECT 28.145 47.840 28.435 47.885 ;
        RECT 32.820 47.840 32.960 48.040 ;
        RECT 33.650 47.980 33.970 48.040 ;
        RECT 36.405 48.180 37.055 48.225 ;
        RECT 39.170 48.180 39.490 48.240 ;
        RECT 40.005 48.180 40.295 48.225 ;
        RECT 36.405 48.040 40.295 48.180 ;
        RECT 36.405 47.995 37.055 48.040 ;
        RECT 39.170 47.980 39.490 48.040 ;
        RECT 39.705 47.995 40.295 48.040 ;
        RECT 43.770 48.180 44.090 48.240 ;
        RECT 44.245 48.180 44.535 48.225 ;
        RECT 43.770 48.040 44.535 48.180 ;
        RECT 28.145 47.700 32.960 47.840 ;
        RECT 33.210 47.840 33.500 47.885 ;
        RECT 35.045 47.840 35.335 47.885 ;
        RECT 38.625 47.840 38.915 47.885 ;
        RECT 33.210 47.700 38.915 47.840 ;
        RECT 28.145 47.655 28.435 47.700 ;
        RECT 33.210 47.655 33.500 47.700 ;
        RECT 35.045 47.655 35.335 47.700 ;
        RECT 38.625 47.655 38.915 47.700 ;
        RECT 39.705 47.680 39.995 47.995 ;
        RECT 43.770 47.980 44.090 48.040 ;
        RECT 44.245 47.995 44.535 48.040 ;
        RECT 46.525 48.180 47.175 48.225 ;
        RECT 50.125 48.180 50.415 48.225 ;
        RECT 53.980 48.180 54.120 48.320 ;
        RECT 46.525 48.040 50.415 48.180 ;
        RECT 46.525 47.995 47.175 48.040 ;
        RECT 49.825 47.995 50.415 48.040 ;
        RECT 53.520 48.040 54.120 48.180 ;
        RECT 43.330 47.840 43.620 47.885 ;
        RECT 45.165 47.840 45.455 47.885 ;
        RECT 48.745 47.840 49.035 47.885 ;
        RECT 43.330 47.700 49.035 47.840 ;
        RECT 43.330 47.655 43.620 47.700 ;
        RECT 45.165 47.655 45.455 47.700 ;
        RECT 48.745 47.655 49.035 47.700 ;
        RECT 49.825 47.680 50.115 47.995 ;
        RECT 52.065 47.840 52.355 47.885 ;
        RECT 52.510 47.840 52.830 47.900 ;
        RECT 52.065 47.700 52.830 47.840 ;
        RECT 20.325 47.500 20.615 47.545 ;
        RECT 22.150 47.500 22.470 47.560 ;
        RECT 20.325 47.360 22.470 47.500 ;
        RECT 20.325 47.315 20.615 47.360 ;
        RECT 22.150 47.300 22.470 47.360 ;
        RECT 23.070 47.500 23.390 47.560 ;
        RECT 24.005 47.500 24.295 47.545 ;
        RECT 26.750 47.500 27.070 47.560 ;
        RECT 27.225 47.500 27.515 47.545 ;
        RECT 23.070 47.360 27.515 47.500 ;
        RECT 23.070 47.300 23.390 47.360 ;
        RECT 24.005 47.315 24.295 47.360 ;
        RECT 26.750 47.300 27.070 47.360 ;
        RECT 27.225 47.315 27.515 47.360 ;
        RECT 32.745 47.500 33.035 47.545 ;
        RECT 32.745 47.360 33.420 47.500 ;
        RECT 32.745 47.315 33.035 47.360 ;
        RECT 12.455 47.160 12.745 47.205 ;
        RECT 14.345 47.160 14.635 47.205 ;
        RECT 17.465 47.160 17.755 47.205 ;
        RECT 12.455 47.020 17.755 47.160 ;
        RECT 12.455 46.975 12.745 47.020 ;
        RECT 14.345 46.975 14.635 47.020 ;
        RECT 17.465 46.975 17.755 47.020 ;
        RECT 33.280 46.820 33.420 47.360 ;
        RECT 34.110 47.300 34.430 47.560 ;
        RECT 42.865 47.500 43.155 47.545 ;
        RECT 49.840 47.500 49.980 47.680 ;
        RECT 52.065 47.655 52.355 47.700 ;
        RECT 52.510 47.640 52.830 47.700 ;
        RECT 52.970 47.640 53.290 47.900 ;
        RECT 53.520 47.885 53.660 48.040 ;
        RECT 55.270 47.980 55.590 48.240 ;
        RECT 64.470 48.180 64.790 48.240 ;
        RECT 64.945 48.180 65.235 48.225 ;
        RECT 64.470 48.040 65.235 48.180 ;
        RECT 64.470 47.980 64.790 48.040 ;
        RECT 64.945 47.995 65.235 48.040 ;
        RECT 53.445 47.655 53.735 47.885 ;
        RECT 53.905 47.840 54.195 47.885 ;
        RECT 54.810 47.840 55.130 47.900 ;
        RECT 53.905 47.700 55.130 47.840 ;
        RECT 53.905 47.655 54.195 47.700 ;
        RECT 54.810 47.640 55.130 47.700 ;
        RECT 55.745 47.840 56.035 47.885 ;
        RECT 62.170 47.840 62.490 47.900 ;
        RECT 63.550 47.840 63.870 47.900 ;
        RECT 66.770 47.840 67.090 47.900 ;
        RECT 55.745 47.700 56.880 47.840 ;
        RECT 55.745 47.655 56.035 47.700 ;
        RECT 56.205 47.500 56.495 47.545 ;
        RECT 42.865 47.360 43.540 47.500 ;
        RECT 49.840 47.360 56.495 47.500 ;
        RECT 42.865 47.315 43.155 47.360 ;
        RECT 33.615 47.160 33.905 47.205 ;
        RECT 35.505 47.160 35.795 47.205 ;
        RECT 38.625 47.160 38.915 47.205 ;
        RECT 42.390 47.160 42.710 47.220 ;
        RECT 43.400 47.160 43.540 47.360 ;
        RECT 56.205 47.315 56.495 47.360 ;
        RECT 33.615 47.020 38.915 47.160 ;
        RECT 33.615 46.975 33.905 47.020 ;
        RECT 35.505 46.975 35.795 47.020 ;
        RECT 38.625 46.975 38.915 47.020 ;
        RECT 39.260 47.020 43.540 47.160 ;
        RECT 39.260 46.820 39.400 47.020 ;
        RECT 42.390 46.960 42.710 47.020 ;
        RECT 33.280 46.680 39.400 46.820 ;
        RECT 43.400 46.820 43.540 47.020 ;
        RECT 43.735 47.160 44.025 47.205 ;
        RECT 45.625 47.160 45.915 47.205 ;
        RECT 48.745 47.160 49.035 47.205 ;
        RECT 43.735 47.020 49.035 47.160 ;
        RECT 43.735 46.975 44.025 47.020 ;
        RECT 45.625 46.975 45.915 47.020 ;
        RECT 48.745 46.975 49.035 47.020 ;
        RECT 50.210 47.160 50.530 47.220 ;
        RECT 56.740 47.160 56.880 47.700 ;
        RECT 62.170 47.700 67.090 47.840 ;
        RECT 62.170 47.640 62.490 47.700 ;
        RECT 63.550 47.640 63.870 47.700 ;
        RECT 66.770 47.640 67.090 47.700 ;
        RECT 76.430 47.640 76.750 47.900 ;
        RECT 77.810 47.840 78.130 47.900 ;
        RECT 78.745 47.840 79.035 47.885 ;
        RECT 77.810 47.700 79.035 47.840 ;
        RECT 82.960 47.840 83.100 48.380 ;
        RECT 89.310 48.320 89.630 48.380 ;
        RECT 89.770 48.320 90.090 48.580 ;
        RECT 108.185 48.520 108.475 48.565 ;
        RECT 109.090 48.520 109.410 48.580 ;
        RECT 108.185 48.380 109.410 48.520 ;
        RECT 108.185 48.335 108.475 48.380 ;
        RECT 109.090 48.320 109.410 48.380 ;
        RECT 83.790 48.180 84.110 48.240 ;
        RECT 88.390 48.180 88.710 48.240 ;
        RECT 83.790 48.040 88.710 48.180 ;
        RECT 83.790 47.980 84.110 48.040 ;
        RECT 84.710 47.840 85.030 47.900 ;
        RECT 85.260 47.885 85.400 48.040 ;
        RECT 88.390 47.980 88.710 48.040 ;
        RECT 92.085 48.180 92.375 48.225 ;
        RECT 99.890 48.180 100.210 48.240 ;
        RECT 101.285 48.180 101.575 48.225 ;
        RECT 92.085 48.040 101.575 48.180 ;
        RECT 92.085 47.995 92.375 48.040 ;
        RECT 99.890 47.980 100.210 48.040 ;
        RECT 101.285 47.995 101.575 48.040 ;
        RECT 82.960 47.700 85.030 47.840 ;
        RECT 77.810 47.640 78.130 47.700 ;
        RECT 78.745 47.655 79.035 47.700 ;
        RECT 84.710 47.640 85.030 47.700 ;
        RECT 85.185 47.655 85.475 47.885 ;
        RECT 85.645 47.655 85.935 47.885 ;
        RECT 86.565 47.840 86.855 47.885 ;
        RECT 87.470 47.840 87.790 47.900 ;
        RECT 91.150 47.840 91.470 47.900 ;
        RECT 86.565 47.700 91.470 47.840 ;
        RECT 86.565 47.655 86.855 47.700 ;
        RECT 62.630 47.300 62.950 47.560 ;
        RECT 63.105 47.315 63.395 47.545 ;
        RECT 64.025 47.500 64.315 47.545 ;
        RECT 65.390 47.500 65.710 47.560 ;
        RECT 64.025 47.360 65.710 47.500 ;
        RECT 64.025 47.315 64.315 47.360 ;
        RECT 50.210 47.020 56.880 47.160 ;
        RECT 63.180 47.160 63.320 47.315 ;
        RECT 65.390 47.300 65.710 47.360 ;
        RECT 75.970 47.500 76.290 47.560 ;
        RECT 77.365 47.500 77.655 47.545 ;
        RECT 75.970 47.360 77.655 47.500 ;
        RECT 75.970 47.300 76.290 47.360 ;
        RECT 77.365 47.315 77.655 47.360 ;
        RECT 78.285 47.500 78.575 47.545 ;
        RECT 82.410 47.500 82.730 47.560 ;
        RECT 78.285 47.360 82.730 47.500 ;
        RECT 85.720 47.500 85.860 47.655 ;
        RECT 87.470 47.640 87.790 47.700 ;
        RECT 91.150 47.640 91.470 47.700 ;
        RECT 91.625 47.655 91.915 47.885 ;
        RECT 95.290 47.840 95.610 47.900 ;
        RECT 98.065 47.840 98.355 47.885 ;
        RECT 95.290 47.700 98.355 47.840 ;
        RECT 90.230 47.500 90.550 47.560 ;
        RECT 85.720 47.360 90.550 47.500 ;
        RECT 91.700 47.500 91.840 47.655 ;
        RECT 95.290 47.640 95.610 47.700 ;
        RECT 98.065 47.655 98.355 47.700 ;
        RECT 107.265 47.840 107.555 47.885 ;
        RECT 109.105 47.840 109.395 47.885 ;
        RECT 107.265 47.700 109.395 47.840 ;
        RECT 107.265 47.655 107.555 47.700 ;
        RECT 109.105 47.655 109.395 47.700 ;
        RECT 110.930 47.840 111.250 47.900 ;
        RECT 111.865 47.840 112.155 47.885 ;
        RECT 110.930 47.700 112.155 47.840 ;
        RECT 110.930 47.640 111.250 47.700 ;
        RECT 111.865 47.655 112.155 47.700 ;
        RECT 114.150 47.840 114.470 47.900 ;
        RECT 115.545 47.840 115.835 47.885 ;
        RECT 114.150 47.700 115.835 47.840 ;
        RECT 114.150 47.640 114.470 47.700 ;
        RECT 115.545 47.655 115.835 47.700 ;
        RECT 92.070 47.500 92.390 47.560 ;
        RECT 91.700 47.360 92.390 47.500 ;
        RECT 78.285 47.315 78.575 47.360 ;
        RECT 63.180 47.020 64.240 47.160 ;
        RECT 50.210 46.960 50.530 47.020 ;
        RECT 64.100 46.880 64.240 47.020 ;
        RECT 44.690 46.820 45.010 46.880 ;
        RECT 43.400 46.680 45.010 46.820 ;
        RECT 44.690 46.620 45.010 46.680 ;
        RECT 51.605 46.820 51.895 46.865 ;
        RECT 53.430 46.820 53.750 46.880 ;
        RECT 51.605 46.680 53.750 46.820 ;
        RECT 51.605 46.635 51.895 46.680 ;
        RECT 53.430 46.620 53.750 46.680 ;
        RECT 64.010 46.620 64.330 46.880 ;
        RECT 75.050 46.820 75.370 46.880 ;
        RECT 75.525 46.820 75.815 46.865 ;
        RECT 75.050 46.680 75.815 46.820 ;
        RECT 77.440 46.820 77.580 47.315 ;
        RECT 82.410 47.300 82.730 47.360 ;
        RECT 90.230 47.300 90.550 47.360 ;
        RECT 92.070 47.300 92.390 47.360 ;
        RECT 92.545 47.315 92.835 47.545 ;
        RECT 80.585 47.160 80.875 47.205 ;
        RECT 82.870 47.160 83.190 47.220 ;
        RECT 80.585 47.020 83.190 47.160 ;
        RECT 80.585 46.975 80.875 47.020 ;
        RECT 82.870 46.960 83.190 47.020 ;
        RECT 83.345 47.160 83.635 47.205 ;
        RECT 86.550 47.160 86.870 47.220 ;
        RECT 92.620 47.160 92.760 47.315 ;
        RECT 83.345 47.020 86.870 47.160 ;
        RECT 83.345 46.975 83.635 47.020 ;
        RECT 86.550 46.960 86.870 47.020 ;
        RECT 92.160 47.020 92.760 47.160 ;
        RECT 92.160 46.820 92.300 47.020 ;
        RECT 77.440 46.680 92.300 46.820 ;
        RECT 105.410 46.820 105.730 46.880 ;
        RECT 112.785 46.820 113.075 46.865 ;
        RECT 105.410 46.680 113.075 46.820 ;
        RECT 75.050 46.620 75.370 46.680 ;
        RECT 75.525 46.635 75.815 46.680 ;
        RECT 105.410 46.620 105.730 46.680 ;
        RECT 112.785 46.635 113.075 46.680 ;
        RECT 5.520 46.000 125.580 46.480 ;
        RECT 13.870 45.800 14.190 45.860 ;
        RECT 18.945 45.800 19.235 45.845 ;
        RECT 13.870 45.660 19.235 45.800 ;
        RECT 13.870 45.600 14.190 45.660 ;
        RECT 18.945 45.615 19.235 45.660 ;
        RECT 33.650 45.800 33.970 45.860 ;
        RECT 34.585 45.800 34.875 45.845 ;
        RECT 33.650 45.660 34.875 45.800 ;
        RECT 33.650 45.600 33.970 45.660 ;
        RECT 34.585 45.615 34.875 45.660 ;
        RECT 39.170 45.800 39.490 45.860 ;
        RECT 40.105 45.800 40.395 45.845 ;
        RECT 39.170 45.660 40.395 45.800 ;
        RECT 10.155 45.460 10.445 45.505 ;
        RECT 12.045 45.460 12.335 45.505 ;
        RECT 15.165 45.460 15.455 45.505 ;
        RECT 10.155 45.320 15.455 45.460 ;
        RECT 10.155 45.275 10.445 45.320 ;
        RECT 12.045 45.275 12.335 45.320 ;
        RECT 15.165 45.275 15.455 45.320 ;
        RECT 18.025 45.460 18.315 45.505 ;
        RECT 20.310 45.460 20.630 45.520 ;
        RECT 18.025 45.320 20.630 45.460 ;
        RECT 18.025 45.275 18.315 45.320 ;
        RECT 20.310 45.260 20.630 45.320 ;
        RECT 26.715 45.460 27.005 45.505 ;
        RECT 28.605 45.460 28.895 45.505 ;
        RECT 31.725 45.460 32.015 45.505 ;
        RECT 26.715 45.320 32.015 45.460 ;
        RECT 26.715 45.275 27.005 45.320 ;
        RECT 28.605 45.275 28.895 45.320 ;
        RECT 31.725 45.275 32.015 45.320 ;
        RECT 7.430 45.120 7.750 45.180 ;
        RECT 9.285 45.120 9.575 45.165 ;
        RECT 22.165 45.120 22.455 45.165 ;
        RECT 23.070 45.120 23.390 45.180 ;
        RECT 29.510 45.120 29.830 45.180 ;
        RECT 7.430 44.980 18.700 45.120 ;
        RECT 7.430 44.920 7.750 44.980 ;
        RECT 9.285 44.935 9.575 44.980 ;
        RECT 9.750 44.780 10.040 44.825 ;
        RECT 11.585 44.780 11.875 44.825 ;
        RECT 15.165 44.780 15.455 44.825 ;
        RECT 9.750 44.640 15.455 44.780 ;
        RECT 9.750 44.595 10.040 44.640 ;
        RECT 11.585 44.595 11.875 44.640 ;
        RECT 15.165 44.595 15.455 44.640 ;
        RECT 10.665 44.440 10.955 44.485 ;
        RECT 12.030 44.440 12.350 44.500 ;
        RECT 16.245 44.485 16.535 44.800 ;
        RECT 18.560 44.500 18.700 44.980 ;
        RECT 22.165 44.980 23.390 45.120 ;
        RECT 22.165 44.935 22.455 44.980 ;
        RECT 23.070 44.920 23.390 44.980 ;
        RECT 24.540 44.980 29.830 45.120 ;
        RECT 34.660 45.120 34.800 45.615 ;
        RECT 39.170 45.600 39.490 45.660 ;
        RECT 40.105 45.615 40.395 45.660 ;
        RECT 45.625 45.800 45.915 45.845 ;
        RECT 48.370 45.800 48.690 45.860 ;
        RECT 45.625 45.660 48.690 45.800 ;
        RECT 45.625 45.615 45.915 45.660 ;
        RECT 48.370 45.600 48.690 45.660 ;
        RECT 82.410 45.600 82.730 45.860 ;
        RECT 86.565 45.800 86.855 45.845 ;
        RECT 87.930 45.800 88.250 45.860 ;
        RECT 86.565 45.660 88.250 45.800 ;
        RECT 86.565 45.615 86.855 45.660 ;
        RECT 87.930 45.600 88.250 45.660 ;
        RECT 111.850 45.600 112.170 45.860 ;
        RECT 74.555 45.460 74.845 45.505 ;
        RECT 76.445 45.460 76.735 45.505 ;
        RECT 79.565 45.460 79.855 45.505 ;
        RECT 74.555 45.320 79.855 45.460 ;
        RECT 82.500 45.460 82.640 45.600 ;
        RECT 107.265 45.460 107.555 45.505 ;
        RECT 82.500 45.320 89.080 45.460 ;
        RECT 74.555 45.275 74.845 45.320 ;
        RECT 76.445 45.275 76.735 45.320 ;
        RECT 79.565 45.275 79.855 45.320 ;
        RECT 35.965 45.120 36.255 45.165 ;
        RECT 34.660 44.980 36.255 45.120 ;
        RECT 24.540 44.825 24.680 44.980 ;
        RECT 29.510 44.920 29.830 44.980 ;
        RECT 35.965 44.935 36.255 44.980 ;
        RECT 36.410 45.120 36.730 45.180 ;
        RECT 39.185 45.120 39.475 45.165 ;
        RECT 36.410 44.980 39.475 45.120 ;
        RECT 36.410 44.920 36.730 44.980 ;
        RECT 39.185 44.935 39.475 44.980 ;
        RECT 47.910 45.120 48.230 45.180 ;
        RECT 48.385 45.120 48.675 45.165 ;
        RECT 52.525 45.120 52.815 45.165 ;
        RECT 47.910 44.980 52.815 45.120 ;
        RECT 47.910 44.920 48.230 44.980 ;
        RECT 48.385 44.935 48.675 44.980 ;
        RECT 52.525 44.935 52.815 44.980 ;
        RECT 53.430 45.120 53.750 45.180 ;
        RECT 56.665 45.120 56.955 45.165 ;
        RECT 53.430 44.980 56.955 45.120 ;
        RECT 53.430 44.920 53.750 44.980 ;
        RECT 56.665 44.935 56.955 44.980 ;
        RECT 75.050 44.920 75.370 45.180 ;
        RECT 77.810 45.120 78.130 45.180 ;
        RECT 82.885 45.120 83.175 45.165 ;
        RECT 77.810 44.980 83.175 45.120 ;
        RECT 77.810 44.920 78.130 44.980 ;
        RECT 82.885 44.935 83.175 44.980 ;
        RECT 84.710 45.120 85.030 45.180 ;
        RECT 84.710 44.980 88.160 45.120 ;
        RECT 84.710 44.920 85.030 44.980 ;
        RECT 24.465 44.595 24.755 44.825 ;
        RECT 25.845 44.595 26.135 44.825 ;
        RECT 26.310 44.780 26.600 44.825 ;
        RECT 28.145 44.780 28.435 44.825 ;
        RECT 31.725 44.780 32.015 44.825 ;
        RECT 26.310 44.640 32.015 44.780 ;
        RECT 26.310 44.595 26.600 44.640 ;
        RECT 28.145 44.595 28.435 44.640 ;
        RECT 31.725 44.595 32.015 44.640 ;
        RECT 10.665 44.300 12.350 44.440 ;
        RECT 10.665 44.255 10.955 44.300 ;
        RECT 12.030 44.240 12.350 44.300 ;
        RECT 12.945 44.440 13.595 44.485 ;
        RECT 16.245 44.440 16.835 44.485 ;
        RECT 17.090 44.440 17.410 44.500 ;
        RECT 12.945 44.300 17.410 44.440 ;
        RECT 12.945 44.255 13.595 44.300 ;
        RECT 16.545 44.255 16.835 44.300 ;
        RECT 17.090 44.240 17.410 44.300 ;
        RECT 18.470 44.440 18.790 44.500 ;
        RECT 25.920 44.440 26.060 44.595 ;
        RECT 18.470 44.300 26.060 44.440 ;
        RECT 18.470 44.240 18.790 44.300 ;
        RECT 27.225 44.255 27.515 44.485 ;
        RECT 29.505 44.440 30.155 44.485 ;
        RECT 32.270 44.440 32.590 44.500 ;
        RECT 32.805 44.485 33.095 44.800 ;
        RECT 38.250 44.780 38.570 44.840 ;
        RECT 40.565 44.780 40.855 44.825 ;
        RECT 38.250 44.640 40.855 44.780 ;
        RECT 38.250 44.580 38.570 44.640 ;
        RECT 40.565 44.595 40.855 44.640 ;
        RECT 47.450 44.580 47.770 44.840 ;
        RECT 72.750 44.780 73.070 44.840 ;
        RECT 88.020 44.825 88.160 44.980 ;
        RECT 88.940 44.840 89.080 45.320 ;
        RECT 107.265 45.320 110.700 45.460 ;
        RECT 107.265 45.275 107.555 45.320 ;
        RECT 103.570 45.120 103.890 45.180 ;
        RECT 110.560 45.165 110.700 45.320 ;
        RECT 104.045 45.120 104.335 45.165 ;
        RECT 103.570 44.980 104.335 45.120 ;
        RECT 103.570 44.920 103.890 44.980 ;
        RECT 104.045 44.935 104.335 44.980 ;
        RECT 110.485 44.935 110.775 45.165 ;
        RECT 73.685 44.780 73.975 44.825 ;
        RECT 72.750 44.640 73.975 44.780 ;
        RECT 72.750 44.580 73.070 44.640 ;
        RECT 73.685 44.595 73.975 44.640 ;
        RECT 74.150 44.780 74.440 44.825 ;
        RECT 75.985 44.780 76.275 44.825 ;
        RECT 79.565 44.780 79.855 44.825 ;
        RECT 74.150 44.640 79.855 44.780 ;
        RECT 74.150 44.595 74.440 44.640 ;
        RECT 75.985 44.595 76.275 44.640 ;
        RECT 79.565 44.595 79.855 44.640 ;
        RECT 32.805 44.440 33.395 44.485 ;
        RECT 29.505 44.300 33.395 44.440 ;
        RECT 29.505 44.255 30.155 44.300 ;
        RECT 20.770 43.900 21.090 44.160 ;
        RECT 21.230 43.900 21.550 44.160 ;
        RECT 25.385 44.100 25.675 44.145 ;
        RECT 27.300 44.100 27.440 44.255 ;
        RECT 32.270 44.240 32.590 44.300 ;
        RECT 33.105 44.255 33.395 44.300 ;
        RECT 47.925 44.440 48.215 44.485 ;
        RECT 51.605 44.440 51.895 44.485 ;
        RECT 53.905 44.440 54.195 44.485 ;
        RECT 47.925 44.300 54.195 44.440 ;
        RECT 47.925 44.255 48.215 44.300 ;
        RECT 51.605 44.255 51.895 44.300 ;
        RECT 53.905 44.255 54.195 44.300 ;
        RECT 77.345 44.440 77.995 44.485 ;
        RECT 78.730 44.440 79.050 44.500 ;
        RECT 80.645 44.485 80.935 44.800 ;
        RECT 85.645 44.595 85.935 44.825 ;
        RECT 87.945 44.595 88.235 44.825 ;
        RECT 80.645 44.440 81.235 44.485 ;
        RECT 77.345 44.300 81.235 44.440 ;
        RECT 77.345 44.255 77.995 44.300 ;
        RECT 78.730 44.240 79.050 44.300 ;
        RECT 80.945 44.255 81.235 44.300 ;
        RECT 25.385 43.960 27.440 44.100 ;
        RECT 43.770 44.100 44.090 44.160 ;
        RECT 49.765 44.100 50.055 44.145 ;
        RECT 43.770 43.960 50.055 44.100 ;
        RECT 25.385 43.915 25.675 43.960 ;
        RECT 43.770 43.900 44.090 43.960 ;
        RECT 49.765 43.915 50.055 43.960 ;
        RECT 51.130 44.100 51.450 44.160 ;
        RECT 52.065 44.100 52.355 44.145 ;
        RECT 52.970 44.100 53.290 44.160 ;
        RECT 51.130 43.960 53.290 44.100 ;
        RECT 51.130 43.900 51.450 43.960 ;
        RECT 52.065 43.915 52.355 43.960 ;
        RECT 52.970 43.900 53.290 43.960 ;
        RECT 79.650 44.100 79.970 44.160 ;
        RECT 85.720 44.100 85.860 44.595 ;
        RECT 88.390 44.580 88.710 44.840 ;
        RECT 88.850 44.580 89.170 44.840 ;
        RECT 89.785 44.780 90.075 44.825 ;
        RECT 91.150 44.780 91.470 44.840 ;
        RECT 89.785 44.640 91.470 44.780 ;
        RECT 89.785 44.595 90.075 44.640 ;
        RECT 91.150 44.580 91.470 44.640 ;
        RECT 93.005 44.595 93.295 44.825 ;
        RECT 102.190 44.780 102.510 44.840 ;
        RECT 104.965 44.780 105.255 44.825 ;
        RECT 102.190 44.640 105.255 44.780 ;
        RECT 87.010 44.440 87.330 44.500 ;
        RECT 92.070 44.440 92.390 44.500 ;
        RECT 93.080 44.440 93.220 44.595 ;
        RECT 102.190 44.580 102.510 44.640 ;
        RECT 104.965 44.595 105.255 44.640 ;
        RECT 87.010 44.300 93.220 44.440 ;
        RECT 105.040 44.440 105.180 44.595 ;
        RECT 105.410 44.580 105.730 44.840 ;
        RECT 111.390 44.580 111.710 44.840 ;
        RECT 111.850 44.440 112.170 44.500 ;
        RECT 105.040 44.300 112.170 44.440 ;
        RECT 87.010 44.240 87.330 44.300 ;
        RECT 92.070 44.240 92.390 44.300 ;
        RECT 111.850 44.240 112.170 44.300 ;
        RECT 79.650 43.960 85.860 44.100 ;
        RECT 89.770 44.100 90.090 44.160 ;
        RECT 90.245 44.100 90.535 44.145 ;
        RECT 89.770 43.960 90.535 44.100 ;
        RECT 79.650 43.900 79.970 43.960 ;
        RECT 89.770 43.900 90.090 43.960 ;
        RECT 90.245 43.915 90.535 43.960 ;
        RECT 105.870 44.100 106.190 44.160 ;
        RECT 107.725 44.100 108.015 44.145 ;
        RECT 105.870 43.960 108.015 44.100 ;
        RECT 105.870 43.900 106.190 43.960 ;
        RECT 107.725 43.915 108.015 43.960 ;
        RECT 5.520 43.280 125.580 43.760 ;
        RECT 17.565 43.080 17.855 43.125 ;
        RECT 18.010 43.080 18.330 43.140 ;
        RECT 17.565 42.940 18.330 43.080 ;
        RECT 17.565 42.895 17.855 42.940 ;
        RECT 18.010 42.880 18.330 42.940 ;
        RECT 20.770 43.080 21.090 43.140 ;
        RECT 24.465 43.080 24.755 43.125 ;
        RECT 20.770 42.940 24.755 43.080 ;
        RECT 20.770 42.880 21.090 42.940 ;
        RECT 24.465 42.895 24.755 42.940 ;
        RECT 32.270 42.880 32.590 43.140 ;
        RECT 34.110 43.080 34.430 43.140 ;
        RECT 35.045 43.080 35.335 43.125 ;
        RECT 34.110 42.940 35.335 43.080 ;
        RECT 34.110 42.880 34.430 42.940 ;
        RECT 35.045 42.895 35.335 42.940 ;
        RECT 65.850 42.880 66.170 43.140 ;
        RECT 78.730 42.880 79.050 43.140 ;
        RECT 85.645 43.080 85.935 43.125 ;
        RECT 87.010 43.080 87.330 43.140 ;
        RECT 85.645 42.940 87.330 43.080 ;
        RECT 85.645 42.895 85.935 42.940 ;
        RECT 87.010 42.880 87.330 42.940 ;
        RECT 98.065 43.080 98.355 43.125 ;
        RECT 103.125 43.080 103.415 43.125 ;
        RECT 104.950 43.080 105.270 43.140 ;
        RECT 98.065 42.940 105.270 43.080 ;
        RECT 98.065 42.895 98.355 42.940 ;
        RECT 103.125 42.895 103.415 42.940 ;
        RECT 104.950 42.880 105.270 42.940 ;
        RECT 17.090 42.740 17.410 42.800 ;
        RECT 18.945 42.740 19.235 42.785 ;
        RECT 17.090 42.600 19.235 42.740 ;
        RECT 17.090 42.540 17.410 42.600 ;
        RECT 18.945 42.555 19.235 42.600 ;
        RECT 21.230 42.740 21.550 42.800 ;
        RECT 24.005 42.740 24.295 42.785 ;
        RECT 38.250 42.740 38.570 42.800 ;
        RECT 39.170 42.740 39.490 42.800 ;
        RECT 62.185 42.740 62.475 42.785 ;
        RECT 65.390 42.740 65.710 42.800 ;
        RECT 96.210 42.740 96.530 42.800 ;
        RECT 21.230 42.600 24.295 42.740 ;
        RECT 21.230 42.540 21.550 42.600 ;
        RECT 24.005 42.555 24.295 42.600 ;
        RECT 32.820 42.600 44.460 42.740 ;
        RECT 18.010 42.400 18.330 42.460 ;
        RECT 19.405 42.400 19.695 42.445 ;
        RECT 18.010 42.260 19.695 42.400 ;
        RECT 18.010 42.200 18.330 42.260 ;
        RECT 19.405 42.215 19.695 42.260 ;
        RECT 20.310 42.400 20.630 42.460 ;
        RECT 32.820 42.445 32.960 42.600 ;
        RECT 38.250 42.540 38.570 42.600 ;
        RECT 39.170 42.540 39.490 42.600 ;
        RECT 20.785 42.400 21.075 42.445 ;
        RECT 20.310 42.260 21.075 42.400 ;
        RECT 20.310 42.200 20.630 42.260 ;
        RECT 20.785 42.215 21.075 42.260 ;
        RECT 32.745 42.215 33.035 42.445 ;
        RECT 35.965 42.400 36.255 42.445 ;
        RECT 38.710 42.400 39.030 42.460 ;
        RECT 35.965 42.260 39.030 42.400 ;
        RECT 35.965 42.215 36.255 42.260 ;
        RECT 38.710 42.200 39.030 42.260 ;
        RECT 43.770 42.200 44.090 42.460 ;
        RECT 44.320 42.400 44.460 42.600 ;
        RECT 62.185 42.600 65.710 42.740 ;
        RECT 62.185 42.555 62.475 42.600 ;
        RECT 65.390 42.540 65.710 42.600 ;
        RECT 80.660 42.600 96.530 42.740 ;
        RECT 80.660 42.460 80.800 42.600 ;
        RECT 46.085 42.400 46.375 42.445 ;
        RECT 50.210 42.400 50.530 42.460 ;
        RECT 44.320 42.260 50.530 42.400 ;
        RECT 46.085 42.215 46.375 42.260 ;
        RECT 50.210 42.200 50.530 42.260 ;
        RECT 67.245 42.400 67.535 42.445 ;
        RECT 67.690 42.400 68.010 42.460 ;
        RECT 67.245 42.260 68.010 42.400 ;
        RECT 67.245 42.215 67.535 42.260 ;
        RECT 67.690 42.200 68.010 42.260 ;
        RECT 77.350 42.400 77.670 42.460 ;
        RECT 78.285 42.400 78.575 42.445 ;
        RECT 80.570 42.400 80.890 42.460 ;
        RECT 77.350 42.260 80.890 42.400 ;
        RECT 77.350 42.200 77.670 42.260 ;
        RECT 78.285 42.215 78.575 42.260 ;
        RECT 80.570 42.200 80.890 42.260 ;
        RECT 85.185 42.400 85.475 42.445 ;
        RECT 87.485 42.400 87.775 42.445 ;
        RECT 85.185 42.260 87.775 42.400 ;
        RECT 85.185 42.215 85.475 42.260 ;
        RECT 87.485 42.215 87.775 42.260 ;
        RECT 88.850 42.400 89.170 42.460 ;
        RECT 91.240 42.445 91.380 42.600 ;
        RECT 96.210 42.540 96.530 42.600 ;
        RECT 102.665 42.740 102.955 42.785 ;
        RECT 109.105 42.740 109.395 42.785 ;
        RECT 102.665 42.600 109.395 42.740 ;
        RECT 102.665 42.555 102.955 42.600 ;
        RECT 109.105 42.555 109.395 42.600 ;
        RECT 111.390 42.740 111.710 42.800 ;
        RECT 111.390 42.600 113.000 42.740 ;
        RECT 111.390 42.540 111.710 42.600 ;
        RECT 90.245 42.400 90.535 42.445 ;
        RECT 88.850 42.260 90.535 42.400 ;
        RECT 88.850 42.200 89.170 42.260 ;
        RECT 90.245 42.215 90.535 42.260 ;
        RECT 91.165 42.215 91.455 42.445 ;
        RECT 92.990 42.400 93.310 42.460 ;
        RECT 95.305 42.400 95.595 42.445 ;
        RECT 104.965 42.400 105.255 42.445 ;
        RECT 105.870 42.400 106.190 42.460 ;
        RECT 92.990 42.260 95.595 42.400 ;
        RECT 92.990 42.200 93.310 42.260 ;
        RECT 95.305 42.215 95.595 42.260 ;
        RECT 98.140 42.260 99.200 42.400 ;
        RECT 23.990 42.060 24.310 42.120 ;
        RECT 27.685 42.060 27.975 42.105 ;
        RECT 47.910 42.060 48.230 42.120 ;
        RECT 23.990 41.920 27.975 42.060 ;
        RECT 23.990 41.860 24.310 41.920 ;
        RECT 27.685 41.875 27.975 41.920 ;
        RECT 33.280 41.920 48.230 42.060 ;
        RECT 26.750 41.720 27.070 41.780 ;
        RECT 32.730 41.720 33.050 41.780 ;
        RECT 33.280 41.720 33.420 41.920 ;
        RECT 47.910 41.860 48.230 41.920 ;
        RECT 64.470 41.860 64.790 42.120 ;
        RECT 64.930 41.860 65.250 42.120 ;
        RECT 75.970 42.060 76.290 42.120 ;
        RECT 86.105 42.060 86.395 42.105 ;
        RECT 86.550 42.060 86.870 42.120 ;
        RECT 98.140 42.060 98.280 42.260 ;
        RECT 75.970 41.920 98.280 42.060 ;
        RECT 75.970 41.860 76.290 41.920 ;
        RECT 86.105 41.875 86.395 41.920 ;
        RECT 86.550 41.860 86.870 41.920 ;
        RECT 98.510 41.860 98.830 42.120 ;
        RECT 99.060 42.105 99.200 42.260 ;
        RECT 104.965 42.260 106.190 42.400 ;
        RECT 104.965 42.215 105.255 42.260 ;
        RECT 105.870 42.200 106.190 42.260 ;
        RECT 111.850 42.200 112.170 42.460 ;
        RECT 112.860 42.445 113.000 42.600 ;
        RECT 112.785 42.215 113.075 42.445 ;
        RECT 98.985 42.060 99.275 42.105 ;
        RECT 103.570 42.060 103.890 42.120 ;
        RECT 98.985 41.920 103.890 42.060 ;
        RECT 98.985 41.875 99.275 41.920 ;
        RECT 103.570 41.860 103.890 41.920 ;
        RECT 26.750 41.580 33.420 41.720 ;
        RECT 46.545 41.720 46.835 41.765 ;
        RECT 48.370 41.720 48.690 41.780 ;
        RECT 46.545 41.580 48.690 41.720 ;
        RECT 26.750 41.520 27.070 41.580 ;
        RECT 32.730 41.520 33.050 41.580 ;
        RECT 46.545 41.535 46.835 41.580 ;
        RECT 48.370 41.520 48.690 41.580 ;
        RECT 62.170 41.520 62.490 41.780 ;
        RECT 91.610 41.520 91.930 41.780 ;
        RECT 92.530 41.520 92.850 41.780 ;
        RECT 93.910 41.720 94.230 41.780 ;
        RECT 96.225 41.720 96.515 41.765 ;
        RECT 93.910 41.580 96.515 41.720 ;
        RECT 93.910 41.520 94.230 41.580 ;
        RECT 96.225 41.535 96.515 41.580 ;
        RECT 97.130 41.720 97.450 41.780 ;
        RECT 100.825 41.720 101.115 41.765 ;
        RECT 97.130 41.580 101.115 41.720 ;
        RECT 97.130 41.520 97.450 41.580 ;
        RECT 100.825 41.535 101.115 41.580 ;
        RECT 105.885 41.720 106.175 41.765 ;
        RECT 109.550 41.720 109.870 41.780 ;
        RECT 105.885 41.580 109.870 41.720 ;
        RECT 105.885 41.535 106.175 41.580 ;
        RECT 109.550 41.520 109.870 41.580 ;
        RECT 113.230 41.520 113.550 41.780 ;
        RECT 44.705 41.380 44.995 41.425 ;
        RECT 46.070 41.380 46.390 41.440 ;
        RECT 44.705 41.240 46.390 41.380 ;
        RECT 44.705 41.195 44.995 41.240 ;
        RECT 46.070 41.180 46.390 41.240 ;
        RECT 66.310 41.380 66.630 41.440 ;
        RECT 66.785 41.380 67.075 41.425 ;
        RECT 66.310 41.240 67.075 41.380 ;
        RECT 66.310 41.180 66.630 41.240 ;
        RECT 66.785 41.195 67.075 41.240 ;
        RECT 83.345 41.380 83.635 41.425 ;
        RECT 85.170 41.380 85.490 41.440 ;
        RECT 83.345 41.240 85.490 41.380 ;
        RECT 83.345 41.195 83.635 41.240 ;
        RECT 85.170 41.180 85.490 41.240 ;
        RECT 5.520 40.560 125.580 41.040 ;
        RECT 51.130 40.360 51.450 40.420 ;
        RECT 53.675 40.360 53.965 40.405 ;
        RECT 51.130 40.220 53.965 40.360 ;
        RECT 51.130 40.160 51.450 40.220 ;
        RECT 53.675 40.175 53.965 40.220 ;
        RECT 64.930 40.360 65.250 40.420 ;
        RECT 66.785 40.360 67.075 40.405 ;
        RECT 67.230 40.360 67.550 40.420 ;
        RECT 64.930 40.220 67.550 40.360 ;
        RECT 64.930 40.160 65.250 40.220 ;
        RECT 66.785 40.175 67.075 40.220 ;
        RECT 67.230 40.160 67.550 40.220 ;
        RECT 79.650 40.160 79.970 40.420 ;
        RECT 104.950 40.360 105.270 40.420 ;
        RECT 107.495 40.360 107.785 40.405 ;
        RECT 104.950 40.220 107.785 40.360 ;
        RECT 104.950 40.160 105.270 40.220 ;
        RECT 107.495 40.175 107.785 40.220 ;
        RECT 111.850 40.360 112.170 40.420 ;
        RECT 116.925 40.360 117.215 40.405 ;
        RECT 111.850 40.220 117.215 40.360 ;
        RECT 111.850 40.160 112.170 40.220 ;
        RECT 116.925 40.175 117.215 40.220 ;
        RECT 45.170 40.020 45.460 40.065 ;
        RECT 47.030 40.020 47.320 40.065 ;
        RECT 49.810 40.020 50.100 40.065 ;
        RECT 45.170 39.880 50.100 40.020 ;
        RECT 45.170 39.835 45.460 39.880 ;
        RECT 47.030 39.835 47.320 39.880 ;
        RECT 49.810 39.835 50.100 39.880 ;
        RECT 58.915 40.020 59.205 40.065 ;
        RECT 60.805 40.020 61.095 40.065 ;
        RECT 63.925 40.020 64.215 40.065 ;
        RECT 58.915 39.880 64.215 40.020 ;
        RECT 58.915 39.835 59.205 39.880 ;
        RECT 60.805 39.835 61.095 39.880 ;
        RECT 63.925 39.835 64.215 39.880 ;
        RECT 71.795 40.020 72.085 40.065 ;
        RECT 73.685 40.020 73.975 40.065 ;
        RECT 76.805 40.020 77.095 40.065 ;
        RECT 71.795 39.880 77.095 40.020 ;
        RECT 71.795 39.835 72.085 39.880 ;
        RECT 73.685 39.835 73.975 39.880 ;
        RECT 76.805 39.835 77.095 39.880 ;
        RECT 98.990 40.020 99.280 40.065 ;
        RECT 100.850 40.020 101.140 40.065 ;
        RECT 103.630 40.020 103.920 40.065 ;
        RECT 98.990 39.880 103.920 40.020 ;
        RECT 98.990 39.835 99.280 39.880 ;
        RECT 100.850 39.835 101.140 39.880 ;
        RECT 103.630 39.835 103.920 39.880 ;
        RECT 109.055 40.020 109.345 40.065 ;
        RECT 110.945 40.020 111.235 40.065 ;
        RECT 114.065 40.020 114.355 40.065 ;
        RECT 109.055 39.880 114.355 40.020 ;
        RECT 109.055 39.835 109.345 39.880 ;
        RECT 110.945 39.835 111.235 39.880 ;
        RECT 114.065 39.835 114.355 39.880 ;
        RECT 27.670 39.680 27.990 39.740 ;
        RECT 30.905 39.680 31.195 39.725 ;
        RECT 27.670 39.540 31.195 39.680 ;
        RECT 27.670 39.480 27.990 39.540 ;
        RECT 30.905 39.495 31.195 39.540 ;
        RECT 44.690 39.680 45.010 39.740 ;
        RECT 52.050 39.680 52.370 39.740 ;
        RECT 58.045 39.680 58.335 39.725 ;
        RECT 44.690 39.540 58.335 39.680 ;
        RECT 44.690 39.480 45.010 39.540 ;
        RECT 52.050 39.480 52.370 39.540 ;
        RECT 58.045 39.495 58.335 39.540 ;
        RECT 70.925 39.680 71.215 39.725 ;
        RECT 72.750 39.680 73.070 39.740 ;
        RECT 83.330 39.680 83.650 39.740 ;
        RECT 70.925 39.540 83.650 39.680 ;
        RECT 70.925 39.495 71.215 39.540 ;
        RECT 72.750 39.480 73.070 39.540 ;
        RECT 83.330 39.480 83.650 39.540 ;
        RECT 85.170 39.480 85.490 39.740 ;
        RECT 86.550 39.480 86.870 39.740 ;
        RECT 87.485 39.680 87.775 39.725 ;
        RECT 92.530 39.680 92.850 39.740 ;
        RECT 87.485 39.540 92.850 39.680 ;
        RECT 87.485 39.495 87.775 39.540 ;
        RECT 92.530 39.480 92.850 39.540 ;
        RECT 98.525 39.680 98.815 39.725 ;
        RECT 104.030 39.680 104.350 39.740 ;
        RECT 107.710 39.680 108.030 39.740 ;
        RECT 108.185 39.680 108.475 39.725 ;
        RECT 98.525 39.540 108.475 39.680 ;
        RECT 98.525 39.495 98.815 39.540 ;
        RECT 104.030 39.480 104.350 39.540 ;
        RECT 107.710 39.480 108.030 39.540 ;
        RECT 108.185 39.495 108.475 39.540 ;
        RECT 109.550 39.480 109.870 39.740 ;
        RECT 40.550 39.140 40.870 39.400 ;
        RECT 46.070 39.340 46.390 39.400 ;
        RECT 46.545 39.340 46.835 39.385 ;
        RECT 49.810 39.340 50.100 39.385 ;
        RECT 46.070 39.200 46.835 39.340 ;
        RECT 46.070 39.140 46.390 39.200 ;
        RECT 46.545 39.155 46.835 39.200 ;
        RECT 47.565 39.200 50.100 39.340 ;
        RECT 47.565 39.045 47.780 39.200 ;
        RECT 49.810 39.155 50.100 39.200 ;
        RECT 58.510 39.340 58.800 39.385 ;
        RECT 60.345 39.340 60.635 39.385 ;
        RECT 63.925 39.340 64.215 39.385 ;
        RECT 58.510 39.200 64.215 39.340 ;
        RECT 58.510 39.155 58.800 39.200 ;
        RECT 60.345 39.155 60.635 39.200 ;
        RECT 63.925 39.155 64.215 39.200 ;
        RECT 45.630 39.000 45.920 39.045 ;
        RECT 47.490 39.000 47.780 39.045 ;
        RECT 45.630 38.860 47.780 39.000 ;
        RECT 45.630 38.815 45.920 38.860 ;
        RECT 47.490 38.815 47.780 38.860 ;
        RECT 48.370 39.045 48.690 39.060 ;
        RECT 48.370 39.000 48.700 39.045 ;
        RECT 51.670 39.000 51.960 39.045 ;
        RECT 48.370 38.860 51.960 39.000 ;
        RECT 48.370 38.815 48.700 38.860 ;
        RECT 51.670 38.815 51.960 38.860 ;
        RECT 59.425 39.000 59.715 39.045 ;
        RECT 59.870 39.000 60.190 39.060 ;
        RECT 65.005 39.045 65.295 39.360 ;
        RECT 68.625 39.340 68.915 39.385 ;
        RECT 70.450 39.340 70.770 39.400 ;
        RECT 68.625 39.200 70.770 39.340 ;
        RECT 68.625 39.155 68.915 39.200 ;
        RECT 70.450 39.140 70.770 39.200 ;
        RECT 71.390 39.340 71.680 39.385 ;
        RECT 73.225 39.340 73.515 39.385 ;
        RECT 76.805 39.340 77.095 39.385 ;
        RECT 71.390 39.200 77.095 39.340 ;
        RECT 71.390 39.155 71.680 39.200 ;
        RECT 73.225 39.155 73.515 39.200 ;
        RECT 76.805 39.155 77.095 39.200 ;
        RECT 59.425 38.860 60.190 39.000 ;
        RECT 59.425 38.815 59.715 38.860 ;
        RECT 48.370 38.800 48.690 38.815 ;
        RECT 59.870 38.800 60.190 38.860 ;
        RECT 61.705 39.000 62.355 39.045 ;
        RECT 65.005 39.000 65.595 39.045 ;
        RECT 66.310 39.000 66.630 39.060 ;
        RECT 61.705 38.860 66.630 39.000 ;
        RECT 61.705 38.815 62.355 38.860 ;
        RECT 65.305 38.815 65.595 38.860 ;
        RECT 66.310 38.800 66.630 38.860 ;
        RECT 72.305 39.000 72.595 39.045 ;
        RECT 73.670 39.000 73.990 39.060 ;
        RECT 77.885 39.045 78.175 39.360 ;
        RECT 81.045 39.340 81.335 39.385 ;
        RECT 82.425 39.340 82.715 39.385 ;
        RECT 81.045 39.200 82.715 39.340 ;
        RECT 81.045 39.155 81.335 39.200 ;
        RECT 82.425 39.155 82.715 39.200 ;
        RECT 87.945 39.340 88.235 39.385 ;
        RECT 89.770 39.340 90.090 39.400 ;
        RECT 87.945 39.200 90.090 39.340 ;
        RECT 87.945 39.155 88.235 39.200 ;
        RECT 89.770 39.140 90.090 39.200 ;
        RECT 90.230 39.140 90.550 39.400 ;
        RECT 94.845 39.155 95.135 39.385 ;
        RECT 72.305 38.860 73.990 39.000 ;
        RECT 72.305 38.815 72.595 38.860 ;
        RECT 73.670 38.800 73.990 38.860 ;
        RECT 74.585 39.000 75.235 39.045 ;
        RECT 77.885 39.000 78.475 39.045 ;
        RECT 80.110 39.000 80.430 39.060 ;
        RECT 94.920 39.000 95.060 39.155 ;
        RECT 96.210 39.140 96.530 39.400 ;
        RECT 98.050 39.340 98.370 39.400 ;
        RECT 100.365 39.340 100.655 39.385 ;
        RECT 103.630 39.340 103.920 39.385 ;
        RECT 98.050 39.200 100.655 39.340 ;
        RECT 98.050 39.140 98.370 39.200 ;
        RECT 100.365 39.155 100.655 39.200 ;
        RECT 101.385 39.200 103.920 39.340 ;
        RECT 101.385 39.045 101.600 39.200 ;
        RECT 103.630 39.155 103.920 39.200 ;
        RECT 108.650 39.340 108.940 39.385 ;
        RECT 110.485 39.340 110.775 39.385 ;
        RECT 114.065 39.340 114.355 39.385 ;
        RECT 108.650 39.200 114.355 39.340 ;
        RECT 108.650 39.155 108.940 39.200 ;
        RECT 110.485 39.155 110.775 39.200 ;
        RECT 114.065 39.155 114.355 39.200 ;
        RECT 74.585 38.860 80.430 39.000 ;
        RECT 74.585 38.815 75.235 38.860 ;
        RECT 78.185 38.815 78.475 38.860 ;
        RECT 80.110 38.800 80.430 38.860 ;
        RECT 89.860 38.860 95.060 39.000 ;
        RECT 99.450 39.000 99.740 39.045 ;
        RECT 101.310 39.000 101.600 39.045 ;
        RECT 99.450 38.860 101.600 39.000 ;
        RECT 33.190 38.660 33.510 38.720 ;
        RECT 34.125 38.660 34.415 38.705 ;
        RECT 33.190 38.520 34.415 38.660 ;
        RECT 33.190 38.460 33.510 38.520 ;
        RECT 34.125 38.475 34.415 38.520 ;
        RECT 38.250 38.660 38.570 38.720 ;
        RECT 39.645 38.660 39.935 38.705 ;
        RECT 38.250 38.520 39.935 38.660 ;
        RECT 38.250 38.460 38.570 38.520 ;
        RECT 39.645 38.475 39.935 38.520 ;
        RECT 60.330 38.660 60.650 38.720 ;
        RECT 62.630 38.660 62.950 38.720 ;
        RECT 67.705 38.660 67.995 38.705 ;
        RECT 60.330 38.520 67.995 38.660 ;
        RECT 60.330 38.460 60.650 38.520 ;
        RECT 62.630 38.460 62.950 38.520 ;
        RECT 67.705 38.475 67.995 38.520 ;
        RECT 81.950 38.460 82.270 38.720 ;
        RECT 89.860 38.705 90.000 38.860 ;
        RECT 99.450 38.815 99.740 38.860 ;
        RECT 101.310 38.815 101.600 38.860 ;
        RECT 102.230 39.000 102.520 39.045 ;
        RECT 104.490 39.000 104.810 39.060 ;
        RECT 105.490 39.000 105.780 39.045 ;
        RECT 102.230 38.860 105.780 39.000 ;
        RECT 102.230 38.815 102.520 38.860 ;
        RECT 104.490 38.800 104.810 38.860 ;
        RECT 105.490 38.815 105.780 38.860 ;
        RECT 111.845 39.000 112.495 39.045 ;
        RECT 113.230 39.000 113.550 39.060 ;
        RECT 115.145 39.045 115.435 39.360 ;
        RECT 115.145 39.000 115.735 39.045 ;
        RECT 111.845 38.860 115.735 39.000 ;
        RECT 111.845 38.815 112.495 38.860 ;
        RECT 113.230 38.800 113.550 38.860 ;
        RECT 115.445 38.815 115.735 38.860 ;
        RECT 89.785 38.475 90.075 38.705 ;
        RECT 93.450 38.460 93.770 38.720 ;
        RECT 93.925 38.660 94.215 38.705 ;
        RECT 94.370 38.660 94.690 38.720 ;
        RECT 93.925 38.520 94.690 38.660 ;
        RECT 93.925 38.475 94.215 38.520 ;
        RECT 94.370 38.460 94.690 38.520 ;
        RECT 96.685 38.660 96.975 38.705 ;
        RECT 97.590 38.660 97.910 38.720 ;
        RECT 96.685 38.520 97.910 38.660 ;
        RECT 96.685 38.475 96.975 38.520 ;
        RECT 97.590 38.460 97.910 38.520 ;
        RECT 5.520 37.840 125.580 38.320 ;
        RECT 23.085 37.640 23.375 37.685 ;
        RECT 23.990 37.640 24.310 37.700 ;
        RECT 23.085 37.500 24.310 37.640 ;
        RECT 23.085 37.455 23.375 37.500 ;
        RECT 23.990 37.440 24.310 37.500 ;
        RECT 25.385 37.640 25.675 37.685 ;
        RECT 33.190 37.640 33.510 37.700 ;
        RECT 25.385 37.500 33.510 37.640 ;
        RECT 25.385 37.455 25.675 37.500 ;
        RECT 33.190 37.440 33.510 37.500 ;
        RECT 40.550 37.640 40.870 37.700 ;
        RECT 46.085 37.640 46.375 37.685 ;
        RECT 40.550 37.500 46.375 37.640 ;
        RECT 40.550 37.440 40.870 37.500 ;
        RECT 46.085 37.455 46.375 37.500 ;
        RECT 47.925 37.640 48.215 37.685 ;
        RECT 51.130 37.640 51.450 37.700 ;
        RECT 47.925 37.500 51.450 37.640 ;
        RECT 47.925 37.455 48.215 37.500 ;
        RECT 51.130 37.440 51.450 37.500 ;
        RECT 58.490 37.440 58.810 37.700 ;
        RECT 59.870 37.440 60.190 37.700 ;
        RECT 63.550 37.640 63.870 37.700 ;
        RECT 64.485 37.640 64.775 37.685 ;
        RECT 62.030 37.500 62.860 37.640 ;
        RECT 18.005 37.300 18.655 37.345 ;
        RECT 20.770 37.300 21.090 37.360 ;
        RECT 21.605 37.300 21.895 37.345 ;
        RECT 18.005 37.160 21.895 37.300 ;
        RECT 18.005 37.115 18.655 37.160 ;
        RECT 20.770 37.100 21.090 37.160 ;
        RECT 21.305 37.115 21.895 37.160 ;
        RECT 37.350 37.300 37.640 37.345 ;
        RECT 39.210 37.300 39.500 37.345 ;
        RECT 37.350 37.160 39.500 37.300 ;
        RECT 37.350 37.115 37.640 37.160 ;
        RECT 39.210 37.115 39.500 37.160 ;
        RECT 40.130 37.300 40.420 37.345 ;
        RECT 41.930 37.300 42.250 37.360 ;
        RECT 43.390 37.300 43.680 37.345 ;
        RECT 48.385 37.300 48.675 37.345 ;
        RECT 58.580 37.300 58.720 37.440 ;
        RECT 62.030 37.300 62.170 37.500 ;
        RECT 40.130 37.160 43.680 37.300 ;
        RECT 40.130 37.115 40.420 37.160 ;
        RECT 14.810 36.960 15.100 37.005 ;
        RECT 16.645 36.960 16.935 37.005 ;
        RECT 20.225 36.960 20.515 37.005 ;
        RECT 14.810 36.820 20.515 36.960 ;
        RECT 14.810 36.775 15.100 36.820 ;
        RECT 16.645 36.775 16.935 36.820 ;
        RECT 20.225 36.775 20.515 36.820 ;
        RECT 21.305 36.800 21.595 37.115 ;
        RECT 25.845 36.960 26.135 37.005 ;
        RECT 26.750 36.960 27.070 37.020 ;
        RECT 25.845 36.820 27.070 36.960 ;
        RECT 25.845 36.775 26.135 36.820 ;
        RECT 26.750 36.760 27.070 36.820 ;
        RECT 33.665 36.775 33.955 37.005 ;
        RECT 36.425 36.960 36.715 37.005 ;
        RECT 39.285 36.960 39.500 37.115 ;
        RECT 41.930 37.100 42.250 37.160 ;
        RECT 43.390 37.115 43.680 37.160 ;
        RECT 45.700 37.160 58.720 37.300 ;
        RECT 59.960 37.160 62.170 37.300 ;
        RECT 41.530 36.960 41.820 37.005 ;
        RECT 36.425 36.820 38.940 36.960 ;
        RECT 39.285 36.820 41.820 36.960 ;
        RECT 36.425 36.775 36.715 36.820 ;
        RECT 14.345 36.435 14.635 36.665 ;
        RECT 14.420 35.940 14.560 36.435 ;
        RECT 15.710 36.420 16.030 36.680 ;
        RECT 22.610 36.620 22.930 36.680 ;
        RECT 26.305 36.620 26.595 36.665 ;
        RECT 32.730 36.620 33.050 36.680 ;
        RECT 22.610 36.480 33.050 36.620 ;
        RECT 22.610 36.420 22.930 36.480 ;
        RECT 26.305 36.435 26.595 36.480 ;
        RECT 32.730 36.420 33.050 36.480 ;
        RECT 15.215 36.280 15.505 36.325 ;
        RECT 17.105 36.280 17.395 36.325 ;
        RECT 20.225 36.280 20.515 36.325 ;
        RECT 15.215 36.140 20.515 36.280 ;
        RECT 33.740 36.280 33.880 36.775 ;
        RECT 38.250 36.420 38.570 36.680 ;
        RECT 38.800 36.620 38.940 36.820 ;
        RECT 41.530 36.775 41.820 36.820 ;
        RECT 44.690 36.620 45.010 36.680 ;
        RECT 38.800 36.480 45.010 36.620 ;
        RECT 44.690 36.420 45.010 36.480 ;
        RECT 36.890 36.280 37.180 36.325 ;
        RECT 38.750 36.280 39.040 36.325 ;
        RECT 41.530 36.280 41.820 36.325 ;
        RECT 45.700 36.280 45.840 37.160 ;
        RECT 48.385 37.115 48.675 37.160 ;
        RECT 46.990 36.960 47.310 37.020 ;
        RECT 57.110 36.960 57.430 37.020 ;
        RECT 58.505 36.960 58.795 37.005 ;
        RECT 59.960 36.960 60.100 37.160 ;
        RECT 46.990 36.820 60.100 36.960 ;
        RECT 46.990 36.760 47.310 36.820 ;
        RECT 57.110 36.760 57.430 36.820 ;
        RECT 58.505 36.775 58.795 36.820 ;
        RECT 60.330 36.760 60.650 37.020 ;
        RECT 62.720 36.960 62.860 37.500 ;
        RECT 63.550 37.500 64.775 37.640 ;
        RECT 63.550 37.440 63.870 37.500 ;
        RECT 64.485 37.455 64.775 37.500 ;
        RECT 70.450 37.440 70.770 37.700 ;
        RECT 73.670 37.440 73.990 37.700 ;
        RECT 77.810 37.440 78.130 37.700 ;
        RECT 80.110 37.440 80.430 37.700 ;
        RECT 93.450 37.640 93.770 37.700 ;
        RECT 98.510 37.640 98.830 37.700 ;
        RECT 81.580 37.500 98.830 37.640 ;
        RECT 63.105 37.300 63.395 37.345 ;
        RECT 77.365 37.300 77.655 37.345 ;
        RECT 81.580 37.300 81.720 37.500 ;
        RECT 93.450 37.440 93.770 37.500 ;
        RECT 98.510 37.440 98.830 37.500 ;
        RECT 104.490 37.440 104.810 37.700 ;
        RECT 63.105 37.160 67.460 37.300 ;
        RECT 63.105 37.115 63.395 37.160 ;
        RECT 67.320 37.020 67.460 37.160 ;
        RECT 77.365 37.160 81.720 37.300 ;
        RECT 81.950 37.300 82.270 37.360 ;
        RECT 84.725 37.300 85.015 37.345 ;
        RECT 81.950 37.160 85.015 37.300 ;
        RECT 77.365 37.115 77.655 37.160 ;
        RECT 81.950 37.100 82.270 37.160 ;
        RECT 84.725 37.115 85.015 37.160 ;
        RECT 87.005 37.300 87.655 37.345 ;
        RECT 90.605 37.300 90.895 37.345 ;
        RECT 87.005 37.160 90.895 37.300 ;
        RECT 87.005 37.115 87.655 37.160 ;
        RECT 90.305 37.115 90.895 37.160 ;
        RECT 91.610 37.300 91.930 37.360 ;
        RECT 94.025 37.300 94.315 37.345 ;
        RECT 97.265 37.300 97.915 37.345 ;
        RECT 91.610 37.160 97.915 37.300 ;
        RECT 63.690 36.960 63.980 37.005 ;
        RECT 64.470 36.960 64.790 37.020 ;
        RECT 65.405 36.960 65.695 37.005 ;
        RECT 62.720 36.820 63.320 36.960 ;
        RECT 47.910 36.620 48.230 36.680 ;
        RECT 48.845 36.620 49.135 36.665 ;
        RECT 47.910 36.480 49.135 36.620 ;
        RECT 47.910 36.420 48.230 36.480 ;
        RECT 48.845 36.435 49.135 36.480 ;
        RECT 61.265 36.620 61.555 36.665 ;
        RECT 61.265 36.480 62.170 36.620 ;
        RECT 61.265 36.435 61.555 36.480 ;
        RECT 33.740 36.140 36.640 36.280 ;
        RECT 15.215 36.095 15.505 36.140 ;
        RECT 17.105 36.095 17.395 36.140 ;
        RECT 20.225 36.095 20.515 36.140 ;
        RECT 18.470 35.940 18.790 36.000 ;
        RECT 14.420 35.800 18.790 35.940 ;
        RECT 18.470 35.740 18.790 35.800 ;
        RECT 23.545 35.940 23.835 35.985 ;
        RECT 24.910 35.940 25.230 36.000 ;
        RECT 23.545 35.800 25.230 35.940 ;
        RECT 23.545 35.755 23.835 35.800 ;
        RECT 24.910 35.740 25.230 35.800 ;
        RECT 35.490 35.740 35.810 36.000 ;
        RECT 36.500 35.940 36.640 36.140 ;
        RECT 36.890 36.140 41.820 36.280 ;
        RECT 36.890 36.095 37.180 36.140 ;
        RECT 38.750 36.095 39.040 36.140 ;
        RECT 41.530 36.095 41.820 36.140 ;
        RECT 45.470 36.140 45.840 36.280 ;
        RECT 62.030 36.280 62.170 36.480 ;
        RECT 62.630 36.420 62.950 36.680 ;
        RECT 63.180 36.620 63.320 36.820 ;
        RECT 63.690 36.820 65.695 36.960 ;
        RECT 63.690 36.775 63.980 36.820 ;
        RECT 64.470 36.760 64.790 36.820 ;
        RECT 65.405 36.775 65.695 36.820 ;
        RECT 67.230 36.760 67.550 37.020 ;
        RECT 74.605 36.960 74.895 37.005 ;
        RECT 80.570 36.960 80.890 37.020 ;
        RECT 81.505 36.960 81.795 37.005 ;
        RECT 74.605 36.820 75.740 36.960 ;
        RECT 74.605 36.775 74.895 36.820 ;
        RECT 67.690 36.620 68.010 36.680 ;
        RECT 63.180 36.480 68.010 36.620 ;
        RECT 67.690 36.420 68.010 36.480 ;
        RECT 63.090 36.280 63.410 36.340 ;
        RECT 65.390 36.280 65.710 36.340 ;
        RECT 75.600 36.325 75.740 36.820 ;
        RECT 80.570 36.820 81.795 36.960 ;
        RECT 80.570 36.760 80.890 36.820 ;
        RECT 81.505 36.775 81.795 36.820 ;
        RECT 83.810 36.960 84.100 37.005 ;
        RECT 85.645 36.960 85.935 37.005 ;
        RECT 89.225 36.960 89.515 37.005 ;
        RECT 83.810 36.820 89.515 36.960 ;
        RECT 83.810 36.775 84.100 36.820 ;
        RECT 85.645 36.775 85.935 36.820 ;
        RECT 89.225 36.775 89.515 36.820 ;
        RECT 90.305 36.800 90.595 37.115 ;
        RECT 91.610 37.100 91.930 37.160 ;
        RECT 94.025 37.115 94.615 37.160 ;
        RECT 97.265 37.115 97.915 37.160 ;
        RECT 94.325 36.800 94.615 37.115 ;
        RECT 95.405 36.960 95.695 37.005 ;
        RECT 98.985 36.960 99.275 37.005 ;
        RECT 100.820 36.960 101.110 37.005 ;
        RECT 95.405 36.820 101.110 36.960 ;
        RECT 75.970 36.620 76.290 36.680 ;
        RECT 78.285 36.620 78.575 36.665 ;
        RECT 75.970 36.480 78.575 36.620 ;
        RECT 75.970 36.420 76.290 36.480 ;
        RECT 78.285 36.435 78.575 36.480 ;
        RECT 83.330 36.420 83.650 36.680 ;
        RECT 90.320 36.620 90.460 36.800 ;
        RECT 95.405 36.775 95.695 36.820 ;
        RECT 98.985 36.775 99.275 36.820 ;
        RECT 100.820 36.775 101.110 36.820 ;
        RECT 101.285 36.960 101.575 37.005 ;
        RECT 104.030 36.960 104.350 37.020 ;
        RECT 101.285 36.820 104.350 36.960 ;
        RECT 101.285 36.775 101.575 36.820 ;
        RECT 104.030 36.760 104.350 36.820 ;
        RECT 104.965 36.960 105.255 37.005 ;
        RECT 111.390 36.960 111.710 37.020 ;
        RECT 104.965 36.820 111.710 36.960 ;
        RECT 104.965 36.775 105.255 36.820 ;
        RECT 111.390 36.760 111.710 36.820 ;
        RECT 83.880 36.480 90.460 36.620 ;
        RECT 62.030 36.140 65.710 36.280 ;
        RECT 45.470 35.985 45.610 36.140 ;
        RECT 63.090 36.080 63.410 36.140 ;
        RECT 65.390 36.080 65.710 36.140 ;
        RECT 75.525 36.095 75.815 36.325 ;
        RECT 81.965 36.280 82.255 36.325 ;
        RECT 83.880 36.280 84.020 36.480 ;
        RECT 92.070 36.420 92.390 36.680 ;
        RECT 96.670 36.620 96.990 36.680 ;
        RECT 99.905 36.620 100.195 36.665 ;
        RECT 96.670 36.480 100.195 36.620 ;
        RECT 96.670 36.420 96.990 36.480 ;
        RECT 99.905 36.435 100.195 36.480 ;
        RECT 81.965 36.140 84.020 36.280 ;
        RECT 84.215 36.280 84.505 36.325 ;
        RECT 86.105 36.280 86.395 36.325 ;
        RECT 89.225 36.280 89.515 36.325 ;
        RECT 84.215 36.140 89.515 36.280 ;
        RECT 81.965 36.095 82.255 36.140 ;
        RECT 84.215 36.095 84.505 36.140 ;
        RECT 86.105 36.095 86.395 36.140 ;
        RECT 89.225 36.095 89.515 36.140 ;
        RECT 90.230 36.280 90.550 36.340 ;
        RECT 92.545 36.280 92.835 36.325 ;
        RECT 90.230 36.140 92.835 36.280 ;
        RECT 90.230 36.080 90.550 36.140 ;
        RECT 92.545 36.095 92.835 36.140 ;
        RECT 95.405 36.280 95.695 36.325 ;
        RECT 98.525 36.280 98.815 36.325 ;
        RECT 100.415 36.280 100.705 36.325 ;
        RECT 95.405 36.140 100.705 36.280 ;
        RECT 95.405 36.095 95.695 36.140 ;
        RECT 98.525 36.095 98.815 36.140 ;
        RECT 100.415 36.095 100.705 36.140 ;
        RECT 45.395 35.940 45.685 35.985 ;
        RECT 36.500 35.800 45.685 35.940 ;
        RECT 45.395 35.755 45.685 35.800 ;
        RECT 58.045 35.940 58.335 35.985 ;
        RECT 58.490 35.940 58.810 36.000 ;
        RECT 58.045 35.800 58.810 35.940 ;
        RECT 58.045 35.755 58.335 35.800 ;
        RECT 58.490 35.740 58.810 35.800 ;
        RECT 63.550 35.940 63.870 36.000 ;
        RECT 65.865 35.940 66.155 35.985 ;
        RECT 63.550 35.800 66.155 35.940 ;
        RECT 63.550 35.740 63.870 35.800 ;
        RECT 65.865 35.755 66.155 35.800 ;
        RECT 5.520 35.120 125.580 35.600 ;
        RECT 14.345 34.920 14.635 34.965 ;
        RECT 15.710 34.920 16.030 34.980 ;
        RECT 14.345 34.780 16.030 34.920 ;
        RECT 14.345 34.735 14.635 34.780 ;
        RECT 15.710 34.720 16.030 34.780 ;
        RECT 27.225 34.920 27.515 34.965 ;
        RECT 27.670 34.920 27.990 34.980 ;
        RECT 27.225 34.780 27.990 34.920 ;
        RECT 27.225 34.735 27.515 34.780 ;
        RECT 27.670 34.720 27.990 34.780 ;
        RECT 85.580 34.920 85.870 34.965 ;
        RECT 94.370 34.920 94.690 34.980 ;
        RECT 85.580 34.780 94.690 34.920 ;
        RECT 85.580 34.735 85.870 34.780 ;
        RECT 94.370 34.720 94.690 34.780 ;
        RECT 98.050 34.720 98.370 34.980 ;
        RECT 23.990 34.580 24.310 34.640 ;
        RECT 22.240 34.440 24.310 34.580 ;
        RECT 22.240 34.285 22.380 34.440 ;
        RECT 23.990 34.380 24.310 34.440 ;
        RECT 30.085 34.580 30.375 34.625 ;
        RECT 33.205 34.580 33.495 34.625 ;
        RECT 35.095 34.580 35.385 34.625 ;
        RECT 30.085 34.440 35.385 34.580 ;
        RECT 30.085 34.395 30.375 34.440 ;
        RECT 33.205 34.395 33.495 34.440 ;
        RECT 35.095 34.395 35.385 34.440 ;
        RECT 52.935 34.580 53.225 34.625 ;
        RECT 54.825 34.580 55.115 34.625 ;
        RECT 57.945 34.580 58.235 34.625 ;
        RECT 52.935 34.440 58.235 34.580 ;
        RECT 52.935 34.395 53.225 34.440 ;
        RECT 54.825 34.395 55.115 34.440 ;
        RECT 57.945 34.395 58.235 34.440 ;
        RECT 67.690 34.380 68.010 34.640 ;
        RECT 85.135 34.580 85.425 34.625 ;
        RECT 87.025 34.580 87.315 34.625 ;
        RECT 90.145 34.580 90.435 34.625 ;
        RECT 85.135 34.440 90.435 34.580 ;
        RECT 85.135 34.395 85.425 34.440 ;
        RECT 87.025 34.395 87.315 34.440 ;
        RECT 90.145 34.395 90.435 34.440 ;
        RECT 22.165 34.055 22.455 34.285 ;
        RECT 22.610 34.040 22.930 34.300 ;
        RECT 35.965 34.240 36.255 34.285 ;
        RECT 23.160 34.100 36.255 34.240 ;
        RECT 13.425 33.900 13.715 33.945 ;
        RECT 14.805 33.900 15.095 33.945 ;
        RECT 13.425 33.760 15.095 33.900 ;
        RECT 13.425 33.715 13.715 33.760 ;
        RECT 14.805 33.715 15.095 33.760 ;
        RECT 18.025 33.715 18.315 33.945 ;
        RECT 18.470 33.900 18.790 33.960 ;
        RECT 23.160 33.900 23.300 34.100 ;
        RECT 35.965 34.055 36.255 34.100 ;
        RECT 41.025 34.240 41.315 34.285 ;
        RECT 41.930 34.240 42.250 34.300 ;
        RECT 41.025 34.100 42.250 34.240 ;
        RECT 41.025 34.055 41.315 34.100 ;
        RECT 41.930 34.040 42.250 34.100 ;
        RECT 53.445 34.240 53.735 34.285 ;
        RECT 56.650 34.240 56.970 34.300 ;
        RECT 53.445 34.100 56.970 34.240 ;
        RECT 53.445 34.055 53.735 34.100 ;
        RECT 56.650 34.040 56.970 34.100 ;
        RECT 60.805 34.240 61.095 34.285 ;
        RECT 64.470 34.240 64.790 34.300 ;
        RECT 60.805 34.100 64.790 34.240 ;
        RECT 67.780 34.240 67.920 34.380 ;
        RECT 72.750 34.240 73.070 34.300 ;
        RECT 67.780 34.100 73.070 34.240 ;
        RECT 60.805 34.055 61.095 34.100 ;
        RECT 64.470 34.040 64.790 34.100 ;
        RECT 72.750 34.040 73.070 34.100 ;
        RECT 92.990 34.040 93.310 34.300 ;
        RECT 18.470 33.760 23.300 33.900 ;
        RECT 18.100 33.560 18.240 33.715 ;
        RECT 18.470 33.700 18.790 33.760 ;
        RECT 24.910 33.700 25.230 33.960 ;
        RECT 21.705 33.560 21.995 33.605 ;
        RECT 26.750 33.560 27.070 33.620 ;
        RECT 29.005 33.605 29.295 33.920 ;
        RECT 30.085 33.900 30.375 33.945 ;
        RECT 33.665 33.900 33.955 33.945 ;
        RECT 35.500 33.900 35.790 33.945 ;
        RECT 30.085 33.760 35.790 33.900 ;
        RECT 30.085 33.715 30.375 33.760 ;
        RECT 33.665 33.715 33.955 33.760 ;
        RECT 35.500 33.715 35.790 33.760 ;
        RECT 39.170 33.900 39.490 33.960 ;
        RECT 40.565 33.900 40.855 33.945 ;
        RECT 39.170 33.760 40.855 33.900 ;
        RECT 39.170 33.700 39.490 33.760 ;
        RECT 40.565 33.715 40.855 33.760 ;
        RECT 49.290 33.900 49.610 33.960 ;
        RECT 52.050 33.900 52.370 33.960 ;
        RECT 49.290 33.760 52.370 33.900 ;
        RECT 49.290 33.700 49.610 33.760 ;
        RECT 52.050 33.700 52.370 33.760 ;
        RECT 52.530 33.900 52.820 33.945 ;
        RECT 54.365 33.900 54.655 33.945 ;
        RECT 57.945 33.900 58.235 33.945 ;
        RECT 52.530 33.760 58.235 33.900 ;
        RECT 52.530 33.715 52.820 33.760 ;
        RECT 54.365 33.715 54.655 33.760 ;
        RECT 57.945 33.715 58.235 33.760 ;
        RECT 32.270 33.605 32.590 33.620 ;
        RECT 18.100 33.420 20.080 33.560 ;
        RECT 19.940 33.265 20.080 33.420 ;
        RECT 21.705 33.420 27.070 33.560 ;
        RECT 21.705 33.375 21.995 33.420 ;
        RECT 26.750 33.360 27.070 33.420 ;
        RECT 28.705 33.560 29.295 33.605 ;
        RECT 31.945 33.560 32.595 33.605 ;
        RECT 28.705 33.420 32.595 33.560 ;
        RECT 28.705 33.375 28.995 33.420 ;
        RECT 31.945 33.375 32.595 33.420 ;
        RECT 32.270 33.360 32.590 33.375 ;
        RECT 34.570 33.360 34.890 33.620 ;
        RECT 55.725 33.560 56.375 33.605 ;
        RECT 58.490 33.560 58.810 33.620 ;
        RECT 59.025 33.605 59.315 33.920 ;
        RECT 61.265 33.900 61.555 33.945 ;
        RECT 62.630 33.900 62.950 33.960 ;
        RECT 61.265 33.760 62.950 33.900 ;
        RECT 61.265 33.715 61.555 33.760 ;
        RECT 62.630 33.700 62.950 33.760 ;
        RECT 83.790 33.900 84.110 33.960 ;
        RECT 84.265 33.900 84.555 33.945 ;
        RECT 83.790 33.760 84.555 33.900 ;
        RECT 83.790 33.700 84.110 33.760 ;
        RECT 84.265 33.715 84.555 33.760 ;
        RECT 84.730 33.900 85.020 33.945 ;
        RECT 86.565 33.900 86.855 33.945 ;
        RECT 90.145 33.900 90.435 33.945 ;
        RECT 84.730 33.760 90.435 33.900 ;
        RECT 84.730 33.715 85.020 33.760 ;
        RECT 86.565 33.715 86.855 33.760 ;
        RECT 90.145 33.715 90.435 33.760 ;
        RECT 91.225 33.605 91.515 33.920 ;
        RECT 93.910 33.700 94.230 33.960 ;
        RECT 97.130 33.700 97.450 33.960 ;
        RECT 59.025 33.560 59.615 33.605 ;
        RECT 55.725 33.420 59.615 33.560 ;
        RECT 55.725 33.375 56.375 33.420 ;
        RECT 58.490 33.360 58.810 33.420 ;
        RECT 59.325 33.375 59.615 33.420 ;
        RECT 87.925 33.560 88.575 33.605 ;
        RECT 91.225 33.560 91.815 33.605 ;
        RECT 97.590 33.560 97.910 33.620 ;
        RECT 87.925 33.420 97.910 33.560 ;
        RECT 87.925 33.375 88.575 33.420 ;
        RECT 91.525 33.375 91.815 33.420 ;
        RECT 97.590 33.360 97.910 33.420 ;
        RECT 19.865 33.035 20.155 33.265 ;
        RECT 23.990 33.020 24.310 33.280 ;
        RECT 62.170 33.220 62.490 33.280 ;
        RECT 64.010 33.220 64.330 33.280 ;
        RECT 62.170 33.080 64.330 33.220 ;
        RECT 62.170 33.020 62.490 33.080 ;
        RECT 64.010 33.020 64.330 33.080 ;
        RECT 94.845 33.220 95.135 33.265 ;
        RECT 96.670 33.220 96.990 33.280 ;
        RECT 94.845 33.080 96.990 33.220 ;
        RECT 94.845 33.035 95.135 33.080 ;
        RECT 96.670 33.020 96.990 33.080 ;
        RECT 5.520 32.400 125.580 32.880 ;
        RECT 23.990 32.200 24.310 32.260 ;
        RECT 19.940 32.060 24.310 32.200 ;
        RECT 19.940 31.905 20.080 32.060 ;
        RECT 23.990 32.000 24.310 32.060 ;
        RECT 26.750 32.200 27.070 32.260 ;
        RECT 27.685 32.200 27.975 32.245 ;
        RECT 26.750 32.060 27.975 32.200 ;
        RECT 26.750 32.000 27.070 32.060 ;
        RECT 27.685 32.015 27.975 32.060 ;
        RECT 32.270 32.000 32.590 32.260 ;
        RECT 34.125 32.200 34.415 32.245 ;
        RECT 34.570 32.200 34.890 32.260 ;
        RECT 34.125 32.060 34.890 32.200 ;
        RECT 34.125 32.015 34.415 32.060 ;
        RECT 34.570 32.000 34.890 32.060 ;
        RECT 55.285 32.200 55.575 32.245 ;
        RECT 56.650 32.200 56.970 32.260 ;
        RECT 55.285 32.060 56.970 32.200 ;
        RECT 55.285 32.015 55.575 32.060 ;
        RECT 56.650 32.000 56.970 32.060 ;
        RECT 57.585 32.015 57.875 32.245 ;
        RECT 58.425 32.200 58.715 32.245 ;
        RECT 61.855 32.200 62.145 32.245 ;
        RECT 63.105 32.200 63.395 32.245 ;
        RECT 58.425 32.060 61.020 32.200 ;
        RECT 58.425 32.015 58.715 32.060 ;
        RECT 19.865 31.675 20.155 31.905 ;
        RECT 22.145 31.860 22.795 31.905 ;
        RECT 25.745 31.860 26.035 31.905 ;
        RECT 57.110 31.860 57.430 31.920 ;
        RECT 22.145 31.720 26.035 31.860 ;
        RECT 22.145 31.675 22.795 31.720 ;
        RECT 25.445 31.675 26.035 31.720 ;
        RECT 32.820 31.720 57.430 31.860 ;
        RECT 18.010 31.320 18.330 31.580 ;
        RECT 18.470 31.320 18.790 31.580 ;
        RECT 18.950 31.520 19.240 31.565 ;
        RECT 20.785 31.520 21.075 31.565 ;
        RECT 24.365 31.520 24.655 31.565 ;
        RECT 18.950 31.380 24.655 31.520 ;
        RECT 18.950 31.335 19.240 31.380 ;
        RECT 20.785 31.335 21.075 31.380 ;
        RECT 24.365 31.335 24.655 31.380 ;
        RECT 25.445 31.520 25.735 31.675 ;
        RECT 28.130 31.520 28.450 31.580 ;
        RECT 25.445 31.380 28.450 31.520 ;
        RECT 25.445 31.360 25.735 31.380 ;
        RECT 28.130 31.320 28.450 31.380 ;
        RECT 28.590 31.520 28.910 31.580 ;
        RECT 32.820 31.565 32.960 31.720 ;
        RECT 32.745 31.520 33.035 31.565 ;
        RECT 28.590 31.380 33.035 31.520 ;
        RECT 28.590 31.320 28.910 31.380 ;
        RECT 32.745 31.335 33.035 31.380 ;
        RECT 33.205 31.520 33.495 31.565 ;
        RECT 35.490 31.520 35.810 31.580 ;
        RECT 53.520 31.565 53.660 31.720 ;
        RECT 57.110 31.660 57.430 31.720 ;
        RECT 33.205 31.380 35.810 31.520 ;
        RECT 33.205 31.335 33.495 31.380 ;
        RECT 35.490 31.320 35.810 31.380 ;
        RECT 53.445 31.335 53.735 31.565 ;
        RECT 56.205 31.520 56.495 31.565 ;
        RECT 57.660 31.520 57.800 32.015 ;
        RECT 60.880 31.905 61.020 32.060 ;
        RECT 61.855 32.060 63.395 32.200 ;
        RECT 61.855 32.015 62.145 32.060 ;
        RECT 63.105 32.015 63.395 32.060 ;
        RECT 59.425 31.675 59.715 31.905 ;
        RECT 60.805 31.860 61.095 31.905 ;
        RECT 61.250 31.860 61.570 31.920 ;
        RECT 60.805 31.720 61.570 31.860 ;
        RECT 60.805 31.675 61.095 31.720 ;
        RECT 56.205 31.380 57.800 31.520 ;
        RECT 58.030 31.520 58.350 31.580 ;
        RECT 59.500 31.520 59.640 31.675 ;
        RECT 61.250 31.660 61.570 31.720 ;
        RECT 58.030 31.380 59.640 31.520 ;
        RECT 60.330 31.520 60.650 31.580 ;
        RECT 64.485 31.520 64.775 31.565 ;
        RECT 60.330 31.380 64.775 31.520 ;
        RECT 56.205 31.335 56.495 31.380 ;
        RECT 58.030 31.320 58.350 31.380 ;
        RECT 60.330 31.320 60.650 31.380 ;
        RECT 64.485 31.335 64.775 31.380 ;
        RECT 69.070 31.520 69.390 31.580 ;
        RECT 71.845 31.520 72.135 31.565 ;
        RECT 69.070 31.380 72.135 31.520 ;
        RECT 69.070 31.320 69.390 31.380 ;
        RECT 71.845 31.335 72.135 31.380 ;
        RECT 72.750 31.320 73.070 31.580 ;
        RECT 18.100 31.180 18.240 31.320 ;
        RECT 18.100 31.040 25.600 31.180 ;
        RECT 19.355 30.840 19.645 30.885 ;
        RECT 21.245 30.840 21.535 30.885 ;
        RECT 24.365 30.840 24.655 30.885 ;
        RECT 19.355 30.700 24.655 30.840 ;
        RECT 25.460 30.840 25.600 31.040 ;
        RECT 30.445 30.995 30.735 31.225 ;
        RECT 28.590 30.840 28.910 30.900 ;
        RECT 25.460 30.700 28.910 30.840 ;
        RECT 19.355 30.655 19.645 30.700 ;
        RECT 21.245 30.655 21.535 30.700 ;
        RECT 24.365 30.655 24.655 30.700 ;
        RECT 28.590 30.640 28.910 30.700 ;
        RECT 17.565 30.500 17.855 30.545 ;
        RECT 20.770 30.500 21.090 30.560 ;
        RECT 17.565 30.360 21.090 30.500 ;
        RECT 17.565 30.315 17.855 30.360 ;
        RECT 20.770 30.300 21.090 30.360 ;
        RECT 23.530 30.500 23.850 30.560 ;
        RECT 27.225 30.500 27.515 30.545 ;
        RECT 30.520 30.500 30.660 30.995 ;
        RECT 64.010 30.980 64.330 31.240 ;
        RECT 64.945 30.995 65.235 31.225 ;
        RECT 60.330 30.840 60.650 30.900 ;
        RECT 63.550 30.840 63.870 30.900 ;
        RECT 65.020 30.840 65.160 30.995 ;
        RECT 65.390 30.980 65.710 31.240 ;
        RECT 60.330 30.700 65.160 30.840 ;
        RECT 60.330 30.640 60.650 30.700 ;
        RECT 63.550 30.640 63.870 30.700 ;
        RECT 23.530 30.360 30.660 30.500 ;
        RECT 23.530 30.300 23.850 30.360 ;
        RECT 27.225 30.315 27.515 30.360 ;
        RECT 53.890 30.300 54.210 30.560 ;
        RECT 58.490 30.300 58.810 30.560 ;
        RECT 61.710 30.300 62.030 30.560 ;
        RECT 62.645 30.500 62.935 30.545 ;
        RECT 66.310 30.500 66.630 30.560 ;
        RECT 62.645 30.360 66.630 30.500 ;
        RECT 62.645 30.315 62.935 30.360 ;
        RECT 66.310 30.300 66.630 30.360 ;
        RECT 66.770 30.500 67.090 30.560 ;
        RECT 69.085 30.500 69.375 30.545 ;
        RECT 66.770 30.360 69.375 30.500 ;
        RECT 66.770 30.300 67.090 30.360 ;
        RECT 69.085 30.315 69.375 30.360 ;
        RECT 73.210 30.300 73.530 30.560 ;
        RECT 5.520 29.680 125.580 30.160 ;
        RECT 28.130 29.280 28.450 29.540 ;
        RECT 58.045 29.480 58.335 29.525 ;
        RECT 62.630 29.480 62.950 29.540 ;
        RECT 58.045 29.340 62.950 29.480 ;
        RECT 58.045 29.295 58.335 29.340 ;
        RECT 62.630 29.280 62.950 29.340 ;
        RECT 64.945 29.480 65.235 29.525 ;
        RECT 69.070 29.480 69.390 29.540 ;
        RECT 70.925 29.480 71.215 29.525 ;
        RECT 64.945 29.340 71.215 29.480 ;
        RECT 64.945 29.295 65.235 29.340 ;
        RECT 69.070 29.280 69.390 29.340 ;
        RECT 70.925 29.295 71.215 29.340 ;
        RECT 50.175 29.140 50.465 29.185 ;
        RECT 52.065 29.140 52.355 29.185 ;
        RECT 55.185 29.140 55.475 29.185 ;
        RECT 50.175 29.000 55.475 29.140 ;
        RECT 50.175 28.955 50.465 29.000 ;
        RECT 52.065 28.955 52.355 29.000 ;
        RECT 55.185 28.955 55.475 29.000 ;
        RECT 61.710 28.940 62.030 29.200 ;
        RECT 63.090 29.140 63.410 29.200 ;
        RECT 65.390 29.140 65.710 29.200 ;
        RECT 63.090 29.000 65.710 29.140 ;
        RECT 63.090 28.940 63.410 29.000 ;
        RECT 65.390 28.940 65.710 29.000 ;
        RECT 68.625 28.955 68.915 29.185 ;
        RECT 73.785 29.140 74.075 29.185 ;
        RECT 76.905 29.140 77.195 29.185 ;
        RECT 78.795 29.140 79.085 29.185 ;
        RECT 73.785 29.000 79.085 29.140 ;
        RECT 73.785 28.955 74.075 29.000 ;
        RECT 76.905 28.955 77.195 29.000 ;
        RECT 78.795 28.955 79.085 29.000 ;
        RECT 60.330 28.800 60.650 28.860 ;
        RECT 58.580 28.660 60.650 28.800 ;
        RECT 61.800 28.800 61.940 28.940 ;
        RECT 66.325 28.800 66.615 28.845 ;
        RECT 61.800 28.660 66.615 28.800 ;
        RECT 68.700 28.800 68.840 28.955 ;
        RECT 78.285 28.800 78.575 28.845 ;
        RECT 68.700 28.660 78.575 28.800 ;
        RECT 28.590 28.260 28.910 28.520 ;
        RECT 49.290 28.260 49.610 28.520 ;
        RECT 58.580 28.505 58.720 28.660 ;
        RECT 60.330 28.600 60.650 28.660 ;
        RECT 66.325 28.615 66.615 28.660 ;
        RECT 78.285 28.615 78.575 28.660 ;
        RECT 79.665 28.800 79.955 28.845 ;
        RECT 83.790 28.800 84.110 28.860 ;
        RECT 79.665 28.660 84.110 28.800 ;
        RECT 79.665 28.615 79.955 28.660 ;
        RECT 83.790 28.600 84.110 28.660 ;
        RECT 49.770 28.460 50.060 28.505 ;
        RECT 51.605 28.460 51.895 28.505 ;
        RECT 55.185 28.460 55.475 28.505 ;
        RECT 49.770 28.320 55.475 28.460 ;
        RECT 49.770 28.275 50.060 28.320 ;
        RECT 51.605 28.275 51.895 28.320 ;
        RECT 55.185 28.275 55.475 28.320 ;
        RECT 50.670 27.920 50.990 28.180 ;
        RECT 52.965 28.120 53.615 28.165 ;
        RECT 53.890 28.120 54.210 28.180 ;
        RECT 56.265 28.165 56.555 28.480 ;
        RECT 58.505 28.275 58.795 28.505 ;
        RECT 59.425 28.275 59.715 28.505 ;
        RECT 62.185 28.460 62.475 28.505 ;
        RECT 63.090 28.460 63.410 28.520 ;
        RECT 62.185 28.320 63.410 28.460 ;
        RECT 62.185 28.275 62.475 28.320 ;
        RECT 56.265 28.120 56.855 28.165 ;
        RECT 52.965 27.980 56.855 28.120 ;
        RECT 59.500 28.120 59.640 28.275 ;
        RECT 63.090 28.260 63.410 28.320 ;
        RECT 63.550 28.260 63.870 28.520 ;
        RECT 65.405 28.275 65.695 28.505 ;
        RECT 65.480 28.120 65.620 28.275 ;
        RECT 66.770 28.260 67.090 28.520 ;
        RECT 72.705 28.165 72.995 28.480 ;
        RECT 73.785 28.460 74.075 28.505 ;
        RECT 77.365 28.460 77.655 28.505 ;
        RECT 79.200 28.460 79.490 28.505 ;
        RECT 73.785 28.320 79.490 28.460 ;
        RECT 73.785 28.275 74.075 28.320 ;
        RECT 77.365 28.275 77.655 28.320 ;
        RECT 79.200 28.275 79.490 28.320 ;
        RECT 59.500 27.980 65.620 28.120 ;
        RECT 72.405 28.120 72.995 28.165 ;
        RECT 73.210 28.120 73.530 28.180 ;
        RECT 75.645 28.120 76.295 28.165 ;
        RECT 72.405 27.980 76.295 28.120 ;
        RECT 52.965 27.935 53.615 27.980 ;
        RECT 53.890 27.920 54.210 27.980 ;
        RECT 56.565 27.935 56.855 27.980 ;
        RECT 58.030 27.780 58.350 27.840 ;
        RECT 58.505 27.780 58.795 27.825 ;
        RECT 58.030 27.640 58.795 27.780 ;
        RECT 58.030 27.580 58.350 27.640 ;
        RECT 58.505 27.595 58.795 27.640 ;
        RECT 60.790 27.780 61.110 27.840 ;
        RECT 61.340 27.825 61.480 27.980 ;
        RECT 72.405 27.935 72.695 27.980 ;
        RECT 73.210 27.920 73.530 27.980 ;
        RECT 75.645 27.935 76.295 27.980 ;
        RECT 61.265 27.780 61.555 27.825 ;
        RECT 60.790 27.640 61.555 27.780 ;
        RECT 60.790 27.580 61.110 27.640 ;
        RECT 61.265 27.595 61.555 27.640 ;
        RECT 61.710 27.580 62.030 27.840 ;
        RECT 62.630 27.580 62.950 27.840 ;
        RECT 5.520 26.960 125.580 27.440 ;
        RECT 50.670 26.760 50.990 26.820 ;
        RECT 52.525 26.760 52.815 26.805 ;
        RECT 50.670 26.620 52.815 26.760 ;
        RECT 50.670 26.560 50.990 26.620 ;
        RECT 52.525 26.575 52.815 26.620 ;
        RECT 58.490 26.560 58.810 26.820 ;
        RECT 61.250 26.560 61.570 26.820 ;
        RECT 49.290 26.420 49.610 26.480 ;
        RECT 68.145 26.420 68.795 26.465 ;
        RECT 71.745 26.420 72.035 26.465 ;
        RECT 49.290 26.280 64.700 26.420 ;
        RECT 49.290 26.220 49.610 26.280 ;
        RECT 54.365 25.895 54.655 26.125 ;
        RECT 59.425 26.080 59.715 26.125 ;
        RECT 59.870 26.080 60.190 26.140 ;
        RECT 59.425 25.940 60.190 26.080 ;
        RECT 59.425 25.895 59.715 25.940 ;
        RECT 54.440 25.060 54.580 25.895 ;
        RECT 59.870 25.880 60.190 25.940 ;
        RECT 60.345 26.080 60.635 26.125 ;
        RECT 60.790 26.080 61.110 26.140 ;
        RECT 60.345 25.940 61.110 26.080 ;
        RECT 60.345 25.895 60.635 25.940 ;
        RECT 60.790 25.880 61.110 25.940 ;
        RECT 62.630 25.880 62.950 26.140 ;
        RECT 63.090 26.080 63.410 26.140 ;
        RECT 64.560 26.125 64.700 26.280 ;
        RECT 68.145 26.280 72.035 26.420 ;
        RECT 68.145 26.235 68.795 26.280 ;
        RECT 71.445 26.235 72.035 26.280 ;
        RECT 64.025 26.080 64.315 26.125 ;
        RECT 63.090 25.940 64.315 26.080 ;
        RECT 63.090 25.880 63.410 25.940 ;
        RECT 64.025 25.895 64.315 25.940 ;
        RECT 64.485 25.895 64.775 26.125 ;
        RECT 64.950 26.080 65.240 26.125 ;
        RECT 66.785 26.080 67.075 26.125 ;
        RECT 70.365 26.080 70.655 26.125 ;
        RECT 64.950 25.940 70.655 26.080 ;
        RECT 64.950 25.895 65.240 25.940 ;
        RECT 66.785 25.895 67.075 25.940 ;
        RECT 70.365 25.895 70.655 25.940 ;
        RECT 71.445 26.080 71.735 26.235 ;
        RECT 71.445 25.940 72.060 26.080 ;
        RECT 71.445 25.920 71.735 25.940 ;
        RECT 54.825 25.740 55.115 25.785 ;
        RECT 58.030 25.740 58.350 25.800 ;
        RECT 54.825 25.600 58.350 25.740 ;
        RECT 64.100 25.740 64.240 25.895 ;
        RECT 71.920 25.800 72.060 25.940 ;
        RECT 64.100 25.600 64.700 25.740 ;
        RECT 54.825 25.555 55.115 25.600 ;
        RECT 58.030 25.540 58.350 25.600 ;
        RECT 61.710 25.060 62.030 25.120 ;
        RECT 62.185 25.060 62.475 25.105 ;
        RECT 64.010 25.060 64.330 25.120 ;
        RECT 54.440 24.920 64.330 25.060 ;
        RECT 64.560 25.060 64.700 25.600 ;
        RECT 65.850 25.540 66.170 25.800 ;
        RECT 71.830 25.540 72.150 25.800 ;
        RECT 74.605 25.555 74.895 25.785 ;
        RECT 65.355 25.400 65.645 25.445 ;
        RECT 67.245 25.400 67.535 25.445 ;
        RECT 70.365 25.400 70.655 25.445 ;
        RECT 65.355 25.260 70.655 25.400 ;
        RECT 65.355 25.215 65.645 25.260 ;
        RECT 67.245 25.215 67.535 25.260 ;
        RECT 70.365 25.215 70.655 25.260 ;
        RECT 74.680 25.060 74.820 25.555 ;
        RECT 64.560 24.920 74.820 25.060 ;
        RECT 61.710 24.860 62.030 24.920 ;
        RECT 62.185 24.875 62.475 24.920 ;
        RECT 64.010 24.860 64.330 24.920 ;
        RECT 5.520 24.240 125.580 24.720 ;
        RECT 65.850 24.040 66.170 24.100 ;
        RECT 67.245 24.040 67.535 24.085 ;
        RECT 65.850 23.900 67.535 24.040 ;
        RECT 65.850 23.840 66.170 23.900 ;
        RECT 67.245 23.855 67.535 23.900 ;
        RECT 70.925 24.040 71.215 24.085 ;
        RECT 71.830 24.040 72.150 24.100 ;
        RECT 70.925 23.900 72.150 24.040 ;
        RECT 70.925 23.855 71.215 23.900 ;
        RECT 71.830 23.840 72.150 23.900 ;
        RECT 66.310 23.020 66.630 23.080 ;
        RECT 68.165 23.020 68.455 23.065 ;
        RECT 66.310 22.880 68.455 23.020 ;
        RECT 66.310 22.820 66.630 22.880 ;
        RECT 68.165 22.835 68.455 22.880 ;
        RECT 71.385 23.020 71.675 23.065 ;
        RECT 72.750 23.020 73.070 23.080 ;
        RECT 71.385 22.880 73.070 23.020 ;
        RECT 71.385 22.835 71.675 22.880 ;
        RECT 72.750 22.820 73.070 22.880 ;
        RECT 5.520 21.520 125.580 22.000 ;
        RECT 5.520 18.800 125.580 19.280 ;
        RECT 5.520 16.080 125.580 16.560 ;
        RECT 5.520 13.360 125.580 13.840 ;
        RECT 5.520 10.640 125.580 11.120 ;
      LAYER met2 ;
        RECT 8.900 140.350 10.670 140.490 ;
        RECT 30.270 140.350 31.580 140.490 ;
        RECT 49.590 140.350 49.980 140.490 ;
        RECT 56.030 140.350 57.340 140.490 ;
        RECT 101.110 140.350 102.880 140.490 ;
        RECT 1.930 122.555 2.210 122.925 ;
        RECT 2.000 118.650 2.140 122.555 ;
        RECT 4.300 121.370 4.440 139.870 ;
        RECT 8.900 124.090 9.040 140.350 ;
        RECT 13.440 128.190 13.700 128.510 ;
        RECT 9.580 127.655 11.460 128.025 ;
        RECT 12.060 126.490 12.320 126.810 ;
        RECT 8.840 123.770 9.100 124.090 ;
        RECT 9.580 122.215 11.460 122.585 ;
        RECT 12.120 121.370 12.260 126.490 ;
        RECT 13.500 124.430 13.640 128.190 ;
        RECT 17.180 126.470 17.320 139.870 ;
        RECT 18.500 129.210 18.760 129.530 ;
        RECT 17.120 126.150 17.380 126.470 ;
        RECT 17.580 125.810 17.840 126.130 ;
        RECT 13.440 124.110 13.700 124.430 ;
        RECT 17.640 124.090 17.780 125.810 ;
        RECT 18.560 124.090 18.700 129.210 ;
        RECT 20.340 125.470 20.600 125.790 ;
        RECT 17.580 123.770 17.840 124.090 ;
        RECT 18.500 123.770 18.760 124.090 ;
        RECT 12.520 123.430 12.780 123.750 ;
        RECT 17.120 123.430 17.380 123.750 ;
        RECT 4.240 121.050 4.500 121.370 ;
        RECT 12.060 121.050 12.320 121.370 ;
        RECT 12.120 120.770 12.260 121.050 ;
        RECT 11.660 120.630 12.260 120.770 ;
        RECT 11.140 120.030 11.400 120.350 ;
        RECT 11.200 119.330 11.340 120.030 ;
        RECT 11.140 119.010 11.400 119.330 ;
        RECT 1.940 118.330 2.200 118.650 ;
        RECT 9.580 116.775 11.460 117.145 ;
        RECT 11.660 113.210 11.800 120.630 ;
        RECT 12.580 119.330 12.720 123.430 ;
        RECT 17.180 121.370 17.320 123.430 ;
        RECT 18.560 121.370 18.700 123.770 ;
        RECT 20.400 122.050 20.540 125.470 ;
        RECT 23.620 124.170 23.760 139.870 ;
        RECT 24.580 130.375 26.460 130.745 ;
        RECT 31.440 126.470 31.580 140.350 ;
        RECT 34.600 129.550 34.860 129.870 ;
        RECT 35.980 129.550 36.240 129.870 ;
        RECT 31.840 128.870 32.100 129.190 ;
        RECT 31.900 126.810 32.040 128.870 ;
        RECT 31.840 126.490 32.100 126.810 ;
        RECT 30.000 126.150 30.260 126.470 ;
        RECT 31.380 126.150 31.640 126.470 ;
        RECT 33.680 126.150 33.940 126.470 ;
        RECT 27.700 125.470 27.960 125.790 ;
        RECT 24.580 124.935 26.460 125.305 ;
        RECT 23.620 124.030 24.220 124.170 ;
        RECT 24.080 123.750 24.220 124.030 ;
        RECT 26.320 123.770 26.580 124.090 ;
        RECT 23.560 123.430 23.820 123.750 ;
        RECT 24.020 123.430 24.280 123.750 ;
        RECT 23.620 122.050 23.760 123.430 ;
        RECT 26.380 122.050 26.520 123.770 ;
        RECT 27.760 122.050 27.900 125.470 ;
        RECT 30.060 124.090 30.200 126.150 ;
        RECT 33.740 124.430 33.880 126.150 ;
        RECT 33.680 124.110 33.940 124.430 ;
        RECT 30.000 123.770 30.260 124.090 ;
        RECT 30.920 123.770 31.180 124.090 ;
        RECT 20.340 121.730 20.600 122.050 ;
        RECT 23.560 121.730 23.820 122.050 ;
        RECT 26.320 121.730 26.580 122.050 ;
        RECT 27.700 121.730 27.960 122.050 ;
        RECT 30.980 121.370 31.120 123.770 ;
        RECT 34.660 122.050 34.800 129.550 ;
        RECT 35.060 125.810 35.320 126.130 ;
        RECT 35.120 122.050 35.260 125.810 ;
        RECT 36.040 124.090 36.180 129.550 ;
        RECT 36.500 129.190 36.640 139.870 ;
        RECT 36.440 128.870 36.700 129.190 ;
        RECT 39.580 127.655 41.460 128.025 ;
        RECT 42.940 126.810 43.080 139.870 ;
        RECT 42.880 126.490 43.140 126.810 ;
        RECT 48.400 126.490 48.660 126.810 ;
        RECT 40.580 126.150 40.840 126.470 ;
        RECT 46.560 126.150 46.820 126.470 ;
        RECT 40.640 124.090 40.780 126.150 ;
        RECT 35.980 123.770 36.240 124.090 ;
        RECT 40.580 123.770 40.840 124.090 ;
        RECT 46.620 123.750 46.760 126.150 ;
        RECT 48.460 124.850 48.600 126.490 ;
        RECT 49.320 125.470 49.580 125.790 ;
        RECT 48.000 124.770 49.060 124.850 ;
        RECT 47.940 124.710 49.060 124.770 ;
        RECT 47.940 124.450 48.200 124.710 ;
        RECT 45.640 123.430 45.900 123.750 ;
        RECT 46.560 123.430 46.820 123.750 ;
        RECT 39.580 122.215 41.460 122.585 ;
        RECT 45.700 122.050 45.840 123.430 ;
        RECT 46.620 123.070 46.760 123.430 ;
        RECT 46.560 122.750 46.820 123.070 ;
        RECT 34.600 121.730 34.860 122.050 ;
        RECT 35.060 121.730 35.320 122.050 ;
        RECT 45.640 121.730 45.900 122.050 ;
        RECT 17.120 121.050 17.380 121.370 ;
        RECT 18.500 121.050 18.760 121.370 ;
        RECT 30.920 121.050 31.180 121.370 ;
        RECT 13.440 120.370 13.700 120.690 ;
        RECT 13.500 119.330 13.640 120.370 ;
        RECT 12.520 119.010 12.780 119.330 ;
        RECT 13.440 119.010 13.700 119.330 ;
        RECT 18.560 118.650 18.700 121.050 ;
        RECT 22.180 120.710 22.440 121.030 ;
        RECT 28.620 120.710 28.880 121.030 ;
        RECT 35.520 120.710 35.780 121.030 ;
        RECT 46.560 120.710 46.820 121.030 ;
        RECT 12.060 118.330 12.320 118.650 ;
        RECT 18.500 118.330 18.760 118.650 ;
        RECT 11.600 112.890 11.860 113.210 ;
        RECT 9.580 111.335 11.460 111.705 ;
        RECT 8.840 106.430 9.100 106.750 ;
        RECT 8.900 104.710 9.040 106.430 ;
        RECT 9.580 105.895 11.460 106.265 ;
        RECT 11.660 105.050 11.800 112.890 ;
        RECT 11.600 104.730 11.860 105.050 ;
        RECT 8.840 104.390 9.100 104.710 ;
        RECT 11.660 102.330 11.800 104.730 ;
        RECT 11.600 102.010 11.860 102.330 ;
        RECT 9.580 100.455 11.460 100.825 ;
        RECT 9.580 95.015 11.460 95.385 ;
        RECT 11.660 94.170 11.800 102.010 ;
        RECT 12.120 101.050 12.260 118.330 ;
        RECT 16.200 115.270 16.460 115.590 ;
        RECT 13.440 114.590 13.700 114.910 ;
        RECT 13.500 112.870 13.640 114.590 ;
        RECT 13.440 112.550 13.700 112.870 ;
        RECT 16.260 111.170 16.400 115.270 ;
        RECT 17.120 113.230 17.380 113.550 ;
        RECT 16.200 110.850 16.460 111.170 ;
        RECT 17.180 110.490 17.320 113.230 ;
        RECT 21.720 111.870 21.980 112.190 ;
        RECT 17.120 110.170 17.380 110.490 ;
        RECT 20.800 110.170 21.060 110.490 ;
        RECT 16.200 109.830 16.460 110.150 ;
        RECT 20.860 109.890 21.000 110.170 ;
        RECT 16.260 107.770 16.400 109.830 ;
        RECT 20.860 109.750 21.460 109.890 ;
        RECT 12.980 107.450 13.240 107.770 ;
        RECT 16.200 107.450 16.460 107.770 ;
        RECT 18.500 107.450 18.760 107.770 ;
        RECT 20.800 107.450 21.060 107.770 ;
        RECT 12.520 106.430 12.780 106.750 ;
        RECT 12.580 102.330 12.720 106.430 ;
        RECT 13.040 105.730 13.180 107.450 ;
        RECT 15.740 106.430 16.000 106.750 ;
        RECT 12.980 105.410 13.240 105.730 ;
        RECT 14.820 104.050 15.080 104.370 ;
        RECT 12.520 102.010 12.780 102.330 ;
        RECT 12.120 100.910 12.720 101.050 ;
        RECT 12.060 95.550 12.320 95.870 ;
        RECT 7.460 93.850 7.720 94.170 ;
        RECT 11.600 93.850 11.860 94.170 ;
        RECT 7.520 91.450 7.660 93.850 ;
        RECT 11.140 93.570 11.400 93.830 ;
        RECT 12.120 93.570 12.260 95.550 ;
        RECT 11.140 93.510 12.260 93.570 ;
        RECT 11.200 93.430 12.260 93.510 ;
        RECT 7.460 91.130 7.720 91.450 ;
        RECT 8.840 90.790 9.100 91.110 ;
        RECT 8.900 89.410 9.040 90.790 ;
        RECT 9.580 89.575 11.460 89.945 ;
        RECT 8.840 89.090 9.100 89.410 ;
        RECT 9.580 84.135 11.460 84.505 ;
        RECT 8.380 79.570 8.640 79.890 ;
        RECT 7.460 77.190 7.720 77.510 ;
        RECT 7.520 75.130 7.660 77.190 ;
        RECT 8.440 75.810 8.580 79.570 ;
        RECT 12.580 79.550 12.720 100.910 ;
        RECT 14.880 100.290 15.020 104.050 ;
        RECT 15.800 102.670 15.940 106.430 ;
        RECT 15.740 102.350 16.000 102.670 ;
        RECT 14.820 99.970 15.080 100.290 ;
        RECT 16.260 99.270 16.400 107.450 ;
        RECT 18.560 103.010 18.700 107.450 ;
        RECT 20.860 104.030 21.000 107.450 ;
        RECT 21.320 107.430 21.460 109.750 ;
        RECT 21.780 109.470 21.920 111.870 ;
        RECT 21.720 109.150 21.980 109.470 ;
        RECT 21.260 107.110 21.520 107.430 ;
        RECT 21.320 105.730 21.460 107.110 ;
        RECT 21.260 105.410 21.520 105.730 ;
        RECT 21.780 104.030 21.920 109.150 ;
        RECT 20.800 103.710 21.060 104.030 ;
        RECT 21.720 103.710 21.980 104.030 ;
        RECT 18.500 102.690 18.760 103.010 ;
        RECT 16.200 98.950 16.460 99.270 ;
        RECT 12.980 91.470 13.240 91.790 ;
        RECT 13.040 89.410 13.180 91.470 ;
        RECT 12.980 89.090 13.240 89.410 ;
        RECT 15.740 87.390 16.000 87.710 ;
        RECT 15.800 82.610 15.940 87.390 ;
        RECT 15.740 82.290 16.000 82.610 ;
        RECT 15.800 81.250 15.940 82.290 ;
        RECT 15.740 80.930 16.000 81.250 ;
        RECT 8.840 79.230 9.100 79.550 ;
        RECT 12.520 79.230 12.780 79.550 ;
        RECT 8.900 77.850 9.040 79.230 ;
        RECT 9.580 78.695 11.460 79.065 ;
        RECT 15.800 78.530 15.940 80.930 ;
        RECT 15.740 78.210 16.000 78.530 ;
        RECT 8.840 77.530 9.100 77.850 ;
        RECT 8.380 75.490 8.640 75.810 ;
        RECT 16.260 75.130 16.400 98.950 ;
        RECT 18.560 98.930 18.700 102.690 ;
        RECT 20.860 99.610 21.000 103.710 ;
        RECT 21.780 99.950 21.920 103.710 ;
        RECT 21.720 99.630 21.980 99.950 ;
        RECT 20.800 99.290 21.060 99.610 ;
        RECT 18.500 98.610 18.760 98.930 ;
        RECT 17.120 96.570 17.380 96.890 ;
        RECT 17.180 92.130 17.320 96.570 ;
        RECT 21.720 93.170 21.980 93.490 ;
        RECT 20.800 92.830 21.060 93.150 ;
        RECT 20.860 92.130 21.000 92.830 ;
        RECT 21.780 92.130 21.920 93.170 ;
        RECT 17.120 91.810 17.380 92.130 ;
        RECT 20.800 91.810 21.060 92.130 ;
        RECT 21.720 91.810 21.980 92.130 ;
        RECT 18.960 91.130 19.220 91.450 ;
        RECT 20.340 91.130 20.600 91.450 ;
        RECT 17.120 90.790 17.380 91.110 ;
        RECT 17.180 88.730 17.320 90.790 ;
        RECT 17.120 88.410 17.380 88.730 ;
        RECT 17.180 80.230 17.320 88.410 ;
        RECT 18.040 88.070 18.300 88.390 ;
        RECT 17.120 79.910 17.380 80.230 ;
        RECT 18.100 77.510 18.240 88.070 ;
        RECT 19.020 88.050 19.160 91.130 ;
        RECT 20.400 88.390 20.540 91.130 ;
        RECT 20.860 88.730 21.000 91.810 ;
        RECT 20.800 88.410 21.060 88.730 ;
        RECT 20.340 88.070 20.600 88.390 ;
        RECT 21.720 88.070 21.980 88.390 ;
        RECT 18.960 87.730 19.220 88.050 ;
        RECT 21.780 87.710 21.920 88.070 ;
        RECT 21.720 87.390 21.980 87.710 ;
        RECT 22.240 86.690 22.380 120.710 ;
        RECT 26.780 120.370 27.040 120.690 ;
        RECT 24.580 119.495 26.460 119.865 ;
        RECT 24.580 114.055 26.460 114.425 ;
        RECT 23.560 112.550 23.820 112.870 ;
        RECT 23.620 111.170 23.760 112.550 ;
        RECT 23.560 110.850 23.820 111.170 ;
        RECT 24.580 108.615 26.460 108.985 ;
        RECT 23.560 107.450 23.820 107.770 ;
        RECT 23.620 103.010 23.760 107.450 ;
        RECT 26.840 107.170 26.980 120.370 ;
        RECT 27.240 113.230 27.500 113.550 ;
        RECT 27.300 108.450 27.440 113.230 ;
        RECT 27.700 112.550 27.960 112.870 ;
        RECT 27.760 109.470 27.900 112.550 ;
        RECT 27.700 109.150 27.960 109.470 ;
        RECT 27.240 108.130 27.500 108.450 ;
        RECT 27.760 107.770 27.900 109.150 ;
        RECT 27.700 107.450 27.960 107.770 ;
        RECT 26.840 107.030 27.440 107.170 ;
        RECT 26.780 106.430 27.040 106.750 ;
        RECT 24.020 105.410 24.280 105.730 ;
        RECT 23.560 102.690 23.820 103.010 ;
        RECT 24.080 101.990 24.220 105.410 ;
        RECT 26.840 104.710 26.980 106.430 ;
        RECT 26.780 104.390 27.040 104.710 ;
        RECT 24.580 103.175 26.460 103.545 ;
        RECT 24.020 101.670 24.280 101.990 ;
        RECT 23.560 98.270 23.820 98.590 ;
        RECT 24.020 98.270 24.280 98.590 ;
        RECT 26.780 98.270 27.040 98.590 ;
        RECT 22.630 90.595 22.910 90.965 ;
        RECT 22.180 86.370 22.440 86.690 ;
        RECT 22.180 85.350 22.440 85.670 ;
        RECT 20.800 82.690 21.060 82.950 ;
        RECT 20.400 82.630 21.060 82.690 ;
        RECT 20.400 82.550 21.000 82.630 ;
        RECT 18.960 80.590 19.220 80.910 ;
        RECT 19.020 78.530 19.160 80.590 ;
        RECT 20.400 80.570 20.540 82.550 ;
        RECT 20.800 81.950 21.060 82.270 ;
        RECT 20.860 80.910 21.000 81.950 ;
        RECT 20.800 80.590 21.060 80.910 ;
        RECT 20.340 80.250 20.600 80.570 ;
        RECT 21.720 80.250 21.980 80.570 ;
        RECT 18.960 78.210 19.220 78.530 ;
        RECT 21.780 77.510 21.920 80.250 ;
        RECT 18.040 77.420 18.300 77.510 ;
        RECT 17.640 77.280 18.300 77.420 ;
        RECT 7.460 74.810 7.720 75.130 ;
        RECT 16.200 74.810 16.460 75.130 ;
        RECT 7.520 63.910 7.660 74.810 ;
        RECT 16.200 74.130 16.460 74.450 ;
        RECT 9.580 73.255 11.460 73.625 ;
        RECT 13.900 69.370 14.160 69.690 ;
        RECT 9.580 67.815 11.460 68.185 ;
        RECT 11.140 65.970 11.400 66.290 ;
        RECT 10.680 65.630 10.940 65.950 ;
        RECT 10.740 64.250 10.880 65.630 ;
        RECT 11.200 64.250 11.340 65.970 ;
        RECT 10.680 63.930 10.940 64.250 ;
        RECT 11.140 63.930 11.400 64.250 ;
        RECT 7.460 63.590 7.720 63.910 ;
        RECT 7.520 61.530 7.660 63.590 ;
        RECT 8.840 62.910 9.100 63.230 ;
        RECT 8.900 62.210 9.040 62.910 ;
        RECT 9.580 62.375 11.460 62.745 ;
        RECT 8.840 61.890 9.100 62.210 ;
        RECT 7.460 61.210 7.720 61.530 ;
        RECT 7.520 56.090 7.660 61.210 ;
        RECT 12.520 60.530 12.780 60.850 ;
        RECT 12.580 59.490 12.720 60.530 ;
        RECT 12.520 59.170 12.780 59.490 ;
        RECT 11.600 57.470 11.860 57.790 ;
        RECT 9.580 56.935 11.460 57.305 ;
        RECT 11.660 56.090 11.800 57.470 ;
        RECT 7.460 55.770 7.720 56.090 ;
        RECT 11.600 55.770 11.860 56.090 ;
        RECT 5.620 53.050 5.880 53.370 ;
        RECT 5.680 52.205 5.820 53.050 ;
        RECT 5.610 51.835 5.890 52.205 ;
        RECT 7.520 47.930 7.660 55.770 ;
        RECT 13.960 53.710 14.100 69.370 ;
        RECT 16.260 66.630 16.400 74.130 ;
        RECT 17.640 70.030 17.780 77.280 ;
        RECT 18.040 77.190 18.300 77.280 ;
        RECT 21.720 77.190 21.980 77.510 ;
        RECT 21.780 75.810 21.920 77.190 ;
        RECT 21.720 75.490 21.980 75.810 ;
        RECT 19.880 74.810 20.140 75.130 ;
        RECT 20.340 74.810 20.600 75.130 ;
        RECT 18.040 71.410 18.300 71.730 ;
        RECT 17.580 69.710 17.840 70.030 ;
        RECT 16.200 66.310 16.460 66.630 ;
        RECT 17.580 66.370 17.840 66.630 ;
        RECT 17.180 66.310 17.840 66.370 ;
        RECT 15.280 58.490 15.540 58.810 ;
        RECT 14.820 55.090 15.080 55.410 ;
        RECT 14.880 54.050 15.020 55.090 ;
        RECT 14.820 53.730 15.080 54.050 ;
        RECT 13.900 53.390 14.160 53.710 ;
        RECT 15.340 53.370 15.480 58.490 ;
        RECT 16.260 56.770 16.400 66.310 ;
        RECT 17.180 66.230 17.780 66.310 ;
        RECT 17.180 65.950 17.320 66.230 ;
        RECT 17.120 65.630 17.380 65.950 ;
        RECT 17.180 59.490 17.320 65.630 ;
        RECT 18.100 62.170 18.240 71.410 ;
        RECT 19.940 69.690 20.080 74.810 ;
        RECT 20.400 74.110 20.540 74.810 ;
        RECT 20.340 73.790 20.600 74.110 ;
        RECT 20.400 72.070 20.540 73.790 ;
        RECT 20.340 71.750 20.600 72.070 ;
        RECT 20.800 71.070 21.060 71.390 ;
        RECT 19.880 69.370 20.140 69.690 ;
        RECT 19.940 62.210 20.080 69.370 ;
        RECT 20.340 66.650 20.600 66.970 ;
        RECT 17.640 62.030 18.240 62.170 ;
        RECT 17.640 60.510 17.780 62.030 ;
        RECT 19.880 61.890 20.140 62.210 ;
        RECT 20.400 61.530 20.540 66.650 ;
        RECT 20.340 61.210 20.600 61.530 ;
        RECT 20.860 60.850 21.000 71.070 ;
        RECT 21.260 64.270 21.520 64.590 ;
        RECT 20.800 60.530 21.060 60.850 ;
        RECT 17.580 60.190 17.840 60.510 ;
        RECT 18.960 60.190 19.220 60.510 ;
        RECT 17.120 59.170 17.380 59.490 ;
        RECT 17.640 58.470 17.780 60.190 ;
        RECT 19.020 58.810 19.160 60.190 ;
        RECT 21.320 59.490 21.460 64.270 ;
        RECT 21.260 59.170 21.520 59.490 ;
        RECT 18.960 58.490 19.220 58.810 ;
        RECT 17.580 58.150 17.840 58.470 ;
        RECT 16.200 56.450 16.460 56.770 ;
        RECT 22.240 56.430 22.380 85.350 ;
        RECT 22.700 69.770 22.840 90.595 ;
        RECT 23.100 87.390 23.360 87.710 ;
        RECT 23.160 83.630 23.300 87.390 ;
        RECT 23.620 84.990 23.760 98.270 ;
        RECT 24.080 92.130 24.220 98.270 ;
        RECT 24.580 97.735 26.460 98.105 ;
        RECT 24.580 92.295 26.460 92.665 ;
        RECT 24.020 91.810 24.280 92.130 ;
        RECT 25.400 91.810 25.660 92.130 ;
        RECT 24.480 91.130 24.740 91.450 ;
        RECT 24.540 89.410 24.680 91.130 ;
        RECT 24.940 90.965 25.200 91.110 ;
        RECT 24.930 90.595 25.210 90.965 ;
        RECT 25.460 90.770 25.600 91.810 ;
        RECT 25.400 90.450 25.660 90.770 ;
        RECT 26.320 90.450 26.580 90.770 ;
        RECT 24.940 90.170 25.200 90.430 ;
        RECT 26.380 90.170 26.520 90.450 ;
        RECT 24.940 90.110 26.520 90.170 ;
        RECT 25.000 90.030 26.520 90.110 ;
        RECT 24.480 89.090 24.740 89.410 ;
        RECT 24.020 88.070 24.280 88.390 ;
        RECT 25.860 88.070 26.120 88.390 ;
        RECT 24.080 86.600 24.220 88.070 ;
        RECT 25.920 87.710 26.060 88.070 ;
        RECT 25.860 87.390 26.120 87.710 ;
        RECT 24.580 86.855 26.460 87.225 ;
        RECT 24.080 86.460 24.680 86.600 ;
        RECT 24.020 85.690 24.280 86.010 ;
        RECT 23.560 84.670 23.820 84.990 ;
        RECT 23.100 83.310 23.360 83.630 ;
        RECT 23.160 82.950 23.300 83.310 ;
        RECT 23.100 82.630 23.360 82.950 ;
        RECT 23.100 81.950 23.360 82.270 ;
        RECT 23.160 80.570 23.300 81.950 ;
        RECT 23.100 80.250 23.360 80.570 ;
        RECT 23.560 80.250 23.820 80.570 ;
        RECT 23.100 76.510 23.360 76.830 ;
        RECT 23.160 75.470 23.300 76.510 ;
        RECT 23.620 75.810 23.760 80.250 ;
        RECT 23.560 75.490 23.820 75.810 ;
        RECT 23.100 75.150 23.360 75.470 ;
        RECT 23.100 74.470 23.360 74.790 ;
        RECT 23.160 72.410 23.300 74.470 ;
        RECT 23.560 74.130 23.820 74.450 ;
        RECT 23.100 72.090 23.360 72.410 ;
        RECT 23.620 72.070 23.760 74.130 ;
        RECT 24.080 73.090 24.220 85.690 ;
        RECT 24.540 83.630 24.680 86.460 ;
        RECT 25.400 85.690 25.660 86.010 ;
        RECT 25.460 83.970 25.600 85.690 ;
        RECT 25.400 83.650 25.660 83.970 ;
        RECT 24.480 83.310 24.740 83.630 ;
        RECT 24.540 82.610 24.680 83.310 ;
        RECT 24.480 82.290 24.740 82.610 ;
        RECT 24.580 81.415 26.460 81.785 ;
        RECT 26.840 79.550 26.980 98.270 ;
        RECT 27.300 92.130 27.440 107.030 ;
        RECT 27.760 105.050 27.900 107.450 ;
        RECT 27.700 104.730 27.960 105.050 ;
        RECT 27.760 93.830 27.900 104.730 ;
        RECT 28.160 102.690 28.420 103.010 ;
        RECT 28.220 99.610 28.360 102.690 ;
        RECT 28.160 99.290 28.420 99.610 ;
        RECT 27.700 93.510 27.960 93.830 ;
        RECT 27.240 91.810 27.500 92.130 ;
        RECT 27.240 91.130 27.500 91.450 ;
        RECT 27.300 83.370 27.440 91.130 ;
        RECT 27.760 86.690 27.900 93.510 ;
        RECT 28.680 92.130 28.820 120.710 ;
        RECT 31.380 117.990 31.640 118.310 ;
        RECT 29.080 107.450 29.340 107.770 ;
        RECT 30.000 107.450 30.260 107.770 ;
        RECT 29.140 96.890 29.280 107.450 ;
        RECT 29.540 106.430 29.800 106.750 ;
        RECT 29.600 104.370 29.740 106.430 ;
        RECT 29.540 104.050 29.800 104.370 ;
        RECT 30.060 104.030 30.200 107.450 ;
        RECT 30.000 103.710 30.260 104.030 ;
        RECT 30.060 103.010 30.200 103.710 ;
        RECT 30.000 102.690 30.260 103.010 ;
        RECT 31.440 99.010 31.580 117.990 ;
        RECT 34.600 112.550 34.860 112.870 ;
        RECT 32.300 112.210 32.560 112.530 ;
        RECT 31.840 111.870 32.100 112.190 ;
        RECT 31.900 110.150 32.040 111.870 ;
        RECT 32.360 110.830 32.500 112.210 ;
        RECT 32.300 110.510 32.560 110.830 ;
        RECT 31.840 109.830 32.100 110.150 ;
        RECT 32.360 99.610 32.500 110.510 ;
        RECT 33.670 109.635 33.950 110.005 ;
        RECT 33.680 109.490 33.940 109.635 ;
        RECT 34.660 107.430 34.800 112.550 ;
        RECT 34.600 107.110 34.860 107.430 ;
        RECT 34.660 105.390 34.800 107.110 ;
        RECT 34.600 105.070 34.860 105.390 ;
        RECT 32.300 99.290 32.560 99.610 ;
        RECT 31.440 98.870 32.500 99.010 ;
        RECT 30.000 98.270 30.260 98.590 ;
        RECT 31.380 98.270 31.640 98.590 ;
        RECT 29.080 96.570 29.340 96.890 ;
        RECT 28.620 91.810 28.880 92.130 ;
        RECT 29.540 91.130 29.800 91.450 ;
        RECT 28.620 88.070 28.880 88.390 ;
        RECT 27.700 86.370 27.960 86.690 ;
        RECT 28.680 83.970 28.820 88.070 ;
        RECT 29.080 87.730 29.340 88.050 ;
        RECT 28.620 83.650 28.880 83.970 ;
        RECT 27.300 83.230 27.900 83.370 ;
        RECT 27.240 80.250 27.500 80.570 ;
        RECT 26.780 79.230 27.040 79.550 ;
        RECT 24.580 75.975 26.460 76.345 ;
        RECT 25.400 75.490 25.660 75.810 ;
        RECT 24.480 75.150 24.740 75.470 ;
        RECT 24.540 74.790 24.680 75.150 ;
        RECT 25.460 75.130 25.600 75.490 ;
        RECT 24.940 74.810 25.200 75.130 ;
        RECT 25.400 74.810 25.660 75.130 ;
        RECT 24.480 74.470 24.740 74.790 ;
        RECT 24.020 72.770 24.280 73.090 ;
        RECT 24.540 72.750 24.680 74.470 ;
        RECT 24.480 72.430 24.740 72.750 ;
        RECT 23.560 71.750 23.820 72.070 ;
        RECT 24.480 71.980 24.740 72.070 ;
        RECT 24.080 71.840 24.740 71.980 ;
        RECT 22.700 69.630 23.300 69.770 ;
        RECT 22.640 69.030 22.900 69.350 ;
        RECT 22.700 64.250 22.840 69.030 ;
        RECT 22.640 63.930 22.900 64.250 ;
        RECT 22.640 60.190 22.900 60.510 ;
        RECT 22.700 56.770 22.840 60.190 ;
        RECT 22.640 56.450 22.900 56.770 ;
        RECT 22.180 56.110 22.440 56.430 ;
        RECT 23.160 56.170 23.300 69.630 ;
        RECT 24.080 66.970 24.220 71.840 ;
        RECT 24.480 71.750 24.740 71.840 ;
        RECT 25.000 71.390 25.140 74.810 ;
        RECT 25.460 72.070 25.600 74.810 ;
        RECT 25.400 71.750 25.660 72.070 ;
        RECT 24.940 71.070 25.200 71.390 ;
        RECT 24.580 70.535 26.460 70.905 ;
        RECT 24.020 66.650 24.280 66.970 ;
        RECT 24.080 64.840 24.220 66.650 ;
        RECT 26.780 65.630 27.040 65.950 ;
        RECT 24.580 65.095 26.460 65.465 ;
        RECT 26.840 64.930 26.980 65.630 ;
        RECT 23.620 64.700 24.220 64.840 ;
        RECT 23.620 63.570 23.760 64.700 ;
        RECT 26.780 64.610 27.040 64.930 ;
        RECT 24.020 63.930 24.280 64.250 ;
        RECT 23.560 63.250 23.820 63.570 ;
        RECT 24.080 61.190 24.220 63.930 ;
        RECT 24.020 60.870 24.280 61.190 ;
        RECT 24.080 59.490 24.220 60.870 ;
        RECT 26.780 60.530 27.040 60.850 ;
        RECT 24.580 59.655 26.460 60.025 ;
        RECT 26.840 59.490 26.980 60.530 ;
        RECT 24.020 59.170 24.280 59.490 ;
        RECT 26.780 59.170 27.040 59.490 ;
        RECT 22.700 56.030 23.300 56.170 ;
        RECT 22.700 54.050 22.840 56.030 ;
        RECT 23.100 55.430 23.360 55.750 ;
        RECT 24.020 55.430 24.280 55.750 ;
        RECT 22.640 53.730 22.900 54.050 ;
        RECT 23.160 53.370 23.300 55.430 ;
        RECT 23.560 55.090 23.820 55.410 ;
        RECT 23.620 53.710 23.760 55.090 ;
        RECT 23.560 53.390 23.820 53.710 ;
        RECT 15.280 53.050 15.540 53.370 ;
        RECT 20.340 53.050 20.600 53.370 ;
        RECT 23.100 53.050 23.360 53.370 ;
        RECT 9.580 51.495 11.460 51.865 ;
        RECT 13.900 49.990 14.160 50.310 ;
        RECT 12.060 49.310 12.320 49.630 ;
        RECT 7.460 47.610 7.720 47.930 ;
        RECT 7.520 45.210 7.660 47.610 ;
        RECT 9.580 46.055 11.460 46.425 ;
        RECT 7.460 44.890 7.720 45.210 ;
        RECT 12.120 44.530 12.260 49.310 ;
        RECT 13.960 45.890 14.100 49.990 ;
        RECT 14.360 49.310 14.620 49.630 ;
        RECT 14.420 48.270 14.560 49.310 ;
        RECT 14.360 47.950 14.620 48.270 ;
        RECT 18.040 47.950 18.300 48.270 ;
        RECT 13.900 45.570 14.160 45.890 ;
        RECT 12.060 44.210 12.320 44.530 ;
        RECT 17.120 44.210 17.380 44.530 ;
        RECT 17.180 42.830 17.320 44.210 ;
        RECT 18.100 43.170 18.240 47.950 ;
        RECT 20.400 45.550 20.540 53.050 ;
        RECT 23.160 52.350 23.300 53.050 ;
        RECT 23.560 52.710 23.820 53.030 ;
        RECT 23.100 52.030 23.360 52.350 ;
        RECT 20.800 49.990 21.060 50.310 ;
        RECT 22.180 49.990 22.440 50.310 ;
        RECT 20.860 48.610 21.000 49.990 ;
        RECT 20.800 48.290 21.060 48.610 ;
        RECT 21.260 47.610 21.520 47.930 ;
        RECT 20.340 45.230 20.600 45.550 ;
        RECT 18.500 44.210 18.760 44.530 ;
        RECT 18.040 42.850 18.300 43.170 ;
        RECT 17.120 42.510 17.380 42.830 ;
        RECT 18.040 42.170 18.300 42.490 ;
        RECT 9.580 40.615 11.460 40.985 ;
        RECT 15.740 36.390 16.000 36.710 ;
        RECT 9.580 35.175 11.460 35.545 ;
        RECT 15.800 35.010 15.940 36.390 ;
        RECT 15.740 34.690 16.000 35.010 ;
        RECT 18.100 31.610 18.240 42.170 ;
        RECT 18.560 36.030 18.700 44.210 ;
        RECT 20.400 42.490 20.540 45.230 ;
        RECT 21.320 44.190 21.460 47.610 ;
        RECT 22.240 47.590 22.380 49.990 ;
        RECT 23.100 49.310 23.360 49.630 ;
        RECT 23.160 48.610 23.300 49.310 ;
        RECT 23.100 48.290 23.360 48.610 ;
        RECT 22.180 47.270 22.440 47.590 ;
        RECT 23.100 47.270 23.360 47.590 ;
        RECT 23.160 45.210 23.300 47.270 ;
        RECT 23.100 44.890 23.360 45.210 ;
        RECT 20.800 43.870 21.060 44.190 ;
        RECT 21.260 43.870 21.520 44.190 ;
        RECT 20.860 43.170 21.000 43.870 ;
        RECT 20.800 42.850 21.060 43.170 ;
        RECT 21.320 42.830 21.460 43.870 ;
        RECT 21.260 42.510 21.520 42.830 ;
        RECT 20.340 42.170 20.600 42.490 ;
        RECT 20.800 37.070 21.060 37.390 ;
        RECT 18.500 35.710 18.760 36.030 ;
        RECT 18.560 33.990 18.700 35.710 ;
        RECT 18.500 33.670 18.760 33.990 ;
        RECT 18.560 31.610 18.700 33.670 ;
        RECT 18.040 31.290 18.300 31.610 ;
        RECT 18.500 31.290 18.760 31.610 ;
        RECT 20.860 30.590 21.000 37.070 ;
        RECT 22.640 36.390 22.900 36.710 ;
        RECT 22.700 34.330 22.840 36.390 ;
        RECT 22.640 34.010 22.900 34.330 ;
        RECT 23.620 30.590 23.760 52.710 ;
        RECT 24.080 42.150 24.220 55.430 ;
        RECT 24.580 54.215 26.460 54.585 ;
        RECT 27.300 54.050 27.440 80.250 ;
        RECT 27.760 73.090 27.900 83.230 ;
        RECT 28.160 83.200 28.420 83.290 ;
        RECT 29.140 83.200 29.280 87.730 ;
        RECT 28.160 83.060 29.280 83.200 ;
        RECT 28.160 82.970 28.420 83.060 ;
        RECT 28.620 81.950 28.880 82.270 ;
        RECT 28.680 81.250 28.820 81.950 ;
        RECT 28.620 80.930 28.880 81.250 ;
        RECT 28.620 80.250 28.880 80.570 ;
        RECT 28.680 75.810 28.820 80.250 ;
        RECT 29.080 79.910 29.340 80.230 ;
        RECT 28.620 75.490 28.880 75.810 ;
        RECT 28.620 74.810 28.880 75.130 ;
        RECT 27.700 72.770 27.960 73.090 ;
        RECT 28.160 66.310 28.420 66.630 ;
        RECT 28.220 64.930 28.360 66.310 ;
        RECT 28.160 64.610 28.420 64.930 ;
        RECT 28.680 64.590 28.820 74.810 ;
        RECT 28.620 64.270 28.880 64.590 ;
        RECT 28.620 62.910 28.880 63.230 ;
        RECT 28.680 61.530 28.820 62.910 ;
        RECT 28.620 61.210 28.880 61.530 ;
        RECT 28.620 55.430 28.880 55.750 ;
        RECT 27.240 53.730 27.500 54.050 ;
        RECT 28.680 53.370 28.820 55.430 ;
        RECT 29.140 54.050 29.280 79.910 ;
        RECT 29.600 75.810 29.740 91.130 ;
        RECT 30.060 90.430 30.200 98.270 ;
        RECT 30.920 91.130 31.180 91.450 ;
        RECT 30.460 90.790 30.720 91.110 ;
        RECT 30.000 90.110 30.260 90.430 ;
        RECT 29.540 75.490 29.800 75.810 ;
        RECT 30.000 69.370 30.260 69.690 ;
        RECT 30.060 67.650 30.200 69.370 ;
        RECT 30.000 67.330 30.260 67.650 ;
        RECT 29.540 65.630 29.800 65.950 ;
        RECT 29.600 64.250 29.740 65.630 ;
        RECT 29.540 63.930 29.800 64.250 ;
        RECT 29.080 53.730 29.340 54.050 ;
        RECT 27.240 53.050 27.500 53.370 ;
        RECT 27.700 53.050 27.960 53.370 ;
        RECT 28.620 53.050 28.880 53.370 ;
        RECT 25.860 52.710 26.120 53.030 ;
        RECT 25.920 52.350 26.060 52.710 ;
        RECT 25.860 52.030 26.120 52.350 ;
        RECT 25.920 50.310 26.060 52.030 ;
        RECT 27.300 50.310 27.440 53.050 ;
        RECT 25.860 49.990 26.120 50.310 ;
        RECT 27.240 49.990 27.500 50.310 ;
        RECT 24.580 48.775 26.460 49.145 ;
        RECT 26.780 47.270 27.040 47.590 ;
        RECT 24.580 43.335 26.460 43.705 ;
        RECT 24.020 41.830 24.280 42.150 ;
        RECT 24.080 37.730 24.220 41.830 ;
        RECT 26.840 41.810 26.980 47.270 ;
        RECT 26.780 41.490 27.040 41.810 ;
        RECT 27.760 39.770 27.900 53.050 ;
        RECT 28.680 52.350 28.820 53.050 ;
        RECT 28.620 52.030 28.880 52.350 ;
        RECT 28.680 50.310 28.820 52.030 ;
        RECT 30.520 51.330 30.660 90.790 ;
        RECT 30.980 89.410 31.120 91.130 ;
        RECT 30.920 89.090 31.180 89.410 ;
        RECT 30.920 81.950 31.180 82.270 ;
        RECT 30.980 80.910 31.120 81.950 ;
        RECT 30.920 80.590 31.180 80.910 ;
        RECT 31.440 79.550 31.580 98.270 ;
        RECT 31.840 92.830 32.100 93.150 ;
        RECT 31.900 92.130 32.040 92.830 ;
        RECT 31.840 91.810 32.100 92.130 ;
        RECT 32.360 79.890 32.500 98.870 ;
        RECT 33.220 95.550 33.480 95.870 ;
        RECT 33.280 93.490 33.420 95.550 ;
        RECT 35.580 93.570 35.720 120.710 ;
        RECT 39.580 116.775 41.460 117.145 ;
        RECT 36.900 112.890 37.160 113.210 ;
        RECT 41.040 112.890 41.300 113.210 ;
        RECT 35.980 111.870 36.240 112.190 ;
        RECT 36.040 110.150 36.180 111.870 ;
        RECT 35.980 109.830 36.240 110.150 ;
        RECT 36.440 109.150 36.700 109.470 ;
        RECT 36.500 107.770 36.640 109.150 ;
        RECT 36.960 108.450 37.100 112.890 ;
        RECT 38.740 112.210 39.000 112.530 ;
        RECT 38.800 109.810 38.940 112.210 ;
        RECT 41.100 112.190 41.240 112.890 ;
        RECT 41.960 112.550 42.220 112.870 ;
        RECT 39.200 111.870 39.460 112.190 ;
        RECT 41.040 111.870 41.300 112.190 ;
        RECT 38.740 109.490 39.000 109.810 ;
        RECT 36.900 108.130 37.160 108.450 ;
        RECT 36.440 107.450 36.700 107.770 ;
        RECT 36.500 105.050 36.640 107.450 ;
        RECT 39.260 107.430 39.400 111.870 ;
        RECT 39.580 111.335 41.460 111.705 ;
        RECT 39.200 107.110 39.460 107.430 ;
        RECT 39.580 105.895 41.460 106.265 ;
        RECT 42.020 105.730 42.160 112.550 ;
        RECT 44.720 107.110 44.980 107.430 ;
        RECT 41.960 105.410 42.220 105.730 ;
        RECT 36.440 104.730 36.700 105.050 ;
        RECT 36.500 99.610 36.640 104.730 ;
        RECT 43.340 102.010 43.600 102.330 ;
        RECT 39.580 100.455 41.460 100.825 ;
        RECT 36.440 99.290 36.700 99.610 ;
        RECT 41.500 99.290 41.760 99.610 ;
        RECT 38.740 98.950 39.000 99.270 ;
        RECT 38.280 98.270 38.540 98.590 ;
        RECT 33.220 93.170 33.480 93.490 ;
        RECT 35.580 93.430 36.180 93.570 ;
        RECT 35.520 92.830 35.780 93.150 ;
        RECT 35.580 92.130 35.720 92.830 ;
        RECT 34.600 91.810 34.860 92.130 ;
        RECT 35.520 91.810 35.780 92.130 ;
        RECT 34.660 88.390 34.800 91.810 ;
        RECT 36.040 89.070 36.180 93.430 ;
        RECT 38.340 89.410 38.480 98.270 ;
        RECT 38.800 94.850 38.940 98.950 ;
        RECT 39.200 98.270 39.460 98.590 ;
        RECT 39.260 96.890 39.400 98.270 ;
        RECT 41.560 97.570 41.700 99.290 ;
        RECT 41.500 97.250 41.760 97.570 ;
        RECT 42.880 96.910 43.140 97.230 ;
        RECT 39.200 96.570 39.460 96.890 ;
        RECT 41.960 95.550 42.220 95.870 ;
        RECT 39.580 95.015 41.460 95.385 ;
        RECT 38.740 94.530 39.000 94.850 ;
        RECT 39.200 93.850 39.460 94.170 ;
        RECT 39.260 90.770 39.400 93.850 ;
        RECT 42.020 93.830 42.160 95.550 ;
        RECT 42.940 94.850 43.080 96.910 ;
        RECT 43.400 96.550 43.540 102.010 ;
        RECT 44.780 99.610 44.920 107.110 ;
        RECT 44.720 99.290 44.980 99.610 ;
        RECT 43.340 96.230 43.600 96.550 ;
        RECT 42.880 94.530 43.140 94.850 ;
        RECT 43.400 93.830 43.540 96.230 ;
        RECT 41.960 93.510 42.220 93.830 ;
        RECT 43.340 93.510 43.600 93.830 ;
        RECT 39.200 90.450 39.460 90.770 ;
        RECT 38.280 89.090 38.540 89.410 ;
        RECT 35.980 88.750 36.240 89.070 ;
        RECT 36.440 88.410 36.700 88.730 ;
        RECT 33.680 88.070 33.940 88.390 ;
        RECT 34.600 88.070 34.860 88.390 ;
        RECT 35.520 88.070 35.780 88.390 ;
        RECT 33.740 87.710 33.880 88.070 ;
        RECT 33.680 87.390 33.940 87.710 ;
        RECT 32.760 86.370 33.020 86.690 ;
        RECT 32.820 83.290 32.960 86.370 ;
        RECT 33.740 85.670 33.880 87.390 ;
        RECT 33.680 85.350 33.940 85.670 ;
        RECT 35.060 83.880 35.320 83.970 ;
        RECT 35.580 83.880 35.720 88.070 ;
        RECT 35.060 83.740 35.720 83.880 ;
        RECT 35.060 83.650 35.320 83.740 ;
        RECT 32.760 82.970 33.020 83.290 ;
        RECT 34.600 82.970 34.860 83.290 ;
        RECT 34.660 81.250 34.800 82.970 ;
        RECT 34.600 80.930 34.860 81.250 ;
        RECT 32.300 79.570 32.560 79.890 ;
        RECT 35.580 79.550 35.720 83.740 ;
        RECT 31.380 79.230 31.640 79.550 ;
        RECT 35.520 79.230 35.780 79.550 ;
        RECT 34.600 76.510 34.860 76.830 ;
        RECT 34.660 75.130 34.800 76.510 ;
        RECT 35.980 75.490 36.240 75.810 ;
        RECT 36.040 75.130 36.180 75.490 ;
        RECT 34.600 74.810 34.860 75.130 ;
        RECT 35.060 74.810 35.320 75.130 ;
        RECT 35.980 74.810 36.240 75.130 ;
        RECT 30.920 74.470 31.180 74.790 ;
        RECT 30.980 72.070 31.120 74.470 ;
        RECT 34.660 74.450 34.800 74.810 ;
        RECT 34.600 74.130 34.860 74.450 ;
        RECT 33.220 73.790 33.480 74.110 ;
        RECT 33.280 72.070 33.420 73.790 ;
        RECT 30.920 71.750 31.180 72.070 ;
        RECT 33.220 71.750 33.480 72.070 ;
        RECT 35.120 69.350 35.260 74.810 ;
        RECT 36.040 74.645 36.180 74.810 ;
        RECT 35.970 74.275 36.250 74.645 ;
        RECT 35.980 70.050 36.240 70.370 ;
        RECT 35.520 69.710 35.780 70.030 ;
        RECT 35.060 69.030 35.320 69.350 ;
        RECT 35.120 66.630 35.260 69.030 ;
        RECT 35.580 67.650 35.720 69.710 ;
        RECT 35.520 67.330 35.780 67.650 ;
        RECT 36.040 66.630 36.180 70.050 ;
        RECT 35.060 66.310 35.320 66.630 ;
        RECT 35.980 66.310 36.240 66.630 ;
        RECT 33.220 65.630 33.480 65.950 ;
        RECT 33.280 64.930 33.420 65.630 ;
        RECT 33.220 64.610 33.480 64.930 ;
        RECT 32.760 64.270 33.020 64.590 ;
        RECT 32.820 62.210 32.960 64.270 ;
        RECT 32.760 61.890 33.020 62.210 ;
        RECT 34.600 60.870 34.860 61.190 ;
        RECT 34.660 59.150 34.800 60.870 ;
        RECT 30.910 58.635 31.190 59.005 ;
        RECT 34.600 58.890 34.860 59.150 ;
        RECT 34.600 58.830 35.260 58.890 ;
        RECT 34.660 58.750 35.260 58.830 ;
        RECT 30.920 58.490 31.180 58.635 ;
        RECT 34.600 58.150 34.860 58.470 ;
        RECT 34.660 56.770 34.800 58.150 ;
        RECT 34.600 56.450 34.860 56.770 ;
        RECT 35.120 56.090 35.260 58.750 ;
        RECT 35.060 55.770 35.320 56.090 ;
        RECT 36.500 54.050 36.640 88.410 ;
        RECT 38.740 88.070 39.000 88.390 ;
        RECT 38.800 75.810 38.940 88.070 ;
        RECT 39.260 80.230 39.400 90.450 ;
        RECT 39.580 89.575 41.460 89.945 ;
        RECT 41.960 87.390 42.220 87.710 ;
        RECT 39.580 84.135 41.460 84.505 ;
        RECT 42.020 80.910 42.160 87.390 ;
        RECT 43.400 86.010 43.540 93.510 ;
        RECT 44.780 86.010 44.920 99.290 ;
        RECT 46.620 94.850 46.760 120.710 ;
        RECT 48.400 115.270 48.660 115.590 ;
        RECT 47.940 114.590 48.200 114.910 ;
        RECT 48.000 113.550 48.140 114.590 ;
        RECT 47.940 113.230 48.200 113.550 ;
        RECT 48.460 112.190 48.600 115.270 ;
        RECT 48.920 112.870 49.060 124.710 ;
        RECT 49.380 124.430 49.520 125.470 ;
        RECT 49.320 124.110 49.580 124.430 ;
        RECT 49.840 124.090 49.980 140.350 ;
        RECT 54.580 130.375 56.460 130.745 ;
        RECT 57.200 126.470 57.340 140.350 ;
        RECT 62.260 129.190 62.400 139.870 ;
        RECT 62.660 129.550 62.920 129.870 ;
        RECT 57.600 128.870 57.860 129.190 ;
        RECT 58.980 128.870 59.240 129.190 ;
        RECT 62.200 128.870 62.460 129.190 ;
        RECT 57.660 126.810 57.800 128.870 ;
        RECT 57.600 126.490 57.860 126.810 ;
        RECT 57.140 126.150 57.400 126.470 ;
        RECT 50.240 125.810 50.500 126.130 ;
        RECT 56.680 125.810 56.940 126.130 ;
        RECT 50.300 124.770 50.440 125.810 ;
        RECT 54.580 124.935 56.460 125.305 ;
        RECT 50.240 124.450 50.500 124.770 ;
        RECT 49.780 123.770 50.040 124.090 ;
        RECT 53.460 123.770 53.720 124.090 ;
        RECT 53.000 122.750 53.260 123.070 ;
        RECT 52.540 113.570 52.800 113.890 ;
        RECT 48.860 112.550 49.120 112.870 ;
        RECT 50.700 112.550 50.960 112.870 ;
        RECT 48.400 111.870 48.660 112.190 ;
        RECT 47.020 110.170 47.280 110.490 ;
        RECT 48.460 110.470 48.600 111.870 ;
        RECT 48.920 111.170 49.060 112.550 ;
        RECT 48.860 110.850 49.120 111.170 ;
        RECT 48.460 110.330 49.060 110.470 ;
        RECT 47.080 107.430 47.220 110.170 ;
        RECT 48.920 107.770 49.060 110.330 ;
        RECT 50.760 108.450 50.900 112.550 ;
        RECT 50.700 108.130 50.960 108.450 ;
        RECT 52.600 107.770 52.740 113.570 ;
        RECT 48.860 107.450 49.120 107.770 ;
        RECT 52.540 107.450 52.800 107.770 ;
        RECT 47.020 107.110 47.280 107.430 ;
        RECT 48.400 106.430 48.660 106.750 ;
        RECT 48.460 104.710 48.600 106.430 ;
        RECT 52.600 105.390 52.740 107.450 ;
        RECT 52.540 105.070 52.800 105.390 ;
        RECT 48.400 104.390 48.660 104.710 ;
        RECT 48.400 100.990 48.660 101.310 ;
        RECT 47.020 98.950 47.280 99.270 ;
        RECT 47.080 97.570 47.220 98.950 ;
        RECT 48.460 98.930 48.600 100.990 ;
        RECT 48.400 98.610 48.660 98.930 ;
        RECT 50.700 98.270 50.960 98.590 ;
        RECT 50.760 97.570 50.900 98.270 ;
        RECT 47.020 97.250 47.280 97.570 ;
        RECT 50.700 97.250 50.960 97.570 ;
        RECT 52.080 96.230 52.340 96.550 ;
        RECT 46.560 94.530 46.820 94.850 ;
        RECT 52.140 90.770 52.280 96.230 ;
        RECT 52.080 90.450 52.340 90.770 ;
        RECT 52.140 88.730 52.280 90.450 ;
        RECT 47.940 88.410 48.200 88.730 ;
        RECT 52.080 88.410 52.340 88.730 ;
        RECT 47.020 87.390 47.280 87.710 ;
        RECT 47.480 87.390 47.740 87.710 ;
        RECT 47.080 86.010 47.220 87.390 ;
        RECT 43.340 85.690 43.600 86.010 ;
        RECT 44.720 85.690 44.980 86.010 ;
        RECT 47.020 85.690 47.280 86.010 ;
        RECT 41.960 80.590 42.220 80.910 ;
        RECT 43.400 80.570 43.540 85.690 ;
        RECT 44.780 83.290 44.920 85.690 ;
        RECT 47.540 83.290 47.680 87.390 ;
        RECT 48.000 83.290 48.140 88.410 ;
        RECT 52.140 83.630 52.280 88.410 ;
        RECT 52.080 83.310 52.340 83.630 ;
        RECT 43.800 82.970 44.060 83.290 ;
        RECT 44.720 82.970 44.980 83.290 ;
        RECT 47.480 82.970 47.740 83.290 ;
        RECT 47.940 82.970 48.200 83.290 ;
        RECT 43.340 80.250 43.600 80.570 ;
        RECT 39.200 79.910 39.460 80.230 ;
        RECT 39.580 78.695 41.460 79.065 ;
        RECT 38.740 75.490 39.000 75.810 ;
        RECT 43.860 75.130 44.000 82.970 ;
        RECT 48.000 81.250 48.140 82.970 ;
        RECT 53.060 82.610 53.200 122.750 ;
        RECT 53.520 121.370 53.660 123.770 ;
        RECT 56.740 123.750 56.880 125.810 ;
        RECT 59.040 124.770 59.180 128.870 ;
        RECT 62.200 125.810 62.460 126.130 ;
        RECT 58.980 124.450 59.240 124.770 ;
        RECT 57.600 124.000 57.860 124.090 ;
        RECT 57.600 123.860 58.260 124.000 ;
        RECT 57.600 123.770 57.860 123.860 ;
        RECT 56.680 123.430 56.940 123.750 ;
        RECT 53.460 121.050 53.720 121.370 ;
        RECT 54.580 119.495 56.460 119.865 ;
        RECT 57.600 115.270 57.860 115.590 ;
        RECT 56.680 114.590 56.940 114.910 ;
        RECT 54.580 114.055 56.460 114.425 ;
        RECT 56.740 112.870 56.880 114.590 ;
        RECT 53.920 112.550 54.180 112.870 ;
        RECT 56.680 112.550 56.940 112.870 ;
        RECT 53.450 109.635 53.730 110.005 ;
        RECT 53.460 109.490 53.720 109.635 ;
        RECT 53.980 106.750 54.120 112.550 ;
        RECT 56.680 111.870 56.940 112.190 ;
        RECT 54.580 108.615 56.460 108.985 ;
        RECT 56.740 107.770 56.880 111.870 ;
        RECT 57.140 110.170 57.400 110.490 ;
        RECT 57.200 108.450 57.340 110.170 ;
        RECT 57.660 108.450 57.800 115.270 ;
        RECT 57.140 108.130 57.400 108.450 ;
        RECT 57.600 108.130 57.860 108.450 ;
        RECT 56.680 107.450 56.940 107.770 ;
        RECT 55.300 107.110 55.560 107.430 ;
        RECT 53.920 106.430 54.180 106.750 ;
        RECT 53.980 102.330 54.120 106.430 ;
        RECT 55.360 105.050 55.500 107.110 ;
        RECT 55.300 104.730 55.560 105.050 ;
        RECT 54.580 103.175 56.460 103.545 ;
        RECT 53.920 102.010 54.180 102.330 ;
        RECT 56.680 100.990 56.940 101.310 ;
        RECT 57.600 100.990 57.860 101.310 ;
        RECT 56.740 100.290 56.880 100.990 ;
        RECT 56.680 99.970 56.940 100.290 ;
        RECT 53.920 99.290 54.180 99.610 ;
        RECT 53.460 98.950 53.720 99.270 ;
        RECT 53.520 97.570 53.660 98.950 ;
        RECT 53.460 97.250 53.720 97.570 ;
        RECT 53.980 88.810 54.120 99.290 ;
        RECT 57.140 98.950 57.400 99.270 ;
        RECT 56.680 98.270 56.940 98.590 ;
        RECT 54.580 97.735 56.460 98.105 ;
        RECT 56.740 97.570 56.880 98.270 ;
        RECT 56.680 97.250 56.940 97.570 ;
        RECT 56.220 96.570 56.480 96.890 ;
        RECT 56.280 93.150 56.420 96.570 ;
        RECT 56.220 92.830 56.480 93.150 ;
        RECT 54.580 92.295 56.460 92.665 ;
        RECT 53.520 88.670 54.120 88.810 ;
        RECT 48.400 82.290 48.660 82.610 ;
        RECT 53.000 82.290 53.260 82.610 ;
        RECT 48.460 81.250 48.600 82.290 ;
        RECT 47.940 80.930 48.200 81.250 ;
        RECT 48.400 80.930 48.660 81.250 ;
        RECT 52.080 75.150 52.340 75.470 ;
        RECT 43.800 74.810 44.060 75.130 ;
        RECT 47.480 74.810 47.740 75.130 ;
        RECT 39.200 74.470 39.460 74.790 ;
        RECT 39.260 69.010 39.400 74.470 ;
        RECT 47.010 74.275 47.290 74.645 ;
        RECT 39.580 73.255 41.460 73.625 ;
        RECT 47.080 72.410 47.220 74.275 ;
        RECT 44.720 72.090 44.980 72.410 ;
        RECT 47.020 72.090 47.280 72.410 ;
        RECT 39.200 68.690 39.460 69.010 ;
        RECT 39.260 66.970 39.400 68.690 ;
        RECT 39.580 67.815 41.460 68.185 ;
        RECT 39.200 66.650 39.460 66.970 ;
        RECT 39.260 63.910 39.400 66.650 ;
        RECT 44.780 64.250 44.920 72.090 ;
        RECT 47.540 72.070 47.680 74.810 ;
        RECT 49.780 73.790 50.040 74.110 ;
        RECT 47.480 71.750 47.740 72.070 ;
        RECT 47.940 71.750 48.200 72.070 ;
        RECT 47.540 66.630 47.680 71.750 ;
        RECT 48.000 70.370 48.140 71.750 ;
        RECT 49.840 71.730 49.980 73.790 ;
        RECT 52.140 73.090 52.280 75.150 ;
        RECT 52.080 72.770 52.340 73.090 ;
        RECT 49.780 71.410 50.040 71.730 ;
        RECT 52.140 70.370 52.280 72.770 ;
        RECT 52.540 72.430 52.800 72.750 ;
        RECT 52.600 70.370 52.740 72.430 ;
        RECT 47.940 70.050 48.200 70.370 ;
        RECT 52.080 70.050 52.340 70.370 ;
        RECT 52.540 70.050 52.800 70.370 ;
        RECT 51.150 66.795 51.430 67.165 ;
        RECT 47.480 66.310 47.740 66.630 ;
        RECT 49.320 65.970 49.580 66.290 ;
        RECT 45.180 65.630 45.440 65.950 ;
        RECT 48.400 65.630 48.660 65.950 ;
        RECT 45.240 64.930 45.380 65.630 ;
        RECT 45.180 64.610 45.440 64.930 ;
        RECT 48.460 64.250 48.600 65.630 ;
        RECT 44.720 63.930 44.980 64.250 ;
        RECT 48.400 63.930 48.660 64.250 ;
        RECT 39.200 63.590 39.460 63.910 ;
        RECT 44.260 63.590 44.520 63.910 ;
        RECT 39.260 61.530 39.400 63.590 ;
        RECT 41.960 62.910 42.220 63.230 ;
        RECT 39.580 62.375 41.460 62.745 ;
        RECT 39.200 61.210 39.460 61.530 ;
        RECT 42.020 61.190 42.160 62.910 ;
        RECT 41.960 60.870 42.220 61.190 ;
        RECT 36.900 60.190 37.160 60.510 ;
        RECT 36.960 55.750 37.100 60.190 ;
        RECT 44.320 59.490 44.460 63.590 ;
        RECT 44.780 61.190 44.920 63.930 ;
        RECT 44.720 60.870 44.980 61.190 ;
        RECT 47.020 60.870 47.280 61.190 ;
        RECT 44.260 59.170 44.520 59.490 ;
        RECT 38.280 58.830 38.540 59.150 ;
        RECT 38.340 56.770 38.480 58.830 ;
        RECT 44.780 57.790 44.920 60.870 ;
        RECT 47.080 59.490 47.220 60.870 ;
        RECT 49.380 60.850 49.520 65.970 ;
        RECT 50.700 61.550 50.960 61.870 ;
        RECT 49.320 60.530 49.580 60.850 ;
        RECT 47.020 59.170 47.280 59.490 ;
        RECT 48.850 58.635 49.130 59.005 ;
        RECT 41.960 57.470 42.220 57.790 ;
        RECT 44.720 57.470 44.980 57.790 ;
        RECT 39.580 56.935 41.460 57.305 ;
        RECT 38.280 56.450 38.540 56.770 ;
        RECT 42.020 55.750 42.160 57.470 ;
        RECT 48.400 56.450 48.660 56.770 ;
        RECT 47.940 55.770 48.200 56.090 ;
        RECT 36.900 55.430 37.160 55.750 ;
        RECT 38.280 55.430 38.540 55.750 ;
        RECT 41.960 55.430 42.220 55.750 ;
        RECT 42.880 55.430 43.140 55.750 ;
        RECT 35.060 53.730 35.320 54.050 ;
        RECT 36.440 53.730 36.700 54.050 ;
        RECT 31.380 53.620 31.640 53.710 ;
        RECT 32.300 53.620 32.560 53.710 ;
        RECT 31.380 53.480 32.560 53.620 ;
        RECT 31.380 53.390 31.640 53.480 ;
        RECT 32.300 53.390 32.560 53.480 ;
        RECT 35.120 53.370 35.260 53.730 ;
        RECT 33.680 53.050 33.940 53.370 ;
        RECT 35.060 53.050 35.320 53.370 ;
        RECT 30.460 51.010 30.720 51.330 ;
        RECT 28.620 49.990 28.880 50.310 ;
        RECT 32.300 49.990 32.560 50.310 ;
        RECT 29.540 49.310 29.800 49.630 ;
        RECT 29.600 45.210 29.740 49.310 ;
        RECT 32.360 48.610 32.500 49.990 ;
        RECT 32.300 48.290 32.560 48.610 ;
        RECT 33.740 48.270 33.880 53.050 ;
        RECT 36.440 49.310 36.700 49.630 ;
        RECT 33.680 47.950 33.940 48.270 ;
        RECT 33.740 45.890 33.880 47.950 ;
        RECT 34.140 47.270 34.400 47.590 ;
        RECT 33.680 45.570 33.940 45.890 ;
        RECT 29.540 44.890 29.800 45.210 ;
        RECT 32.300 44.210 32.560 44.530 ;
        RECT 32.360 43.170 32.500 44.210 ;
        RECT 34.200 43.170 34.340 47.270 ;
        RECT 36.500 45.210 36.640 49.310 ;
        RECT 36.440 44.890 36.700 45.210 ;
        RECT 38.340 44.870 38.480 55.430 ;
        RECT 42.020 53.710 42.160 55.430 ;
        RECT 41.960 53.390 42.220 53.710 ;
        RECT 39.580 51.495 41.460 51.865 ;
        RECT 41.500 49.650 41.760 49.970 ;
        RECT 38.740 49.310 39.000 49.630 ;
        RECT 38.280 44.550 38.540 44.870 ;
        RECT 32.300 42.850 32.560 43.170 ;
        RECT 34.140 42.850 34.400 43.170 ;
        RECT 38.340 42.830 38.480 44.550 ;
        RECT 38.280 42.510 38.540 42.830 ;
        RECT 38.800 42.490 38.940 49.310 ;
        RECT 41.560 48.610 41.700 49.650 ;
        RECT 41.500 48.290 41.760 48.610 ;
        RECT 42.020 48.370 42.160 53.390 ;
        RECT 42.940 53.370 43.080 55.430 ;
        RECT 47.020 55.090 47.280 55.410 ;
        RECT 42.880 53.050 43.140 53.370 ;
        RECT 43.800 49.310 44.060 49.630 ;
        RECT 39.200 47.950 39.460 48.270 ;
        RECT 42.020 48.230 42.620 48.370 ;
        RECT 43.860 48.270 44.000 49.310 ;
        RECT 39.260 45.890 39.400 47.950 ;
        RECT 42.480 47.250 42.620 48.230 ;
        RECT 43.800 47.950 44.060 48.270 ;
        RECT 42.420 46.930 42.680 47.250 ;
        RECT 44.720 46.590 44.980 46.910 ;
        RECT 39.580 46.055 41.460 46.425 ;
        RECT 39.200 45.570 39.460 45.890 ;
        RECT 43.800 43.870 44.060 44.190 ;
        RECT 39.200 42.510 39.460 42.830 ;
        RECT 38.740 42.170 39.000 42.490 ;
        RECT 32.760 41.490 33.020 41.810 ;
        RECT 27.700 39.450 27.960 39.770 ;
        RECT 24.580 37.895 26.460 38.265 ;
        RECT 24.020 37.410 24.280 37.730 ;
        RECT 24.080 34.670 24.220 37.410 ;
        RECT 26.780 36.730 27.040 37.050 ;
        RECT 24.940 35.710 25.200 36.030 ;
        RECT 24.020 34.350 24.280 34.670 ;
        RECT 25.000 33.990 25.140 35.710 ;
        RECT 24.940 33.670 25.200 33.990 ;
        RECT 26.840 33.650 26.980 36.730 ;
        RECT 27.760 35.010 27.900 39.450 ;
        RECT 32.820 36.710 32.960 41.490 ;
        RECT 33.220 38.430 33.480 38.750 ;
        RECT 38.280 38.430 38.540 38.750 ;
        RECT 33.280 37.730 33.420 38.430 ;
        RECT 33.220 37.410 33.480 37.730 ;
        RECT 38.340 36.710 38.480 38.430 ;
        RECT 32.760 36.390 33.020 36.710 ;
        RECT 38.280 36.390 38.540 36.710 ;
        RECT 35.520 35.710 35.780 36.030 ;
        RECT 27.700 34.690 27.960 35.010 ;
        RECT 26.780 33.330 27.040 33.650 ;
        RECT 32.300 33.330 32.560 33.650 ;
        RECT 34.600 33.330 34.860 33.650 ;
        RECT 24.020 32.990 24.280 33.310 ;
        RECT 24.080 32.290 24.220 32.990 ;
        RECT 24.580 32.455 26.460 32.825 ;
        RECT 26.840 32.290 26.980 33.330 ;
        RECT 32.360 32.290 32.500 33.330 ;
        RECT 34.660 32.290 34.800 33.330 ;
        RECT 24.020 31.970 24.280 32.290 ;
        RECT 26.780 31.970 27.040 32.290 ;
        RECT 32.300 31.970 32.560 32.290 ;
        RECT 34.600 31.970 34.860 32.290 ;
        RECT 35.580 31.610 35.720 35.710 ;
        RECT 39.260 33.990 39.400 42.510 ;
        RECT 43.860 42.490 44.000 43.870 ;
        RECT 43.800 42.170 44.060 42.490 ;
        RECT 39.580 40.615 41.460 40.985 ;
        RECT 44.780 39.770 44.920 46.590 ;
        RECT 46.100 41.150 46.360 41.470 ;
        RECT 44.720 39.450 44.980 39.770 ;
        RECT 40.580 39.110 40.840 39.430 ;
        RECT 40.640 37.730 40.780 39.110 ;
        RECT 40.580 37.410 40.840 37.730 ;
        RECT 41.960 37.070 42.220 37.390 ;
        RECT 39.580 35.175 41.460 35.545 ;
        RECT 42.020 34.330 42.160 37.070 ;
        RECT 44.780 36.710 44.920 39.450 ;
        RECT 46.160 39.430 46.300 41.150 ;
        RECT 46.100 39.110 46.360 39.430 ;
        RECT 47.080 37.050 47.220 55.090 ;
        RECT 47.480 53.050 47.740 53.370 ;
        RECT 47.540 48.610 47.680 53.050 ;
        RECT 48.000 51.330 48.140 55.770 ;
        RECT 48.460 55.750 48.600 56.450 ;
        RECT 48.400 55.430 48.660 55.750 ;
        RECT 48.920 53.710 49.060 58.635 ;
        RECT 50.760 55.750 50.900 61.550 ;
        RECT 50.700 55.430 50.960 55.750 ;
        RECT 48.860 53.390 49.120 53.710 ;
        RECT 47.940 51.010 48.200 51.330 ;
        RECT 47.480 48.290 47.740 48.610 ;
        RECT 47.540 44.870 47.680 48.290 ;
        RECT 48.000 45.210 48.140 51.010 ;
        RECT 50.760 50.310 50.900 55.430 ;
        RECT 51.220 53.030 51.360 66.795 ;
        RECT 52.600 66.630 52.740 70.050 ;
        RECT 52.540 66.310 52.800 66.630 ;
        RECT 52.080 63.250 52.340 63.570 ;
        RECT 52.140 58.810 52.280 63.250 ;
        RECT 52.080 58.490 52.340 58.810 ;
        RECT 51.620 55.430 51.880 55.750 ;
        RECT 51.680 55.070 51.820 55.430 ;
        RECT 51.620 54.750 51.880 55.070 ;
        RECT 53.520 54.050 53.660 88.670 ;
        RECT 56.740 88.390 56.880 97.250 ;
        RECT 56.680 88.070 56.940 88.390 ;
        RECT 53.920 87.730 54.180 88.050 ;
        RECT 53.980 86.690 54.120 87.730 ;
        RECT 54.580 86.855 56.460 87.225 ;
        RECT 53.920 86.370 54.180 86.690 ;
        RECT 55.760 85.690 56.020 86.010 ;
        RECT 55.820 83.290 55.960 85.690 ;
        RECT 55.760 82.970 56.020 83.290 ;
        RECT 56.220 82.970 56.480 83.290 ;
        RECT 56.280 82.690 56.420 82.970 ;
        RECT 56.280 82.550 56.880 82.690 ;
        RECT 54.580 81.415 56.460 81.785 ;
        RECT 54.580 75.975 56.460 76.345 ;
        RECT 53.910 74.955 54.190 75.325 ;
        RECT 53.920 74.810 54.180 74.955 ;
        RECT 53.980 72.070 54.120 74.810 ;
        RECT 53.920 71.750 54.180 72.070 ;
        RECT 54.580 70.535 56.460 70.905 ;
        RECT 55.300 68.690 55.560 69.010 ;
        RECT 55.360 66.970 55.500 68.690 ;
        RECT 55.300 66.650 55.560 66.970 ;
        RECT 54.580 65.095 56.460 65.465 ;
        RECT 54.580 59.655 56.460 60.025 ;
        RECT 54.580 54.215 56.460 54.585 ;
        RECT 53.460 53.730 53.720 54.050 ;
        RECT 51.160 52.710 51.420 53.030 ;
        RECT 53.920 52.710 54.180 53.030 ;
        RECT 52.540 52.370 52.800 52.690 ;
        RECT 52.600 50.310 52.740 52.370 ;
        RECT 53.980 50.310 54.120 52.710 ;
        RECT 56.740 51.330 56.880 82.550 ;
        RECT 57.200 75.810 57.340 98.950 ;
        RECT 57.660 94.850 57.800 100.990 ;
        RECT 57.600 94.530 57.860 94.850 ;
        RECT 57.600 93.510 57.860 93.830 ;
        RECT 57.660 92.210 57.800 93.510 ;
        RECT 58.120 92.890 58.260 123.860 ;
        RECT 62.260 122.050 62.400 125.810 ;
        RECT 62.720 124.090 62.860 129.550 ;
        RECT 68.700 126.810 68.840 139.870 ;
        RECT 69.580 127.655 71.460 128.025 ;
        RECT 68.640 126.490 68.900 126.810 ;
        RECT 67.720 126.150 67.980 126.470 ;
        RECT 62.660 123.770 62.920 124.090 ;
        RECT 67.780 123.750 67.920 126.150 ;
        RECT 68.640 125.810 68.900 126.130 ;
        RECT 67.720 123.430 67.980 123.750 ;
        RECT 62.200 121.730 62.460 122.050 ;
        RECT 58.980 121.390 59.240 121.710 ;
        RECT 58.520 120.710 58.780 121.030 ;
        RECT 58.580 117.970 58.720 120.710 ;
        RECT 58.520 117.650 58.780 117.970 ;
        RECT 59.040 113.800 59.180 121.390 ;
        RECT 63.120 120.030 63.380 120.350 ;
        RECT 61.740 115.270 62.000 115.590 ;
        RECT 61.280 114.590 61.540 114.910 ;
        RECT 58.580 113.660 59.180 113.800 ;
        RECT 58.580 100.290 58.720 113.660 ;
        RECT 61.340 113.550 61.480 114.590 ;
        RECT 61.280 113.230 61.540 113.550 ;
        RECT 58.980 112.890 59.240 113.210 ;
        RECT 59.040 109.470 59.180 112.890 ;
        RECT 60.820 112.210 61.080 112.530 ;
        RECT 59.440 111.870 59.700 112.190 ;
        RECT 58.980 109.150 59.240 109.470 ;
        RECT 59.040 107.430 59.180 109.150 ;
        RECT 59.500 108.450 59.640 111.870 ;
        RECT 59.440 108.130 59.700 108.450 ;
        RECT 58.980 107.110 59.240 107.430 ;
        RECT 59.500 105.050 59.640 108.130 ;
        RECT 60.880 107.430 61.020 112.210 ;
        RECT 61.800 110.490 61.940 115.270 ;
        RECT 61.740 110.170 62.000 110.490 ;
        RECT 59.900 107.110 60.160 107.430 ;
        RECT 60.820 107.110 61.080 107.430 ;
        RECT 59.440 104.730 59.700 105.050 ;
        RECT 58.980 104.390 59.240 104.710 ;
        RECT 59.040 102.330 59.180 104.390 ;
        RECT 59.440 104.050 59.700 104.370 ;
        RECT 58.980 102.010 59.240 102.330 ;
        RECT 58.520 99.970 58.780 100.290 ;
        RECT 58.520 98.270 58.780 98.590 ;
        RECT 58.580 93.570 58.720 98.270 ;
        RECT 59.040 94.510 59.180 102.010 ;
        RECT 58.980 94.190 59.240 94.510 ;
        RECT 58.580 93.430 59.180 93.570 ;
        RECT 59.040 93.150 59.180 93.430 ;
        RECT 58.120 92.750 58.720 92.890 ;
        RECT 58.980 92.830 59.240 93.150 ;
        RECT 57.660 92.070 58.260 92.210 ;
        RECT 58.580 92.130 58.720 92.750 ;
        RECT 57.600 91.130 57.860 91.450 ;
        RECT 57.660 89.410 57.800 91.130 ;
        RECT 57.600 89.090 57.860 89.410 ;
        RECT 57.600 84.670 57.860 84.990 ;
        RECT 57.660 82.950 57.800 84.670 ;
        RECT 57.600 82.630 57.860 82.950 ;
        RECT 58.120 75.810 58.260 92.070 ;
        RECT 58.520 91.810 58.780 92.130 ;
        RECT 58.980 91.130 59.240 91.450 ;
        RECT 58.520 90.790 58.780 91.110 ;
        RECT 58.580 90.285 58.720 90.790 ;
        RECT 58.510 89.915 58.790 90.285 ;
        RECT 58.520 88.070 58.780 88.390 ;
        RECT 58.580 86.350 58.720 88.070 ;
        RECT 58.520 86.030 58.780 86.350 ;
        RECT 57.140 75.490 57.400 75.810 ;
        RECT 58.060 75.490 58.320 75.810 ;
        RECT 58.520 74.810 58.780 75.130 ;
        RECT 58.580 72.070 58.720 74.810 ;
        RECT 59.040 73.090 59.180 91.130 ;
        RECT 59.500 90.430 59.640 104.050 ;
        RECT 59.960 102.330 60.100 107.110 ;
        RECT 60.360 103.710 60.620 104.030 ;
        RECT 59.900 102.010 60.160 102.330 ;
        RECT 60.420 94.930 60.560 103.710 ;
        RECT 60.880 102.670 61.020 107.110 ;
        RECT 61.800 107.090 61.940 110.170 ;
        RECT 61.740 106.770 62.000 107.090 ;
        RECT 60.820 102.350 61.080 102.670 ;
        RECT 61.280 96.910 61.540 97.230 ;
        RECT 60.820 95.550 61.080 95.870 ;
        RECT 59.960 94.790 60.560 94.930 ;
        RECT 59.440 90.110 59.700 90.430 ;
        RECT 59.960 83.970 60.100 94.790 ;
        RECT 60.360 93.850 60.620 94.170 ;
        RECT 59.900 83.650 60.160 83.970 ;
        RECT 59.440 82.290 59.700 82.610 ;
        RECT 59.500 73.090 59.640 82.290 ;
        RECT 59.900 75.490 60.160 75.810 ;
        RECT 58.980 72.770 59.240 73.090 ;
        RECT 59.440 72.770 59.700 73.090 ;
        RECT 59.440 72.090 59.700 72.410 ;
        RECT 58.520 71.750 58.780 72.070 ;
        RECT 57.140 71.070 57.400 71.390 ;
        RECT 57.200 66.630 57.340 71.070 ;
        RECT 59.500 68.670 59.640 72.090 ;
        RECT 59.960 71.730 60.100 75.490 ;
        RECT 59.900 71.410 60.160 71.730 ;
        RECT 59.440 68.350 59.700 68.670 ;
        RECT 57.140 66.310 57.400 66.630 ;
        RECT 57.200 64.930 57.340 66.310 ;
        RECT 57.140 64.610 57.400 64.930 ;
        RECT 59.440 64.610 59.700 64.930 ;
        RECT 59.500 60.510 59.640 64.610 ;
        RECT 59.440 60.190 59.700 60.510 ;
        RECT 59.900 55.770 60.160 56.090 ;
        RECT 57.600 54.750 57.860 55.070 ;
        RECT 57.660 53.370 57.800 54.750 ;
        RECT 59.960 53.370 60.100 55.770 ;
        RECT 57.600 53.050 57.860 53.370 ;
        RECT 59.900 53.050 60.160 53.370 ;
        RECT 56.680 51.010 56.940 51.330 ;
        RECT 57.660 50.310 57.800 53.050 ;
        RECT 60.420 50.990 60.560 93.850 ;
        RECT 60.880 93.830 61.020 95.550 ;
        RECT 60.820 93.510 61.080 93.830 ;
        RECT 60.820 92.830 61.080 93.150 ;
        RECT 60.880 88.390 61.020 92.830 ;
        RECT 61.340 88.730 61.480 96.910 ;
        RECT 61.740 96.570 62.000 96.890 ;
        RECT 61.800 89.070 61.940 96.570 ;
        RECT 63.180 96.550 63.320 120.030 ;
        RECT 67.780 112.870 67.920 123.430 ;
        RECT 68.700 121.710 68.840 125.810 ;
        RECT 75.140 123.750 75.280 139.870 ;
        RECT 81.580 126.810 81.720 139.870 ;
        RECT 84.580 130.375 86.460 130.745 ;
        RECT 88.020 126.810 88.160 139.870 ;
        RECT 81.520 126.490 81.780 126.810 ;
        RECT 87.960 126.490 88.220 126.810 ;
        RECT 86.180 126.130 86.780 126.210 ;
        RECT 76.460 125.810 76.720 126.130 ;
        RECT 80.140 125.810 80.400 126.130 ;
        RECT 86.120 126.070 86.780 126.130 ;
        RECT 86.120 125.810 86.380 126.070 ;
        RECT 69.100 123.430 69.360 123.750 ;
        RECT 75.080 123.430 75.340 123.750 ;
        RECT 69.160 122.050 69.300 123.430 ;
        RECT 69.580 122.215 71.460 122.585 ;
        RECT 76.520 122.050 76.660 125.810 ;
        RECT 80.200 123.750 80.340 125.810 ;
        RECT 84.580 124.935 86.460 125.305 ;
        RECT 82.900 123.770 83.160 124.090 ;
        RECT 80.140 123.430 80.400 123.750 ;
        RECT 69.100 121.730 69.360 122.050 ;
        RECT 76.460 121.730 76.720 122.050 ;
        RECT 68.640 121.390 68.900 121.710 ;
        RECT 82.960 121.370 83.100 123.770 ;
        RECT 86.640 122.050 86.780 126.070 ;
        RECT 90.720 125.810 90.980 126.130 ;
        RECT 87.040 125.470 87.300 125.790 ;
        RECT 87.100 123.750 87.240 125.470 ;
        RECT 87.040 123.430 87.300 123.750 ;
        RECT 88.420 123.430 88.680 123.750 ;
        RECT 86.580 121.730 86.840 122.050 ;
        RECT 82.900 121.050 83.160 121.370 ;
        RECT 68.180 120.710 68.440 121.030 ;
        RECT 75.080 120.710 75.340 121.030 ;
        RECT 76.460 120.710 76.720 121.030 ;
        RECT 81.520 120.710 81.780 121.030 ;
        RECT 65.420 112.550 65.680 112.870 ;
        RECT 67.720 112.550 67.980 112.870 ;
        RECT 65.480 110.490 65.620 112.550 ;
        RECT 65.420 110.170 65.680 110.490 ;
        RECT 64.960 102.010 65.220 102.330 ;
        RECT 63.580 99.630 63.840 99.950 ;
        RECT 63.120 96.230 63.380 96.550 ;
        RECT 63.640 95.870 63.780 99.630 ;
        RECT 65.020 98.930 65.160 102.010 ;
        RECT 64.960 98.610 65.220 98.930 ;
        RECT 65.020 97.570 65.160 98.610 ;
        RECT 64.960 97.250 65.220 97.570 ;
        RECT 64.500 96.570 64.760 96.890 ;
        RECT 64.040 95.890 64.300 96.210 ;
        RECT 63.580 95.550 63.840 95.870 ;
        RECT 63.640 91.790 63.780 95.550 ;
        RECT 63.580 91.470 63.840 91.790 ;
        RECT 61.740 88.750 62.000 89.070 ;
        RECT 61.280 88.410 61.540 88.730 ;
        RECT 60.820 88.070 61.080 88.390 ;
        RECT 60.880 86.010 61.020 88.070 ;
        RECT 61.340 86.690 61.480 88.410 ;
        RECT 61.280 86.370 61.540 86.690 ;
        RECT 61.800 86.350 61.940 88.750 ;
        RECT 61.740 86.030 62.000 86.350 ;
        RECT 60.820 85.690 61.080 86.010 ;
        RECT 60.880 82.270 61.020 85.690 ;
        RECT 63.120 82.630 63.380 82.950 ;
        RECT 61.280 82.290 61.540 82.610 ;
        RECT 60.820 81.950 61.080 82.270 ;
        RECT 61.340 81.250 61.480 82.290 ;
        RECT 61.280 80.930 61.540 81.250 ;
        RECT 62.660 80.480 62.920 80.570 ;
        RECT 63.180 80.480 63.320 82.630 ;
        RECT 64.100 82.180 64.240 95.890 ;
        RECT 64.560 93.490 64.700 96.570 ;
        RECT 65.480 96.550 65.620 110.170 ;
        RECT 66.340 109.830 66.600 110.150 ;
        RECT 65.420 96.230 65.680 96.550 ;
        RECT 64.500 93.170 64.760 93.490 ;
        RECT 64.560 91.790 64.700 93.170 ;
        RECT 64.500 91.470 64.760 91.790 ;
        RECT 65.480 91.450 65.620 96.230 ;
        RECT 65.420 91.130 65.680 91.450 ;
        RECT 65.880 85.690 66.140 86.010 ;
        RECT 65.420 82.630 65.680 82.950 ;
        RECT 64.500 82.180 64.760 82.270 ;
        RECT 64.100 82.040 64.760 82.180 ;
        RECT 64.500 81.950 64.760 82.040 ;
        RECT 62.660 80.340 63.320 80.480 ;
        RECT 62.660 80.250 62.920 80.340 ;
        RECT 63.180 77.510 63.320 80.340 ;
        RECT 64.040 79.800 64.300 79.890 ;
        RECT 64.560 79.800 64.700 81.950 ;
        RECT 65.480 80.570 65.620 82.630 ;
        RECT 65.940 80.570 66.080 85.690 ;
        RECT 65.420 80.250 65.680 80.570 ;
        RECT 65.880 80.250 66.140 80.570 ;
        RECT 65.480 80.085 65.620 80.250 ;
        RECT 64.040 79.660 64.700 79.800 ;
        RECT 65.410 79.715 65.690 80.085 ;
        RECT 64.040 79.570 64.300 79.660 ;
        RECT 63.120 77.190 63.380 77.510 ;
        RECT 60.810 74.955 61.090 75.325 ;
        RECT 61.280 75.150 61.540 75.470 ;
        RECT 60.820 74.810 61.080 74.955 ;
        RECT 61.340 72.750 61.480 75.150 ;
        RECT 62.200 74.810 62.460 75.130 ;
        RECT 61.280 72.430 61.540 72.750 ;
        RECT 62.260 72.070 62.400 74.810 ;
        RECT 63.180 72.070 63.320 77.190 ;
        RECT 64.040 75.490 64.300 75.810 ;
        RECT 64.100 74.110 64.240 75.490 ;
        RECT 64.040 73.790 64.300 74.110 ;
        RECT 61.740 71.750 62.000 72.070 ;
        RECT 62.200 71.750 62.460 72.070 ;
        RECT 63.120 71.980 63.380 72.070 ;
        RECT 62.720 71.840 63.380 71.980 ;
        RECT 60.820 66.650 61.080 66.970 ;
        RECT 60.880 63.910 61.020 66.650 ;
        RECT 61.280 66.310 61.540 66.630 ;
        RECT 60.820 63.590 61.080 63.910 ;
        RECT 61.340 63.820 61.480 66.310 ;
        RECT 61.800 64.930 61.940 71.750 ;
        RECT 62.200 67.165 62.460 67.310 ;
        RECT 62.190 66.795 62.470 67.165 ;
        RECT 62.720 66.630 62.860 71.840 ;
        RECT 63.120 71.750 63.380 71.840 ;
        RECT 63.120 71.070 63.380 71.390 ;
        RECT 63.180 70.370 63.320 71.070 ;
        RECT 64.100 70.370 64.240 73.790 ;
        RECT 63.120 70.050 63.380 70.370 ;
        RECT 64.040 70.050 64.300 70.370 ;
        RECT 63.120 69.370 63.380 69.690 ;
        RECT 64.040 69.370 64.300 69.690 ;
        RECT 62.660 66.310 62.920 66.630 ;
        RECT 61.740 64.610 62.000 64.930 ;
        RECT 62.200 64.610 62.460 64.930 ;
        RECT 61.740 63.820 62.000 63.910 ;
        RECT 61.340 63.680 62.000 63.820 ;
        RECT 61.740 63.590 62.000 63.680 ;
        RECT 60.880 62.210 61.020 63.590 ;
        RECT 60.820 61.890 61.080 62.210 ;
        RECT 61.800 58.720 61.940 63.590 ;
        RECT 62.260 61.190 62.400 64.610 ;
        RECT 63.180 63.230 63.320 69.370 ;
        RECT 64.100 64.250 64.240 69.370 ;
        RECT 64.040 63.930 64.300 64.250 ;
        RECT 63.120 62.910 63.380 63.230 ;
        RECT 62.200 60.870 62.460 61.190 ;
        RECT 62.200 58.720 62.460 58.810 ;
        RECT 61.800 58.580 62.460 58.720 ;
        RECT 62.200 58.490 62.460 58.580 ;
        RECT 62.260 56.090 62.400 58.490 ;
        RECT 62.200 55.770 62.460 56.090 ;
        RECT 61.280 52.370 61.540 52.690 ;
        RECT 60.360 50.670 60.620 50.990 ;
        RECT 61.340 50.310 61.480 52.370 ;
        RECT 61.730 50.475 62.010 50.845 ;
        RECT 61.740 50.330 62.000 50.475 ;
        RECT 48.400 49.990 48.660 50.310 ;
        RECT 50.700 49.990 50.960 50.310 ;
        RECT 52.540 49.990 52.800 50.310 ;
        RECT 53.460 49.990 53.720 50.310 ;
        RECT 53.920 49.990 54.180 50.310 ;
        RECT 57.600 49.990 57.860 50.310 ;
        RECT 58.520 49.990 58.780 50.310 ;
        RECT 61.280 50.165 61.540 50.310 ;
        RECT 48.460 45.890 48.600 49.990 ;
        RECT 50.240 49.650 50.500 49.970 ;
        RECT 50.300 47.250 50.440 49.650 ;
        RECT 52.600 47.930 52.740 49.990 ;
        RECT 52.540 47.610 52.800 47.930 ;
        RECT 53.000 47.610 53.260 47.930 ;
        RECT 50.240 46.930 50.500 47.250 ;
        RECT 48.400 45.570 48.660 45.890 ;
        RECT 47.940 44.890 48.200 45.210 ;
        RECT 47.480 44.550 47.740 44.870 ;
        RECT 48.000 42.150 48.140 44.890 ;
        RECT 50.300 42.490 50.440 46.930 ;
        RECT 53.060 44.190 53.200 47.610 ;
        RECT 53.520 46.910 53.660 49.990 ;
        RECT 53.980 48.610 54.120 49.990 ;
        RECT 54.580 48.775 56.460 49.145 ;
        RECT 57.660 48.610 57.800 49.990 ;
        RECT 53.920 48.290 54.180 48.610 ;
        RECT 54.840 48.290 55.100 48.610 ;
        RECT 57.600 48.290 57.860 48.610 ;
        RECT 54.900 47.930 55.040 48.290 ;
        RECT 55.300 48.125 55.560 48.270 ;
        RECT 54.840 47.610 55.100 47.930 ;
        RECT 55.290 47.755 55.570 48.125 ;
        RECT 53.460 46.590 53.720 46.910 ;
        RECT 53.520 45.210 53.660 46.590 ;
        RECT 53.460 44.890 53.720 45.210 ;
        RECT 51.160 43.870 51.420 44.190 ;
        RECT 53.000 43.870 53.260 44.190 ;
        RECT 50.240 42.170 50.500 42.490 ;
        RECT 47.940 41.830 48.200 42.150 ;
        RECT 47.020 36.730 47.280 37.050 ;
        RECT 48.000 36.710 48.140 41.830 ;
        RECT 48.400 41.490 48.660 41.810 ;
        RECT 48.460 39.090 48.600 41.490 ;
        RECT 51.220 40.450 51.360 43.870 ;
        RECT 54.580 43.335 56.460 43.705 ;
        RECT 51.160 40.130 51.420 40.450 ;
        RECT 48.400 38.770 48.660 39.090 ;
        RECT 51.220 37.730 51.360 40.130 ;
        RECT 52.080 39.450 52.340 39.770 ;
        RECT 51.160 37.410 51.420 37.730 ;
        RECT 44.720 36.390 44.980 36.710 ;
        RECT 47.940 36.390 48.200 36.710 ;
        RECT 41.960 34.010 42.220 34.330 ;
        RECT 52.140 33.990 52.280 39.450 ;
        RECT 54.580 37.895 56.460 38.265 ;
        RECT 58.580 37.730 58.720 49.990 ;
        RECT 61.270 49.795 61.550 50.165 ;
        RECT 62.260 49.630 62.400 55.770 ;
        RECT 62.660 52.370 62.920 52.690 ;
        RECT 62.720 50.650 62.860 52.370 ;
        RECT 62.660 50.330 62.920 50.650 ;
        RECT 61.740 49.310 62.000 49.630 ;
        RECT 62.200 49.310 62.460 49.630 ;
        RECT 61.800 48.610 61.940 49.310 ;
        RECT 61.740 48.290 62.000 48.610 ;
        RECT 62.200 47.610 62.460 47.930 ;
        RECT 62.260 41.810 62.400 47.610 ;
        RECT 62.720 47.590 62.860 50.330 ;
        RECT 62.660 47.270 62.920 47.590 ;
        RECT 62.200 41.490 62.460 41.810 ;
        RECT 59.900 38.770 60.160 39.090 ;
        RECT 59.960 37.730 60.100 38.770 ;
        RECT 60.360 38.430 60.620 38.750 ;
        RECT 58.520 37.410 58.780 37.730 ;
        RECT 59.900 37.410 60.160 37.730 ;
        RECT 60.420 37.050 60.560 38.430 ;
        RECT 57.140 36.730 57.400 37.050 ;
        RECT 60.360 36.730 60.620 37.050 ;
        RECT 56.680 34.010 56.940 34.330 ;
        RECT 39.200 33.670 39.460 33.990 ;
        RECT 49.320 33.670 49.580 33.990 ;
        RECT 52.080 33.670 52.340 33.990 ;
        RECT 28.160 31.290 28.420 31.610 ;
        RECT 28.620 31.290 28.880 31.610 ;
        RECT 35.520 31.290 35.780 31.610 ;
        RECT 20.800 30.270 21.060 30.590 ;
        RECT 23.560 30.270 23.820 30.590 ;
        RECT 9.580 29.735 11.460 30.105 ;
        RECT 28.220 29.570 28.360 31.290 ;
        RECT 28.680 30.930 28.820 31.290 ;
        RECT 28.620 30.610 28.880 30.930 ;
        RECT 28.160 29.250 28.420 29.570 ;
        RECT 28.680 28.550 28.820 30.610 ;
        RECT 39.580 29.735 41.460 30.105 ;
        RECT 49.380 28.550 49.520 33.670 ;
        RECT 54.580 32.455 56.460 32.825 ;
        RECT 56.740 32.290 56.880 34.010 ;
        RECT 56.680 31.970 56.940 32.290 ;
        RECT 57.200 31.950 57.340 36.730 ;
        RECT 58.520 35.710 58.780 36.030 ;
        RECT 58.580 33.650 58.720 35.710 ;
        RECT 58.520 33.330 58.780 33.650 ;
        RECT 57.140 31.630 57.400 31.950 ;
        RECT 60.420 31.690 60.560 36.730 ;
        RECT 62.260 33.310 62.400 41.490 ;
        RECT 62.720 38.750 62.860 47.270 ;
        RECT 62.660 38.430 62.920 38.750 ;
        RECT 63.180 37.640 63.320 62.910 ;
        RECT 63.580 56.110 63.840 56.430 ;
        RECT 63.640 53.370 63.780 56.110 ;
        RECT 63.580 53.050 63.840 53.370 ;
        RECT 64.100 50.990 64.240 63.930 ;
        RECT 64.560 63.910 64.700 79.660 ;
        RECT 64.950 75.635 65.230 76.005 ;
        RECT 65.020 75.470 65.160 75.635 ;
        RECT 64.960 75.150 65.220 75.470 ;
        RECT 64.960 66.650 65.220 66.970 ;
        RECT 64.500 63.590 64.760 63.910 ;
        RECT 64.560 56.430 64.700 63.590 ;
        RECT 65.020 61.190 65.160 66.650 ;
        RECT 64.960 60.870 65.220 61.190 ;
        RECT 64.500 56.110 64.760 56.430 ;
        RECT 64.500 55.430 64.760 55.750 ;
        RECT 63.570 50.475 63.850 50.845 ;
        RECT 64.040 50.670 64.300 50.990 ;
        RECT 63.640 49.880 63.780 50.475 ;
        RECT 64.040 49.880 64.300 49.970 ;
        RECT 63.640 49.740 64.300 49.880 ;
        RECT 64.040 49.650 64.300 49.740 ;
        RECT 63.580 48.290 63.840 48.610 ;
        RECT 63.640 47.930 63.780 48.290 ;
        RECT 63.580 47.610 63.840 47.930 ;
        RECT 64.100 46.910 64.240 49.650 ;
        RECT 64.560 48.270 64.700 55.430 ;
        RECT 65.940 53.450 66.080 80.250 ;
        RECT 66.400 68.410 66.540 109.830 ;
        RECT 67.720 99.630 67.980 99.950 ;
        RECT 67.260 98.270 67.520 98.590 ;
        RECT 67.320 97.570 67.460 98.270 ;
        RECT 67.260 97.250 67.520 97.570 ;
        RECT 67.780 96.890 67.920 99.630 ;
        RECT 67.720 96.570 67.980 96.890 ;
        RECT 68.240 92.210 68.380 120.710 ;
        RECT 75.140 118.650 75.280 120.710 ;
        RECT 75.080 118.330 75.340 118.650 ;
        RECT 69.580 116.775 71.460 117.145 ;
        RECT 75.540 113.230 75.800 113.550 ;
        RECT 71.860 112.550 72.120 112.870 ;
        RECT 69.580 111.335 71.460 111.705 ;
        RECT 71.920 111.170 72.060 112.550 ;
        RECT 71.860 110.850 72.120 111.170 ;
        RECT 68.640 109.830 68.900 110.150 ;
        RECT 70.940 109.830 71.200 110.150 ;
        RECT 68.700 107.090 68.840 109.830 ;
        RECT 71.000 108.450 71.140 109.830 ;
        RECT 74.160 109.490 74.420 109.810 ;
        RECT 74.220 108.450 74.360 109.490 ;
        RECT 75.600 108.450 75.740 113.230 ;
        RECT 76.000 109.150 76.260 109.470 ;
        RECT 70.940 108.130 71.200 108.450 ;
        RECT 74.160 108.130 74.420 108.450 ;
        RECT 75.540 108.130 75.800 108.450 ;
        RECT 76.060 108.110 76.200 109.150 ;
        RECT 76.000 107.790 76.260 108.110 ;
        RECT 69.100 107.450 69.360 107.770 ;
        RECT 71.860 107.450 72.120 107.770 ;
        RECT 68.640 106.770 68.900 107.090 ;
        RECT 69.160 105.730 69.300 107.450 ;
        RECT 69.580 105.895 71.460 106.265 ;
        RECT 69.100 105.410 69.360 105.730 ;
        RECT 69.100 101.330 69.360 101.650 ;
        RECT 69.160 100.290 69.300 101.330 ;
        RECT 69.580 100.455 71.460 100.825 ;
        RECT 69.100 99.970 69.360 100.290 ;
        RECT 71.920 99.270 72.060 107.450 ;
        RECT 74.620 107.110 74.880 107.430 ;
        RECT 74.680 105.050 74.820 107.110 ;
        RECT 74.620 104.730 74.880 105.050 ;
        RECT 71.860 98.950 72.120 99.270 ;
        RECT 73.240 98.950 73.500 99.270 ;
        RECT 71.400 98.270 71.660 98.590 ;
        RECT 71.460 97.230 71.600 98.270 ;
        RECT 71.400 96.910 71.660 97.230 ;
        RECT 69.580 95.015 71.460 95.385 ;
        RECT 73.300 94.850 73.440 98.950 ;
        RECT 74.160 98.610 74.420 98.930 ;
        RECT 73.240 94.530 73.500 94.850 ;
        RECT 68.240 92.070 68.840 92.210 ;
        RECT 68.180 91.470 68.440 91.790 ;
        RECT 66.800 90.790 67.060 91.110 ;
        RECT 66.860 89.410 67.000 90.790 ;
        RECT 66.800 89.090 67.060 89.410 ;
        RECT 67.720 74.470 67.980 74.790 ;
        RECT 67.780 68.670 67.920 74.470 ;
        RECT 66.400 68.270 67.000 68.410 ;
        RECT 67.720 68.350 67.980 68.670 ;
        RECT 66.860 66.630 67.000 68.270 ;
        RECT 66.800 66.310 67.060 66.630 ;
        RECT 66.340 65.970 66.600 66.290 ;
        RECT 66.400 64.930 66.540 65.970 ;
        RECT 66.340 64.610 66.600 64.930 ;
        RECT 66.860 63.230 67.000 66.310 ;
        RECT 66.800 62.910 67.060 63.230 ;
        RECT 66.340 60.870 66.600 61.190 ;
        RECT 66.400 58.810 66.540 60.870 ;
        RECT 66.340 58.490 66.600 58.810 ;
        RECT 68.240 53.710 68.380 91.470 ;
        RECT 68.700 90.430 68.840 92.070 ;
        RECT 68.640 90.110 68.900 90.430 ;
        RECT 69.580 89.575 71.460 89.945 ;
        RECT 72.320 88.410 72.580 88.730 ;
        RECT 69.100 86.030 69.360 86.350 ;
        RECT 69.160 83.970 69.300 86.030 ;
        RECT 69.580 84.135 71.460 84.505 ;
        RECT 69.100 83.650 69.360 83.970 ;
        RECT 72.380 82.950 72.520 88.410 ;
        RECT 74.220 87.450 74.360 98.610 ;
        RECT 74.680 94.510 74.820 104.730 ;
        RECT 76.060 104.710 76.200 107.790 ;
        RECT 76.000 104.390 76.260 104.710 ;
        RECT 75.080 104.050 75.340 104.370 ;
        RECT 75.140 97.230 75.280 104.050 ;
        RECT 76.060 99.610 76.200 104.390 ;
        RECT 76.000 99.290 76.260 99.610 ;
        RECT 76.000 98.610 76.260 98.930 ;
        RECT 75.080 96.910 75.340 97.230 ;
        RECT 74.620 94.190 74.880 94.510 ;
        RECT 74.680 93.570 74.820 94.190 ;
        RECT 75.140 94.170 75.280 96.910 ;
        RECT 76.060 96.890 76.200 98.610 ;
        RECT 76.000 96.570 76.260 96.890 ;
        RECT 75.080 93.850 75.340 94.170 ;
        RECT 74.680 93.430 75.740 93.570 ;
        RECT 74.620 92.830 74.880 93.150 ;
        RECT 74.680 92.130 74.820 92.830 ;
        RECT 74.620 91.810 74.880 92.130 ;
        RECT 74.680 88.390 74.820 91.810 ;
        RECT 75.080 91.470 75.340 91.790 ;
        RECT 75.140 89.410 75.280 91.470 ;
        RECT 75.600 90.770 75.740 93.430 ;
        RECT 76.060 91.450 76.200 96.570 ;
        RECT 76.520 94.850 76.660 120.710 ;
        RECT 76.920 111.870 77.180 112.190 ;
        RECT 76.980 108.110 77.120 111.870 ;
        RECT 80.600 109.830 80.860 110.150 ;
        RECT 80.660 108.450 80.800 109.830 ;
        RECT 80.600 108.130 80.860 108.450 ;
        RECT 76.920 107.790 77.180 108.110 ;
        RECT 76.980 104.710 77.120 107.790 ;
        RECT 79.680 107.450 79.940 107.770 ;
        RECT 79.740 105.730 79.880 107.450 ;
        RECT 79.680 105.410 79.940 105.730 ;
        RECT 76.920 104.390 77.180 104.710 ;
        RECT 79.220 99.630 79.480 99.950 ;
        RECT 79.280 99.270 79.420 99.630 ;
        RECT 78.760 98.950 79.020 99.270 ;
        RECT 79.220 98.950 79.480 99.270 ;
        RECT 78.820 96.550 78.960 98.950 ;
        RECT 79.280 96.890 79.420 98.950 ;
        RECT 80.600 98.270 80.860 98.590 ;
        RECT 80.660 97.230 80.800 98.270 ;
        RECT 81.580 97.570 81.720 120.710 ;
        RECT 84.580 119.495 86.460 119.865 ;
        RECT 83.360 114.590 83.620 114.910 ;
        RECT 83.420 113.890 83.560 114.590 ;
        RECT 84.580 114.055 86.460 114.425 ;
        RECT 83.360 113.570 83.620 113.890 ;
        RECT 82.900 112.890 83.160 113.210 ;
        RECT 82.960 108.110 83.100 112.890 ;
        RECT 86.580 112.210 86.840 112.530 ;
        RECT 83.820 111.870 84.080 112.190 ;
        RECT 83.350 109.635 83.630 110.005 ;
        RECT 83.880 109.810 84.020 111.870 ;
        RECT 82.900 107.790 83.160 108.110 ;
        RECT 83.420 107.770 83.560 109.635 ;
        RECT 83.820 109.490 84.080 109.810 ;
        RECT 84.580 108.615 86.460 108.985 ;
        RECT 83.360 107.450 83.620 107.770 ;
        RECT 83.420 107.285 83.560 107.450 ;
        RECT 86.640 107.430 86.780 112.210 ;
        RECT 87.100 110.490 87.240 123.430 ;
        RECT 88.480 122.050 88.620 123.430 ;
        RECT 90.780 123.070 90.920 125.810 ;
        RECT 93.940 123.770 94.200 124.090 ;
        RECT 90.720 122.750 90.980 123.070 ;
        RECT 94.000 122.050 94.140 123.770 ;
        RECT 94.460 123.750 94.600 139.870 ;
        RECT 99.580 127.655 101.460 128.025 ;
        RECT 97.620 125.810 97.880 126.130 ;
        RECT 98.080 125.810 98.340 126.130 ;
        RECT 94.400 123.430 94.660 123.750 ;
        RECT 94.860 123.090 95.120 123.410 ;
        RECT 88.420 121.730 88.680 122.050 ;
        RECT 93.940 121.730 94.200 122.050 ;
        RECT 94.920 121.030 95.060 123.090 ;
        RECT 97.680 121.710 97.820 125.810 ;
        RECT 98.140 124.090 98.280 125.810 ;
        RECT 102.740 125.790 102.880 140.350 ;
        RECT 107.340 127.490 107.480 139.870 ;
        RECT 110.040 128.870 110.300 129.190 ;
        RECT 111.880 128.870 112.140 129.190 ;
        RECT 107.280 127.170 107.540 127.490 ;
        RECT 110.100 126.810 110.240 128.870 ;
        RECT 110.040 126.490 110.300 126.810 ;
        RECT 106.820 125.810 107.080 126.130 ;
        RECT 102.680 125.470 102.940 125.790 ;
        RECT 98.080 123.770 98.340 124.090 ;
        RECT 99.580 122.215 101.460 122.585 ;
        RECT 106.880 122.050 107.020 125.810 ;
        RECT 110.100 124.430 110.240 126.490 ;
        RECT 110.500 125.810 110.760 126.130 ;
        RECT 110.560 124.770 110.700 125.810 ;
        RECT 110.500 124.450 110.760 124.770 ;
        RECT 110.040 124.110 110.300 124.430 ;
        RECT 107.280 123.770 107.540 124.090 ;
        RECT 106.820 121.730 107.080 122.050 ;
        RECT 107.340 121.710 107.480 123.770 ;
        RECT 108.200 123.430 108.460 123.750 ;
        RECT 108.260 122.050 108.400 123.430 ;
        RECT 108.200 121.730 108.460 122.050 ;
        RECT 97.620 121.390 97.880 121.710 ;
        RECT 107.280 121.390 107.540 121.710 ;
        RECT 108.200 121.050 108.460 121.370 ;
        RECT 88.420 120.710 88.680 121.030 ;
        RECT 90.260 120.710 90.520 121.030 ;
        RECT 92.100 120.710 92.360 121.030 ;
        RECT 94.860 120.710 95.120 121.030 ;
        RECT 104.520 120.710 104.780 121.030 ;
        RECT 87.500 112.890 87.760 113.210 ;
        RECT 87.560 110.830 87.700 112.890 ;
        RECT 87.500 110.510 87.760 110.830 ;
        RECT 87.040 110.170 87.300 110.490 ;
        RECT 83.350 106.915 83.630 107.285 ;
        RECT 86.580 107.110 86.840 107.430 ;
        RECT 86.640 105.390 86.780 107.110 ;
        RECT 87.100 106.750 87.240 110.170 ;
        RECT 87.040 106.430 87.300 106.750 ;
        RECT 86.580 105.070 86.840 105.390 ;
        RECT 81.980 104.390 82.240 104.710 ;
        RECT 86.580 104.390 86.840 104.710 ;
        RECT 82.040 99.270 82.180 104.390 ;
        RECT 84.580 103.175 86.460 103.545 ;
        RECT 84.280 102.010 84.540 102.330 ;
        RECT 84.340 100.290 84.480 102.010 ;
        RECT 84.280 99.970 84.540 100.290 ;
        RECT 86.640 99.950 86.780 104.390 ;
        RECT 82.440 99.690 82.700 99.950 ;
        RECT 82.440 99.630 83.100 99.690 ;
        RECT 86.580 99.630 86.840 99.950 ;
        RECT 82.500 99.550 83.100 99.630 ;
        RECT 82.960 99.270 83.100 99.550 ;
        RECT 81.980 98.950 82.240 99.270 ;
        RECT 82.900 98.950 83.160 99.270 ;
        RECT 82.440 98.270 82.700 98.590 ;
        RECT 82.900 98.270 83.160 98.590 ;
        RECT 81.520 97.250 81.780 97.570 ;
        RECT 80.600 96.910 80.860 97.230 ;
        RECT 79.220 96.570 79.480 96.890 ;
        RECT 81.060 96.570 81.320 96.890 ;
        RECT 78.760 96.230 79.020 96.550 ;
        RECT 76.460 94.530 76.720 94.850 ;
        RECT 78.820 91.790 78.960 96.230 ;
        RECT 80.600 95.550 80.860 95.870 ;
        RECT 80.140 93.850 80.400 94.170 ;
        RECT 79.220 93.510 79.480 93.830 ;
        RECT 78.760 91.470 79.020 91.790 ;
        RECT 76.000 91.130 76.260 91.450 ;
        RECT 75.540 90.450 75.800 90.770 ;
        RECT 75.080 89.090 75.340 89.410 ;
        RECT 75.600 89.070 75.740 90.450 ;
        RECT 75.540 88.750 75.800 89.070 ;
        RECT 74.620 88.070 74.880 88.390 ;
        RECT 75.080 88.070 75.340 88.390 ;
        RECT 75.140 87.450 75.280 88.070 ;
        RECT 74.220 87.310 75.280 87.450 ;
        RECT 77.840 87.390 78.100 87.710 ;
        RECT 72.780 82.970 73.040 83.290 ;
        RECT 71.400 82.630 71.660 82.950 ;
        RECT 72.320 82.630 72.580 82.950 ;
        RECT 70.480 81.950 70.740 82.270 ;
        RECT 70.540 80.570 70.680 81.950 ;
        RECT 70.480 80.250 70.740 80.570 ;
        RECT 71.460 80.230 71.600 82.630 ;
        RECT 68.640 79.910 68.900 80.230 ;
        RECT 71.400 79.910 71.660 80.230 ;
        RECT 68.700 77.850 68.840 79.910 ;
        RECT 69.580 78.695 71.460 79.065 ;
        RECT 72.380 78.530 72.520 82.630 ;
        RECT 72.320 78.210 72.580 78.530 ;
        RECT 68.640 77.530 68.900 77.850 ;
        RECT 71.860 73.790 72.120 74.110 ;
        RECT 69.580 73.255 71.460 73.625 ;
        RECT 68.640 72.770 68.900 73.090 ;
        RECT 68.700 70.370 68.840 72.770 ;
        RECT 71.920 72.070 72.060 73.790 ;
        RECT 69.100 71.750 69.360 72.070 ;
        RECT 71.860 71.750 72.120 72.070 ;
        RECT 68.640 70.050 68.900 70.370 ;
        RECT 69.160 69.090 69.300 71.750 ;
        RECT 68.700 68.950 69.300 69.090 ;
        RECT 68.700 67.310 68.840 68.950 ;
        RECT 69.100 68.350 69.360 68.670 ;
        RECT 68.640 66.990 68.900 67.310 ;
        RECT 69.160 66.630 69.300 68.350 ;
        RECT 69.580 67.815 71.460 68.185 ;
        RECT 72.320 66.650 72.580 66.970 ;
        RECT 69.100 66.310 69.360 66.630 ;
        RECT 72.380 64.250 72.520 66.650 ;
        RECT 71.860 63.930 72.120 64.250 ;
        RECT 72.320 63.930 72.580 64.250 ;
        RECT 69.580 62.375 71.460 62.745 ;
        RECT 71.920 62.170 72.060 63.930 ;
        RECT 71.920 62.030 72.520 62.170 ;
        RECT 72.380 60.510 72.520 62.030 ;
        RECT 72.840 61.530 72.980 82.970 ;
        RECT 74.160 81.950 74.420 82.270 ;
        RECT 74.220 80.910 74.360 81.950 ;
        RECT 74.160 80.590 74.420 80.910 ;
        RECT 73.690 75.635 73.970 76.005 ;
        RECT 73.760 75.470 73.900 75.635 ;
        RECT 73.700 75.150 73.960 75.470 ;
        RECT 74.680 74.110 74.820 87.310 ;
        RECT 76.460 85.350 76.720 85.670 ;
        RECT 76.000 84.670 76.260 84.990 ;
        RECT 75.080 77.420 75.340 77.510 ;
        RECT 76.060 77.420 76.200 84.670 ;
        RECT 75.080 77.280 76.200 77.420 ;
        RECT 75.080 77.190 75.340 77.280 ;
        RECT 74.620 73.790 74.880 74.110 ;
        RECT 75.540 69.030 75.800 69.350 ;
        RECT 75.600 67.650 75.740 69.030 ;
        RECT 75.540 67.330 75.800 67.650 ;
        RECT 74.160 65.970 74.420 66.290 ;
        RECT 74.220 64.930 74.360 65.970 ;
        RECT 74.160 64.610 74.420 64.930 ;
        RECT 73.700 63.590 73.960 63.910 ;
        RECT 73.760 62.210 73.900 63.590 ;
        RECT 76.000 62.910 76.260 63.230 ;
        RECT 73.700 61.890 73.960 62.210 ;
        RECT 72.780 61.210 73.040 61.530 ;
        RECT 72.320 60.190 72.580 60.510 ;
        RECT 72.380 59.150 72.520 60.190 ;
        RECT 72.320 58.830 72.580 59.150 ;
        RECT 69.580 56.935 71.460 57.305 ;
        RECT 74.620 55.090 74.880 55.410 ;
        RECT 70.480 54.750 70.740 55.070 ;
        RECT 70.540 53.710 70.680 54.750 ;
        RECT 65.940 53.310 66.540 53.450 ;
        RECT 66.800 53.390 67.060 53.710 ;
        RECT 67.720 53.390 67.980 53.710 ;
        RECT 68.180 53.390 68.440 53.710 ;
        RECT 70.480 53.390 70.740 53.710 ;
        RECT 66.400 53.030 66.540 53.310 ;
        RECT 66.860 53.030 67.000 53.390 ;
        RECT 64.960 52.940 65.220 53.030 ;
        RECT 64.960 52.800 65.620 52.940 ;
        RECT 64.960 52.710 65.220 52.800 ;
        RECT 65.480 50.650 65.620 52.800 ;
        RECT 65.880 52.710 66.140 53.030 ;
        RECT 66.340 52.710 66.600 53.030 ;
        RECT 66.800 52.710 67.060 53.030 ;
        RECT 65.420 50.330 65.680 50.650 ;
        RECT 64.500 47.950 64.760 48.270 ;
        RECT 65.480 47.590 65.620 50.330 ;
        RECT 65.940 50.310 66.080 52.710 ;
        RECT 66.340 52.030 66.600 52.350 ;
        RECT 66.400 50.650 66.540 52.030 ;
        RECT 66.340 50.330 66.600 50.650 ;
        RECT 66.860 50.310 67.000 52.710 ;
        RECT 67.260 52.030 67.520 52.350 ;
        RECT 67.320 51.330 67.460 52.030 ;
        RECT 67.260 51.010 67.520 51.330 ;
        RECT 67.780 50.990 67.920 53.390 ;
        RECT 68.180 52.710 68.440 53.030 ;
        RECT 69.100 52.710 69.360 53.030 ;
        RECT 67.720 50.670 67.980 50.990 ;
        RECT 68.240 50.650 68.380 52.710 ;
        RECT 68.180 50.330 68.440 50.650 ;
        RECT 69.160 50.310 69.300 52.710 ;
        RECT 69.580 51.495 71.460 51.865 ;
        RECT 74.680 50.310 74.820 55.090 ;
        RECT 76.060 54.130 76.200 62.910 ;
        RECT 76.520 57.790 76.660 85.350 ;
        RECT 77.900 83.290 78.040 87.390 ;
        RECT 78.760 85.690 79.020 86.010 ;
        RECT 78.300 84.670 78.560 84.990 ;
        RECT 77.840 82.970 78.100 83.290 ;
        RECT 77.900 81.250 78.040 82.970 ;
        RECT 77.840 80.930 78.100 81.250 ;
        RECT 78.360 77.170 78.500 84.670 ;
        RECT 78.820 83.630 78.960 85.690 ;
        RECT 78.760 83.310 79.020 83.630 ;
        RECT 78.300 76.850 78.560 77.170 ;
        RECT 79.280 73.090 79.420 93.510 ;
        RECT 79.680 85.010 79.940 85.330 ;
        RECT 79.740 82.950 79.880 85.010 ;
        RECT 79.680 82.630 79.940 82.950 ;
        RECT 79.220 72.770 79.480 73.090 ;
        RECT 77.840 71.750 78.100 72.070 ;
        RECT 78.300 71.750 78.560 72.070 ;
        RECT 77.900 71.390 78.040 71.750 ;
        RECT 77.840 71.070 78.100 71.390 ;
        RECT 78.360 70.370 78.500 71.750 ;
        RECT 78.760 71.410 79.020 71.730 ;
        RECT 78.300 70.050 78.560 70.370 ;
        RECT 78.820 69.010 78.960 71.410 ;
        RECT 78.760 68.690 79.020 69.010 ;
        RECT 76.920 67.330 77.180 67.650 ;
        RECT 76.980 61.190 77.120 67.330 ;
        RECT 78.820 66.970 78.960 68.690 ;
        RECT 78.760 66.650 79.020 66.970 ;
        RECT 77.380 64.270 77.640 64.590 ;
        RECT 77.440 62.210 77.580 64.270 ;
        RECT 79.220 63.250 79.480 63.570 ;
        RECT 77.380 61.890 77.640 62.210 ;
        RECT 79.280 61.530 79.420 63.250 ;
        RECT 79.220 61.210 79.480 61.530 ;
        RECT 76.920 60.870 77.180 61.190 ;
        RECT 76.460 57.470 76.720 57.790 ;
        RECT 76.060 53.990 77.580 54.130 ;
        RECT 76.920 53.050 77.180 53.370 ;
        RECT 76.980 50.310 77.120 53.050 ;
        RECT 65.880 49.990 66.140 50.310 ;
        RECT 66.330 49.795 66.610 50.165 ;
        RECT 66.800 49.990 67.060 50.310 ;
        RECT 69.100 49.990 69.360 50.310 ;
        RECT 74.620 49.990 74.880 50.310 ;
        RECT 76.920 49.990 77.180 50.310 ;
        RECT 66.340 49.650 66.600 49.795 ;
        RECT 66.860 47.930 67.000 49.990 ;
        RECT 66.800 47.610 67.060 47.930 ;
        RECT 65.420 47.270 65.680 47.590 ;
        RECT 64.040 46.590 64.300 46.910 ;
        RECT 63.580 37.640 63.840 37.730 ;
        RECT 63.180 37.500 63.840 37.640 ;
        RECT 63.580 37.410 63.840 37.500 ;
        RECT 64.100 37.130 64.240 46.590 ;
        RECT 65.480 42.830 65.620 47.270 ;
        RECT 65.870 42.995 66.150 43.365 ;
        RECT 65.880 42.850 66.140 42.995 ;
        RECT 65.420 42.510 65.680 42.830 ;
        RECT 64.500 41.830 64.760 42.150 ;
        RECT 64.960 41.830 65.220 42.150 ;
        RECT 63.640 36.990 64.240 37.130 ;
        RECT 64.560 37.050 64.700 41.830 ;
        RECT 65.020 40.450 65.160 41.830 ;
        RECT 64.960 40.130 65.220 40.450 ;
        RECT 62.660 36.390 62.920 36.710 ;
        RECT 62.720 33.990 62.860 36.390 ;
        RECT 63.120 36.050 63.380 36.370 ;
        RECT 62.660 33.670 62.920 33.990 ;
        RECT 62.200 32.990 62.460 33.310 ;
        RECT 60.420 31.610 61.020 31.690 ;
        RECT 61.280 31.630 61.540 31.950 ;
        RECT 58.060 31.290 58.320 31.610 ;
        RECT 60.360 31.550 61.020 31.610 ;
        RECT 60.360 31.290 60.620 31.550 ;
        RECT 53.920 30.270 54.180 30.590 ;
        RECT 28.620 28.230 28.880 28.550 ;
        RECT 49.320 28.230 49.580 28.550 ;
        RECT 24.580 27.015 26.460 27.385 ;
        RECT 49.380 26.510 49.520 28.230 ;
        RECT 53.980 28.210 54.120 30.270 ;
        RECT 50.700 27.890 50.960 28.210 ;
        RECT 53.920 27.890 54.180 28.210 ;
        RECT 50.760 26.850 50.900 27.890 ;
        RECT 58.120 27.870 58.260 31.290 ;
        RECT 60.360 30.610 60.620 30.930 ;
        RECT 58.520 30.270 58.780 30.590 ;
        RECT 58.060 27.550 58.320 27.870 ;
        RECT 54.580 27.015 56.460 27.385 ;
        RECT 50.700 26.530 50.960 26.850 ;
        RECT 49.320 26.190 49.580 26.510 ;
        RECT 58.120 25.830 58.260 27.550 ;
        RECT 58.580 26.850 58.720 30.270 ;
        RECT 60.420 28.890 60.560 30.610 ;
        RECT 60.360 28.570 60.620 28.890 ;
        RECT 58.520 26.530 58.780 26.850 ;
        RECT 59.900 26.080 60.160 26.170 ;
        RECT 60.420 26.080 60.560 28.570 ;
        RECT 60.880 27.870 61.020 31.550 ;
        RECT 60.820 27.550 61.080 27.870 ;
        RECT 60.880 26.170 61.020 27.550 ;
        RECT 61.340 26.850 61.480 31.630 ;
        RECT 61.740 30.270 62.000 30.590 ;
        RECT 61.800 29.230 61.940 30.270 ;
        RECT 62.720 29.570 62.860 33.670 ;
        RECT 62.660 29.250 62.920 29.570 ;
        RECT 63.180 29.230 63.320 36.050 ;
        RECT 63.640 36.030 63.780 36.990 ;
        RECT 64.500 36.730 64.760 37.050 ;
        RECT 63.580 35.710 63.840 36.030 ;
        RECT 63.640 30.930 63.780 35.710 ;
        RECT 64.560 34.330 64.700 36.730 ;
        RECT 65.480 36.370 65.620 42.510 ;
        RECT 67.720 42.170 67.980 42.490 ;
        RECT 66.340 41.150 66.600 41.470 ;
        RECT 66.400 39.090 66.540 41.150 ;
        RECT 67.260 40.130 67.520 40.450 ;
        RECT 66.340 38.770 66.600 39.090 ;
        RECT 67.320 37.050 67.460 40.130 ;
        RECT 67.260 36.730 67.520 37.050 ;
        RECT 67.780 36.710 67.920 42.170 ;
        RECT 67.720 36.390 67.980 36.710 ;
        RECT 65.420 36.050 65.680 36.370 ;
        RECT 67.780 34.670 67.920 36.390 ;
        RECT 67.720 34.350 67.980 34.670 ;
        RECT 64.500 34.010 64.760 34.330 ;
        RECT 64.040 32.990 64.300 33.310 ;
        RECT 64.100 31.270 64.240 32.990 ;
        RECT 69.160 31.610 69.300 49.990 ;
        RECT 76.000 49.310 76.260 49.630 ;
        RECT 76.460 49.310 76.720 49.630 ;
        RECT 76.060 47.590 76.200 49.310 ;
        RECT 76.520 47.930 76.660 49.310 ;
        RECT 76.460 47.610 76.720 47.930 ;
        RECT 76.000 47.270 76.260 47.590 ;
        RECT 75.080 46.590 75.340 46.910 ;
        RECT 69.580 46.055 71.460 46.425 ;
        RECT 75.140 45.210 75.280 46.590 ;
        RECT 75.080 44.890 75.340 45.210 ;
        RECT 72.780 44.550 73.040 44.870 ;
        RECT 69.580 40.615 71.460 40.985 ;
        RECT 72.840 39.770 72.980 44.550 ;
        RECT 76.060 42.150 76.200 47.270 ;
        RECT 77.440 42.490 77.580 53.990 ;
        RECT 78.760 53.390 79.020 53.710 ;
        RECT 78.300 52.030 78.560 52.350 ;
        RECT 78.360 50.990 78.500 52.030 ;
        RECT 78.300 50.670 78.560 50.990 ;
        RECT 78.820 50.320 78.960 53.390 ;
        RECT 80.200 51.330 80.340 93.850 ;
        RECT 80.660 93.830 80.800 95.550 ;
        RECT 81.120 94.170 81.260 96.570 ;
        RECT 81.060 93.850 81.320 94.170 ;
        RECT 80.600 93.510 80.860 93.830 ;
        RECT 81.120 93.060 81.260 93.850 ;
        RECT 82.500 93.830 82.640 98.270 ;
        RECT 82.960 94.850 83.100 98.270 ;
        RECT 84.580 97.735 86.460 98.105 ;
        RECT 83.820 96.570 84.080 96.890 ;
        RECT 82.900 94.530 83.160 94.850 ;
        RECT 82.440 93.510 82.700 93.830 ;
        RECT 80.660 92.920 81.260 93.060 ;
        RECT 80.660 91.450 80.800 92.920 ;
        RECT 80.600 91.130 80.860 91.450 ;
        RECT 83.360 91.130 83.620 91.450 ;
        RECT 80.660 86.350 80.800 91.130 ;
        RECT 80.600 86.030 80.860 86.350 ;
        RECT 82.900 85.350 83.160 85.670 ;
        RECT 82.960 83.370 83.100 85.350 ;
        RECT 82.500 83.230 83.100 83.370 ;
        RECT 81.520 82.630 81.780 82.950 ;
        RECT 80.600 82.290 80.860 82.610 ;
        RECT 80.660 80.570 80.800 82.290 ;
        RECT 81.580 81.250 81.720 82.630 ;
        RECT 82.500 81.250 82.640 83.230 ;
        RECT 82.900 82.630 83.160 82.950 ;
        RECT 81.520 80.930 81.780 81.250 ;
        RECT 82.440 80.930 82.700 81.250 ;
        RECT 80.600 80.250 80.860 80.570 ;
        RECT 82.440 80.250 82.700 80.570 ;
        RECT 80.660 79.550 80.800 80.250 ;
        RECT 81.980 79.910 82.240 80.230 ;
        RECT 80.600 79.230 80.860 79.550 ;
        RECT 82.040 78.530 82.180 79.910 ;
        RECT 81.980 78.210 82.240 78.530 ;
        RECT 82.500 77.510 82.640 80.250 ;
        RECT 82.960 77.850 83.100 82.630 ;
        RECT 82.900 77.530 83.160 77.850 ;
        RECT 82.440 77.190 82.700 77.510 ;
        RECT 82.500 76.830 82.640 77.190 ;
        RECT 82.440 76.510 82.700 76.830 ;
        RECT 81.060 74.130 81.320 74.450 ;
        RECT 81.120 72.070 81.260 74.130 ;
        RECT 81.060 71.750 81.320 72.070 ;
        RECT 81.520 71.750 81.780 72.070 ;
        RECT 81.580 71.390 81.720 71.750 ;
        RECT 81.520 71.070 81.780 71.390 ;
        RECT 81.520 69.370 81.780 69.690 ;
        RECT 81.060 69.030 81.320 69.350 ;
        RECT 80.600 67.330 80.860 67.650 ;
        RECT 80.660 67.165 80.800 67.330 ;
        RECT 80.590 66.795 80.870 67.165 ;
        RECT 81.120 66.970 81.260 69.030 ;
        RECT 81.060 66.650 81.320 66.970 ;
        RECT 81.120 66.370 81.260 66.650 ;
        RECT 81.580 66.630 81.720 69.370 ;
        RECT 81.980 67.050 82.240 67.310 ;
        RECT 82.960 67.050 83.100 77.530 ;
        RECT 83.420 73.090 83.560 91.130 ;
        RECT 83.880 73.090 84.020 96.570 ;
        RECT 85.660 96.230 85.920 96.550 ;
        RECT 85.720 93.830 85.860 96.230 ;
        RECT 85.660 93.510 85.920 93.830 ;
        RECT 86.580 93.170 86.840 93.490 ;
        RECT 84.580 92.295 86.460 92.665 ;
        RECT 86.640 92.130 86.780 93.170 ;
        RECT 86.580 91.810 86.840 92.130 ;
        RECT 86.580 90.790 86.840 91.110 ;
        RECT 84.580 86.855 86.460 87.225 ;
        RECT 84.580 81.415 86.460 81.785 ;
        RECT 86.120 79.910 86.380 80.230 ;
        RECT 86.180 78.190 86.320 79.910 ;
        RECT 86.120 77.870 86.380 78.190 ;
        RECT 84.580 75.975 86.460 76.345 ;
        RECT 83.360 72.770 83.620 73.090 ;
        RECT 83.820 72.770 84.080 73.090 ;
        RECT 85.200 72.430 85.460 72.750 ;
        RECT 85.260 72.070 85.400 72.430 ;
        RECT 85.200 71.750 85.460 72.070 ;
        RECT 83.820 71.410 84.080 71.730 ;
        RECT 83.880 70.280 84.020 71.410 ;
        RECT 84.580 70.535 86.460 70.905 ;
        RECT 83.880 70.140 84.480 70.280 ;
        RECT 84.340 69.690 84.480 70.140 ;
        RECT 84.280 69.370 84.540 69.690 ;
        RECT 83.820 69.030 84.080 69.350 ;
        RECT 83.360 68.350 83.620 68.670 ;
        RECT 81.980 66.990 83.100 67.050 ;
        RECT 82.040 66.910 83.100 66.990 ;
        RECT 80.660 66.230 81.260 66.370 ;
        RECT 81.520 66.310 81.780 66.630 ;
        RECT 80.660 63.910 80.800 66.230 ;
        RECT 81.060 65.630 81.320 65.950 ;
        RECT 81.120 64.930 81.260 65.630 ;
        RECT 81.060 64.610 81.320 64.930 ;
        RECT 82.960 64.590 83.100 66.910 ;
        RECT 82.900 64.270 83.160 64.590 ;
        RECT 80.600 63.590 80.860 63.910 ;
        RECT 82.960 63.570 83.100 64.270 ;
        RECT 83.420 64.250 83.560 68.350 ;
        RECT 83.880 64.930 84.020 69.030 ;
        RECT 84.340 65.950 84.480 69.370 ;
        RECT 85.660 68.690 85.920 69.010 ;
        RECT 85.720 66.970 85.860 68.690 ;
        RECT 85.660 66.650 85.920 66.970 ;
        RECT 84.280 65.630 84.540 65.950 ;
        RECT 84.580 65.095 86.460 65.465 ;
        RECT 83.820 64.610 84.080 64.930 ;
        RECT 83.360 63.930 83.620 64.250 ;
        RECT 82.900 63.250 83.160 63.570 ;
        RECT 81.520 62.910 81.780 63.230 ;
        RECT 81.580 62.170 81.720 62.910 ;
        RECT 81.120 62.030 81.720 62.170 ;
        RECT 81.120 60.850 81.260 62.030 ;
        RECT 83.360 61.210 83.620 61.530 ;
        RECT 81.060 60.530 81.320 60.850 ;
        RECT 83.420 58.470 83.560 61.210 ;
        RECT 84.580 59.655 86.460 60.025 ;
        RECT 83.360 58.150 83.620 58.470 ;
        RECT 80.140 51.010 80.400 51.330 ;
        RECT 78.760 50.000 79.020 50.320 ;
        RECT 82.900 49.990 83.160 50.310 ;
        RECT 79.680 49.650 79.940 49.970 ;
        RECT 77.840 47.610 78.100 47.930 ;
        RECT 77.900 45.210 78.040 47.610 ;
        RECT 77.840 44.890 78.100 45.210 ;
        RECT 77.380 42.170 77.640 42.490 ;
        RECT 76.000 41.830 76.260 42.150 ;
        RECT 72.780 39.450 73.040 39.770 ;
        RECT 70.480 39.110 70.740 39.430 ;
        RECT 70.540 37.730 70.680 39.110 ;
        RECT 73.700 38.770 73.960 39.090 ;
        RECT 73.760 37.730 73.900 38.770 ;
        RECT 70.480 37.410 70.740 37.730 ;
        RECT 73.700 37.410 73.960 37.730 ;
        RECT 76.060 36.710 76.200 41.830 ;
        RECT 77.900 37.730 78.040 44.890 ;
        RECT 78.760 44.210 79.020 44.530 ;
        RECT 78.820 43.170 78.960 44.210 ;
        RECT 79.740 44.190 79.880 49.650 ;
        RECT 82.440 47.270 82.700 47.590 ;
        RECT 82.500 45.890 82.640 47.270 ;
        RECT 82.960 47.250 83.100 49.990 ;
        RECT 83.420 49.630 83.560 58.150 ;
        RECT 84.580 54.215 86.460 54.585 ;
        RECT 86.120 53.050 86.380 53.370 ;
        RECT 86.180 52.690 86.320 53.050 ;
        RECT 86.120 52.370 86.380 52.690 ;
        RECT 83.820 52.030 84.080 52.350 ;
        RECT 83.880 51.330 84.020 52.030 ;
        RECT 86.180 51.330 86.320 52.370 ;
        RECT 83.820 51.010 84.080 51.330 ;
        RECT 86.120 51.010 86.380 51.330 ;
        RECT 83.360 49.310 83.620 49.630 ;
        RECT 82.900 46.930 83.160 47.250 ;
        RECT 82.440 45.570 82.700 45.890 ;
        RECT 79.680 43.870 79.940 44.190 ;
        RECT 78.760 42.850 79.020 43.170 ;
        RECT 79.740 40.450 79.880 43.870 ;
        RECT 80.600 42.170 80.860 42.490 ;
        RECT 79.680 40.130 79.940 40.450 ;
        RECT 80.140 38.770 80.400 39.090 ;
        RECT 80.200 37.730 80.340 38.770 ;
        RECT 77.840 37.410 78.100 37.730 ;
        RECT 80.140 37.410 80.400 37.730 ;
        RECT 80.660 37.050 80.800 42.170 ;
        RECT 83.420 39.770 83.560 49.310 ;
        RECT 83.880 48.270 84.020 51.010 ;
        RECT 84.580 48.775 86.460 49.145 ;
        RECT 83.820 47.950 84.080 48.270 ;
        RECT 84.740 47.610 85.000 47.930 ;
        RECT 84.800 45.210 84.940 47.610 ;
        RECT 86.640 47.250 86.780 90.790 ;
        RECT 87.100 88.730 87.240 106.430 ;
        RECT 87.560 104.710 87.700 110.510 ;
        RECT 87.500 104.390 87.760 104.710 ;
        RECT 88.480 103.010 88.620 120.710 ;
        RECT 88.880 117.310 89.140 117.630 ;
        RECT 88.940 115.250 89.080 117.310 ;
        RECT 88.880 114.930 89.140 115.250 ;
        RECT 88.880 113.570 89.140 113.890 ;
        RECT 88.940 110.470 89.080 113.570 ;
        RECT 88.940 110.330 89.540 110.470 ;
        RECT 88.880 103.710 89.140 104.030 ;
        RECT 88.420 102.690 88.680 103.010 ;
        RECT 87.500 102.010 87.760 102.330 ;
        RECT 87.960 102.010 88.220 102.330 ;
        RECT 87.040 88.410 87.300 88.730 ;
        RECT 87.560 73.090 87.700 102.010 ;
        RECT 88.020 100.290 88.160 102.010 ;
        RECT 88.420 101.670 88.680 101.990 ;
        RECT 87.960 99.970 88.220 100.290 ;
        RECT 87.960 92.830 88.220 93.150 ;
        RECT 88.020 90.430 88.160 92.830 ;
        RECT 87.960 90.110 88.220 90.430 ;
        RECT 87.960 84.670 88.220 84.990 ;
        RECT 88.020 83.290 88.160 84.670 ;
        RECT 87.960 82.970 88.220 83.290 ;
        RECT 87.960 79.230 88.220 79.550 ;
        RECT 87.040 72.770 87.300 73.090 ;
        RECT 87.500 72.770 87.760 73.090 ;
        RECT 87.100 72.070 87.240 72.770 ;
        RECT 87.040 71.750 87.300 72.070 ;
        RECT 87.500 71.410 87.760 71.730 ;
        RECT 87.040 68.350 87.300 68.670 ;
        RECT 87.100 66.290 87.240 68.350 ;
        RECT 87.040 65.970 87.300 66.290 ;
        RECT 87.100 64.930 87.240 65.970 ;
        RECT 87.560 64.930 87.700 71.410 ;
        RECT 87.040 64.610 87.300 64.930 ;
        RECT 87.500 64.610 87.760 64.930 ;
        RECT 87.560 64.250 87.700 64.610 ;
        RECT 87.500 63.930 87.760 64.250 ;
        RECT 87.040 52.710 87.300 53.030 ;
        RECT 86.580 46.930 86.840 47.250 ;
        RECT 84.740 44.890 85.000 45.210 ;
        RECT 87.100 44.530 87.240 52.710 ;
        RECT 87.500 52.030 87.760 52.350 ;
        RECT 87.560 47.930 87.700 52.030 ;
        RECT 87.500 47.610 87.760 47.930 ;
        RECT 88.020 45.890 88.160 79.230 ;
        RECT 88.480 54.050 88.620 101.670 ;
        RECT 88.940 101.310 89.080 103.710 ;
        RECT 88.880 100.990 89.140 101.310 ;
        RECT 88.880 96.570 89.140 96.890 ;
        RECT 88.940 86.770 89.080 96.570 ;
        RECT 89.400 92.130 89.540 110.330 ;
        RECT 90.320 103.010 90.460 120.710 ;
        RECT 90.720 115.270 90.980 115.590 ;
        RECT 90.780 113.890 90.920 115.270 ;
        RECT 90.720 113.570 90.980 113.890 ;
        RECT 91.640 103.710 91.900 104.030 ;
        RECT 90.260 102.690 90.520 103.010 ;
        RECT 90.260 102.010 90.520 102.330 ;
        RECT 89.800 101.670 90.060 101.990 ;
        RECT 89.340 91.810 89.600 92.130 ;
        RECT 88.940 86.630 89.540 86.770 ;
        RECT 88.880 85.690 89.140 86.010 ;
        RECT 88.940 81.250 89.080 85.690 ;
        RECT 88.880 80.930 89.140 81.250 ;
        RECT 89.400 79.550 89.540 86.630 ;
        RECT 89.340 79.230 89.600 79.550 ;
        RECT 88.880 72.430 89.140 72.750 ;
        RECT 88.940 72.070 89.080 72.430 ;
        RECT 88.880 71.750 89.140 72.070 ;
        RECT 88.880 69.710 89.140 70.030 ;
        RECT 88.940 68.670 89.080 69.710 ;
        RECT 88.880 68.350 89.140 68.670 ;
        RECT 89.340 65.630 89.600 65.950 ;
        RECT 88.880 64.610 89.140 64.930 ;
        RECT 88.940 61.530 89.080 64.610 ;
        RECT 89.400 62.210 89.540 65.630 ;
        RECT 89.340 61.890 89.600 62.210 ;
        RECT 88.880 61.210 89.140 61.530 ;
        RECT 88.420 53.730 88.680 54.050 ;
        RECT 89.340 53.050 89.600 53.370 ;
        RECT 89.400 52.350 89.540 53.050 ;
        RECT 89.860 52.690 90.000 101.670 ;
        RECT 90.320 73.090 90.460 102.010 ;
        RECT 90.720 101.330 90.980 101.650 ;
        RECT 90.780 95.870 90.920 101.330 ;
        RECT 91.700 101.310 91.840 103.710 ;
        RECT 91.640 100.990 91.900 101.310 ;
        RECT 92.160 97.570 92.300 120.710 ;
        RECT 104.060 120.370 104.320 120.690 ;
        RECT 96.240 118.330 96.500 118.650 ;
        RECT 96.300 115.590 96.440 118.330 ;
        RECT 99.580 116.775 101.460 117.145 ;
        RECT 95.320 115.270 95.580 115.590 ;
        RECT 96.240 115.270 96.500 115.590 ;
        RECT 102.220 115.270 102.480 115.590 ;
        RECT 103.600 115.270 103.860 115.590 ;
        RECT 92.560 112.890 92.820 113.210 ;
        RECT 92.620 111.170 92.760 112.890 ;
        RECT 95.380 112.870 95.520 115.270 ;
        RECT 95.320 112.610 95.580 112.870 ;
        RECT 95.320 112.550 95.980 112.610 ;
        RECT 95.380 112.470 95.980 112.550 ;
        RECT 92.560 110.850 92.820 111.170 ;
        RECT 95.840 107.430 95.980 112.470 ;
        RECT 95.780 107.110 96.040 107.430 ;
        RECT 92.560 104.390 92.820 104.710 ;
        RECT 92.620 102.330 92.760 104.390 ;
        RECT 92.560 102.010 92.820 102.330 ;
        RECT 94.860 101.670 95.120 101.990 ;
        RECT 94.400 100.990 94.660 101.310 ;
        RECT 92.100 97.250 92.360 97.570 ;
        RECT 93.480 96.910 93.740 97.230 ;
        RECT 90.720 95.550 90.980 95.870 ;
        RECT 90.720 90.790 90.980 91.110 ;
        RECT 90.780 89.410 90.920 90.790 ;
        RECT 91.640 90.110 91.900 90.430 ;
        RECT 93.020 90.110 93.280 90.430 ;
        RECT 90.720 89.090 90.980 89.410 ;
        RECT 91.700 88.730 91.840 90.110 ;
        RECT 92.560 89.090 92.820 89.410 ;
        RECT 91.640 88.410 91.900 88.730 ;
        RECT 92.620 86.010 92.760 89.090 ;
        RECT 93.080 88.050 93.220 90.110 ;
        RECT 93.020 87.730 93.280 88.050 ;
        RECT 92.560 85.920 92.820 86.010 ;
        RECT 92.160 85.780 92.820 85.920 ;
        RECT 91.640 85.350 91.900 85.670 ;
        RECT 90.720 85.010 90.980 85.330 ;
        RECT 90.780 83.290 90.920 85.010 ;
        RECT 91.700 83.290 91.840 85.350 ;
        RECT 90.720 82.970 90.980 83.290 ;
        RECT 91.640 82.970 91.900 83.290 ;
        RECT 91.700 80.570 91.840 82.970 ;
        RECT 92.160 81.250 92.300 85.780 ;
        RECT 92.560 85.690 92.820 85.780 ;
        RECT 92.560 82.290 92.820 82.610 ;
        RECT 92.620 81.250 92.760 82.290 ;
        RECT 92.100 80.930 92.360 81.250 ;
        RECT 92.560 80.930 92.820 81.250 ;
        RECT 91.640 80.250 91.900 80.570 ;
        RECT 91.180 74.810 91.440 75.130 ;
        RECT 92.100 74.810 92.360 75.130 ;
        RECT 90.260 72.770 90.520 73.090 ;
        RECT 91.240 72.070 91.380 74.810 ;
        RECT 91.180 71.750 91.440 72.070 ;
        RECT 92.160 70.370 92.300 74.810 ;
        RECT 92.100 70.050 92.360 70.370 ;
        RECT 90.720 69.030 90.980 69.350 ;
        RECT 90.780 67.310 90.920 69.030 ;
        RECT 90.720 66.990 90.980 67.310 ;
        RECT 93.020 63.590 93.280 63.910 ;
        RECT 93.080 62.210 93.220 63.590 ;
        RECT 93.020 61.890 93.280 62.210 ;
        RECT 92.090 59.315 92.370 59.685 ;
        RECT 92.160 59.150 92.300 59.315 ;
        RECT 92.100 58.830 92.360 59.150 ;
        RECT 91.180 57.470 91.440 57.790 ;
        RECT 90.720 55.430 90.980 55.750 ;
        RECT 90.260 55.090 90.520 55.410 ;
        RECT 90.320 54.050 90.460 55.090 ;
        RECT 90.260 53.730 90.520 54.050 ;
        RECT 89.800 52.370 90.060 52.690 ;
        RECT 89.340 52.030 89.600 52.350 ;
        RECT 89.400 48.610 89.540 52.030 ;
        RECT 90.780 51.330 90.920 55.430 ;
        RECT 91.240 53.710 91.380 57.470 ;
        RECT 93.540 56.770 93.680 96.910 ;
        RECT 93.940 96.570 94.200 96.890 ;
        RECT 94.000 75.810 94.140 96.570 ;
        RECT 94.460 95.870 94.600 100.990 ;
        RECT 94.920 99.270 95.060 101.670 ;
        RECT 95.840 99.610 95.980 107.110 ;
        RECT 95.780 99.290 96.040 99.610 ;
        RECT 94.860 98.950 95.120 99.270 ;
        RECT 94.400 95.550 94.660 95.870 ;
        RECT 94.920 93.830 95.060 98.950 ;
        RECT 95.840 96.890 95.980 99.290 ;
        RECT 95.320 96.570 95.580 96.890 ;
        RECT 95.780 96.570 96.040 96.890 ;
        RECT 95.380 94.850 95.520 96.570 ;
        RECT 95.320 94.530 95.580 94.850 ;
        RECT 94.860 93.510 95.120 93.830 ;
        RECT 96.300 91.450 96.440 115.270 ;
        RECT 99.920 114.590 100.180 114.910 ;
        RECT 99.980 113.550 100.120 114.590 ;
        RECT 99.920 113.230 100.180 113.550 ;
        RECT 96.700 112.550 96.960 112.870 ;
        RECT 96.760 109.470 96.900 112.550 ;
        RECT 99.580 111.335 101.460 111.705 ;
        RECT 98.540 110.170 98.800 110.490 ;
        RECT 102.280 110.470 102.420 115.270 ;
        RECT 103.660 113.890 103.800 115.270 ;
        RECT 103.600 113.570 103.860 113.890 ;
        RECT 103.600 112.210 103.860 112.530 ;
        RECT 103.660 111.930 103.800 112.210 ;
        RECT 103.200 111.790 103.800 111.930 ;
        RECT 103.200 110.490 103.340 111.790 ;
        RECT 101.820 110.330 102.420 110.470 ;
        RECT 96.700 109.150 96.960 109.470 ;
        RECT 96.760 105.050 96.900 109.150 ;
        RECT 97.160 107.110 97.420 107.430 ;
        RECT 97.220 105.730 97.360 107.110 ;
        RECT 97.160 105.410 97.420 105.730 ;
        RECT 98.600 105.050 98.740 110.170 ;
        RECT 99.000 109.150 99.260 109.470 ;
        RECT 99.060 106.750 99.200 109.150 ;
        RECT 101.820 107.770 101.960 110.330 ;
        RECT 103.140 110.170 103.400 110.490 ;
        RECT 101.760 107.450 102.020 107.770 ;
        RECT 99.000 106.430 99.260 106.750 ;
        RECT 96.700 104.730 96.960 105.050 ;
        RECT 98.540 104.730 98.800 105.050 ;
        RECT 99.060 103.940 99.200 106.430 ;
        RECT 99.580 105.895 101.460 106.265 ;
        RECT 100.380 104.730 100.640 105.050 ;
        RECT 99.460 103.940 99.720 104.030 ;
        RECT 99.060 103.800 99.720 103.940 ;
        RECT 99.460 103.710 99.720 103.800 ;
        RECT 99.520 102.670 99.660 103.710 ;
        RECT 99.460 102.350 99.720 102.670 ;
        RECT 100.440 101.650 100.580 104.730 ;
        RECT 101.820 102.330 101.960 107.450 ;
        RECT 103.130 106.915 103.410 107.285 ;
        RECT 103.200 104.710 103.340 106.915 ;
        RECT 103.140 104.390 103.400 104.710 ;
        RECT 102.680 103.710 102.940 104.030 ;
        RECT 101.760 102.010 102.020 102.330 ;
        RECT 99.000 101.330 99.260 101.650 ;
        RECT 100.380 101.330 100.640 101.650 ;
        RECT 98.080 98.950 98.340 99.270 ;
        RECT 97.620 98.270 97.880 98.590 ;
        RECT 97.680 96.890 97.820 98.270 ;
        RECT 97.620 96.570 97.880 96.890 ;
        RECT 98.140 94.850 98.280 98.950 ;
        RECT 98.080 94.530 98.340 94.850 ;
        RECT 99.060 94.170 99.200 101.330 ;
        RECT 99.580 100.455 101.460 100.825 ;
        RECT 101.820 99.270 101.960 102.010 ;
        RECT 101.760 98.950 102.020 99.270 ;
        RECT 102.740 98.930 102.880 103.710 ;
        RECT 102.680 98.610 102.940 98.930 ;
        RECT 101.300 98.270 101.560 98.590 ;
        RECT 101.760 98.270 102.020 98.590 ;
        RECT 101.360 97.230 101.500 98.270 ;
        RECT 101.300 96.910 101.560 97.230 ;
        RECT 99.580 95.015 101.460 95.385 ;
        RECT 99.000 93.850 99.260 94.170 ;
        RECT 101.820 93.830 101.960 98.270 ;
        RECT 102.220 96.570 102.480 96.890 ;
        RECT 101.760 93.510 102.020 93.830 ;
        RECT 94.400 91.130 94.660 91.450 ;
        RECT 96.240 91.130 96.500 91.450 ;
        RECT 94.460 86.350 94.600 91.130 ;
        RECT 99.580 89.575 101.460 89.945 ;
        RECT 94.400 86.030 94.660 86.350 ;
        RECT 94.460 80.570 94.600 86.030 ;
        RECT 94.860 85.010 95.120 85.330 ;
        RECT 94.920 83.630 95.060 85.010 ;
        RECT 102.280 84.990 102.420 96.570 ;
        RECT 102.740 95.870 102.880 98.610 ;
        RECT 102.680 95.550 102.940 95.870 ;
        RECT 102.740 93.490 102.880 95.550 ;
        RECT 102.680 93.170 102.940 93.490 ;
        RECT 104.120 86.090 104.260 120.370 ;
        RECT 104.580 86.690 104.720 120.710 ;
        RECT 105.900 114.590 106.160 114.910 ;
        RECT 105.440 112.890 105.700 113.210 ;
        RECT 105.500 109.470 105.640 112.890 ;
        RECT 105.960 110.150 106.100 114.590 ;
        RECT 105.900 109.830 106.160 110.150 ;
        RECT 105.440 109.150 105.700 109.470 ;
        RECT 105.500 104.370 105.640 109.150 ;
        RECT 105.440 104.050 105.700 104.370 ;
        RECT 107.280 98.950 107.540 99.270 ;
        RECT 105.900 96.230 106.160 96.550 ;
        RECT 105.960 88.390 106.100 96.230 ;
        RECT 107.340 94.850 107.480 98.950 ;
        RECT 107.740 95.550 108.000 95.870 ;
        RECT 107.280 94.530 107.540 94.850 ;
        RECT 107.800 93.830 107.940 95.550 ;
        RECT 107.740 93.510 108.000 93.830 ;
        RECT 105.900 88.070 106.160 88.390 ;
        RECT 104.980 87.390 105.240 87.710 ;
        RECT 104.520 86.370 104.780 86.690 ;
        RECT 103.600 85.690 103.860 86.010 ;
        RECT 104.120 85.950 104.720 86.090 ;
        RECT 102.680 85.350 102.940 85.670 ;
        RECT 95.780 84.670 96.040 84.990 ;
        RECT 102.220 84.670 102.480 84.990 ;
        RECT 94.860 83.310 95.120 83.630 ;
        RECT 95.840 82.950 95.980 84.670 ;
        RECT 99.580 84.135 101.460 84.505 ;
        RECT 95.780 82.630 96.040 82.950 ;
        RECT 96.700 82.690 96.960 82.950 ;
        RECT 96.300 82.630 96.960 82.690 ;
        RECT 96.300 82.550 96.900 82.630 ;
        RECT 96.300 82.270 96.440 82.550 ;
        RECT 96.240 81.950 96.500 82.270 ;
        RECT 96.300 80.910 96.440 81.950 ;
        RECT 96.240 80.590 96.500 80.910 ;
        RECT 94.400 80.250 94.660 80.570 ;
        RECT 96.700 80.250 96.960 80.570 ;
        RECT 93.940 75.490 94.200 75.810 ;
        RECT 96.240 75.490 96.500 75.810 ;
        RECT 93.940 74.470 94.200 74.790 ;
        RECT 94.000 72.070 94.140 74.470 ;
        RECT 93.940 71.750 94.200 72.070 ;
        RECT 94.400 71.750 94.660 72.070 ;
        RECT 94.460 71.390 94.600 71.750 ;
        RECT 94.400 71.070 94.660 71.390 ;
        RECT 96.300 70.370 96.440 75.490 ;
        RECT 96.240 70.050 96.500 70.370 ;
        RECT 96.760 66.370 96.900 80.250 ;
        RECT 97.160 79.910 97.420 80.230 ;
        RECT 97.220 73.090 97.360 79.910 ;
        RECT 99.580 78.695 101.460 79.065 ;
        RECT 101.300 77.190 101.560 77.510 ;
        RECT 102.220 77.190 102.480 77.510 ;
        RECT 100.840 76.850 101.100 77.170 ;
        RECT 100.900 75.130 101.040 76.850 ;
        RECT 101.360 75.130 101.500 77.190 ;
        RECT 100.840 74.810 101.100 75.130 ;
        RECT 101.300 74.810 101.560 75.130 ;
        RECT 97.620 74.470 97.880 74.790 ;
        RECT 97.160 72.770 97.420 73.090 ;
        RECT 97.160 72.090 97.420 72.410 ;
        RECT 97.220 66.970 97.360 72.090 ;
        RECT 97.160 66.650 97.420 66.970 ;
        RECT 97.680 66.630 97.820 74.470 ;
        RECT 102.280 74.450 102.420 77.190 ;
        RECT 99.000 74.130 99.260 74.450 ;
        RECT 102.220 74.130 102.480 74.450 ;
        RECT 98.080 68.350 98.340 68.670 ;
        RECT 98.540 68.350 98.800 68.670 ;
        RECT 96.760 66.230 97.360 66.370 ;
        RECT 97.620 66.310 97.880 66.630 ;
        RECT 94.400 65.630 94.660 65.950 ;
        RECT 94.460 61.190 94.600 65.630 ;
        RECT 96.700 64.270 96.960 64.590 ;
        RECT 96.760 62.210 96.900 64.270 ;
        RECT 96.700 61.890 96.960 62.210 ;
        RECT 94.400 60.870 94.660 61.190 ;
        RECT 93.480 56.450 93.740 56.770 ;
        RECT 91.640 56.110 91.900 56.430 ;
        RECT 91.180 53.390 91.440 53.710 ;
        RECT 91.700 53.370 91.840 56.110 ;
        RECT 97.220 54.050 97.360 66.230 ;
        RECT 97.680 63.570 97.820 66.310 ;
        RECT 98.140 64.930 98.280 68.350 ;
        RECT 98.600 66.630 98.740 68.350 ;
        RECT 98.540 66.310 98.800 66.630 ;
        RECT 98.080 64.610 98.340 64.930 ;
        RECT 99.060 64.250 99.200 74.130 ;
        RECT 99.580 73.255 101.460 73.625 ;
        RECT 99.920 71.750 100.180 72.070 ;
        RECT 99.460 71.070 99.720 71.390 ;
        RECT 99.520 68.670 99.660 71.070 ;
        RECT 99.980 70.370 100.120 71.750 ;
        RECT 100.380 71.410 100.640 71.730 ;
        RECT 99.920 70.050 100.180 70.370 ;
        RECT 100.440 68.920 100.580 71.410 ;
        RECT 102.220 69.030 102.480 69.350 ;
        RECT 100.440 68.780 101.960 68.920 ;
        RECT 99.460 68.350 99.720 68.670 ;
        RECT 99.580 67.815 101.460 68.185 ;
        RECT 101.820 67.650 101.960 68.780 ;
        RECT 102.280 67.650 102.420 69.030 ;
        RECT 101.760 67.330 102.020 67.650 ;
        RECT 102.220 67.330 102.480 67.650 ;
        RECT 100.840 65.970 101.100 66.290 ;
        RECT 100.900 64.930 101.040 65.970 ;
        RECT 100.840 64.610 101.100 64.930 ;
        RECT 99.000 63.930 99.260 64.250 ;
        RECT 97.620 63.250 97.880 63.570 ;
        RECT 99.580 62.375 101.460 62.745 ;
        RECT 97.620 60.870 97.880 61.190 ;
        RECT 97.160 53.730 97.420 54.050 ;
        RECT 91.640 53.050 91.900 53.370 ;
        RECT 90.720 51.010 90.980 51.330 ;
        RECT 89.800 50.330 90.060 50.650 ;
        RECT 89.860 48.610 90.000 50.330 ;
        RECT 89.340 48.290 89.600 48.610 ;
        RECT 89.800 48.290 90.060 48.610 ;
        RECT 88.420 47.950 88.680 48.270 ;
        RECT 87.960 45.570 88.220 45.890 ;
        RECT 88.480 44.870 88.620 47.950 ;
        RECT 91.180 47.840 91.440 47.930 ;
        RECT 91.700 47.840 91.840 53.050 ;
        RECT 92.560 52.710 92.820 53.030 ;
        RECT 91.180 47.700 91.840 47.840 ;
        RECT 92.620 47.840 92.760 52.710 ;
        RECT 95.320 51.010 95.580 51.330 ;
        RECT 95.380 47.930 95.520 51.010 ;
        RECT 97.680 50.310 97.820 60.870 ;
        RECT 101.820 58.810 101.960 67.330 ;
        RECT 98.540 58.490 98.800 58.810 ;
        RECT 101.760 58.490 102.020 58.810 ;
        RECT 98.600 55.750 98.740 58.490 ;
        RECT 102.220 58.150 102.480 58.470 ;
        RECT 99.580 56.935 101.460 57.305 ;
        RECT 98.540 55.430 98.800 55.750 ;
        RECT 99.000 55.430 99.260 55.750 ;
        RECT 99.060 54.050 99.200 55.430 ;
        RECT 102.280 55.410 102.420 58.150 ;
        RECT 102.740 56.770 102.880 85.350 ;
        RECT 103.660 78.530 103.800 85.690 ;
        RECT 104.060 82.630 104.320 82.950 ;
        RECT 103.600 78.210 103.860 78.530 ;
        RECT 104.120 78.190 104.260 82.630 ;
        RECT 104.580 82.270 104.720 85.950 ;
        RECT 105.040 83.970 105.180 87.390 ;
        RECT 105.960 86.010 106.100 88.070 ;
        RECT 106.360 87.390 106.620 87.710 ;
        RECT 105.900 85.690 106.160 86.010 ;
        RECT 105.440 84.670 105.700 84.990 ;
        RECT 104.980 83.650 105.240 83.970 ;
        RECT 104.520 81.950 104.780 82.270 ;
        RECT 105.500 79.890 105.640 84.670 ;
        RECT 106.420 83.970 106.560 87.390 ;
        RECT 106.360 83.650 106.620 83.970 ;
        RECT 105.900 82.970 106.160 83.290 ;
        RECT 105.440 79.570 105.700 79.890 ;
        RECT 104.060 77.870 104.320 78.190 ;
        RECT 103.140 77.190 103.400 77.510 ;
        RECT 104.520 77.190 104.780 77.510 ;
        RECT 103.200 75.810 103.340 77.190 ;
        RECT 104.060 76.850 104.320 77.170 ;
        RECT 103.140 75.490 103.400 75.810 ;
        RECT 104.120 75.130 104.260 76.850 ;
        RECT 104.580 75.130 104.720 77.190 ;
        RECT 104.060 74.810 104.320 75.130 ;
        RECT 104.520 74.810 104.780 75.130 ;
        RECT 103.600 74.130 103.860 74.450 ;
        RECT 103.140 73.790 103.400 74.110 ;
        RECT 103.200 69.770 103.340 73.790 ;
        RECT 103.660 71.390 103.800 74.130 ;
        RECT 103.600 71.070 103.860 71.390 ;
        RECT 103.660 70.370 103.800 71.070 ;
        RECT 103.600 70.050 103.860 70.370 ;
        RECT 103.200 69.690 103.800 69.770 ;
        RECT 103.200 69.630 103.860 69.690 ;
        RECT 103.600 69.370 103.860 69.630 ;
        RECT 103.660 67.050 103.800 69.370 ;
        RECT 103.200 66.910 103.800 67.050 ;
        RECT 103.200 64.250 103.340 66.910 ;
        RECT 103.140 63.930 103.400 64.250 ;
        RECT 104.520 60.870 104.780 61.190 ;
        RECT 104.580 58.130 104.720 60.870 ;
        RECT 105.960 59.490 106.100 82.970 ;
        RECT 106.360 82.630 106.620 82.950 ;
        RECT 106.420 75.810 106.560 82.630 ;
        RECT 108.260 81.250 108.400 121.050 ;
        RECT 110.100 121.030 110.240 124.110 ;
        RECT 108.660 120.710 108.920 121.030 ;
        RECT 110.040 120.710 110.300 121.030 ;
        RECT 108.720 82.270 108.860 120.710 ;
        RECT 110.100 115.590 110.240 120.710 ;
        RECT 111.940 120.690 112.080 128.870 ;
        RECT 112.800 124.110 113.060 124.430 ;
        RECT 112.860 123.070 113.000 124.110 ;
        RECT 113.780 123.750 113.920 139.870 ;
        RECT 114.580 130.375 116.460 130.745 ;
        RECT 120.220 129.870 120.360 139.870 ;
        RECT 119.700 129.550 119.960 129.870 ;
        RECT 120.160 129.550 120.420 129.870 ;
        RECT 114.580 124.935 116.460 125.305 ;
        RECT 119.760 124.090 119.900 129.550 ;
        RECT 119.700 123.770 119.960 124.090 ;
        RECT 120.620 123.770 120.880 124.090 ;
        RECT 113.720 123.430 113.980 123.750 ;
        RECT 112.800 122.750 113.060 123.070 ;
        RECT 118.780 122.750 119.040 123.070 ;
        RECT 118.840 120.690 118.980 122.750 ;
        RECT 120.680 122.050 120.820 123.770 ;
        RECT 120.620 121.730 120.880 122.050 ;
        RECT 126.660 121.370 126.800 139.870 ;
        RECT 126.600 121.050 126.860 121.370 ;
        RECT 111.880 120.370 112.140 120.690 ;
        RECT 118.780 120.370 119.040 120.690 ;
        RECT 114.580 119.495 116.460 119.865 ;
        RECT 119.240 115.610 119.500 115.930 ;
        RECT 110.040 115.270 110.300 115.590 ;
        RECT 110.100 112.870 110.240 115.270 ;
        RECT 118.320 114.590 118.580 114.910 ;
        RECT 114.580 114.055 116.460 114.425 ;
        RECT 117.860 113.230 118.120 113.550 ;
        RECT 110.040 112.550 110.300 112.870 ;
        RECT 112.800 112.550 113.060 112.870 ;
        RECT 110.100 110.490 110.240 112.550 ;
        RECT 110.040 110.170 110.300 110.490 ;
        RECT 109.580 109.490 109.840 109.810 ;
        RECT 109.640 108.450 109.780 109.490 ;
        RECT 109.580 108.130 109.840 108.450 ;
        RECT 110.100 104.030 110.240 110.170 ;
        RECT 112.860 108.450 113.000 112.550 ;
        RECT 117.400 111.870 117.660 112.190 ;
        RECT 114.180 110.170 114.440 110.490 ;
        RECT 117.460 110.470 117.600 111.870 ;
        RECT 117.920 110.490 118.060 113.230 ;
        RECT 117.000 110.330 117.600 110.470 ;
        RECT 113.720 109.150 113.980 109.470 ;
        RECT 112.800 108.130 113.060 108.450 ;
        RECT 113.780 107.770 113.920 109.150 ;
        RECT 114.240 108.360 114.380 110.170 ;
        RECT 117.000 109.470 117.140 110.330 ;
        RECT 117.860 110.170 118.120 110.490 ;
        RECT 116.940 109.150 117.200 109.470 ;
        RECT 114.580 108.615 116.460 108.985 ;
        RECT 114.240 108.220 114.840 108.360 ;
        RECT 113.720 107.450 113.980 107.770 ;
        RECT 114.180 107.450 114.440 107.770 ;
        RECT 114.240 107.170 114.380 107.450 ;
        RECT 114.700 107.430 114.840 108.220 ;
        RECT 117.000 107.430 117.140 109.150 ;
        RECT 118.380 107.770 118.520 114.590 ;
        RECT 119.300 111.170 119.440 115.610 ;
        RECT 122.460 114.930 122.720 115.250 ;
        RECT 119.240 110.850 119.500 111.170 ;
        RECT 122.520 110.490 122.660 114.930 ;
        RECT 122.460 110.170 122.720 110.490 ;
        RECT 118.780 109.830 119.040 110.150 ;
        RECT 119.240 109.830 119.500 110.150 ;
        RECT 118.320 107.450 118.580 107.770 ;
        RECT 113.780 107.030 114.380 107.170 ;
        RECT 114.640 107.110 114.900 107.430 ;
        RECT 116.940 107.110 117.200 107.430 ;
        RECT 110.040 103.710 110.300 104.030 ;
        RECT 110.100 99.610 110.240 103.710 ;
        RECT 110.960 100.990 111.220 101.310 ;
        RECT 110.040 99.290 110.300 99.610 ;
        RECT 110.100 97.230 110.240 99.290 ;
        RECT 111.020 98.930 111.160 100.990 ;
        RECT 113.780 98.930 113.920 107.030 ;
        RECT 114.700 106.490 114.840 107.110 ;
        RECT 114.240 106.350 114.840 106.490 ;
        RECT 114.240 105.050 114.380 106.350 ;
        RECT 114.180 104.730 114.440 105.050 ;
        RECT 114.240 99.610 114.380 104.730 ;
        RECT 114.580 103.175 116.460 103.545 ;
        RECT 117.000 101.990 117.140 107.110 ;
        RECT 118.840 102.330 118.980 109.830 ;
        RECT 119.300 108.450 119.440 109.830 ;
        RECT 119.240 108.130 119.500 108.450 ;
        RECT 118.780 102.010 119.040 102.330 ;
        RECT 116.940 101.670 117.200 101.990 ;
        RECT 118.840 99.610 118.980 102.010 ;
        RECT 114.180 99.290 114.440 99.610 ;
        RECT 118.780 99.290 119.040 99.610 ;
        RECT 110.960 98.610 111.220 98.930 ;
        RECT 113.720 98.610 113.980 98.930 ;
        RECT 111.420 98.270 111.680 98.590 ;
        RECT 111.480 97.570 111.620 98.270 ;
        RECT 111.420 97.250 111.680 97.570 ;
        RECT 110.040 96.910 110.300 97.230 ;
        RECT 110.100 88.730 110.240 96.910 ;
        RECT 111.420 96.570 111.680 96.890 ;
        RECT 110.960 90.790 111.220 91.110 ;
        RECT 110.500 90.110 110.760 90.430 ;
        RECT 110.040 88.410 110.300 88.730 ;
        RECT 110.100 86.010 110.240 88.410 ;
        RECT 110.560 88.390 110.700 90.110 ;
        RECT 110.500 88.070 110.760 88.390 ;
        RECT 111.020 88.050 111.160 90.790 ;
        RECT 111.480 89.410 111.620 96.570 ;
        RECT 113.780 96.210 113.920 98.610 ;
        RECT 114.240 96.290 114.380 99.290 ;
        RECT 116.940 98.270 117.200 98.590 ;
        RECT 114.580 97.735 116.460 98.105 ;
        RECT 114.640 96.290 114.900 96.550 ;
        RECT 114.240 96.230 114.900 96.290 ;
        RECT 113.720 95.890 113.980 96.210 ;
        RECT 114.240 96.150 114.840 96.230 ;
        RECT 114.240 91.530 114.380 96.150 ;
        RECT 117.000 95.870 117.140 98.270 ;
        RECT 116.940 95.550 117.200 95.870 ;
        RECT 114.580 92.295 116.460 92.665 ;
        RECT 117.000 91.530 117.140 95.550 ;
        RECT 118.840 93.830 118.980 99.290 ;
        RECT 119.240 98.270 119.500 98.590 ;
        RECT 122.460 98.270 122.720 98.590 ;
        RECT 119.300 97.570 119.440 98.270 ;
        RECT 119.240 97.250 119.500 97.570 ;
        RECT 122.520 97.230 122.660 98.270 ;
        RECT 122.460 96.910 122.720 97.230 ;
        RECT 118.780 93.510 119.040 93.830 ;
        RECT 118.320 92.830 118.580 93.150 ;
        RECT 114.240 91.390 114.840 91.530 ;
        RECT 114.700 90.770 114.840 91.390 ;
        RECT 116.540 91.390 117.140 91.530 ;
        RECT 116.540 91.110 116.680 91.390 ;
        RECT 117.400 91.130 117.660 91.450 ;
        RECT 116.480 90.790 116.740 91.110 ;
        RECT 114.640 90.450 114.900 90.770 ;
        RECT 111.420 89.090 111.680 89.410 ;
        RECT 110.960 87.730 111.220 88.050 ;
        RECT 117.460 87.710 117.600 91.130 ;
        RECT 117.860 87.730 118.120 88.050 ;
        RECT 117.400 87.390 117.660 87.710 ;
        RECT 114.580 86.855 116.460 87.225 ;
        RECT 117.460 86.690 117.600 87.390 ;
        RECT 117.400 86.370 117.660 86.690 ;
        RECT 110.040 85.690 110.300 86.010 ;
        RECT 112.800 83.310 113.060 83.630 ;
        RECT 108.660 81.950 108.920 82.270 ;
        RECT 108.200 80.930 108.460 81.250 ;
        RECT 110.500 77.190 110.760 77.510 ;
        RECT 112.340 77.190 112.600 77.510 ;
        RECT 110.560 75.810 110.700 77.190 ;
        RECT 106.360 75.490 106.620 75.810 ;
        RECT 110.500 75.490 110.760 75.810 ;
        RECT 111.420 74.810 111.680 75.130 ;
        RECT 110.040 74.470 110.300 74.790 ;
        RECT 110.500 74.470 110.760 74.790 ;
        RECT 106.820 71.410 107.080 71.730 ;
        RECT 106.880 70.370 107.020 71.410 ;
        RECT 106.820 70.050 107.080 70.370 ;
        RECT 110.100 66.630 110.240 74.470 ;
        RECT 110.560 69.010 110.700 74.470 ;
        RECT 111.480 71.390 111.620 74.810 ;
        RECT 112.400 72.070 112.540 77.190 ;
        RECT 112.340 71.750 112.600 72.070 ;
        RECT 111.420 71.070 111.680 71.390 ;
        RECT 110.500 68.690 110.760 69.010 ;
        RECT 110.040 66.310 110.300 66.630 ;
        RECT 110.100 64.930 110.240 66.310 ;
        RECT 110.040 64.610 110.300 64.930 ;
        RECT 110.560 63.910 110.700 68.690 ;
        RECT 112.400 63.910 112.540 71.750 ;
        RECT 106.360 63.590 106.620 63.910 ;
        RECT 110.500 63.590 110.760 63.910 ;
        RECT 112.340 63.590 112.600 63.910 ;
        RECT 106.420 62.210 106.560 63.590 ;
        RECT 106.360 61.890 106.620 62.210 ;
        RECT 112.400 62.170 112.540 63.590 ;
        RECT 111.940 62.030 112.540 62.170 ;
        RECT 111.940 61.530 112.080 62.030 ;
        RECT 111.880 61.210 112.140 61.530 ;
        RECT 110.960 60.530 111.220 60.850 ;
        RECT 111.020 59.490 111.160 60.530 ;
        RECT 105.900 59.170 106.160 59.490 ;
        RECT 110.960 59.170 111.220 59.490 ;
        RECT 107.740 58.830 108.000 59.150 ;
        RECT 104.980 58.490 105.240 58.810 ;
        RECT 105.440 58.490 105.700 58.810 ;
        RECT 105.900 58.490 106.160 58.810 ;
        RECT 104.520 57.810 104.780 58.130 ;
        RECT 102.680 56.450 102.940 56.770 ;
        RECT 102.220 55.090 102.480 55.410 ;
        RECT 99.000 53.730 99.260 54.050 ;
        RECT 98.080 52.710 98.340 53.030 ;
        RECT 99.060 52.770 99.200 53.730 ;
        RECT 102.220 53.390 102.480 53.710 ;
        RECT 98.140 51.330 98.280 52.710 ;
        RECT 98.600 52.630 99.200 52.770 ;
        RECT 98.080 51.010 98.340 51.330 ;
        RECT 98.600 50.650 98.740 52.630 ;
        RECT 99.000 52.030 99.260 52.350 ;
        RECT 98.540 50.330 98.800 50.650 ;
        RECT 99.060 50.310 99.200 52.030 ;
        RECT 99.580 51.495 101.460 51.865 ;
        RECT 97.620 49.990 97.880 50.310 ;
        RECT 99.000 49.990 99.260 50.310 ;
        RECT 99.920 49.310 100.180 49.630 ;
        RECT 99.980 48.270 100.120 49.310 ;
        RECT 99.920 47.950 100.180 48.270 ;
        RECT 92.620 47.700 93.220 47.840 ;
        RECT 91.180 47.610 91.440 47.700 ;
        RECT 90.260 47.270 90.520 47.590 ;
        RECT 88.420 44.550 88.680 44.870 ;
        RECT 88.880 44.550 89.140 44.870 ;
        RECT 87.040 44.210 87.300 44.530 ;
        RECT 84.580 43.335 86.460 43.705 ;
        RECT 87.100 43.170 87.240 44.210 ;
        RECT 87.040 42.850 87.300 43.170 ;
        RECT 88.940 42.490 89.080 44.550 ;
        RECT 89.800 43.870 90.060 44.190 ;
        RECT 88.880 42.170 89.140 42.490 ;
        RECT 86.580 41.830 86.840 42.150 ;
        RECT 85.200 41.150 85.460 41.470 ;
        RECT 85.260 39.770 85.400 41.150 ;
        RECT 86.640 39.770 86.780 41.830 ;
        RECT 83.360 39.450 83.620 39.770 ;
        RECT 85.200 39.450 85.460 39.770 ;
        RECT 86.580 39.450 86.840 39.770 ;
        RECT 81.980 38.430 82.240 38.750 ;
        RECT 82.040 37.390 82.180 38.430 ;
        RECT 81.980 37.070 82.240 37.390 ;
        RECT 80.600 36.730 80.860 37.050 ;
        RECT 83.420 36.710 83.560 39.450 ;
        RECT 89.860 39.430 90.000 43.870 ;
        RECT 90.320 39.430 90.460 47.270 ;
        RECT 91.240 44.870 91.380 47.610 ;
        RECT 92.100 47.330 92.360 47.590 ;
        RECT 92.100 47.270 92.760 47.330 ;
        RECT 92.160 47.190 92.760 47.270 ;
        RECT 91.180 44.550 91.440 44.870 ;
        RECT 92.100 44.210 92.360 44.530 ;
        RECT 91.640 41.490 91.900 41.810 ;
        RECT 89.800 39.110 90.060 39.430 ;
        RECT 90.260 39.110 90.520 39.430 ;
        RECT 84.580 37.895 86.460 38.265 ;
        RECT 76.000 36.390 76.260 36.710 ;
        RECT 83.360 36.450 83.620 36.710 ;
        RECT 83.360 36.390 84.020 36.450 ;
        RECT 83.420 36.310 84.020 36.390 ;
        RECT 90.320 36.370 90.460 39.110 ;
        RECT 91.700 37.390 91.840 41.490 ;
        RECT 91.640 37.070 91.900 37.390 ;
        RECT 92.160 36.710 92.300 44.210 ;
        RECT 92.620 41.810 92.760 47.190 ;
        RECT 93.080 42.490 93.220 47.700 ;
        RECT 95.320 47.610 95.580 47.930 ;
        RECT 99.580 46.055 101.460 46.425 ;
        RECT 102.280 44.870 102.420 53.390 ;
        RECT 102.680 52.710 102.940 53.030 ;
        RECT 102.740 51.330 102.880 52.710 ;
        RECT 102.680 51.010 102.940 51.330 ;
        RECT 103.600 50.330 103.860 50.650 ;
        RECT 103.660 45.210 103.800 50.330 ;
        RECT 103.600 44.890 103.860 45.210 ;
        RECT 102.220 44.550 102.480 44.870 ;
        RECT 96.240 42.510 96.500 42.830 ;
        RECT 93.020 42.170 93.280 42.490 ;
        RECT 92.560 41.490 92.820 41.810 ;
        RECT 92.620 39.770 92.760 41.490 ;
        RECT 92.560 39.450 92.820 39.770 ;
        RECT 92.100 36.390 92.360 36.710 ;
        RECT 69.580 35.175 71.460 35.545 ;
        RECT 72.780 34.010 73.040 34.330 ;
        RECT 72.840 31.610 72.980 34.010 ;
        RECT 83.880 33.990 84.020 36.310 ;
        RECT 90.260 36.050 90.520 36.370 ;
        RECT 93.080 34.330 93.220 42.170 ;
        RECT 93.940 41.490 94.200 41.810 ;
        RECT 93.480 38.430 93.740 38.750 ;
        RECT 93.540 37.730 93.680 38.430 ;
        RECT 93.480 37.410 93.740 37.730 ;
        RECT 93.020 34.010 93.280 34.330 ;
        RECT 94.000 33.990 94.140 41.490 ;
        RECT 96.300 39.430 96.440 42.510 ;
        RECT 103.660 42.150 103.800 44.890 ;
        RECT 105.040 43.170 105.180 58.490 ;
        RECT 105.500 55.070 105.640 58.490 ;
        RECT 105.960 56.090 106.100 58.490 ;
        RECT 107.800 56.090 107.940 58.830 ;
        RECT 111.420 58.490 111.680 58.810 ;
        RECT 111.480 58.130 111.620 58.490 ;
        RECT 111.420 57.810 111.680 58.130 ;
        RECT 105.900 55.770 106.160 56.090 ;
        RECT 107.740 55.770 108.000 56.090 ;
        RECT 105.440 54.750 105.700 55.070 ;
        RECT 105.500 53.280 105.640 54.750 ;
        RECT 105.900 53.280 106.160 53.370 ;
        RECT 105.500 53.140 106.160 53.280 ;
        RECT 105.900 53.050 106.160 53.140 ;
        RECT 105.900 52.370 106.160 52.690 ;
        RECT 105.960 50.310 106.100 52.370 ;
        RECT 107.800 52.350 107.940 55.770 ;
        RECT 111.480 55.750 111.620 57.810 ;
        RECT 111.940 56.090 112.080 61.210 ;
        RECT 111.880 55.770 112.140 56.090 ;
        RECT 111.420 55.430 111.680 55.750 ;
        RECT 107.740 52.030 108.000 52.350 ;
        RECT 107.800 50.650 107.940 52.030 ;
        RECT 107.740 50.330 108.000 50.650 ;
        RECT 105.900 49.990 106.160 50.310 ;
        RECT 105.440 46.590 105.700 46.910 ;
        RECT 105.500 44.870 105.640 46.590 ;
        RECT 105.440 44.550 105.700 44.870 ;
        RECT 105.900 43.870 106.160 44.190 ;
        RECT 104.980 42.850 105.240 43.170 ;
        RECT 98.540 41.830 98.800 42.150 ;
        RECT 103.600 41.830 103.860 42.150 ;
        RECT 97.160 41.490 97.420 41.810 ;
        RECT 96.240 39.110 96.500 39.430 ;
        RECT 94.400 38.430 94.660 38.750 ;
        RECT 94.460 35.010 94.600 38.430 ;
        RECT 96.700 36.390 96.960 36.710 ;
        RECT 94.400 34.690 94.660 35.010 ;
        RECT 83.820 33.670 84.080 33.990 ;
        RECT 93.940 33.670 94.200 33.990 ;
        RECT 69.100 31.290 69.360 31.610 ;
        RECT 72.780 31.290 73.040 31.610 ;
        RECT 64.040 30.950 64.300 31.270 ;
        RECT 65.420 30.950 65.680 31.270 ;
        RECT 63.580 30.610 63.840 30.930 ;
        RECT 61.740 28.910 62.000 29.230 ;
        RECT 63.120 28.910 63.380 29.230 ;
        RECT 63.180 28.550 63.320 28.910 ;
        RECT 63.640 28.550 63.780 30.610 ;
        RECT 63.120 28.230 63.380 28.550 ;
        RECT 63.580 28.230 63.840 28.550 ;
        RECT 61.740 27.550 62.000 27.870 ;
        RECT 62.660 27.550 62.920 27.870 ;
        RECT 61.280 26.530 61.540 26.850 ;
        RECT 59.900 25.940 60.560 26.080 ;
        RECT 59.900 25.850 60.160 25.940 ;
        RECT 60.820 25.850 61.080 26.170 ;
        RECT 58.060 25.510 58.320 25.830 ;
        RECT 61.800 25.150 61.940 27.550 ;
        RECT 62.720 26.170 62.860 27.550 ;
        RECT 63.180 26.170 63.320 28.230 ;
        RECT 62.660 25.850 62.920 26.170 ;
        RECT 63.120 25.850 63.380 26.170 ;
        RECT 64.100 25.150 64.240 30.950 ;
        RECT 65.480 29.230 65.620 30.950 ;
        RECT 66.340 30.270 66.600 30.590 ;
        RECT 66.800 30.270 67.060 30.590 ;
        RECT 65.420 28.910 65.680 29.230 ;
        RECT 65.880 25.510 66.140 25.830 ;
        RECT 61.740 24.830 62.000 25.150 ;
        RECT 64.040 24.830 64.300 25.150 ;
        RECT 9.580 24.295 11.460 24.665 ;
        RECT 39.580 24.295 41.460 24.665 ;
        RECT 65.940 24.130 66.080 25.510 ;
        RECT 65.880 23.810 66.140 24.130 ;
        RECT 66.400 23.110 66.540 30.270 ;
        RECT 66.860 28.550 67.000 30.270 ;
        RECT 69.160 29.570 69.300 31.290 ;
        RECT 69.580 29.735 71.460 30.105 ;
        RECT 69.100 29.250 69.360 29.570 ;
        RECT 66.800 28.230 67.060 28.550 ;
        RECT 71.860 25.510 72.120 25.830 ;
        RECT 69.580 24.295 71.460 24.665 ;
        RECT 71.920 24.130 72.060 25.510 ;
        RECT 71.860 23.810 72.120 24.130 ;
        RECT 72.840 23.110 72.980 31.290 ;
        RECT 73.240 30.270 73.500 30.590 ;
        RECT 73.300 28.210 73.440 30.270 ;
        RECT 83.880 28.890 84.020 33.670 ;
        RECT 96.760 33.310 96.900 36.390 ;
        RECT 97.220 33.990 97.360 41.490 ;
        RECT 98.080 39.110 98.340 39.430 ;
        RECT 97.620 38.430 97.880 38.750 ;
        RECT 97.160 33.670 97.420 33.990 ;
        RECT 97.680 33.650 97.820 38.430 ;
        RECT 98.140 35.010 98.280 39.110 ;
        RECT 98.600 37.730 98.740 41.830 ;
        RECT 99.580 40.615 101.460 40.985 ;
        RECT 105.040 40.450 105.180 42.850 ;
        RECT 105.960 42.490 106.100 43.870 ;
        RECT 105.900 42.170 106.160 42.490 ;
        RECT 104.980 40.130 105.240 40.450 ;
        RECT 107.800 39.770 107.940 50.330 ;
        RECT 109.120 49.650 109.380 49.970 ;
        RECT 109.180 48.610 109.320 49.650 ;
        RECT 110.960 49.310 111.220 49.630 ;
        RECT 109.120 48.290 109.380 48.610 ;
        RECT 111.020 47.930 111.160 49.310 ;
        RECT 110.960 47.610 111.220 47.930 ;
        RECT 111.480 44.870 111.620 55.430 ;
        RECT 111.880 55.090 112.140 55.410 ;
        RECT 111.940 53.710 112.080 55.090 ;
        RECT 112.860 54.050 113.000 83.310 ;
        RECT 117.920 82.950 118.060 87.730 ;
        RECT 118.380 86.350 118.520 92.830 ;
        RECT 118.320 86.030 118.580 86.350 ;
        RECT 118.840 83.290 118.980 93.510 ;
        RECT 120.620 91.130 120.880 91.450 ;
        RECT 120.680 88.730 120.820 91.130 ;
        RECT 122.920 90.110 123.180 90.430 ;
        RECT 120.620 88.410 120.880 88.730 ;
        RECT 120.680 86.690 120.820 88.410 ;
        RECT 122.980 88.390 123.120 90.110 ;
        RECT 122.920 88.070 123.180 88.390 ;
        RECT 122.000 87.390 122.260 87.710 ;
        RECT 120.620 86.370 120.880 86.690 ;
        RECT 122.060 85.670 122.200 87.390 ;
        RECT 122.000 85.350 122.260 85.670 ;
        RECT 118.780 82.970 119.040 83.290 ;
        RECT 117.860 82.630 118.120 82.950 ;
        RECT 114.580 81.415 116.460 81.785 ;
        RECT 117.400 76.850 117.660 77.170 ;
        RECT 114.180 76.510 114.440 76.830 ;
        RECT 114.240 74.790 114.380 76.510 ;
        RECT 114.580 75.975 116.460 76.345 ;
        RECT 117.460 75.810 117.600 76.850 ;
        RECT 117.400 75.490 117.660 75.810 ;
        RECT 117.400 74.810 117.660 75.130 ;
        RECT 118.780 74.810 119.040 75.130 ;
        RECT 114.180 74.470 114.440 74.790 ;
        RECT 113.720 73.790 113.980 74.110 ;
        RECT 113.780 72.410 113.920 73.790 ;
        RECT 113.720 72.090 113.980 72.410 ;
        RECT 114.240 69.690 114.380 74.470 ;
        RECT 117.460 72.410 117.600 74.810 ;
        RECT 117.400 72.090 117.660 72.410 ;
        RECT 116.940 71.070 117.200 71.390 ;
        RECT 114.580 70.535 116.460 70.905 ;
        RECT 114.180 69.370 114.440 69.690 ;
        RECT 115.100 68.690 115.360 69.010 ;
        RECT 115.160 66.970 115.300 68.690 ;
        RECT 116.480 68.580 116.740 68.670 ;
        RECT 117.000 68.580 117.140 71.070 ;
        RECT 117.460 70.030 117.600 72.090 ;
        RECT 118.840 70.370 118.980 74.810 ;
        RECT 121.080 71.750 121.340 72.070 ;
        RECT 118.780 70.050 119.040 70.370 ;
        RECT 117.400 69.710 117.660 70.030 ;
        RECT 116.480 68.440 117.140 68.580 ;
        RECT 116.480 68.350 116.740 68.440 ;
        RECT 115.100 66.650 115.360 66.970 ;
        RECT 116.540 66.630 116.680 68.350 ;
        RECT 121.140 66.630 121.280 71.750 ;
        RECT 116.480 66.310 116.740 66.630 ;
        RECT 121.080 66.310 121.340 66.630 ;
        RECT 118.780 65.630 119.040 65.950 ;
        RECT 120.160 65.630 120.420 65.950 ;
        RECT 114.580 65.095 116.460 65.465 ;
        RECT 118.840 63.910 118.980 65.630 ;
        RECT 120.220 64.590 120.360 65.630 ;
        RECT 120.160 64.270 120.420 64.590 ;
        RECT 118.780 63.590 119.040 63.910 ;
        RECT 113.260 62.910 113.520 63.230 ;
        RECT 113.320 60.850 113.460 62.910 ;
        RECT 113.260 60.530 113.520 60.850 ;
        RECT 114.580 59.655 116.460 60.025 ;
        RECT 114.180 58.150 114.440 58.470 ;
        RECT 113.720 57.470 113.980 57.790 ;
        RECT 112.800 53.730 113.060 54.050 ;
        RECT 113.780 53.710 113.920 57.470 ;
        RECT 111.880 53.390 112.140 53.710 ;
        RECT 113.720 53.390 113.980 53.710 ;
        RECT 114.240 53.370 114.380 58.150 ;
        RECT 114.580 54.215 116.460 54.585 ;
        RECT 114.180 53.050 114.440 53.370 ;
        RECT 115.100 53.050 115.360 53.370 ;
        RECT 115.160 51.330 115.300 53.050 ;
        RECT 114.180 51.010 114.440 51.330 ;
        RECT 115.100 51.010 115.360 51.330 ;
        RECT 111.880 49.650 112.140 49.970 ;
        RECT 111.940 45.890 112.080 49.650 ;
        RECT 114.240 47.930 114.380 51.010 ;
        RECT 114.580 48.775 116.460 49.145 ;
        RECT 114.180 47.610 114.440 47.930 ;
        RECT 111.880 45.570 112.140 45.890 ;
        RECT 111.420 44.550 111.680 44.870 ;
        RECT 111.480 42.830 111.620 44.550 ;
        RECT 111.880 44.210 112.140 44.530 ;
        RECT 111.420 42.510 111.680 42.830 ;
        RECT 109.580 41.490 109.840 41.810 ;
        RECT 109.640 39.770 109.780 41.490 ;
        RECT 104.060 39.450 104.320 39.770 ;
        RECT 107.740 39.450 108.000 39.770 ;
        RECT 109.580 39.450 109.840 39.770 ;
        RECT 98.540 37.410 98.800 37.730 ;
        RECT 104.120 37.050 104.260 39.450 ;
        RECT 104.520 38.770 104.780 39.090 ;
        RECT 104.580 37.730 104.720 38.770 ;
        RECT 104.520 37.410 104.780 37.730 ;
        RECT 111.480 37.050 111.620 42.510 ;
        RECT 111.940 42.490 112.080 44.210 ;
        RECT 114.580 43.335 116.460 43.705 ;
        RECT 111.880 42.170 112.140 42.490 ;
        RECT 111.940 40.450 112.080 42.170 ;
        RECT 113.260 41.490 113.520 41.810 ;
        RECT 111.880 40.130 112.140 40.450 ;
        RECT 113.320 39.090 113.460 41.490 ;
        RECT 113.260 38.770 113.520 39.090 ;
        RECT 114.580 37.895 116.460 38.265 ;
        RECT 104.060 36.730 104.320 37.050 ;
        RECT 111.420 36.730 111.680 37.050 ;
        RECT 99.580 35.175 101.460 35.545 ;
        RECT 98.080 34.690 98.340 35.010 ;
        RECT 97.620 33.330 97.880 33.650 ;
        RECT 96.700 32.990 96.960 33.310 ;
        RECT 84.580 32.455 86.460 32.825 ;
        RECT 114.580 32.455 116.460 32.825 ;
        RECT 99.580 29.735 101.460 30.105 ;
        RECT 83.820 28.570 84.080 28.890 ;
        RECT 73.240 27.890 73.500 28.210 ;
        RECT 84.580 27.015 86.460 27.385 ;
        RECT 114.580 27.015 116.460 27.385 ;
        RECT 99.580 24.295 101.460 24.665 ;
        RECT 66.340 22.790 66.600 23.110 ;
        RECT 72.780 22.790 73.040 23.110 ;
        RECT 24.580 21.575 26.460 21.945 ;
        RECT 54.580 21.575 56.460 21.945 ;
        RECT 84.580 21.575 86.460 21.945 ;
        RECT 114.580 21.575 116.460 21.945 ;
        RECT 9.580 18.855 11.460 19.225 ;
        RECT 39.580 18.855 41.460 19.225 ;
        RECT 69.580 18.855 71.460 19.225 ;
        RECT 99.580 18.855 101.460 19.225 ;
        RECT 24.580 16.135 26.460 16.505 ;
        RECT 54.580 16.135 56.460 16.505 ;
        RECT 84.580 16.135 86.460 16.505 ;
        RECT 114.580 16.135 116.460 16.505 ;
        RECT 9.580 13.415 11.460 13.785 ;
        RECT 39.580 13.415 41.460 13.785 ;
        RECT 69.580 13.415 71.460 13.785 ;
        RECT 99.580 13.415 101.460 13.785 ;
        RECT 24.580 10.695 26.460 11.065 ;
        RECT 54.580 10.695 56.460 11.065 ;
        RECT 84.580 10.695 86.460 11.065 ;
        RECT 114.580 10.695 116.460 11.065 ;
      LAYER met3 ;
        RECT 24.530 130.395 26.510 130.725 ;
        RECT 54.530 130.395 56.510 130.725 ;
        RECT 84.530 130.395 86.510 130.725 ;
        RECT 114.530 130.395 116.510 130.725 ;
        RECT 9.530 127.675 11.510 128.005 ;
        RECT 39.530 127.675 41.510 128.005 ;
        RECT 69.530 127.675 71.510 128.005 ;
        RECT 99.530 127.675 101.510 128.005 ;
        RECT 24.530 124.955 26.510 125.285 ;
        RECT 54.530 124.955 56.510 125.285 ;
        RECT 84.530 124.955 86.510 125.285 ;
        RECT 114.530 124.955 116.510 125.285 ;
        RECT 2.000 122.575 2.235 122.905 ;
        RECT 9.530 122.235 11.510 122.565 ;
        RECT 39.530 122.235 41.510 122.565 ;
        RECT 69.530 122.235 71.510 122.565 ;
        RECT 99.530 122.235 101.510 122.565 ;
        RECT 24.530 119.515 26.510 119.845 ;
        RECT 54.530 119.515 56.510 119.845 ;
        RECT 84.530 119.515 86.510 119.845 ;
        RECT 114.530 119.515 116.510 119.845 ;
        RECT 9.530 116.795 11.510 117.125 ;
        RECT 39.530 116.795 41.510 117.125 ;
        RECT 69.530 116.795 71.510 117.125 ;
        RECT 99.530 116.795 101.510 117.125 ;
        RECT 24.530 114.075 26.510 114.405 ;
        RECT 54.530 114.075 56.510 114.405 ;
        RECT 84.530 114.075 86.510 114.405 ;
        RECT 114.530 114.075 116.510 114.405 ;
        RECT 9.530 111.355 11.510 111.685 ;
        RECT 39.530 111.355 41.510 111.685 ;
        RECT 69.530 111.355 71.510 111.685 ;
        RECT 99.530 111.355 101.510 111.685 ;
        RECT 33.645 109.970 33.975 109.985 ;
        RECT 53.425 109.970 53.755 109.985 ;
        RECT 83.325 109.970 83.655 109.985 ;
        RECT 33.645 109.670 83.655 109.970 ;
        RECT 33.645 109.655 33.975 109.670 ;
        RECT 53.425 109.655 53.755 109.670 ;
        RECT 83.325 109.655 83.655 109.670 ;
        RECT 24.530 108.635 26.510 108.965 ;
        RECT 54.530 108.635 56.510 108.965 ;
        RECT 84.530 108.635 86.510 108.965 ;
        RECT 114.530 108.635 116.510 108.965 ;
        RECT 83.325 107.260 83.655 107.265 ;
        RECT 83.070 107.250 83.655 107.260 ;
        RECT 103.105 107.250 103.435 107.265 ;
        RECT 82.690 106.950 103.435 107.250 ;
        RECT 83.070 106.940 83.655 106.950 ;
        RECT 83.325 106.935 83.655 106.940 ;
        RECT 103.105 106.935 103.435 106.950 ;
        RECT 9.530 105.915 11.510 106.245 ;
        RECT 39.530 105.915 41.510 106.245 ;
        RECT 69.530 105.915 71.510 106.245 ;
        RECT 99.530 105.915 101.510 106.245 ;
        RECT 24.530 103.195 26.510 103.525 ;
        RECT 54.530 103.195 56.510 103.525 ;
        RECT 84.530 103.195 86.510 103.525 ;
        RECT 114.530 103.195 116.510 103.525 ;
        RECT 9.530 100.475 11.510 100.805 ;
        RECT 39.530 100.475 41.510 100.805 ;
        RECT 69.530 100.475 71.510 100.805 ;
        RECT 99.530 100.475 101.510 100.805 ;
        RECT 24.530 97.755 26.510 98.085 ;
        RECT 54.530 97.755 56.510 98.085 ;
        RECT 84.530 97.755 86.510 98.085 ;
        RECT 114.530 97.755 116.510 98.085 ;
        RECT 9.530 95.035 11.510 95.365 ;
        RECT 39.530 95.035 41.510 95.365 ;
        RECT 69.530 95.035 71.510 95.365 ;
        RECT 99.530 95.035 101.510 95.365 ;
        RECT 24.530 92.315 26.510 92.645 ;
        RECT 54.530 92.315 56.510 92.645 ;
        RECT 84.530 92.315 86.510 92.645 ;
        RECT 114.530 92.315 116.510 92.645 ;
        RECT 22.605 90.930 22.935 90.945 ;
        RECT 24.905 90.930 25.235 90.945 ;
        RECT 22.605 90.630 25.235 90.930 ;
        RECT 22.605 90.615 22.935 90.630 ;
        RECT 24.905 90.615 25.235 90.630 ;
        RECT 57.310 90.250 57.690 90.260 ;
        RECT 58.485 90.250 58.815 90.265 ;
        RECT 57.310 89.950 58.815 90.250 ;
        RECT 57.310 89.940 57.690 89.950 ;
        RECT 58.485 89.935 58.815 89.950 ;
        RECT 9.530 89.595 11.510 89.925 ;
        RECT 39.530 89.595 41.510 89.925 ;
        RECT 69.530 89.595 71.510 89.925 ;
        RECT 99.530 89.595 101.510 89.925 ;
        RECT 63.750 88.210 64.130 88.220 ;
        RECT 13.650 87.910 64.130 88.210 ;
        RECT 13.650 87.530 13.950 87.910 ;
        RECT 63.750 87.900 64.130 87.910 ;
        RECT 2.000 87.230 13.950 87.530 ;
        RECT 24.530 86.875 26.510 87.205 ;
        RECT 54.530 86.875 56.510 87.205 ;
        RECT 84.530 86.875 86.510 87.205 ;
        RECT 114.530 86.875 116.510 87.205 ;
        RECT 9.530 84.155 11.510 84.485 ;
        RECT 39.530 84.155 41.510 84.485 ;
        RECT 69.530 84.155 71.510 84.485 ;
        RECT 99.530 84.155 101.510 84.485 ;
        RECT 24.530 81.435 26.510 81.765 ;
        RECT 54.530 81.435 56.510 81.765 ;
        RECT 84.530 81.435 86.510 81.765 ;
        RECT 114.530 81.435 116.510 81.765 ;
        RECT 65.385 80.060 65.715 80.065 ;
        RECT 65.385 80.050 65.970 80.060 ;
        RECT 65.160 79.750 65.970 80.050 ;
        RECT 65.385 79.740 65.970 79.750 ;
        RECT 65.385 79.735 65.715 79.740 ;
        RECT 9.530 78.715 11.510 79.045 ;
        RECT 39.530 78.715 41.510 79.045 ;
        RECT 69.530 78.715 71.510 79.045 ;
        RECT 99.530 78.715 101.510 79.045 ;
        RECT 24.530 75.995 26.510 76.325 ;
        RECT 54.530 75.995 56.510 76.325 ;
        RECT 84.530 75.995 86.510 76.325 ;
        RECT 114.530 75.995 116.510 76.325 ;
        RECT 63.750 75.970 64.130 75.980 ;
        RECT 64.925 75.970 65.255 75.985 ;
        RECT 63.750 75.670 65.255 75.970 ;
        RECT 63.750 75.660 64.130 75.670 ;
        RECT 64.925 75.655 65.255 75.670 ;
        RECT 72.030 75.970 72.410 75.980 ;
        RECT 73.665 75.970 73.995 75.985 ;
        RECT 83.070 75.970 83.450 75.980 ;
        RECT 72.030 75.670 83.450 75.970 ;
        RECT 72.030 75.660 72.410 75.670 ;
        RECT 73.665 75.655 73.995 75.670 ;
        RECT 83.070 75.660 83.450 75.670 ;
        RECT 53.885 75.290 54.215 75.305 ;
        RECT 60.785 75.290 61.115 75.305 ;
        RECT 53.885 74.990 61.115 75.290 ;
        RECT 83.110 75.290 83.410 75.660 ;
        RECT 89.510 75.290 89.890 75.300 ;
        RECT 83.110 74.990 89.890 75.290 ;
        RECT 53.885 74.975 54.215 74.990 ;
        RECT 60.785 74.975 61.115 74.990 ;
        RECT 89.510 74.980 89.890 74.990 ;
        RECT 35.945 74.610 36.275 74.625 ;
        RECT 46.985 74.610 47.315 74.625 ;
        RECT 35.945 74.310 47.315 74.610 ;
        RECT 35.945 74.295 36.275 74.310 ;
        RECT 46.985 74.295 47.315 74.310 ;
        RECT 9.530 73.275 11.510 73.605 ;
        RECT 39.530 73.275 41.510 73.605 ;
        RECT 69.530 73.275 71.510 73.605 ;
        RECT 99.530 73.275 101.510 73.605 ;
        RECT 24.530 70.555 26.510 70.885 ;
        RECT 54.530 70.555 56.510 70.885 ;
        RECT 84.530 70.555 86.510 70.885 ;
        RECT 114.530 70.555 116.510 70.885 ;
        RECT 9.530 67.835 11.510 68.165 ;
        RECT 39.530 67.835 41.510 68.165 ;
        RECT 69.530 67.835 71.510 68.165 ;
        RECT 99.530 67.835 101.510 68.165 ;
        RECT 51.125 67.130 51.455 67.145 ;
        RECT 62.165 67.130 62.495 67.145 ;
        RECT 80.565 67.130 80.895 67.145 ;
        RECT 51.125 66.830 80.895 67.130 ;
        RECT 51.125 66.815 51.455 66.830 ;
        RECT 62.165 66.815 62.495 66.830 ;
        RECT 80.565 66.815 80.895 66.830 ;
        RECT 24.530 65.115 26.510 65.445 ;
        RECT 54.530 65.115 56.510 65.445 ;
        RECT 84.530 65.115 86.510 65.445 ;
        RECT 114.530 65.115 116.510 65.445 ;
        RECT 9.530 62.395 11.510 62.725 ;
        RECT 39.530 62.395 41.510 62.725 ;
        RECT 69.530 62.395 71.510 62.725 ;
        RECT 99.530 62.395 101.510 62.725 ;
        RECT 24.530 59.675 26.510 60.005 ;
        RECT 54.530 59.675 56.510 60.005 ;
        RECT 84.530 59.675 86.510 60.005 ;
        RECT 114.530 59.675 116.510 60.005 ;
        RECT 89.510 59.650 89.890 59.660 ;
        RECT 92.065 59.650 92.395 59.665 ;
        RECT 89.510 59.350 92.395 59.650 ;
        RECT 89.510 59.340 89.890 59.350 ;
        RECT 92.065 59.335 92.395 59.350 ;
        RECT 30.885 58.970 31.215 58.985 ;
        RECT 48.825 58.970 49.155 58.985 ;
        RECT 72.030 58.970 72.410 58.980 ;
        RECT 30.885 58.670 72.410 58.970 ;
        RECT 30.885 58.655 31.215 58.670 ;
        RECT 48.825 58.655 49.155 58.670 ;
        RECT 72.030 58.660 72.410 58.670 ;
        RECT 9.530 56.955 11.510 57.285 ;
        RECT 39.530 56.955 41.510 57.285 ;
        RECT 69.530 56.955 71.510 57.285 ;
        RECT 99.530 56.955 101.510 57.285 ;
        RECT 24.530 54.235 26.510 54.565 ;
        RECT 54.530 54.235 56.510 54.565 ;
        RECT 84.530 54.235 86.510 54.565 ;
        RECT 114.530 54.235 116.510 54.565 ;
        RECT 5.585 52.170 5.915 52.185 ;
        RECT 2.000 51.870 5.915 52.170 ;
        RECT 5.585 51.855 5.915 51.870 ;
        RECT 9.530 51.515 11.510 51.845 ;
        RECT 39.530 51.515 41.510 51.845 ;
        RECT 69.530 51.515 71.510 51.845 ;
        RECT 99.530 51.515 101.510 51.845 ;
        RECT 61.705 50.810 62.035 50.825 ;
        RECT 63.545 50.810 63.875 50.825 ;
        RECT 61.705 50.510 63.875 50.810 ;
        RECT 61.705 50.495 62.035 50.510 ;
        RECT 63.545 50.495 63.875 50.510 ;
        RECT 61.245 50.130 61.575 50.145 ;
        RECT 66.305 50.130 66.635 50.145 ;
        RECT 61.245 49.830 66.635 50.130 ;
        RECT 61.245 49.815 61.575 49.830 ;
        RECT 66.305 49.815 66.635 49.830 ;
        RECT 24.530 48.795 26.510 49.125 ;
        RECT 54.530 48.795 56.510 49.125 ;
        RECT 84.530 48.795 86.510 49.125 ;
        RECT 114.530 48.795 116.510 49.125 ;
        RECT 55.265 48.090 55.595 48.105 ;
        RECT 57.310 48.090 57.690 48.100 ;
        RECT 55.265 47.790 57.690 48.090 ;
        RECT 55.265 47.775 55.595 47.790 ;
        RECT 57.310 47.780 57.690 47.790 ;
        RECT 9.530 46.075 11.510 46.405 ;
        RECT 39.530 46.075 41.510 46.405 ;
        RECT 69.530 46.075 71.510 46.405 ;
        RECT 99.530 46.075 101.510 46.405 ;
        RECT 24.530 43.355 26.510 43.685 ;
        RECT 54.530 43.355 56.510 43.685 ;
        RECT 84.530 43.355 86.510 43.685 ;
        RECT 114.530 43.355 116.510 43.685 ;
        RECT 65.845 43.340 66.175 43.345 ;
        RECT 65.590 43.330 66.175 43.340 ;
        RECT 65.590 43.030 66.400 43.330 ;
        RECT 65.590 43.020 66.175 43.030 ;
        RECT 65.845 43.015 66.175 43.020 ;
        RECT 9.530 40.635 11.510 40.965 ;
        RECT 39.530 40.635 41.510 40.965 ;
        RECT 69.530 40.635 71.510 40.965 ;
        RECT 99.530 40.635 101.510 40.965 ;
        RECT 24.530 37.915 26.510 38.245 ;
        RECT 54.530 37.915 56.510 38.245 ;
        RECT 84.530 37.915 86.510 38.245 ;
        RECT 114.530 37.915 116.510 38.245 ;
        RECT 9.530 35.195 11.510 35.525 ;
        RECT 39.530 35.195 41.510 35.525 ;
        RECT 69.530 35.195 71.510 35.525 ;
        RECT 99.530 35.195 101.510 35.525 ;
        RECT 24.530 32.475 26.510 32.805 ;
        RECT 54.530 32.475 56.510 32.805 ;
        RECT 84.530 32.475 86.510 32.805 ;
        RECT 114.530 32.475 116.510 32.805 ;
        RECT 9.530 29.755 11.510 30.085 ;
        RECT 39.530 29.755 41.510 30.085 ;
        RECT 69.530 29.755 71.510 30.085 ;
        RECT 99.530 29.755 101.510 30.085 ;
        RECT 24.530 27.035 26.510 27.365 ;
        RECT 54.530 27.035 56.510 27.365 ;
        RECT 84.530 27.035 86.510 27.365 ;
        RECT 114.530 27.035 116.510 27.365 ;
        RECT 9.530 24.315 11.510 24.645 ;
        RECT 39.530 24.315 41.510 24.645 ;
        RECT 69.530 24.315 71.510 24.645 ;
        RECT 99.530 24.315 101.510 24.645 ;
        RECT 24.530 21.595 26.510 21.925 ;
        RECT 54.530 21.595 56.510 21.925 ;
        RECT 84.530 21.595 86.510 21.925 ;
        RECT 114.530 21.595 116.510 21.925 ;
        RECT 9.530 18.875 11.510 19.205 ;
        RECT 39.530 18.875 41.510 19.205 ;
        RECT 69.530 18.875 71.510 19.205 ;
        RECT 99.530 18.875 101.510 19.205 ;
        RECT 24.530 16.155 26.510 16.485 ;
        RECT 54.530 16.155 56.510 16.485 ;
        RECT 84.530 16.155 86.510 16.485 ;
        RECT 114.530 16.155 116.510 16.485 ;
        RECT 9.530 13.435 11.510 13.765 ;
        RECT 39.530 13.435 41.510 13.765 ;
        RECT 69.530 13.435 71.510 13.765 ;
        RECT 99.530 13.435 101.510 13.765 ;
        RECT 24.530 10.715 26.510 11.045 ;
        RECT 54.530 10.715 56.510 11.045 ;
        RECT 84.530 10.715 86.510 11.045 ;
        RECT 114.530 10.715 116.510 11.045 ;
      LAYER met4 ;
        RECT 83.095 106.935 83.425 107.265 ;
        RECT 57.335 89.935 57.665 90.265 ;
        RECT 57.350 48.105 57.650 89.935 ;
        RECT 63.775 87.895 64.105 88.225 ;
        RECT 63.790 75.985 64.090 87.895 ;
        RECT 65.615 79.735 65.945 80.065 ;
        RECT 63.775 75.655 64.105 75.985 ;
        RECT 57.335 47.775 57.665 48.105 ;
        RECT 65.630 43.345 65.930 79.735 ;
        RECT 83.110 75.985 83.410 106.935 ;
        RECT 72.055 75.655 72.385 75.985 ;
        RECT 83.095 75.655 83.425 75.985 ;
        RECT 72.070 58.985 72.370 75.655 ;
        RECT 89.535 74.975 89.865 75.305 ;
        RECT 89.550 59.665 89.850 74.975 ;
        RECT 89.535 59.335 89.865 59.665 ;
        RECT 72.055 58.655 72.385 58.985 ;
        RECT 65.615 43.015 65.945 43.345 ;
  END
END digital_top
END LIBRARY

