VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 853.044495 ;
    ANTENNADIFFAREA 1113.359375 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.515 210.815 14.685 211.005 ;
        RECT 18.195 210.815 18.365 211.005 ;
        RECT 23.715 210.815 23.885 211.005 ;
        RECT 25.555 210.815 25.725 211.005 ;
        RECT 31.075 210.815 31.245 211.005 ;
        RECT 36.595 210.815 36.765 211.005 ;
        RECT 38.435 210.815 38.605 211.005 ;
        RECT 43.955 210.815 44.125 211.005 ;
        RECT 49.475 210.815 49.645 211.005 ;
        RECT 51.315 210.815 51.485 211.005 ;
        RECT 56.835 210.815 57.005 211.005 ;
        RECT 62.355 210.815 62.525 211.005 ;
        RECT 64.195 210.815 64.365 211.005 ;
        RECT 69.715 210.815 69.885 211.005 ;
        RECT 75.235 210.815 75.405 211.005 ;
        RECT 77.075 210.815 77.245 211.005 ;
        RECT 82.595 210.815 82.765 211.005 ;
        RECT 88.115 210.815 88.285 211.005 ;
        RECT 89.955 210.815 90.125 211.005 ;
        RECT 95.475 210.815 95.645 211.005 ;
        RECT 100.995 210.815 101.165 211.005 ;
        RECT 102.835 210.815 103.005 211.005 ;
        RECT 108.355 210.815 108.525 211.005 ;
        RECT 113.875 210.815 114.045 211.005 ;
        RECT 114.850 210.865 114.970 210.975 ;
        RECT 120.315 210.815 120.485 211.005 ;
        RECT 125.835 210.815 126.005 211.005 ;
        RECT 127.215 210.815 127.385 211.005 ;
        RECT 14.375 210.005 15.745 210.815 ;
        RECT 15.755 210.005 18.505 210.815 ;
        RECT 18.515 210.005 24.025 210.815 ;
        RECT 24.045 209.945 24.475 210.730 ;
        RECT 24.495 210.005 25.865 210.815 ;
        RECT 25.875 210.005 31.385 210.815 ;
        RECT 31.395 210.005 36.905 210.815 ;
        RECT 36.925 209.945 37.355 210.730 ;
        RECT 37.375 210.005 38.745 210.815 ;
        RECT 38.755 210.005 44.265 210.815 ;
        RECT 44.275 210.005 49.785 210.815 ;
        RECT 49.805 209.945 50.235 210.730 ;
        RECT 50.255 210.005 51.625 210.815 ;
        RECT 51.635 210.005 57.145 210.815 ;
        RECT 57.155 210.005 62.665 210.815 ;
        RECT 62.685 209.945 63.115 210.730 ;
        RECT 63.135 210.005 64.505 210.815 ;
        RECT 64.515 210.005 70.025 210.815 ;
        RECT 70.035 210.005 75.545 210.815 ;
        RECT 75.565 209.945 75.995 210.730 ;
        RECT 76.015 210.005 77.385 210.815 ;
        RECT 77.395 210.005 82.905 210.815 ;
        RECT 82.915 210.005 88.425 210.815 ;
        RECT 88.445 209.945 88.875 210.730 ;
        RECT 88.895 210.005 90.265 210.815 ;
        RECT 90.275 210.005 95.785 210.815 ;
        RECT 95.795 210.005 101.305 210.815 ;
        RECT 101.325 209.945 101.755 210.730 ;
        RECT 101.775 210.005 103.145 210.815 ;
        RECT 103.155 210.005 108.665 210.815 ;
        RECT 108.675 210.005 114.185 210.815 ;
        RECT 114.205 209.945 114.635 210.730 ;
        RECT 115.115 210.005 120.625 210.815 ;
        RECT 120.635 210.005 126.145 210.815 ;
        RECT 126.155 210.005 127.525 210.815 ;
      LAYER nwell ;
        RECT 14.180 206.785 127.720 209.615 ;
      LAYER pwell ;
        RECT 14.375 205.585 15.745 206.395 ;
        RECT 15.755 205.585 18.505 206.395 ;
        RECT 18.515 205.585 24.025 206.395 ;
        RECT 24.045 205.670 24.475 206.455 ;
        RECT 24.955 205.585 27.705 206.395 ;
        RECT 27.715 205.585 33.225 206.395 ;
        RECT 33.235 205.585 38.745 206.395 ;
        RECT 38.755 205.585 44.265 206.395 ;
        RECT 44.275 205.585 49.785 206.395 ;
        RECT 49.805 205.670 50.235 206.455 ;
        RECT 50.255 205.585 55.765 206.395 ;
        RECT 55.775 205.585 61.285 206.395 ;
        RECT 61.295 205.585 66.805 206.395 ;
        RECT 66.815 205.585 72.325 206.395 ;
        RECT 72.345 205.585 73.695 206.495 ;
        RECT 74.200 206.265 75.545 206.495 ;
        RECT 73.715 205.585 75.545 206.265 ;
        RECT 75.565 205.670 75.995 206.455 ;
        RECT 76.935 205.585 80.045 206.495 ;
        RECT 81.075 205.585 84.745 206.395 ;
        RECT 84.755 205.585 90.265 206.395 ;
        RECT 90.275 205.585 95.785 206.395 ;
        RECT 95.795 205.585 101.305 206.395 ;
        RECT 101.325 205.670 101.755 206.455 ;
        RECT 102.235 205.585 104.065 206.395 ;
        RECT 104.075 205.585 109.585 206.395 ;
        RECT 109.595 205.585 115.105 206.395 ;
        RECT 115.115 205.585 120.625 206.395 ;
        RECT 120.635 205.585 126.145 206.395 ;
        RECT 126.155 205.585 127.525 206.395 ;
        RECT 14.515 205.375 14.685 205.585 ;
        RECT 16.355 205.420 16.515 205.530 ;
        RECT 18.195 205.395 18.365 205.585 ;
        RECT 20.035 205.375 20.205 205.565 ;
        RECT 23.715 205.395 23.885 205.585 ;
        RECT 24.690 205.425 24.810 205.535 ;
        RECT 25.555 205.375 25.725 205.565 ;
        RECT 27.395 205.395 27.565 205.585 ;
        RECT 31.075 205.375 31.245 205.565 ;
        RECT 32.915 205.395 33.085 205.585 ;
        RECT 36.595 205.375 36.765 205.565 ;
        RECT 37.570 205.425 37.690 205.535 ;
        RECT 38.435 205.395 38.605 205.585 ;
        RECT 40.275 205.375 40.445 205.565 ;
        RECT 43.955 205.395 44.125 205.585 ;
        RECT 45.795 205.375 45.965 205.565 ;
        RECT 49.475 205.395 49.645 205.585 ;
        RECT 51.315 205.375 51.485 205.565 ;
        RECT 55.455 205.395 55.625 205.585 ;
        RECT 56.835 205.375 57.005 205.565 ;
        RECT 60.975 205.395 61.145 205.585 ;
        RECT 62.355 205.375 62.525 205.565 ;
        RECT 64.195 205.375 64.365 205.565 ;
        RECT 65.575 205.375 65.745 205.565 ;
        RECT 66.495 205.395 66.665 205.585 ;
        RECT 66.955 205.375 67.125 205.565 ;
        RECT 72.015 205.395 72.185 205.585 ;
        RECT 72.475 205.395 72.645 205.585 ;
        RECT 73.855 205.395 74.025 205.585 ;
        RECT 76.615 205.430 76.775 205.540 ;
        RECT 77.075 205.375 77.245 205.565 ;
        RECT 79.835 205.395 80.005 205.585 ;
        RECT 80.755 205.430 80.915 205.540 ;
        RECT 84.435 205.395 84.605 205.585 ;
        RECT 86.275 205.375 86.445 205.565 ;
        RECT 88.115 205.375 88.285 205.565 ;
        RECT 89.090 205.425 89.210 205.535 ;
        RECT 89.955 205.395 90.125 205.585 ;
        RECT 91.795 205.375 91.965 205.565 ;
        RECT 95.475 205.395 95.645 205.585 ;
        RECT 97.315 205.375 97.485 205.565 ;
        RECT 100.995 205.395 101.165 205.585 ;
        RECT 101.970 205.425 102.090 205.535 ;
        RECT 102.835 205.375 103.005 205.565 ;
        RECT 103.755 205.395 103.925 205.585 ;
        RECT 108.355 205.375 108.525 205.565 ;
        RECT 109.275 205.395 109.445 205.585 ;
        RECT 113.875 205.375 114.045 205.565 ;
        RECT 114.795 205.535 114.965 205.585 ;
        RECT 114.795 205.425 114.970 205.535 ;
        RECT 114.795 205.395 114.965 205.425 ;
        RECT 120.315 205.375 120.485 205.585 ;
        RECT 125.835 205.375 126.005 205.585 ;
        RECT 127.215 205.375 127.385 205.585 ;
        RECT 14.375 204.565 15.745 205.375 ;
        RECT 16.675 204.565 20.345 205.375 ;
        RECT 20.355 204.565 25.865 205.375 ;
        RECT 25.875 204.565 31.385 205.375 ;
        RECT 31.395 204.565 36.905 205.375 ;
        RECT 36.925 204.505 37.355 205.290 ;
        RECT 37.835 204.565 40.585 205.375 ;
        RECT 40.595 204.565 46.105 205.375 ;
        RECT 46.115 204.565 51.625 205.375 ;
        RECT 51.635 204.565 57.145 205.375 ;
        RECT 57.155 204.565 62.665 205.375 ;
        RECT 62.685 204.505 63.115 205.290 ;
        RECT 63.135 204.565 64.505 205.375 ;
        RECT 64.525 204.465 65.875 205.375 ;
        RECT 66.825 204.465 68.175 205.375 ;
        RECT 68.195 204.695 77.385 205.375 ;
        RECT 77.395 204.695 86.585 205.375 ;
        RECT 68.195 204.465 69.115 204.695 ;
        RECT 71.945 204.475 72.875 204.695 ;
        RECT 77.395 204.465 78.315 204.695 ;
        RECT 81.145 204.475 82.075 204.695 ;
        RECT 86.595 204.565 88.425 205.375 ;
        RECT 88.445 204.505 88.875 205.290 ;
        RECT 89.355 204.565 92.105 205.375 ;
        RECT 92.115 204.565 97.625 205.375 ;
        RECT 97.635 204.565 103.145 205.375 ;
        RECT 103.155 204.565 108.665 205.375 ;
        RECT 108.675 204.565 114.185 205.375 ;
        RECT 114.205 204.505 114.635 205.290 ;
        RECT 115.115 204.565 120.625 205.375 ;
        RECT 120.635 204.565 126.145 205.375 ;
        RECT 126.155 204.565 127.525 205.375 ;
      LAYER nwell ;
        RECT 14.180 201.345 127.720 204.175 ;
      LAYER pwell ;
        RECT 14.375 200.145 15.745 200.955 ;
        RECT 15.755 200.145 18.505 200.955 ;
        RECT 18.515 200.145 24.025 200.955 ;
        RECT 24.045 200.230 24.475 201.015 ;
        RECT 24.955 200.145 27.705 200.955 ;
        RECT 27.715 200.145 33.225 200.955 ;
        RECT 33.235 200.145 38.745 200.955 ;
        RECT 38.755 200.145 44.265 200.955 ;
        RECT 44.275 200.145 49.785 200.955 ;
        RECT 49.805 200.230 50.235 201.015 ;
        RECT 50.255 200.145 53.925 200.955 ;
        RECT 53.935 200.145 59.445 200.955 ;
        RECT 63.965 200.825 64.895 201.045 ;
        RECT 67.615 200.825 69.825 201.055 ;
        RECT 59.455 200.145 69.825 200.825 ;
        RECT 70.035 200.825 70.965 201.055 ;
        RECT 70.035 200.145 73.705 200.825 ;
        RECT 73.715 200.145 75.545 200.825 ;
        RECT 75.565 200.230 75.995 201.015 ;
        RECT 76.475 200.825 77.395 201.055 ;
        RECT 79.235 200.825 80.155 201.055 ;
        RECT 82.985 200.825 83.915 201.045 ;
        RECT 76.475 200.145 78.765 200.825 ;
        RECT 79.235 200.145 88.425 200.825 ;
        RECT 88.435 200.145 90.265 200.955 ;
        RECT 90.275 200.145 95.785 200.955 ;
        RECT 95.795 200.145 101.305 200.955 ;
        RECT 101.325 200.230 101.755 201.015 ;
        RECT 102.235 200.145 104.065 200.955 ;
        RECT 104.075 200.145 109.585 200.955 ;
        RECT 109.595 200.145 115.105 200.955 ;
        RECT 115.115 200.145 120.625 200.955 ;
        RECT 120.635 200.145 126.145 200.955 ;
        RECT 126.155 200.145 127.525 200.955 ;
        RECT 14.515 199.935 14.685 200.145 ;
        RECT 16.355 199.980 16.515 200.090 ;
        RECT 18.195 199.955 18.365 200.145 ;
        RECT 20.035 199.935 20.205 200.125 ;
        RECT 23.715 199.955 23.885 200.145 ;
        RECT 24.690 199.985 24.810 200.095 ;
        RECT 25.555 199.935 25.725 200.125 ;
        RECT 27.395 199.955 27.565 200.145 ;
        RECT 31.075 199.935 31.245 200.125 ;
        RECT 32.915 199.955 33.085 200.145 ;
        RECT 36.595 199.935 36.765 200.125 ;
        RECT 37.570 199.985 37.690 200.095 ;
        RECT 38.435 199.955 38.605 200.145 ;
        RECT 40.275 199.935 40.445 200.125 ;
        RECT 43.955 199.955 44.125 200.145 ;
        RECT 45.795 199.935 45.965 200.125 ;
        RECT 49.475 199.955 49.645 200.145 ;
        RECT 51.315 199.935 51.485 200.125 ;
        RECT 53.615 199.955 53.785 200.145 ;
        RECT 56.835 199.935 57.005 200.125 ;
        RECT 59.135 199.955 59.305 200.145 ;
        RECT 59.595 199.955 59.765 200.145 ;
        RECT 62.355 199.935 62.525 200.125 ;
        RECT 63.330 199.985 63.450 200.095 ;
        RECT 66.955 199.935 67.125 200.125 ;
        RECT 68.335 199.935 68.505 200.125 ;
        RECT 70.175 199.935 70.345 200.125 ;
        RECT 73.395 199.955 73.565 200.145 ;
        RECT 74.775 199.935 74.945 200.125 ;
        RECT 75.235 199.955 75.405 200.145 ;
        RECT 76.210 199.985 76.330 200.095 ;
        RECT 78.455 199.935 78.625 200.145 ;
        RECT 78.970 199.985 79.090 200.095 ;
        RECT 80.755 199.955 80.925 200.125 ;
        RECT 80.755 199.935 80.920 199.955 ;
        RECT 82.140 199.935 82.310 200.125 ;
        RECT 82.595 199.935 82.765 200.125 ;
        RECT 83.975 199.935 84.145 200.125 ;
        RECT 86.275 199.935 86.445 200.125 ;
        RECT 88.115 199.935 88.285 200.145 ;
        RECT 89.090 199.985 89.210 200.095 ;
        RECT 89.955 199.955 90.125 200.145 ;
        RECT 90.875 199.935 91.045 200.125 ;
        RECT 95.475 199.955 95.645 200.145 ;
        RECT 96.395 199.935 96.565 200.125 ;
        RECT 100.995 199.955 101.165 200.145 ;
        RECT 101.970 199.985 102.090 200.095 ;
        RECT 103.755 199.955 103.925 200.145 ;
        RECT 105.595 199.935 105.765 200.125 ;
        RECT 108.355 199.935 108.525 200.125 ;
        RECT 109.275 199.955 109.445 200.145 ;
        RECT 113.875 199.935 114.045 200.125 ;
        RECT 114.795 200.095 114.965 200.145 ;
        RECT 114.795 199.985 114.970 200.095 ;
        RECT 114.795 199.955 114.965 199.985 ;
        RECT 120.315 199.935 120.485 200.145 ;
        RECT 125.835 199.935 126.005 200.145 ;
        RECT 127.215 199.935 127.385 200.145 ;
        RECT 14.375 199.125 15.745 199.935 ;
        RECT 16.675 199.125 20.345 199.935 ;
        RECT 20.355 199.125 25.865 199.935 ;
        RECT 25.875 199.125 31.385 199.935 ;
        RECT 31.395 199.125 36.905 199.935 ;
        RECT 36.925 199.065 37.355 199.850 ;
        RECT 37.835 199.125 40.585 199.935 ;
        RECT 40.595 199.125 46.105 199.935 ;
        RECT 46.115 199.125 51.625 199.935 ;
        RECT 51.635 199.125 57.145 199.935 ;
        RECT 57.155 199.125 62.665 199.935 ;
        RECT 62.685 199.065 63.115 199.850 ;
        RECT 63.595 199.125 67.265 199.935 ;
        RECT 67.275 199.155 68.645 199.935 ;
        RECT 68.655 199.255 70.485 199.935 ;
        RECT 70.505 199.895 71.425 199.935 ;
        RECT 70.495 199.705 71.425 199.895 ;
        RECT 73.515 199.705 75.085 199.935 ;
        RECT 70.495 199.345 75.085 199.705 ;
        RECT 70.505 199.255 75.085 199.345 ;
        RECT 75.190 199.255 78.655 199.935 ;
        RECT 79.085 199.255 80.920 199.935 ;
        RECT 70.505 199.025 73.505 199.255 ;
        RECT 75.190 199.025 76.110 199.255 ;
        RECT 79.085 199.025 80.015 199.255 ;
        RECT 81.075 199.025 82.425 199.935 ;
        RECT 82.455 199.155 83.825 199.935 ;
        RECT 83.845 199.025 85.195 199.935 ;
        RECT 85.225 199.025 86.575 199.935 ;
        RECT 86.595 199.125 88.425 199.935 ;
        RECT 88.445 199.065 88.875 199.850 ;
        RECT 89.355 199.125 91.185 199.935 ;
        RECT 91.195 199.125 96.705 199.935 ;
        RECT 96.715 199.255 105.905 199.935 ;
        RECT 96.715 199.025 97.635 199.255 ;
        RECT 100.465 199.035 101.395 199.255 ;
        RECT 105.915 199.125 108.665 199.935 ;
        RECT 108.675 199.125 114.185 199.935 ;
        RECT 114.205 199.065 114.635 199.850 ;
        RECT 115.115 199.125 120.625 199.935 ;
        RECT 120.635 199.125 126.145 199.935 ;
        RECT 126.155 199.125 127.525 199.935 ;
      LAYER nwell ;
        RECT 14.180 195.905 127.720 198.735 ;
      LAYER pwell ;
        RECT 14.375 194.705 15.745 195.515 ;
        RECT 15.755 194.705 18.505 195.515 ;
        RECT 18.515 194.705 24.025 195.515 ;
        RECT 24.045 194.790 24.475 195.575 ;
        RECT 24.955 194.705 27.705 195.515 ;
        RECT 27.715 194.705 33.225 195.515 ;
        RECT 33.235 194.705 38.745 195.515 ;
        RECT 38.755 194.705 44.265 195.515 ;
        RECT 44.275 194.705 49.785 195.515 ;
        RECT 49.805 194.790 50.235 195.575 ;
        RECT 50.715 194.705 52.545 195.515 ;
        RECT 52.565 194.705 53.915 195.615 ;
        RECT 56.590 195.385 57.510 195.615 ;
        RECT 54.045 194.705 57.510 195.385 ;
        RECT 57.615 194.705 63.125 195.515 ;
        RECT 63.135 194.705 68.645 195.515 ;
        RECT 68.655 195.385 69.575 195.615 ;
        RECT 68.655 194.705 70.945 195.385 ;
        RECT 70.955 194.705 73.875 195.615 ;
        RECT 74.175 194.705 75.545 195.515 ;
        RECT 75.565 194.790 75.995 195.575 ;
        RECT 76.015 194.705 79.685 195.515 ;
        RECT 79.695 194.705 85.205 195.515 ;
        RECT 85.585 195.505 86.505 195.615 ;
        RECT 85.585 195.385 87.920 195.505 ;
        RECT 92.585 195.385 93.505 195.605 ;
        RECT 85.585 194.705 94.865 195.385 ;
        RECT 94.875 194.705 97.625 195.515 ;
        RECT 100.290 195.385 101.210 195.615 ;
        RECT 97.745 194.705 101.210 195.385 ;
        RECT 101.325 194.790 101.755 195.575 ;
        RECT 101.775 194.705 104.525 195.515 ;
        RECT 104.535 194.705 110.045 195.515 ;
        RECT 110.055 195.385 110.975 195.615 ;
        RECT 113.805 195.385 114.735 195.605 ;
        RECT 110.055 194.705 119.245 195.385 ;
        RECT 119.255 194.705 120.625 195.515 ;
        RECT 120.635 194.705 126.145 195.515 ;
        RECT 126.155 194.705 127.525 195.515 ;
        RECT 14.515 194.495 14.685 194.705 ;
        RECT 16.355 194.540 16.515 194.650 ;
        RECT 18.195 194.515 18.365 194.705 ;
        RECT 20.035 194.495 20.205 194.685 ;
        RECT 23.715 194.515 23.885 194.705 ;
        RECT 24.690 194.545 24.810 194.655 ;
        RECT 25.555 194.495 25.725 194.685 ;
        RECT 27.395 194.515 27.565 194.705 ;
        RECT 31.075 194.495 31.245 194.685 ;
        RECT 32.915 194.515 33.085 194.705 ;
        RECT 36.595 194.495 36.765 194.685 ;
        RECT 37.975 194.540 38.135 194.650 ;
        RECT 38.435 194.515 38.605 194.705 ;
        RECT 41.655 194.495 41.825 194.685 ;
        RECT 43.955 194.515 44.125 194.705 ;
        RECT 47.175 194.495 47.345 194.685 ;
        RECT 48.555 194.495 48.725 194.685 ;
        RECT 49.015 194.495 49.185 194.685 ;
        RECT 49.475 194.515 49.645 194.705 ;
        RECT 50.450 194.545 50.570 194.655 ;
        RECT 52.235 194.515 52.405 194.705 ;
        RECT 53.615 194.515 53.785 194.705 ;
        RECT 54.075 194.515 54.245 194.705 ;
        RECT 58.675 194.540 58.835 194.650 ;
        RECT 62.355 194.495 62.525 194.685 ;
        RECT 62.815 194.515 62.985 194.705 ;
        RECT 64.655 194.495 64.825 194.685 ;
        RECT 66.035 194.495 66.205 194.685 ;
        RECT 66.550 194.545 66.670 194.655 ;
        RECT 68.335 194.495 68.505 194.705 ;
        RECT 14.375 193.685 15.745 194.495 ;
        RECT 16.675 193.685 20.345 194.495 ;
        RECT 20.355 193.685 25.865 194.495 ;
        RECT 25.875 193.685 31.385 194.495 ;
        RECT 31.395 193.685 36.905 194.495 ;
        RECT 36.925 193.625 37.355 194.410 ;
        RECT 38.295 193.685 41.965 194.495 ;
        RECT 41.975 193.685 47.485 194.495 ;
        RECT 47.505 193.585 48.855 194.495 ;
        RECT 48.875 193.815 58.065 194.495 ;
        RECT 53.385 193.595 54.315 193.815 ;
        RECT 57.145 193.585 58.065 193.815 ;
        RECT 58.995 193.685 62.665 194.495 ;
        RECT 62.685 193.625 63.115 194.410 ;
        RECT 63.135 193.685 64.965 194.495 ;
        RECT 64.985 193.585 66.335 194.495 ;
        RECT 66.815 193.685 68.645 194.495 ;
        RECT 68.795 194.465 68.965 194.685 ;
        RECT 70.635 194.515 70.805 194.705 ;
        RECT 71.100 194.515 71.270 194.705 ;
        RECT 70.920 194.465 71.865 194.495 ;
        RECT 68.795 194.265 71.865 194.465 ;
        RECT 68.655 193.785 71.865 194.265 ;
        RECT 68.655 193.585 69.585 193.785 ;
        RECT 70.920 193.585 71.865 193.785 ;
        RECT 71.875 194.465 72.820 194.495 ;
        RECT 74.775 194.465 74.945 194.685 ;
        RECT 75.235 194.515 75.405 194.705 ;
        RECT 78.455 194.495 78.625 194.685 ;
        RECT 79.375 194.515 79.545 194.705 ;
        RECT 83.975 194.495 84.145 194.685 ;
        RECT 84.895 194.515 85.065 194.705 ;
        RECT 87.840 194.495 88.010 194.685 ;
        RECT 89.955 194.495 90.125 194.685 ;
        RECT 92.715 194.495 92.885 194.685 ;
        RECT 93.175 194.495 93.345 194.685 ;
        RECT 94.555 194.495 94.725 194.705 ;
        RECT 97.315 194.515 97.485 194.705 ;
        RECT 97.775 194.515 97.945 194.705 ;
        RECT 104.215 194.515 104.385 194.705 ;
        RECT 104.675 194.495 104.845 194.685 ;
        RECT 108.355 194.495 108.525 194.685 ;
        RECT 108.815 194.495 108.985 194.685 ;
        RECT 109.735 194.515 109.905 194.705 ;
        RECT 113.600 194.495 113.770 194.685 ;
        RECT 115.715 194.495 115.885 194.685 ;
        RECT 116.635 194.540 116.795 194.650 ;
        RECT 118.935 194.515 119.105 194.705 ;
        RECT 120.315 194.495 120.485 194.705 ;
        RECT 125.835 194.495 126.005 194.705 ;
        RECT 127.215 194.495 127.385 194.705 ;
        RECT 71.875 194.265 74.945 194.465 ;
        RECT 71.875 193.785 75.085 194.265 ;
        RECT 71.875 193.585 72.820 193.785 ;
        RECT 74.155 193.585 75.085 193.785 ;
        RECT 75.095 193.685 78.765 194.495 ;
        RECT 78.775 193.685 84.285 194.495 ;
        RECT 84.525 193.815 88.425 194.495 ;
        RECT 87.495 193.585 88.425 193.815 ;
        RECT 88.445 193.625 88.875 194.410 ;
        RECT 88.905 193.585 90.255 194.495 ;
        RECT 90.275 193.685 93.025 194.495 ;
        RECT 93.045 193.585 94.395 194.495 ;
        RECT 94.415 193.815 103.520 194.495 ;
        RECT 103.615 193.685 104.985 194.495 ;
        RECT 104.995 193.685 108.665 194.495 ;
        RECT 108.685 193.585 110.035 194.495 ;
        RECT 110.285 193.815 114.185 194.495 ;
        RECT 113.255 193.585 114.185 193.815 ;
        RECT 114.205 193.625 114.635 194.410 ;
        RECT 114.665 193.585 116.015 194.495 ;
        RECT 116.955 193.685 120.625 194.495 ;
        RECT 120.635 193.685 126.145 194.495 ;
        RECT 126.155 193.685 127.525 194.495 ;
      LAYER nwell ;
        RECT 14.180 190.465 127.720 193.295 ;
      LAYER pwell ;
        RECT 14.375 189.265 15.745 190.075 ;
        RECT 15.755 189.265 18.505 190.075 ;
        RECT 18.515 189.265 24.025 190.075 ;
        RECT 24.045 189.350 24.475 190.135 ;
        RECT 24.955 189.265 30.465 190.075 ;
        RECT 30.475 189.265 35.985 190.075 ;
        RECT 36.365 190.065 37.285 190.175 ;
        RECT 36.365 189.945 38.700 190.065 ;
        RECT 43.365 189.945 44.285 190.165 ;
        RECT 48.855 189.945 49.785 190.175 ;
        RECT 36.365 189.265 45.645 189.945 ;
        RECT 45.885 189.265 49.785 189.945 ;
        RECT 49.805 189.350 50.235 190.135 ;
        RECT 50.715 189.265 52.085 190.045 ;
        RECT 52.095 189.945 53.015 190.175 ;
        RECT 55.845 189.945 56.775 190.165 ;
        RECT 61.335 189.945 62.675 190.175 ;
        RECT 65.505 189.945 66.435 190.165 ;
        RECT 52.095 189.265 61.285 189.945 ;
        RECT 61.335 189.265 70.945 189.945 ;
        RECT 70.955 189.265 74.065 190.175 ;
        RECT 74.175 189.265 75.545 190.075 ;
        RECT 75.565 189.350 75.995 190.135 ;
        RECT 76.015 189.265 78.305 190.175 ;
        RECT 79.235 189.265 82.905 190.075 ;
        RECT 83.285 190.065 84.205 190.175 ;
        RECT 83.285 189.945 85.620 190.065 ;
        RECT 90.285 189.945 91.205 190.165 ;
        RECT 83.285 189.265 92.565 189.945 ;
        RECT 92.575 189.265 93.945 190.045 ;
        RECT 100.375 189.945 101.305 190.175 ;
        RECT 94.335 189.265 96.760 189.945 ;
        RECT 97.405 189.265 101.305 189.945 ;
        RECT 101.325 189.350 101.755 190.135 ;
        RECT 101.775 189.265 103.145 190.045 ;
        RECT 103.155 189.265 104.525 190.075 ;
        RECT 107.735 189.945 108.665 190.175 ;
        RECT 104.765 189.265 108.665 189.945 ;
        RECT 108.675 189.945 109.595 190.175 ;
        RECT 112.425 189.945 113.355 190.165 ;
        RECT 108.675 189.265 117.865 189.945 ;
        RECT 117.875 189.265 119.245 190.045 ;
        RECT 119.255 189.265 120.625 190.075 ;
        RECT 120.635 189.265 126.145 190.075 ;
        RECT 126.155 189.265 127.525 190.075 ;
        RECT 14.515 189.055 14.685 189.265 ;
        RECT 15.950 189.105 16.070 189.215 ;
        RECT 17.735 189.055 17.905 189.245 ;
        RECT 18.195 189.075 18.365 189.265 ;
        RECT 23.255 189.055 23.425 189.245 ;
        RECT 23.715 189.075 23.885 189.265 ;
        RECT 24.690 189.105 24.810 189.215 ;
        RECT 28.775 189.055 28.945 189.245 ;
        RECT 30.155 189.055 30.325 189.265 ;
        RECT 31.535 189.055 31.705 189.245 ;
        RECT 35.215 189.055 35.385 189.245 ;
        RECT 35.675 189.055 35.845 189.265 ;
        RECT 45.335 189.075 45.505 189.265 ;
        RECT 46.255 189.055 46.425 189.245 ;
        RECT 49.200 189.075 49.370 189.265 ;
        RECT 50.450 189.105 50.570 189.215 ;
        RECT 51.775 189.075 51.945 189.265 ;
        RECT 55.455 189.055 55.625 189.245 ;
        RECT 59.320 189.055 59.490 189.245 ;
        RECT 60.975 189.055 61.145 189.265 ;
        RECT 62.355 189.055 62.525 189.245 ;
        RECT 63.330 189.105 63.450 189.215 ;
        RECT 63.735 189.055 63.905 189.245 ;
        RECT 69.715 189.055 69.885 189.245 ;
        RECT 70.635 189.075 70.805 189.265 ;
        RECT 73.855 189.075 74.025 189.265 ;
        RECT 75.235 189.055 75.405 189.265 ;
        RECT 76.160 189.075 76.330 189.265 ;
        RECT 78.915 189.110 79.075 189.220 ;
        RECT 80.755 189.055 80.925 189.245 ;
        RECT 82.595 189.075 82.765 189.265 ;
        RECT 86.275 189.055 86.445 189.245 ;
        RECT 87.655 189.055 87.825 189.245 ;
        RECT 88.170 189.105 88.290 189.215 ;
        RECT 89.035 189.055 89.205 189.245 ;
        RECT 91.795 189.055 91.965 189.245 ;
        RECT 92.255 189.075 92.425 189.265 ;
        RECT 92.715 189.075 92.885 189.265 ;
        RECT 96.855 189.075 97.025 189.245 ;
        RECT 97.315 189.055 97.485 189.245 ;
        RECT 100.720 189.075 100.890 189.265 ;
        RECT 101.915 189.075 102.085 189.265 ;
        RECT 104.215 189.075 104.385 189.265 ;
        RECT 106.515 189.055 106.685 189.245 ;
        RECT 108.080 189.075 108.250 189.265 ;
        RECT 110.195 189.055 110.365 189.245 ;
        RECT 110.710 189.105 110.830 189.215 ;
        RECT 112.495 189.055 112.665 189.245 ;
        RECT 112.955 189.055 113.125 189.245 ;
        RECT 114.850 189.105 114.970 189.215 ;
        RECT 117.555 189.075 117.725 189.265 ;
        RECT 118.935 189.075 119.105 189.265 ;
        RECT 120.315 189.055 120.485 189.265 ;
        RECT 125.835 189.055 126.005 189.265 ;
        RECT 127.215 189.055 127.385 189.265 ;
        RECT 14.375 188.245 15.745 189.055 ;
        RECT 16.215 188.245 18.045 189.055 ;
        RECT 18.055 188.245 23.565 189.055 ;
        RECT 23.575 188.245 29.085 189.055 ;
        RECT 29.105 188.145 30.455 189.055 ;
        RECT 30.475 188.245 31.845 189.055 ;
        RECT 31.855 188.245 35.525 189.055 ;
        RECT 35.545 188.145 36.895 189.055 ;
        RECT 36.925 188.185 37.355 188.970 ;
        RECT 37.375 188.375 46.565 189.055 ;
        RECT 46.660 188.375 55.765 189.055 ;
        RECT 56.005 188.375 59.905 189.055 ;
        RECT 37.375 188.145 38.295 188.375 ;
        RECT 41.125 188.155 42.055 188.375 ;
        RECT 58.975 188.145 59.905 188.375 ;
        RECT 59.915 188.275 61.285 189.055 ;
        RECT 61.295 188.245 62.665 189.055 ;
        RECT 62.685 188.185 63.115 188.970 ;
        RECT 63.705 188.375 67.170 189.055 ;
        RECT 66.250 188.145 67.170 188.375 ;
        RECT 67.275 188.245 70.025 189.055 ;
        RECT 70.035 188.245 75.545 189.055 ;
        RECT 75.555 188.245 81.065 189.055 ;
        RECT 81.075 188.245 86.585 189.055 ;
        RECT 86.605 188.145 87.955 189.055 ;
        RECT 88.445 188.185 88.875 188.970 ;
        RECT 88.895 188.275 90.265 189.055 ;
        RECT 90.275 188.245 92.105 189.055 ;
        RECT 92.115 188.245 97.625 189.055 ;
        RECT 97.635 188.375 106.825 189.055 ;
        RECT 106.930 188.375 110.395 189.055 ;
        RECT 97.635 188.145 98.555 188.375 ;
        RECT 101.385 188.155 102.315 188.375 ;
        RECT 106.930 188.145 107.850 188.375 ;
        RECT 110.975 188.245 112.805 189.055 ;
        RECT 112.815 188.275 114.185 189.055 ;
        RECT 114.205 188.185 114.635 188.970 ;
        RECT 115.115 188.245 120.625 189.055 ;
        RECT 120.635 188.245 126.145 189.055 ;
        RECT 126.155 188.245 127.525 189.055 ;
      LAYER nwell ;
        RECT 14.180 185.025 127.720 187.855 ;
      LAYER pwell ;
        RECT 14.375 183.825 15.745 184.635 ;
        RECT 15.755 183.825 18.505 184.635 ;
        RECT 18.515 183.825 24.025 184.635 ;
        RECT 24.045 183.910 24.475 184.695 ;
        RECT 24.495 183.825 25.865 184.635 ;
        RECT 25.875 184.505 26.795 184.735 ;
        RECT 29.625 184.505 30.555 184.725 ;
        RECT 25.875 183.825 35.065 184.505 ;
        RECT 35.535 183.825 38.285 184.635 ;
        RECT 38.305 183.825 39.655 184.735 ;
        RECT 42.875 184.505 43.805 184.735 ;
        RECT 39.905 183.825 43.805 184.505 ;
        RECT 43.815 184.505 44.745 184.735 ;
        RECT 43.815 183.825 47.715 184.505 ;
        RECT 48.425 183.825 49.775 184.735 ;
        RECT 49.805 183.910 50.235 184.695 ;
        RECT 50.255 184.505 51.175 184.735 ;
        RECT 54.005 184.505 54.935 184.725 ;
        RECT 50.255 183.825 59.445 184.505 ;
        RECT 59.915 183.825 65.425 184.635 ;
        RECT 65.435 183.825 70.945 184.635 ;
        RECT 70.965 184.505 73.965 184.735 ;
        RECT 70.965 184.415 75.545 184.505 ;
        RECT 70.955 184.055 75.545 184.415 ;
        RECT 70.955 183.865 71.885 184.055 ;
        RECT 70.965 183.825 71.885 183.865 ;
        RECT 73.975 183.825 75.545 184.055 ;
        RECT 75.565 183.910 75.995 184.695 ;
        RECT 76.015 183.825 78.765 184.635 ;
        RECT 78.775 183.825 84.285 184.635 ;
        RECT 87.495 184.505 88.425 184.735 ;
        RECT 84.525 183.825 88.425 184.505 ;
        RECT 88.435 183.825 93.945 184.635 ;
        RECT 96.610 184.505 97.530 184.735 ;
        RECT 94.065 183.825 97.530 184.505 ;
        RECT 98.555 183.825 99.925 184.605 ;
        RECT 99.945 183.825 101.295 184.735 ;
        RECT 101.325 183.910 101.755 184.695 ;
        RECT 102.330 184.505 103.250 184.735 ;
        RECT 109.030 184.505 109.950 184.735 ;
        RECT 112.710 184.505 113.630 184.735 ;
        RECT 102.330 183.825 105.795 184.505 ;
        RECT 106.485 183.825 109.950 184.505 ;
        RECT 110.165 183.825 113.630 184.505 ;
        RECT 113.735 183.825 115.105 184.635 ;
        RECT 115.115 183.825 120.625 184.635 ;
        RECT 120.635 183.825 126.145 184.635 ;
        RECT 126.155 183.825 127.525 184.635 ;
        RECT 14.515 183.615 14.685 183.825 ;
        RECT 15.950 183.665 16.070 183.775 ;
        RECT 18.195 183.635 18.365 183.825 ;
        RECT 21.415 183.615 21.585 183.805 ;
        RECT 21.875 183.615 22.045 183.805 ;
        RECT 23.715 183.635 23.885 183.825 ;
        RECT 25.555 183.635 25.725 183.825 ;
        RECT 26.475 183.615 26.645 183.805 ;
        RECT 26.935 183.615 27.105 183.805 ;
        RECT 30.890 183.615 31.060 183.805 ;
        RECT 34.755 183.775 34.925 183.825 ;
        RECT 34.755 183.665 34.930 183.775 ;
        RECT 35.270 183.665 35.390 183.775 ;
        RECT 34.755 183.635 34.925 183.665 ;
        RECT 36.595 183.615 36.765 183.805 ;
        RECT 37.515 183.615 37.685 183.805 ;
        RECT 37.975 183.635 38.145 183.825 ;
        RECT 38.435 183.635 38.605 183.825 ;
        RECT 41.195 183.615 41.365 183.805 ;
        RECT 43.220 183.635 43.390 183.825 ;
        RECT 44.230 183.635 44.400 183.825 ;
        RECT 44.875 183.615 45.045 183.805 ;
        RECT 48.150 183.665 48.270 183.775 ;
        RECT 48.555 183.635 48.725 183.825 ;
        RECT 49.475 183.615 49.645 183.805 ;
        RECT 50.855 183.615 51.025 183.805 ;
        RECT 51.315 183.615 51.485 183.805 ;
        RECT 55.455 183.615 55.625 183.805 ;
        RECT 55.970 183.665 56.090 183.775 ;
        RECT 58.675 183.615 58.845 183.805 ;
        RECT 59.135 183.635 59.305 183.825 ;
        RECT 59.650 183.665 59.770 183.775 ;
        RECT 60.055 183.615 60.225 183.805 ;
        RECT 60.570 183.665 60.690 183.775 ;
        RECT 62.355 183.615 62.525 183.805 ;
        RECT 63.330 183.665 63.450 183.775 ;
        RECT 65.115 183.635 65.285 183.825 ;
        RECT 66.035 183.615 66.205 183.805 ;
        RECT 66.495 183.635 66.665 183.805 ;
        RECT 66.595 183.615 66.665 183.635 ;
        RECT 69.715 183.615 69.885 183.805 ;
        RECT 70.635 183.635 70.805 183.825 ;
        RECT 75.235 183.635 75.405 183.825 ;
        RECT 77.995 183.635 78.165 183.805 ;
        RECT 78.455 183.635 78.625 183.825 ;
        RECT 78.915 183.660 79.075 183.770 ;
        RECT 83.975 183.635 84.145 183.825 ;
        RECT 87.840 183.635 88.010 183.825 ;
        RECT 77.995 183.615 78.065 183.635 ;
        RECT 88.115 183.615 88.285 183.805 ;
        RECT 89.955 183.615 90.125 183.805 ;
        RECT 91.335 183.615 91.505 183.805 ;
        RECT 93.635 183.635 93.805 183.825 ;
        RECT 94.095 183.635 94.265 183.825 ;
        RECT 95.015 183.615 95.185 183.805 ;
        RECT 98.235 183.670 98.395 183.780 ;
        RECT 98.695 183.635 98.865 183.825 ;
        RECT 98.880 183.615 99.050 183.805 ;
        RECT 100.075 183.635 100.245 183.825 ;
        RECT 101.915 183.775 102.085 183.805 ;
        RECT 101.915 183.665 102.090 183.775 ;
        RECT 101.915 183.615 102.085 183.665 ;
        RECT 105.595 183.635 105.765 183.825 ;
        RECT 106.515 183.805 106.685 183.825 ;
        RECT 105.780 183.615 105.950 183.805 ;
        RECT 106.110 183.665 106.230 183.775 ;
        RECT 106.515 183.635 106.690 183.805 ;
        RECT 110.195 183.635 110.365 183.825 ;
        RECT 106.520 183.615 106.690 183.635 ;
        RECT 113.600 183.615 113.770 183.805 ;
        RECT 114.795 183.635 114.965 183.825 ;
        RECT 115.255 183.660 115.415 183.770 ;
        RECT 120.315 183.635 120.485 183.825 ;
        RECT 124.455 183.615 124.625 183.805 ;
        RECT 125.835 183.615 126.005 183.825 ;
        RECT 127.215 183.615 127.385 183.825 ;
        RECT 14.375 182.805 15.745 183.615 ;
        RECT 16.215 182.805 21.725 183.615 ;
        RECT 21.735 182.835 23.105 183.615 ;
        RECT 23.210 182.935 26.675 183.615 ;
        RECT 26.905 182.935 30.370 183.615 ;
        RECT 23.210 182.705 24.130 182.935 ;
        RECT 29.450 182.705 30.370 182.935 ;
        RECT 30.475 182.935 34.375 183.615 ;
        RECT 30.475 182.705 31.405 182.935 ;
        RECT 35.075 182.805 36.905 183.615 ;
        RECT 36.925 182.745 37.355 183.530 ;
        RECT 37.485 182.935 40.950 183.615 ;
        RECT 41.165 182.935 44.630 183.615 ;
        RECT 44.845 182.935 48.310 183.615 ;
        RECT 40.030 182.705 40.950 182.935 ;
        RECT 43.710 182.705 44.630 182.935 ;
        RECT 47.390 182.705 48.310 182.935 ;
        RECT 48.415 182.835 49.785 183.615 ;
        RECT 49.795 182.835 51.165 183.615 ;
        RECT 51.175 182.835 52.545 183.615 ;
        RECT 52.555 182.705 55.715 183.615 ;
        RECT 56.235 182.805 58.985 183.615 ;
        RECT 59.005 182.705 60.355 183.615 ;
        RECT 60.835 182.805 62.665 183.615 ;
        RECT 62.685 182.745 63.115 183.530 ;
        RECT 63.595 182.805 66.345 183.615 ;
        RECT 66.595 183.385 68.865 183.615 ;
        RECT 69.575 183.385 74.000 183.615 ;
        RECT 75.795 183.385 78.065 183.615 ;
        RECT 66.595 182.705 69.350 183.385 ;
        RECT 69.575 182.705 74.940 183.385 ;
        RECT 75.310 182.705 78.065 183.385 ;
        RECT 79.235 182.935 88.425 183.615 ;
        RECT 79.235 182.705 80.155 182.935 ;
        RECT 82.985 182.715 83.915 182.935 ;
        RECT 88.445 182.745 88.875 183.530 ;
        RECT 88.905 182.705 90.255 183.615 ;
        RECT 90.275 182.805 91.645 183.615 ;
        RECT 91.655 182.805 95.325 183.615 ;
        RECT 95.565 182.935 99.465 183.615 ;
        RECT 98.535 182.705 99.465 182.935 ;
        RECT 99.475 182.805 102.225 183.615 ;
        RECT 102.465 182.935 106.365 183.615 ;
        RECT 105.435 182.705 106.365 182.935 ;
        RECT 106.375 182.705 109.850 183.615 ;
        RECT 110.285 182.935 114.185 183.615 ;
        RECT 113.255 182.705 114.185 182.935 ;
        RECT 114.205 182.745 114.635 183.530 ;
        RECT 115.575 182.935 124.765 183.615 ;
        RECT 115.575 182.705 116.495 182.935 ;
        RECT 119.325 182.715 120.255 182.935 ;
        RECT 124.775 182.805 126.145 183.615 ;
        RECT 126.155 182.805 127.525 183.615 ;
      LAYER nwell ;
        RECT 14.180 179.585 127.720 182.415 ;
      LAYER pwell ;
        RECT 14.375 178.385 15.745 179.195 ;
        RECT 15.755 178.385 18.505 179.195 ;
        RECT 18.515 178.385 24.025 179.195 ;
        RECT 24.045 178.470 24.475 179.255 ;
        RECT 29.005 179.065 29.935 179.285 ;
        RECT 32.765 179.065 33.685 179.295 ;
        RECT 24.495 178.385 33.685 179.065 ;
        RECT 33.790 179.065 34.710 179.295 ;
        RECT 33.790 178.385 37.255 179.065 ;
        RECT 37.835 178.385 41.310 179.295 ;
        RECT 41.975 178.385 45.450 179.295 ;
        RECT 48.855 179.065 49.785 179.295 ;
        RECT 45.885 178.385 49.785 179.065 ;
        RECT 49.805 178.470 50.235 179.255 ;
        RECT 52.910 179.065 53.830 179.295 ;
        RECT 50.365 178.385 53.830 179.065 ;
        RECT 53.935 178.385 55.765 179.195 ;
        RECT 55.775 179.065 56.705 179.295 ;
        RECT 55.775 178.385 59.675 179.065 ;
        RECT 59.925 178.385 62.665 179.065 ;
        RECT 62.675 178.385 65.425 179.195 ;
        RECT 65.445 178.385 66.795 179.295 ;
        RECT 66.815 179.065 68.160 179.295 ;
        RECT 66.815 178.385 68.645 179.065 ;
        RECT 68.655 178.385 71.395 179.065 ;
        RECT 71.655 178.615 74.410 179.295 ;
        RECT 71.655 178.385 73.925 178.615 ;
        RECT 75.565 178.470 75.995 179.255 ;
        RECT 78.670 179.065 79.590 179.295 ;
        RECT 76.125 178.385 79.590 179.065 ;
        RECT 79.890 178.385 83.365 179.295 ;
        RECT 83.375 178.385 85.205 179.195 ;
        RECT 88.415 179.065 89.345 179.295 ;
        RECT 85.445 178.385 89.345 179.065 ;
        RECT 89.355 178.385 90.725 179.165 ;
        RECT 90.745 178.385 92.095 179.295 ;
        RECT 92.115 179.065 93.035 179.295 ;
        RECT 95.865 179.065 96.795 179.285 ;
        RECT 92.115 178.385 101.305 179.065 ;
        RECT 101.325 178.470 101.755 179.255 ;
        RECT 101.870 179.065 102.790 179.295 ;
        RECT 105.550 179.065 106.470 179.295 ;
        RECT 101.870 178.385 105.335 179.065 ;
        RECT 105.550 178.385 109.015 179.065 ;
        RECT 109.605 178.385 110.955 179.295 ;
        RECT 110.975 179.065 111.895 179.295 ;
        RECT 114.725 179.065 115.655 179.285 ;
        RECT 110.975 178.385 120.165 179.065 ;
        RECT 120.185 178.385 121.535 179.295 ;
        RECT 121.555 178.385 122.925 179.165 ;
        RECT 123.395 178.385 126.145 179.195 ;
        RECT 126.155 178.385 127.525 179.195 ;
        RECT 14.515 178.175 14.685 178.385 ;
        RECT 18.195 178.195 18.365 178.385 ;
        RECT 19.115 178.175 19.285 178.365 ;
        RECT 23.715 178.195 23.885 178.385 ;
        RECT 24.635 178.175 24.805 178.385 ;
        RECT 26.015 178.175 26.185 178.365 ;
        RECT 26.475 178.175 26.645 178.365 ;
        RECT 36.595 178.175 36.765 178.365 ;
        RECT 37.055 178.195 37.225 178.385 ;
        RECT 37.570 178.225 37.690 178.335 ;
        RECT 37.980 178.195 38.150 178.385 ;
        RECT 40.920 178.175 41.090 178.365 ;
        RECT 41.710 178.225 41.830 178.335 ;
        RECT 42.120 178.330 42.290 178.385 ;
        RECT 42.115 178.220 42.290 178.330 ;
        RECT 42.120 178.195 42.290 178.220 ;
        RECT 42.575 178.175 42.745 178.365 ;
        RECT 49.200 178.195 49.370 178.385 ;
        RECT 49.470 178.175 49.640 178.365 ;
        RECT 49.935 178.175 50.105 178.365 ;
        RECT 50.395 178.195 50.565 178.385 ;
        RECT 55.455 178.195 55.625 178.385 ;
        RECT 56.190 178.195 56.360 178.385 ;
        RECT 62.355 178.175 62.525 178.385 ;
        RECT 64.195 178.175 64.365 178.365 ;
        RECT 65.115 178.195 65.285 178.385 ;
        RECT 65.575 178.195 65.745 178.385 ;
        RECT 66.955 178.175 67.125 178.365 ;
        RECT 68.335 178.195 68.505 178.385 ;
        RECT 68.795 178.175 68.965 178.385 ;
        RECT 71.655 178.365 71.725 178.385 ;
        RECT 69.255 178.175 69.425 178.365 ;
        RECT 71.095 178.175 71.265 178.365 ;
        RECT 71.555 178.195 71.725 178.365 ;
        RECT 75.235 178.175 75.405 178.365 ;
        RECT 75.750 178.225 75.870 178.335 ;
        RECT 76.155 178.195 76.325 178.385 ;
        RECT 79.370 178.175 79.540 178.365 ;
        RECT 79.840 178.175 80.010 178.365 ;
        RECT 83.050 178.195 83.220 178.385 ;
        RECT 84.435 178.175 84.605 178.365 ;
        RECT 84.895 178.175 85.065 178.385 ;
        RECT 88.760 178.195 88.930 178.385 ;
        RECT 90.415 178.195 90.585 178.385 ;
        RECT 90.875 178.195 91.045 178.385 ;
        RECT 92.255 178.175 92.425 178.365 ;
        RECT 97.775 178.175 97.945 178.365 ;
        RECT 100.995 178.195 101.165 178.385 ;
        RECT 101.450 178.175 101.620 178.365 ;
        RECT 102.835 178.175 103.005 178.365 ;
        RECT 104.215 178.175 104.385 178.365 ;
        RECT 104.680 178.175 104.850 178.365 ;
        RECT 105.135 178.195 105.305 178.385 ;
        RECT 108.815 178.195 108.985 178.385 ;
        RECT 109.330 178.225 109.450 178.335 ;
        RECT 109.735 178.175 109.905 178.385 ;
        RECT 113.600 178.175 113.770 178.365 ;
        RECT 116.175 178.175 116.345 178.365 ;
        RECT 116.635 178.175 116.805 178.365 ;
        RECT 119.855 178.195 120.025 178.385 ;
        RECT 120.315 178.175 120.485 178.385 ;
        RECT 121.695 178.195 121.865 178.385 ;
        RECT 123.130 178.225 123.250 178.335 ;
        RECT 125.835 178.175 126.005 178.385 ;
        RECT 127.215 178.175 127.385 178.385 ;
        RECT 14.375 177.365 15.745 178.175 ;
        RECT 15.755 177.365 19.425 178.175 ;
        RECT 19.435 177.365 24.945 178.175 ;
        RECT 24.965 177.265 26.315 178.175 ;
        RECT 26.345 177.265 27.695 178.175 ;
        RECT 27.715 177.495 36.905 178.175 ;
        RECT 27.715 177.265 28.635 177.495 ;
        RECT 31.465 177.275 32.395 177.495 ;
        RECT 36.925 177.305 37.355 178.090 ;
        RECT 37.605 177.495 41.505 178.175 ;
        RECT 42.545 177.495 46.010 178.175 ;
        RECT 40.575 177.265 41.505 177.495 ;
        RECT 45.090 177.265 46.010 177.495 ;
        RECT 46.310 177.265 49.785 178.175 ;
        RECT 49.905 177.495 53.370 178.175 ;
        RECT 52.450 177.265 53.370 177.495 ;
        RECT 53.475 177.495 62.665 178.175 ;
        RECT 53.475 177.265 54.395 177.495 ;
        RECT 57.225 177.275 58.155 177.495 ;
        RECT 62.685 177.305 63.115 178.090 ;
        RECT 63.135 177.395 64.505 178.175 ;
        RECT 64.515 177.365 67.265 178.175 ;
        RECT 67.275 177.495 69.105 178.175 ;
        RECT 69.115 177.495 70.945 178.175 ;
        RECT 70.955 177.495 72.785 178.175 ;
        RECT 67.275 177.265 68.620 177.495 ;
        RECT 69.600 177.265 70.945 177.495 ;
        RECT 71.440 177.265 72.785 177.495 ;
        RECT 72.825 177.265 75.545 178.175 ;
        RECT 76.210 177.265 79.685 178.175 ;
        RECT 79.695 177.265 83.170 178.175 ;
        RECT 83.375 177.365 84.745 178.175 ;
        RECT 84.865 177.495 88.330 178.175 ;
        RECT 87.410 177.265 88.330 177.495 ;
        RECT 88.445 177.305 88.875 178.090 ;
        RECT 88.895 177.365 92.565 178.175 ;
        RECT 92.575 177.365 98.085 178.175 ;
        RECT 98.290 177.265 101.765 178.175 ;
        RECT 101.775 177.395 103.145 178.175 ;
        RECT 103.155 177.365 104.525 178.175 ;
        RECT 104.535 177.265 108.010 178.175 ;
        RECT 108.215 177.365 110.045 178.175 ;
        RECT 110.285 177.495 114.185 178.175 ;
        RECT 113.255 177.265 114.185 177.495 ;
        RECT 114.205 177.305 114.635 178.090 ;
        RECT 114.655 177.365 116.485 178.175 ;
        RECT 116.495 177.395 117.865 178.175 ;
        RECT 117.875 177.365 120.625 178.175 ;
        RECT 120.635 177.365 126.145 178.175 ;
        RECT 126.155 177.365 127.525 178.175 ;
      LAYER nwell ;
        RECT 14.180 174.145 127.720 176.975 ;
      LAYER pwell ;
        RECT 14.375 172.945 15.745 173.755 ;
        RECT 15.755 172.945 18.505 173.755 ;
        RECT 18.515 172.945 24.025 173.755 ;
        RECT 24.045 173.030 24.475 173.815 ;
        RECT 25.415 172.945 26.785 173.725 ;
        RECT 29.450 173.625 30.370 173.855 ;
        RECT 26.905 172.945 30.370 173.625 ;
        RECT 30.475 173.625 31.405 173.855 ;
        RECT 30.475 172.945 34.375 173.625 ;
        RECT 35.270 172.945 38.745 173.855 ;
        RECT 38.755 172.945 42.230 173.855 ;
        RECT 42.630 172.945 46.105 173.855 ;
        RECT 48.770 173.625 49.690 173.855 ;
        RECT 46.225 172.945 49.690 173.625 ;
        RECT 49.805 173.030 50.235 173.815 ;
        RECT 50.255 172.945 53.005 173.755 ;
        RECT 56.215 173.625 57.145 173.855 ;
        RECT 53.245 172.945 57.145 173.625 ;
        RECT 57.155 173.625 58.075 173.855 ;
        RECT 60.905 173.625 61.835 173.845 ;
        RECT 57.155 172.945 66.345 173.625 ;
        RECT 66.355 172.945 68.185 173.755 ;
        RECT 68.195 172.945 70.805 173.855 ;
        RECT 70.955 173.625 72.300 173.855 ;
        RECT 70.955 172.945 72.785 173.625 ;
        RECT 72.795 172.945 75.545 173.755 ;
        RECT 75.565 173.030 75.995 173.815 ;
        RECT 76.935 172.945 80.605 173.755 ;
        RECT 80.615 172.945 84.090 173.855 ;
        RECT 84.755 172.945 90.265 173.755 ;
        RECT 90.275 172.945 95.785 173.755 ;
        RECT 95.795 172.945 101.305 173.755 ;
        RECT 101.325 173.030 101.755 173.815 ;
        RECT 101.775 172.945 103.605 173.755 ;
        RECT 103.810 172.945 107.285 173.855 ;
        RECT 107.295 172.945 110.770 173.855 ;
        RECT 110.975 172.945 112.345 173.755 ;
        RECT 112.355 172.945 117.865 173.755 ;
        RECT 117.885 172.945 119.235 173.855 ;
        RECT 119.255 172.945 120.625 173.755 ;
        RECT 120.635 172.945 126.145 173.755 ;
        RECT 126.155 172.945 127.525 173.755 ;
        RECT 14.515 172.735 14.685 172.945 ;
        RECT 16.355 172.780 16.515 172.890 ;
        RECT 18.195 172.755 18.365 172.945 ;
        RECT 20.035 172.735 20.205 172.925 ;
        RECT 23.715 172.755 23.885 172.945 ;
        RECT 25.095 172.790 25.255 172.900 ;
        RECT 25.555 172.735 25.725 172.925 ;
        RECT 26.475 172.755 26.645 172.945 ;
        RECT 26.935 172.755 27.105 172.945 ;
        RECT 30.890 172.755 31.060 172.945 ;
        RECT 31.075 172.735 31.245 172.925 ;
        RECT 34.810 172.785 34.930 172.895 ;
        RECT 36.595 172.735 36.765 172.925 ;
        RECT 37.520 172.735 37.690 172.925 ;
        RECT 38.430 172.755 38.600 172.945 ;
        RECT 38.900 172.755 39.070 172.945 ;
        RECT 41.250 172.785 41.370 172.895 ;
        RECT 42.575 172.735 42.745 172.925 ;
        RECT 43.495 172.780 43.655 172.890 ;
        RECT 43.960 172.735 44.130 172.925 ;
        RECT 45.790 172.755 45.960 172.945 ;
        RECT 46.255 172.755 46.425 172.945 ;
        RECT 47.640 172.735 47.810 172.925 ;
        RECT 51.320 172.735 51.490 172.925 ;
        RECT 52.695 172.755 52.865 172.945 ;
        RECT 55.915 172.735 56.085 172.925 ;
        RECT 56.560 172.755 56.730 172.945 ;
        RECT 59.595 172.735 59.765 172.925 ;
        RECT 60.975 172.735 61.145 172.925 ;
        RECT 61.435 172.735 61.605 172.925 ;
        RECT 63.330 172.785 63.450 172.895 ;
        RECT 65.115 172.735 65.285 172.925 ;
        RECT 66.035 172.755 66.205 172.945 ;
        RECT 67.875 172.755 68.045 172.945 ;
        RECT 68.340 172.755 68.510 172.945 ;
        RECT 70.635 172.735 70.805 172.925 ;
        RECT 72.475 172.755 72.645 172.945 ;
        RECT 75.235 172.755 75.405 172.945 ;
        RECT 76.155 172.735 76.325 172.925 ;
        RECT 76.615 172.790 76.775 172.900 ;
        RECT 80.295 172.755 80.465 172.945 ;
        RECT 80.760 172.755 80.930 172.945 ;
        RECT 81.675 172.735 81.845 172.925 ;
        RECT 82.140 172.735 82.310 172.925 ;
        RECT 84.490 172.785 84.610 172.895 ;
        RECT 84.895 172.735 85.065 172.925 ;
        RECT 89.090 172.785 89.210 172.895 ;
        RECT 89.495 172.735 89.665 172.925 ;
        RECT 89.955 172.755 90.125 172.945 ;
        RECT 95.475 172.755 95.645 172.945 ;
        RECT 99.615 172.735 99.785 172.925 ;
        RECT 100.535 172.780 100.695 172.890 ;
        RECT 100.995 172.755 101.165 172.945 ;
        RECT 103.295 172.755 103.465 172.945 ;
        RECT 106.055 172.735 106.225 172.925 ;
        RECT 106.970 172.755 107.140 172.945 ;
        RECT 107.440 172.925 107.610 172.945 ;
        RECT 107.435 172.755 107.610 172.925 ;
        RECT 107.435 172.735 107.605 172.755 ;
        RECT 111.110 172.735 111.280 172.925 ;
        RECT 112.035 172.755 112.205 172.945 ;
        RECT 112.495 172.735 112.665 172.925 ;
        RECT 112.955 172.735 113.125 172.925 ;
        RECT 115.255 172.780 115.415 172.890 ;
        RECT 117.555 172.755 117.725 172.945 ;
        RECT 118.015 172.755 118.185 172.945 ;
        RECT 120.315 172.755 120.485 172.945 ;
        RECT 124.455 172.735 124.625 172.925 ;
        RECT 125.835 172.735 126.005 172.945 ;
        RECT 127.215 172.735 127.385 172.945 ;
        RECT 14.375 171.925 15.745 172.735 ;
        RECT 16.675 171.925 20.345 172.735 ;
        RECT 20.355 171.925 25.865 172.735 ;
        RECT 25.875 171.925 31.385 172.735 ;
        RECT 31.395 171.925 36.905 172.735 ;
        RECT 36.925 171.865 37.355 172.650 ;
        RECT 37.375 171.825 40.850 172.735 ;
        RECT 41.515 171.955 42.885 172.735 ;
        RECT 43.815 171.825 47.290 172.735 ;
        RECT 47.495 171.825 50.970 172.735 ;
        RECT 51.175 171.825 54.650 172.735 ;
        RECT 54.855 171.925 56.225 172.735 ;
        RECT 56.235 171.925 59.905 172.735 ;
        RECT 59.925 171.825 61.275 172.735 ;
        RECT 61.295 171.955 62.665 172.735 ;
        RECT 62.685 171.865 63.115 172.650 ;
        RECT 63.595 171.925 65.425 172.735 ;
        RECT 65.435 171.925 70.945 172.735 ;
        RECT 70.955 171.925 76.465 172.735 ;
        RECT 76.475 171.925 81.985 172.735 ;
        RECT 81.995 171.825 84.605 172.735 ;
        RECT 84.865 172.055 88.330 172.735 ;
        RECT 87.410 171.825 88.330 172.055 ;
        RECT 88.445 171.865 88.875 172.650 ;
        RECT 89.365 171.825 90.715 172.735 ;
        RECT 90.735 172.055 99.925 172.735 ;
        RECT 90.735 171.825 91.655 172.055 ;
        RECT 94.485 171.835 95.415 172.055 ;
        RECT 100.855 171.925 106.365 172.735 ;
        RECT 106.385 171.825 107.735 172.735 ;
        RECT 107.950 171.825 111.425 172.735 ;
        RECT 111.435 171.925 112.805 172.735 ;
        RECT 112.825 171.825 114.175 172.735 ;
        RECT 114.205 171.865 114.635 172.650 ;
        RECT 115.575 172.055 124.765 172.735 ;
        RECT 115.575 171.825 116.495 172.055 ;
        RECT 119.325 171.835 120.255 172.055 ;
        RECT 124.775 171.925 126.145 172.735 ;
        RECT 126.155 171.925 127.525 172.735 ;
      LAYER nwell ;
        RECT 14.180 168.705 127.720 171.535 ;
      LAYER pwell ;
        RECT 14.375 167.505 15.745 168.315 ;
        RECT 15.755 167.505 18.505 168.315 ;
        RECT 18.515 167.505 24.025 168.315 ;
        RECT 24.045 167.590 24.475 168.375 ;
        RECT 24.955 167.505 26.785 168.315 ;
        RECT 26.805 167.505 28.155 168.415 ;
        RECT 28.635 167.505 32.305 168.315 ;
        RECT 32.325 167.505 33.675 168.415 ;
        RECT 33.695 167.505 35.065 168.315 ;
        RECT 35.160 167.505 44.265 168.185 ;
        RECT 44.275 167.505 49.785 168.315 ;
        RECT 49.805 167.590 50.235 168.375 ;
        RECT 50.255 167.505 51.625 168.315 ;
        RECT 51.635 167.505 57.145 168.315 ;
        RECT 57.155 167.505 62.665 168.315 ;
        RECT 62.675 167.505 68.185 168.315 ;
        RECT 68.195 168.185 69.540 168.415 ;
        RECT 70.035 168.185 71.380 168.415 ;
        RECT 68.195 167.505 70.025 168.185 ;
        RECT 70.035 167.505 71.865 168.185 ;
        RECT 71.875 167.505 75.545 168.315 ;
        RECT 75.565 167.590 75.995 168.375 ;
        RECT 79.215 168.185 80.145 168.415 ;
        RECT 76.245 167.505 80.145 168.185 ;
        RECT 80.525 168.305 81.445 168.415 ;
        RECT 80.525 168.185 82.860 168.305 ;
        RECT 87.525 168.185 88.445 168.405 ;
        RECT 80.525 167.505 89.805 168.185 ;
        RECT 89.815 167.505 91.185 168.315 ;
        RECT 94.395 168.185 95.325 168.415 ;
        RECT 91.425 167.505 95.325 168.185 ;
        RECT 95.795 167.505 97.165 168.285 ;
        RECT 97.635 167.505 101.305 168.315 ;
        RECT 101.325 167.590 101.755 168.375 ;
        RECT 102.695 168.185 103.615 168.415 ;
        RECT 106.445 168.185 107.375 168.405 ;
        RECT 112.355 168.185 113.285 168.415 ;
        RECT 116.590 168.185 117.510 168.415 ;
        RECT 102.695 167.505 111.885 168.185 ;
        RECT 112.355 167.505 116.255 168.185 ;
        RECT 116.590 167.505 120.055 168.185 ;
        RECT 120.175 167.505 121.545 168.285 ;
        RECT 121.555 167.505 123.385 168.185 ;
        RECT 123.395 167.505 126.145 168.315 ;
        RECT 126.155 167.505 127.525 168.315 ;
        RECT 14.515 167.295 14.685 167.505 ;
        RECT 17.275 167.295 17.445 167.485 ;
        RECT 18.195 167.315 18.365 167.505 ;
        RECT 22.795 167.295 22.965 167.485 ;
        RECT 23.255 167.295 23.425 167.485 ;
        RECT 23.715 167.315 23.885 167.505 ;
        RECT 24.690 167.345 24.810 167.455 ;
        RECT 26.475 167.315 26.645 167.505 ;
        RECT 26.935 167.315 27.105 167.505 ;
        RECT 28.370 167.345 28.490 167.455 ;
        RECT 31.995 167.315 32.165 167.505 ;
        RECT 33.375 167.295 33.545 167.505 ;
        RECT 34.755 167.315 34.925 167.505 ;
        RECT 36.595 167.295 36.765 167.485 ;
        RECT 37.515 167.295 37.685 167.485 ;
        RECT 38.895 167.295 39.065 167.485 ;
        RECT 43.955 167.315 44.125 167.505 ;
        RECT 45.795 167.295 45.965 167.485 ;
        RECT 46.715 167.340 46.875 167.450 ;
        RECT 49.475 167.315 49.645 167.505 ;
        RECT 51.315 167.315 51.485 167.505 ;
        RECT 55.915 167.295 56.085 167.485 ;
        RECT 56.835 167.315 57.005 167.505 ;
        RECT 62.355 167.485 62.525 167.505 ;
        RECT 57.755 167.295 57.925 167.485 ;
        RECT 59.135 167.295 59.305 167.485 ;
        RECT 59.650 167.345 59.770 167.455 ;
        RECT 62.350 167.315 62.525 167.485 ;
        RECT 62.350 167.295 62.520 167.315 ;
        RECT 64.655 167.295 64.825 167.485 ;
        RECT 67.415 167.295 67.585 167.485 ;
        RECT 67.875 167.295 68.045 167.505 ;
        RECT 69.715 167.315 69.885 167.505 ;
        RECT 70.635 167.295 70.805 167.485 ;
        RECT 71.555 167.315 71.725 167.505 ;
        RECT 74.775 167.295 74.945 167.485 ;
        RECT 75.235 167.315 75.405 167.505 ;
        RECT 79.560 167.315 79.730 167.505 ;
        RECT 84.435 167.295 84.605 167.485 ;
        RECT 85.815 167.295 85.985 167.485 ;
        RECT 87.195 167.295 87.365 167.485 ;
        RECT 88.115 167.340 88.275 167.450 ;
        RECT 89.090 167.345 89.210 167.455 ;
        RECT 89.495 167.315 89.665 167.505 ;
        RECT 90.875 167.315 91.045 167.505 ;
        RECT 92.715 167.295 92.885 167.485 ;
        RECT 94.740 167.315 94.910 167.505 ;
        RECT 95.530 167.345 95.650 167.455 ;
        RECT 95.935 167.315 96.105 167.505 ;
        RECT 96.580 167.295 96.750 167.485 ;
        RECT 97.370 167.345 97.490 167.455 ;
        RECT 100.995 167.315 101.165 167.505 ;
        RECT 102.375 167.350 102.535 167.460 ;
        RECT 106.515 167.295 106.685 167.485 ;
        RECT 106.975 167.295 107.145 167.485 ;
        RECT 110.655 167.295 110.825 167.485 ;
        RECT 111.575 167.315 111.745 167.505 ;
        RECT 112.090 167.345 112.210 167.455 ;
        RECT 112.770 167.315 112.940 167.505 ;
        RECT 115.255 167.340 115.415 167.450 ;
        RECT 119.855 167.315 120.025 167.505 ;
        RECT 120.315 167.315 120.485 167.505 ;
        RECT 123.075 167.315 123.245 167.505 ;
        RECT 124.455 167.295 124.625 167.485 ;
        RECT 125.835 167.295 126.005 167.505 ;
        RECT 127.215 167.295 127.385 167.505 ;
        RECT 14.375 166.485 15.745 167.295 ;
        RECT 15.755 166.485 17.585 167.295 ;
        RECT 17.595 166.485 23.105 167.295 ;
        RECT 23.115 166.615 32.305 167.295 ;
        RECT 27.625 166.395 28.555 166.615 ;
        RECT 31.385 166.385 32.305 166.615 ;
        RECT 32.315 166.515 33.685 167.295 ;
        RECT 33.695 166.385 36.855 167.295 ;
        RECT 36.925 166.425 37.355 167.210 ;
        RECT 37.385 166.385 38.735 167.295 ;
        RECT 38.865 166.615 42.330 167.295 ;
        RECT 41.410 166.385 42.330 166.615 ;
        RECT 42.530 166.615 45.995 167.295 ;
        RECT 47.035 166.615 56.225 167.295 ;
        RECT 42.530 166.385 43.450 166.615 ;
        RECT 47.035 166.385 47.955 166.615 ;
        RECT 50.785 166.395 51.715 166.615 ;
        RECT 56.235 166.485 58.065 167.295 ;
        RECT 58.085 166.385 59.435 167.295 ;
        RECT 60.055 166.385 62.665 167.295 ;
        RECT 62.685 166.425 63.115 167.210 ;
        RECT 63.135 166.485 64.965 167.295 ;
        RECT 64.985 166.615 67.725 167.295 ;
        RECT 67.735 166.615 70.475 167.295 ;
        RECT 70.495 166.385 73.215 167.295 ;
        RECT 73.255 166.485 75.085 167.295 ;
        RECT 75.465 166.615 84.745 167.295 ;
        RECT 75.465 166.495 77.800 166.615 ;
        RECT 75.465 166.385 76.385 166.495 ;
        RECT 82.465 166.395 83.385 166.615 ;
        RECT 84.765 166.385 86.115 167.295 ;
        RECT 86.145 166.385 87.495 167.295 ;
        RECT 88.445 166.425 88.875 167.210 ;
        RECT 89.355 166.485 93.025 167.295 ;
        RECT 93.265 166.615 97.165 167.295 ;
        RECT 96.235 166.385 97.165 166.615 ;
        RECT 97.545 166.615 106.825 167.295 ;
        RECT 106.945 166.615 110.410 167.295 ;
        RECT 110.625 166.615 114.090 167.295 ;
        RECT 97.545 166.495 99.880 166.615 ;
        RECT 97.545 166.385 98.465 166.495 ;
        RECT 104.545 166.395 105.465 166.615 ;
        RECT 109.490 166.385 110.410 166.615 ;
        RECT 113.170 166.385 114.090 166.615 ;
        RECT 114.205 166.425 114.635 167.210 ;
        RECT 115.575 166.615 124.765 167.295 ;
        RECT 115.575 166.385 116.495 166.615 ;
        RECT 119.325 166.395 120.255 166.615 ;
        RECT 124.775 166.485 126.145 167.295 ;
        RECT 126.155 166.485 127.525 167.295 ;
      LAYER nwell ;
        RECT 14.180 163.265 127.720 166.095 ;
      LAYER pwell ;
        RECT 14.375 162.065 15.745 162.875 ;
        RECT 15.755 162.065 18.505 162.875 ;
        RECT 18.515 162.065 24.025 162.875 ;
        RECT 24.045 162.150 24.475 162.935 ;
        RECT 25.415 162.065 26.785 162.845 ;
        RECT 31.305 162.745 32.235 162.965 ;
        RECT 35.065 162.745 35.985 162.975 ;
        RECT 26.795 162.065 35.985 162.745 ;
        RECT 35.995 162.745 36.915 162.975 ;
        RECT 39.745 162.745 40.675 162.965 ;
        RECT 48.770 162.745 49.690 162.975 ;
        RECT 35.995 162.065 45.185 162.745 ;
        RECT 46.225 162.065 49.690 162.745 ;
        RECT 49.805 162.150 50.235 162.935 ;
        RECT 50.265 162.065 51.615 162.975 ;
        RECT 51.635 162.065 53.465 162.875 ;
        RECT 53.475 162.065 54.845 162.845 ;
        RECT 54.855 162.745 55.775 162.975 ;
        RECT 58.605 162.745 59.535 162.965 ;
        RECT 54.855 162.065 64.045 162.745 ;
        RECT 64.195 162.065 66.805 162.975 ;
        RECT 66.825 162.065 69.565 162.745 ;
        RECT 70.035 162.065 75.545 162.875 ;
        RECT 75.565 162.150 75.995 162.935 ;
        RECT 76.015 162.065 77.845 162.875 ;
        RECT 81.055 162.745 81.985 162.975 ;
        RECT 78.085 162.065 81.985 162.745 ;
        RECT 81.995 162.065 83.365 162.845 ;
        RECT 83.375 162.065 85.205 162.875 ;
        RECT 85.215 162.065 86.585 162.845 ;
        RECT 86.595 162.065 92.105 162.875 ;
        RECT 92.200 162.065 101.305 162.745 ;
        RECT 101.325 162.150 101.755 162.935 ;
        RECT 104.975 162.745 105.905 162.975 ;
        RECT 102.005 162.065 105.905 162.745 ;
        RECT 106.375 162.745 107.305 162.975 ;
        RECT 106.375 162.065 110.275 162.745 ;
        RECT 110.655 162.065 113.265 162.975 ;
        RECT 113.275 162.745 114.195 162.975 ;
        RECT 117.025 162.745 117.955 162.965 ;
        RECT 113.275 162.065 122.465 162.745 ;
        RECT 122.475 162.065 123.845 162.845 ;
        RECT 124.315 162.065 126.145 162.875 ;
        RECT 126.155 162.065 127.525 162.875 ;
        RECT 14.515 161.855 14.685 162.065 ;
        RECT 17.275 161.855 17.445 162.045 ;
        RECT 18.195 161.875 18.365 162.065 ;
        RECT 23.715 161.875 23.885 162.065 ;
        RECT 25.095 161.910 25.255 162.020 ;
        RECT 26.475 161.875 26.645 162.065 ;
        RECT 26.935 161.855 27.105 162.065 ;
        RECT 27.670 161.855 27.840 162.045 ;
        RECT 32.455 161.855 32.625 162.045 ;
        RECT 33.190 161.855 33.360 162.045 ;
        RECT 37.570 161.905 37.690 162.015 ;
        RECT 39.355 161.855 39.525 162.045 ;
        RECT 39.815 161.855 39.985 162.045 ;
        RECT 43.770 161.855 43.940 162.045 ;
        RECT 44.875 161.875 45.045 162.065 ;
        RECT 45.795 161.910 45.955 162.020 ;
        RECT 46.255 161.875 46.425 162.065 ;
        RECT 48.555 161.855 48.725 162.045 ;
        RECT 49.290 161.855 49.460 162.045 ;
        RECT 51.315 161.875 51.485 162.065 ;
        RECT 53.155 161.875 53.325 162.065 ;
        RECT 53.615 161.875 53.785 162.065 ;
        RECT 56.560 161.855 56.730 162.045 ;
        RECT 57.350 161.905 57.470 162.015 ;
        RECT 59.135 161.855 59.305 162.045 ;
        RECT 59.595 161.855 59.765 162.045 ;
        RECT 62.355 161.855 62.525 162.045 ;
        RECT 63.735 161.875 63.905 162.065 ;
        RECT 64.195 161.855 64.365 162.045 ;
        RECT 66.035 161.855 66.205 162.045 ;
        RECT 66.490 161.875 66.660 162.065 ;
        RECT 67.875 161.855 68.045 162.045 ;
        RECT 68.335 161.855 68.505 162.045 ;
        RECT 69.255 161.875 69.425 162.065 ;
        RECT 69.770 161.905 69.890 162.015 ;
        RECT 70.175 161.855 70.345 162.045 ;
        RECT 72.070 161.905 72.190 162.015 ;
        RECT 74.775 161.855 74.945 162.045 ;
        RECT 75.235 161.875 75.405 162.065 ;
        RECT 77.535 161.875 77.705 162.065 ;
        RECT 80.295 161.855 80.465 162.045 ;
        RECT 81.400 161.875 81.570 162.065 ;
        RECT 81.675 161.855 81.845 162.045 ;
        RECT 82.135 161.875 82.305 162.065 ;
        RECT 84.895 161.875 85.065 162.065 ;
        RECT 85.355 161.875 85.525 162.065 ;
        RECT 85.540 161.855 85.710 162.045 ;
        RECT 86.275 161.855 86.445 162.045 ;
        RECT 88.115 161.900 88.275 162.010 ;
        RECT 89.090 161.905 89.210 162.015 ;
        RECT 91.795 161.875 91.965 162.065 ;
        RECT 98.695 161.855 98.865 162.045 ;
        RECT 100.995 161.875 101.165 162.065 ;
        RECT 101.915 161.855 102.085 162.045 ;
        RECT 102.375 161.855 102.545 162.045 ;
        RECT 105.320 161.875 105.490 162.065 ;
        RECT 106.110 161.905 106.230 162.015 ;
        RECT 106.515 161.855 106.685 162.045 ;
        RECT 106.790 161.875 106.960 162.065 ;
        RECT 112.950 161.875 113.120 162.065 ;
        RECT 113.600 161.855 113.770 162.045 ;
        RECT 118.200 161.855 118.370 162.045 ;
        RECT 118.935 161.855 119.105 162.045 ;
        RECT 120.370 161.905 120.490 162.015 ;
        RECT 120.775 161.855 120.945 162.045 ;
        RECT 122.155 162.015 122.325 162.065 ;
        RECT 122.155 161.905 122.330 162.015 ;
        RECT 122.155 161.875 122.325 161.905 ;
        RECT 123.535 161.875 123.705 162.065 ;
        RECT 124.050 161.905 124.170 162.015 ;
        RECT 125.835 161.855 126.005 162.065 ;
        RECT 127.215 161.855 127.385 162.065 ;
        RECT 14.375 161.045 15.745 161.855 ;
        RECT 15.755 161.045 17.585 161.855 ;
        RECT 17.965 161.175 27.245 161.855 ;
        RECT 27.255 161.175 31.155 161.855 ;
        RECT 17.965 161.055 20.300 161.175 ;
        RECT 17.965 160.945 18.885 161.055 ;
        RECT 24.965 160.955 25.885 161.175 ;
        RECT 27.255 160.945 28.185 161.175 ;
        RECT 31.395 161.045 32.765 161.855 ;
        RECT 32.775 161.175 36.675 161.855 ;
        RECT 32.775 160.945 33.705 161.175 ;
        RECT 36.925 160.985 37.355 161.770 ;
        RECT 37.835 161.045 39.665 161.855 ;
        RECT 39.785 161.175 43.250 161.855 ;
        RECT 42.330 160.945 43.250 161.175 ;
        RECT 43.355 161.175 47.255 161.855 ;
        RECT 43.355 160.945 44.285 161.175 ;
        RECT 47.495 161.075 48.865 161.855 ;
        RECT 48.875 161.175 52.775 161.855 ;
        RECT 53.245 161.175 57.145 161.855 ;
        RECT 48.875 160.945 49.805 161.175 ;
        RECT 56.215 160.945 57.145 161.175 ;
        RECT 57.615 161.045 59.445 161.855 ;
        RECT 59.455 161.075 60.825 161.855 ;
        RECT 60.835 161.045 62.665 161.855 ;
        RECT 62.685 160.985 63.115 161.770 ;
        RECT 63.135 161.045 64.505 161.855 ;
        RECT 64.515 161.175 66.345 161.855 ;
        RECT 66.355 161.175 68.185 161.855 ;
        RECT 68.195 161.175 70.025 161.855 ;
        RECT 70.035 161.175 71.865 161.855 ;
        RECT 64.515 160.945 65.860 161.175 ;
        RECT 66.355 160.945 67.700 161.175 ;
        RECT 68.680 160.945 70.025 161.175 ;
        RECT 70.520 160.945 71.865 161.175 ;
        RECT 72.335 161.045 75.085 161.855 ;
        RECT 75.095 161.045 80.605 161.855 ;
        RECT 80.625 160.945 81.975 161.855 ;
        RECT 82.225 161.175 86.125 161.855 ;
        RECT 85.195 160.945 86.125 161.175 ;
        RECT 86.135 161.075 87.505 161.855 ;
        RECT 88.445 160.985 88.875 161.770 ;
        RECT 89.725 161.175 99.005 161.855 ;
        RECT 89.725 161.055 92.060 161.175 ;
        RECT 89.725 160.945 90.645 161.055 ;
        RECT 96.725 160.955 97.645 161.175 ;
        RECT 99.015 160.945 102.175 161.855 ;
        RECT 102.345 161.175 105.810 161.855 ;
        RECT 106.485 161.175 109.950 161.855 ;
        RECT 110.285 161.175 114.185 161.855 ;
        RECT 104.890 160.945 105.810 161.175 ;
        RECT 109.030 160.945 109.950 161.175 ;
        RECT 113.255 160.945 114.185 161.175 ;
        RECT 114.205 160.985 114.635 161.770 ;
        RECT 114.885 161.175 118.785 161.855 ;
        RECT 117.855 160.945 118.785 161.175 ;
        RECT 118.805 160.945 120.155 161.855 ;
        RECT 120.635 161.075 122.005 161.855 ;
        RECT 122.475 161.045 126.145 161.855 ;
        RECT 126.155 161.045 127.525 161.855 ;
      LAYER nwell ;
        RECT 14.180 157.825 127.720 160.655 ;
      LAYER pwell ;
        RECT 14.375 156.625 15.745 157.435 ;
        RECT 15.755 156.625 17.125 157.435 ;
        RECT 17.145 156.625 18.495 157.535 ;
        RECT 18.525 156.625 19.875 157.535 ;
        RECT 23.095 157.305 24.025 157.535 ;
        RECT 20.125 156.625 24.025 157.305 ;
        RECT 24.045 156.710 24.475 157.495 ;
        RECT 24.495 156.625 25.865 157.405 ;
        RECT 25.875 156.625 27.705 157.435 ;
        RECT 30.370 157.305 31.290 157.535 ;
        RECT 34.050 157.305 34.970 157.535 ;
        RECT 27.825 156.625 31.290 157.305 ;
        RECT 31.505 156.625 34.970 157.305 ;
        RECT 35.075 156.625 38.745 157.435 ;
        RECT 38.950 156.625 42.425 157.535 ;
        RECT 42.630 156.625 46.105 157.535 ;
        RECT 48.770 157.305 49.690 157.535 ;
        RECT 46.225 156.625 49.690 157.305 ;
        RECT 49.805 156.710 50.235 157.495 ;
        RECT 50.255 156.625 53.730 157.535 ;
        RECT 54.395 156.625 59.905 157.435 ;
        RECT 59.925 156.625 61.275 157.535 ;
        RECT 61.435 156.625 64.045 157.535 ;
        RECT 64.515 156.625 68.185 157.435 ;
        RECT 68.680 157.305 70.025 157.535 ;
        RECT 70.520 157.305 71.865 157.535 ;
        RECT 68.195 156.625 70.025 157.305 ;
        RECT 70.035 156.625 71.865 157.305 ;
        RECT 72.070 156.625 75.545 157.535 ;
        RECT 75.565 156.710 75.995 157.495 ;
        RECT 76.670 156.625 80.145 157.535 ;
        RECT 80.985 157.425 81.905 157.535 ;
        RECT 80.985 157.305 83.320 157.425 ;
        RECT 87.985 157.305 88.905 157.525 ;
        RECT 80.985 156.625 90.265 157.305 ;
        RECT 90.735 156.625 92.565 157.435 ;
        RECT 92.585 156.625 93.935 157.535 ;
        RECT 94.415 156.625 96.245 157.435 ;
        RECT 96.255 156.625 97.625 157.405 ;
        RECT 97.635 156.625 99.465 157.435 ;
        RECT 99.485 156.625 100.835 157.535 ;
        RECT 101.325 156.710 101.755 157.495 ;
        RECT 102.235 156.625 104.065 157.435 ;
        RECT 104.075 156.625 105.445 157.405 ;
        RECT 105.455 156.625 106.825 157.405 ;
        RECT 107.755 156.625 111.230 157.535 ;
        RECT 112.355 156.625 116.025 157.435 ;
        RECT 118.690 157.305 119.610 157.535 ;
        RECT 116.145 156.625 119.610 157.305 ;
        RECT 120.635 156.625 126.145 157.435 ;
        RECT 126.155 156.625 127.525 157.435 ;
        RECT 14.515 156.415 14.685 156.625 ;
        RECT 16.355 156.460 16.515 156.570 ;
        RECT 16.815 156.435 16.985 156.625 ;
        RECT 18.195 156.435 18.365 156.625 ;
        RECT 18.655 156.435 18.825 156.625 ;
        RECT 23.440 156.435 23.610 156.625 ;
        RECT 24.635 156.435 24.805 156.625 ;
        RECT 26.015 156.415 26.185 156.605 ;
        RECT 27.395 156.415 27.565 156.625 ;
        RECT 27.855 156.435 28.025 156.625 ;
        RECT 28.775 156.415 28.945 156.605 ;
        RECT 31.535 156.435 31.705 156.625 ;
        RECT 32.455 156.415 32.625 156.605 ;
        RECT 36.320 156.415 36.490 156.605 ;
        RECT 37.570 156.465 37.690 156.575 ;
        RECT 38.435 156.435 38.605 156.625 ;
        RECT 39.355 156.415 39.525 156.605 ;
        RECT 39.820 156.415 39.990 156.605 ;
        RECT 42.110 156.435 42.280 156.625 ;
        RECT 43.500 156.415 43.670 156.605 ;
        RECT 45.790 156.435 45.960 156.625 ;
        RECT 46.255 156.435 46.425 156.625 ;
        RECT 47.180 156.415 47.350 156.605 ;
        RECT 50.400 156.435 50.570 156.625 ;
        RECT 50.910 156.465 51.030 156.575 ;
        RECT 52.695 156.415 52.865 156.605 ;
        RECT 54.130 156.465 54.250 156.575 ;
        RECT 59.595 156.435 59.765 156.625 ;
        RECT 60.975 156.435 61.145 156.625 ;
        RECT 62.355 156.415 62.525 156.605 ;
        RECT 63.330 156.465 63.450 156.575 ;
        RECT 63.730 156.435 63.900 156.625 ;
        RECT 64.250 156.465 64.370 156.575 ;
        RECT 65.115 156.415 65.285 156.605 ;
        RECT 67.875 156.435 68.045 156.625 ;
        RECT 68.335 156.435 68.505 156.625 ;
        RECT 70.175 156.435 70.345 156.625 ;
        RECT 74.315 156.415 74.485 156.605 ;
        RECT 75.230 156.435 75.400 156.625 ;
        RECT 76.155 156.575 76.325 156.605 ;
        RECT 76.155 156.465 76.330 156.575 ;
        RECT 76.155 156.415 76.325 156.465 ;
        RECT 76.620 156.415 76.790 156.605 ;
        RECT 79.830 156.435 80.000 156.625 ;
        RECT 80.300 156.415 80.470 156.605 ;
        RECT 84.435 156.460 84.595 156.570 ;
        RECT 88.115 156.415 88.285 156.605 ;
        RECT 89.955 156.435 90.125 156.625 ;
        RECT 90.470 156.465 90.590 156.575 ;
        RECT 91.335 156.415 91.505 156.605 ;
        RECT 92.255 156.435 92.425 156.625 ;
        RECT 92.715 156.435 92.885 156.625 ;
        RECT 94.150 156.465 94.270 156.575 ;
        RECT 95.935 156.435 96.105 156.625 ;
        RECT 96.395 156.435 96.565 156.625 ;
        RECT 96.855 156.415 97.025 156.605 ;
        RECT 99.155 156.435 99.325 156.625 ;
        RECT 99.615 156.435 99.785 156.625 ;
        RECT 100.530 156.415 100.700 156.605 ;
        RECT 101.050 156.465 101.170 156.575 ;
        RECT 101.970 156.465 102.090 156.575 ;
        RECT 102.835 156.415 103.005 156.605 ;
        RECT 103.300 156.415 103.470 156.605 ;
        RECT 103.755 156.435 103.925 156.625 ;
        RECT 105.135 156.435 105.305 156.625 ;
        RECT 105.595 156.435 105.765 156.625 ;
        RECT 107.435 156.470 107.595 156.580 ;
        RECT 107.900 156.435 108.070 156.625 ;
        RECT 110.190 156.415 110.360 156.605 ;
        RECT 112.035 156.470 112.195 156.580 ;
        RECT 113.875 156.415 114.045 156.605 ;
        RECT 115.715 156.415 115.885 156.625 ;
        RECT 116.175 156.605 116.345 156.625 ;
        RECT 116.175 156.435 116.350 156.605 ;
        RECT 116.180 156.415 116.350 156.435 ;
        RECT 120.315 156.415 120.485 156.605 ;
        RECT 125.835 156.415 126.005 156.625 ;
        RECT 127.215 156.415 127.385 156.625 ;
        RECT 14.375 155.605 15.745 156.415 ;
        RECT 17.045 155.735 26.325 156.415 ;
        RECT 17.045 155.615 19.380 155.735 ;
        RECT 17.045 155.505 17.965 155.615 ;
        RECT 24.045 155.515 24.965 155.735 ;
        RECT 26.335 155.635 27.705 156.415 ;
        RECT 27.715 155.605 29.085 156.415 ;
        RECT 29.095 155.605 32.765 156.415 ;
        RECT 33.005 155.735 36.905 156.415 ;
        RECT 35.975 155.505 36.905 155.735 ;
        RECT 36.925 155.545 37.355 156.330 ;
        RECT 37.835 155.605 39.665 156.415 ;
        RECT 39.675 155.505 43.150 156.415 ;
        RECT 43.355 155.505 46.830 156.415 ;
        RECT 47.035 155.505 50.510 156.415 ;
        RECT 51.175 155.605 53.005 156.415 ;
        RECT 53.385 155.735 62.665 156.415 ;
        RECT 53.385 155.615 55.720 155.735 ;
        RECT 53.385 155.505 54.305 155.615 ;
        RECT 60.385 155.515 61.305 155.735 ;
        RECT 62.685 155.545 63.115 156.330 ;
        RECT 63.595 155.605 65.425 156.415 ;
        RECT 65.520 155.735 74.625 156.415 ;
        RECT 74.635 155.605 76.465 156.415 ;
        RECT 76.475 155.505 79.950 156.415 ;
        RECT 80.155 155.505 83.630 156.415 ;
        RECT 84.755 155.605 88.425 156.415 ;
        RECT 88.445 155.545 88.875 156.330 ;
        RECT 88.895 155.605 91.645 156.415 ;
        RECT 91.655 155.605 97.165 156.415 ;
        RECT 97.370 155.505 100.845 156.415 ;
        RECT 101.315 155.605 103.145 156.415 ;
        RECT 103.155 155.505 106.630 156.415 ;
        RECT 107.030 155.505 110.505 156.415 ;
        RECT 110.515 155.605 114.185 156.415 ;
        RECT 114.205 155.545 114.635 156.330 ;
        RECT 114.655 155.605 116.025 156.415 ;
        RECT 116.035 155.505 118.645 156.415 ;
        RECT 118.795 155.605 120.625 156.415 ;
        RECT 120.635 155.605 126.145 156.415 ;
        RECT 126.155 155.605 127.525 156.415 ;
      LAYER nwell ;
        RECT 14.180 152.385 127.720 155.215 ;
      LAYER pwell ;
        RECT 14.375 151.185 15.745 151.995 ;
        RECT 16.215 151.185 19.885 151.995 ;
        RECT 23.095 151.865 24.025 152.095 ;
        RECT 20.125 151.185 24.025 151.865 ;
        RECT 24.045 151.270 24.475 152.055 ;
        RECT 24.495 151.185 25.865 151.995 ;
        RECT 25.875 151.185 29.545 151.995 ;
        RECT 29.925 151.985 30.845 152.095 ;
        RECT 29.925 151.865 32.260 151.985 ;
        RECT 36.925 151.865 37.845 152.085 ;
        RECT 29.925 151.185 39.205 151.865 ;
        RECT 39.215 151.185 42.690 152.095 ;
        RECT 42.895 151.185 44.265 151.995 ;
        RECT 44.275 151.185 49.785 151.995 ;
        RECT 49.805 151.270 50.235 152.055 ;
        RECT 51.175 151.185 56.685 151.995 ;
        RECT 56.705 151.185 58.055 152.095 ;
        RECT 58.445 151.985 59.365 152.095 ;
        RECT 58.445 151.865 60.780 151.985 ;
        RECT 65.445 151.865 66.365 152.085 ;
        RECT 58.445 151.185 67.725 151.865 ;
        RECT 68.195 151.185 70.945 151.995 ;
        RECT 71.440 151.865 72.785 152.095 ;
        RECT 70.955 151.185 72.785 151.865 ;
        RECT 72.795 151.185 75.515 152.095 ;
        RECT 75.565 151.270 75.995 152.055 ;
        RECT 76.935 151.185 80.605 151.995 ;
        RECT 80.615 151.185 86.125 151.995 ;
        RECT 86.505 151.985 87.425 152.095 ;
        RECT 86.505 151.865 88.840 151.985 ;
        RECT 93.505 151.865 94.425 152.085 ;
        RECT 86.505 151.185 95.785 151.865 ;
        RECT 95.795 151.185 101.305 151.995 ;
        RECT 101.325 151.270 101.755 152.055 ;
        RECT 102.235 151.895 103.180 152.095 ;
        RECT 102.235 151.215 104.985 151.895 ;
        RECT 102.235 151.185 103.180 151.215 ;
        RECT 14.515 150.975 14.685 151.185 ;
        RECT 15.950 151.025 16.070 151.135 ;
        RECT 19.575 150.995 19.745 151.185 ;
        RECT 23.440 150.995 23.610 151.185 ;
        RECT 25.555 150.975 25.725 151.185 ;
        RECT 26.935 150.975 27.105 151.165 ;
        RECT 29.235 150.995 29.405 151.185 ;
        RECT 32.455 150.975 32.625 151.165 ;
        RECT 32.915 150.975 33.085 151.165 ;
        RECT 35.215 150.975 35.385 151.165 ;
        RECT 35.675 150.975 35.845 151.165 ;
        RECT 38.895 150.995 39.065 151.185 ;
        RECT 39.360 150.995 39.530 151.185 ;
        RECT 40.735 150.975 40.905 151.165 ;
        RECT 41.200 150.975 41.370 151.165 ;
        RECT 43.955 150.995 44.125 151.185 ;
        RECT 48.095 150.975 48.265 151.165 ;
        RECT 14.375 150.165 15.745 150.975 ;
        RECT 16.585 150.295 25.865 150.975 ;
        RECT 16.585 150.175 18.920 150.295 ;
        RECT 16.585 150.065 17.505 150.175 ;
        RECT 23.585 150.075 24.505 150.295 ;
        RECT 25.875 150.165 27.245 150.975 ;
        RECT 27.255 150.165 32.765 150.975 ;
        RECT 32.785 150.065 34.135 150.975 ;
        RECT 34.155 150.165 35.525 150.975 ;
        RECT 35.535 150.195 36.905 150.975 ;
        RECT 36.925 150.105 37.355 150.890 ;
        RECT 37.375 150.165 41.045 150.975 ;
        RECT 41.055 150.065 44.530 150.975 ;
        RECT 44.735 150.165 48.405 150.975 ;
        RECT 48.560 150.945 48.730 151.165 ;
        RECT 49.475 150.995 49.645 151.185 ;
        RECT 50.855 151.030 51.015 151.140 ;
        RECT 51.320 150.975 51.490 151.165 ;
        RECT 56.375 150.975 56.545 151.185 ;
        RECT 56.835 150.995 57.005 151.185 ;
        RECT 60.240 150.975 60.410 151.165 ;
        RECT 61.030 151.025 61.150 151.135 ;
        RECT 62.355 150.975 62.525 151.165 ;
        RECT 63.330 151.025 63.450 151.135 ;
        RECT 63.735 150.975 63.905 151.165 ;
        RECT 65.170 151.025 65.290 151.135 ;
        RECT 66.955 150.975 67.125 151.165 ;
        RECT 67.415 150.975 67.585 151.185 ;
        RECT 67.930 151.025 68.050 151.135 ;
        RECT 70.635 150.975 70.805 151.185 ;
        RECT 71.095 150.995 71.265 151.185 ;
        RECT 72.935 150.995 73.105 151.185 ;
        RECT 73.395 150.975 73.565 151.165 ;
        RECT 74.315 151.020 74.475 151.130 ;
        RECT 74.775 150.975 74.945 151.165 ;
        RECT 76.615 151.030 76.775 151.140 ;
        RECT 50.220 150.945 51.165 150.975 ;
        RECT 48.415 150.265 51.165 150.945 ;
        RECT 50.220 150.065 51.165 150.265 ;
        RECT 51.175 150.065 54.650 150.975 ;
        RECT 54.855 150.165 56.685 150.975 ;
        RECT 56.925 150.295 60.825 150.975 ;
        RECT 59.895 150.065 60.825 150.295 ;
        RECT 61.295 150.195 62.665 150.975 ;
        RECT 62.685 150.105 63.115 150.890 ;
        RECT 63.595 150.195 64.965 150.975 ;
        RECT 65.435 150.165 67.265 150.975 ;
        RECT 67.275 150.295 69.105 150.975 ;
        RECT 67.760 150.065 69.105 150.295 ;
        RECT 69.115 150.295 70.945 150.975 ;
        RECT 70.965 150.295 73.705 150.975 ;
        RECT 74.635 150.295 77.375 150.975 ;
        RECT 77.395 150.945 78.340 150.975 ;
        RECT 79.830 150.945 80.000 151.165 ;
        RECT 80.295 151.135 80.465 151.185 ;
        RECT 80.295 151.025 80.470 151.135 ;
        RECT 80.295 150.995 80.465 151.025 ;
        RECT 83.975 150.975 84.145 151.165 ;
        RECT 85.815 150.995 85.985 151.185 ;
        RECT 87.840 150.975 88.010 151.165 ;
        RECT 89.090 151.025 89.210 151.135 ;
        RECT 90.415 150.975 90.585 151.165 ;
        RECT 91.335 151.020 91.495 151.130 ;
        RECT 91.795 150.975 91.965 151.165 ;
        RECT 94.095 150.975 94.265 151.165 ;
        RECT 95.475 150.995 95.645 151.185 ;
        RECT 95.935 150.975 96.105 151.165 ;
        RECT 100.995 150.995 101.165 151.185 ;
        RECT 101.970 151.025 102.090 151.135 ;
        RECT 104.670 150.995 104.840 151.215 ;
        RECT 104.995 151.185 108.470 152.095 ;
        RECT 108.675 151.185 112.150 152.095 ;
        RECT 112.815 151.185 118.325 151.995 ;
        RECT 118.345 151.185 119.695 152.095 ;
        RECT 120.175 151.185 121.545 151.965 ;
        RECT 122.475 151.185 126.145 151.995 ;
        RECT 126.155 151.185 127.525 151.995 ;
        RECT 105.140 151.165 105.310 151.185 ;
        RECT 105.135 150.995 105.310 151.165 ;
        RECT 105.135 150.975 105.305 150.995 ;
        RECT 106.515 150.975 106.685 151.165 ;
        RECT 106.980 150.975 107.150 151.165 ;
        RECT 108.820 150.995 108.990 151.185 ;
        RECT 110.655 150.975 110.825 151.165 ;
        RECT 112.550 151.025 112.670 151.135 ;
        RECT 115.255 151.020 115.415 151.130 ;
        RECT 118.015 150.995 118.185 151.185 ;
        RECT 119.395 150.995 119.565 151.185 ;
        RECT 119.910 151.025 120.030 151.135 ;
        RECT 120.315 150.995 120.485 151.185 ;
        RECT 122.155 151.030 122.315 151.140 ;
        RECT 124.455 150.975 124.625 151.165 ;
        RECT 125.835 150.975 126.005 151.185 ;
        RECT 127.215 150.975 127.385 151.185 ;
        RECT 69.115 150.065 70.460 150.295 ;
        RECT 77.395 150.265 80.145 150.945 ;
        RECT 77.395 150.065 78.340 150.265 ;
        RECT 80.615 150.165 84.285 150.975 ;
        RECT 84.525 150.295 88.425 150.975 ;
        RECT 87.495 150.065 88.425 150.295 ;
        RECT 88.445 150.105 88.875 150.890 ;
        RECT 89.365 150.065 90.715 150.975 ;
        RECT 91.655 150.195 93.025 150.975 ;
        RECT 93.045 150.065 94.395 150.975 ;
        RECT 94.415 150.165 96.245 150.975 ;
        RECT 96.255 150.295 105.445 150.975 ;
        RECT 96.255 150.065 97.175 150.295 ;
        RECT 100.005 150.075 100.935 150.295 ;
        RECT 105.455 150.165 106.825 150.975 ;
        RECT 106.835 150.065 110.310 150.975 ;
        RECT 110.625 150.295 114.090 150.975 ;
        RECT 113.170 150.065 114.090 150.295 ;
        RECT 114.205 150.105 114.635 150.890 ;
        RECT 115.575 150.295 124.765 150.975 ;
        RECT 115.575 150.065 116.495 150.295 ;
        RECT 119.325 150.075 120.255 150.295 ;
        RECT 124.775 150.165 126.145 150.975 ;
        RECT 126.155 150.165 127.525 150.975 ;
      LAYER nwell ;
        RECT 14.180 146.945 127.720 149.775 ;
      LAYER pwell ;
        RECT 14.375 145.745 15.745 146.555 ;
        RECT 16.215 145.745 19.885 146.555 ;
        RECT 23.095 146.425 24.025 146.655 ;
        RECT 20.125 145.745 24.025 146.425 ;
        RECT 24.045 145.830 24.475 146.615 ;
        RECT 24.495 145.745 25.865 146.525 ;
        RECT 25.875 145.745 27.705 146.555 ;
        RECT 27.715 145.745 29.085 146.525 ;
        RECT 29.095 146.425 30.025 146.655 ;
        RECT 29.095 145.745 32.995 146.425 ;
        RECT 33.695 145.745 35.525 146.555 ;
        RECT 35.730 145.745 39.205 146.655 ;
        RECT 39.215 145.745 42.690 146.655 ;
        RECT 43.355 145.745 47.025 146.555 ;
        RECT 48.840 146.455 49.785 146.655 ;
        RECT 47.035 145.775 49.785 146.455 ;
        RECT 49.805 145.830 50.235 146.615 ;
        RECT 14.515 145.535 14.685 145.745 ;
        RECT 15.950 145.585 16.070 145.695 ;
        RECT 19.115 145.535 19.285 145.725 ;
        RECT 19.575 145.535 19.745 145.745 ;
        RECT 20.955 145.535 21.125 145.725 ;
        RECT 23.440 145.555 23.610 145.745 ;
        RECT 25.555 145.555 25.725 145.745 ;
        RECT 27.395 145.555 27.565 145.745 ;
        RECT 27.855 145.555 28.025 145.745 ;
        RECT 29.510 145.555 29.680 145.745 ;
        RECT 31.535 145.535 31.705 145.725 ;
        RECT 32.915 145.535 33.085 145.725 ;
        RECT 33.430 145.585 33.550 145.695 ;
        RECT 35.215 145.555 35.385 145.745 ;
        RECT 36.595 145.535 36.765 145.725 ;
        RECT 37.570 145.585 37.690 145.695 ;
        RECT 38.890 145.555 39.060 145.745 ;
        RECT 39.360 145.555 39.530 145.745 ;
        RECT 40.275 145.535 40.445 145.725 ;
        RECT 40.735 145.535 40.905 145.725 ;
        RECT 43.090 145.585 43.210 145.695 ;
        RECT 46.715 145.555 46.885 145.745 ;
        RECT 47.180 145.555 47.350 145.775 ;
        RECT 48.840 145.745 49.785 145.775 ;
        RECT 50.715 145.745 52.085 146.525 ;
        RECT 53.015 145.745 56.490 146.655 ;
        RECT 56.695 145.745 59.445 146.555 ;
        RECT 62.655 146.425 63.585 146.655 ;
        RECT 59.685 145.745 63.585 146.425 ;
        RECT 63.595 145.745 64.965 146.555 ;
        RECT 64.975 145.745 70.485 146.555 ;
        RECT 70.495 146.425 71.840 146.655 ;
        RECT 72.820 146.425 74.165 146.655 ;
        RECT 70.495 145.745 72.325 146.425 ;
        RECT 72.335 145.745 74.165 146.425 ;
        RECT 74.175 145.745 75.545 146.555 ;
        RECT 75.565 145.830 75.995 146.615 ;
        RECT 76.210 145.745 79.685 146.655 ;
        RECT 79.695 145.745 83.170 146.655 ;
        RECT 83.375 145.745 84.745 146.555 ;
        RECT 85.125 146.545 86.045 146.655 ;
        RECT 85.125 146.425 87.460 146.545 ;
        RECT 92.125 146.425 93.045 146.645 ;
        RECT 85.125 145.745 94.405 146.425 ;
        RECT 94.885 145.745 96.235 146.655 ;
        RECT 99.455 146.425 100.385 146.655 ;
        RECT 96.485 145.745 100.385 146.425 ;
        RECT 101.325 145.830 101.755 146.615 ;
        RECT 101.775 145.745 103.145 146.525 ;
        RECT 103.615 146.455 104.560 146.655 ;
        RECT 103.615 145.775 106.365 146.455 ;
        RECT 103.615 145.745 104.560 145.775 ;
        RECT 50.450 145.585 50.570 145.695 ;
        RECT 51.315 145.535 51.485 145.725 ;
        RECT 51.775 145.555 51.945 145.745 ;
        RECT 52.050 145.535 52.220 145.725 ;
        RECT 52.695 145.590 52.855 145.700 ;
        RECT 53.160 145.555 53.330 145.745 ;
        RECT 55.970 145.585 56.090 145.695 ;
        RECT 57.755 145.535 57.925 145.725 ;
        RECT 58.215 145.535 58.385 145.725 ;
        RECT 59.135 145.555 59.305 145.745 ;
        RECT 59.650 145.585 59.770 145.695 ;
        RECT 62.355 145.535 62.525 145.725 ;
        RECT 63.000 145.555 63.170 145.745 ;
        RECT 63.330 145.585 63.450 145.695 ;
        RECT 64.655 145.555 64.825 145.745 ;
        RECT 67.140 145.535 67.310 145.725 ;
        RECT 67.930 145.585 68.050 145.695 ;
        RECT 70.175 145.555 70.345 145.745 ;
        RECT 72.015 145.555 72.185 145.745 ;
        RECT 72.475 145.555 72.645 145.745 ;
        RECT 73.395 145.535 73.565 145.725 ;
        RECT 75.235 145.555 75.405 145.745 ;
        RECT 79.370 145.725 79.540 145.745 ;
        RECT 78.915 145.535 79.085 145.725 ;
        RECT 79.370 145.555 79.550 145.725 ;
        RECT 79.840 145.555 80.010 145.745 ;
        RECT 82.190 145.585 82.310 145.695 ;
        RECT 14.375 144.725 15.745 145.535 ;
        RECT 15.755 144.725 19.425 145.535 ;
        RECT 19.445 144.625 20.795 145.535 ;
        RECT 20.825 144.625 22.175 145.535 ;
        RECT 22.565 144.855 31.845 145.535 ;
        RECT 22.565 144.735 24.900 144.855 ;
        RECT 22.565 144.625 23.485 144.735 ;
        RECT 29.565 144.635 30.485 144.855 ;
        RECT 31.855 144.725 33.225 145.535 ;
        RECT 33.235 144.725 36.905 145.535 ;
        RECT 36.925 144.665 37.355 145.450 ;
        RECT 37.835 144.725 40.585 145.535 ;
        RECT 40.605 144.625 41.955 145.535 ;
        RECT 42.345 144.855 51.625 145.535 ;
        RECT 51.635 144.855 55.535 145.535 ;
        RECT 42.345 144.735 44.680 144.855 ;
        RECT 42.345 144.625 43.265 144.735 ;
        RECT 49.345 144.635 50.265 144.855 ;
        RECT 51.635 144.625 52.565 144.855 ;
        RECT 56.235 144.725 58.065 145.535 ;
        RECT 58.085 144.625 59.435 145.535 ;
        RECT 59.915 144.725 62.665 145.535 ;
        RECT 62.685 144.665 63.115 145.450 ;
        RECT 63.825 144.855 67.725 145.535 ;
        RECT 66.795 144.625 67.725 144.855 ;
        RECT 68.195 144.725 73.705 145.535 ;
        RECT 73.715 144.725 79.225 145.535 ;
        RECT 79.380 145.505 79.550 145.555 ;
        RECT 83.975 145.535 84.145 145.725 ;
        RECT 84.435 145.555 84.605 145.745 ;
        RECT 87.840 145.535 88.010 145.725 ;
        RECT 89.495 145.580 89.655 145.690 ;
        RECT 89.955 145.535 90.125 145.725 ;
        RECT 91.390 145.585 91.510 145.695 ;
        RECT 93.175 145.535 93.345 145.725 ;
        RECT 93.635 145.535 93.805 145.725 ;
        RECT 94.095 145.555 94.265 145.745 ;
        RECT 94.610 145.585 94.730 145.695 ;
        RECT 95.015 145.555 95.185 145.745 ;
        RECT 97.370 145.585 97.490 145.695 ;
        RECT 99.800 145.555 99.970 145.745 ;
        RECT 100.995 145.535 101.165 145.725 ;
        RECT 101.915 145.555 102.085 145.745 ;
        RECT 103.350 145.585 103.470 145.695 ;
        RECT 106.050 145.555 106.220 145.775 ;
        RECT 106.375 145.745 109.850 146.655 ;
        RECT 110.055 145.745 111.885 146.555 ;
        RECT 115.095 146.425 116.025 146.655 ;
        RECT 112.125 145.745 116.025 146.425 ;
        RECT 116.405 146.545 117.325 146.655 ;
        RECT 116.405 146.425 118.740 146.545 ;
        RECT 123.405 146.425 124.325 146.645 ;
        RECT 116.405 145.745 125.685 146.425 ;
        RECT 126.155 145.745 127.525 146.555 ;
        RECT 106.520 145.725 106.690 145.745 ;
        RECT 106.515 145.555 106.690 145.725 ;
        RECT 106.515 145.535 106.685 145.555 ;
        RECT 81.040 145.505 81.985 145.535 ;
        RECT 79.235 144.825 81.985 145.505 ;
        RECT 81.040 144.625 81.985 144.825 ;
        RECT 82.455 144.725 84.285 145.535 ;
        RECT 84.525 144.855 88.425 145.535 ;
        RECT 87.495 144.625 88.425 144.855 ;
        RECT 88.445 144.665 88.875 145.450 ;
        RECT 89.815 144.755 91.185 145.535 ;
        RECT 91.655 144.725 93.485 145.535 ;
        RECT 93.605 144.855 97.070 145.535 ;
        RECT 96.150 144.625 97.070 144.855 ;
        RECT 97.635 144.725 101.305 145.535 ;
        RECT 101.315 144.725 106.825 145.535 ;
        RECT 106.980 145.505 107.150 145.725 ;
        RECT 109.740 145.535 109.910 145.725 ;
        RECT 111.575 145.555 111.745 145.745 ;
        RECT 113.875 145.580 114.035 145.690 ;
        RECT 114.850 145.585 114.970 145.695 ;
        RECT 115.440 145.555 115.610 145.745 ;
        RECT 118.660 145.535 118.830 145.725 ;
        RECT 119.395 145.535 119.565 145.725 ;
        RECT 120.830 145.585 120.950 145.695 ;
        RECT 121.235 145.535 121.405 145.725 ;
        RECT 125.375 145.555 125.545 145.745 ;
        RECT 125.835 145.695 126.005 145.725 ;
        RECT 125.835 145.585 126.010 145.695 ;
        RECT 125.835 145.535 126.005 145.585 ;
        RECT 127.215 145.535 127.385 145.745 ;
        RECT 108.640 145.505 109.585 145.535 ;
        RECT 106.835 144.825 109.585 145.505 ;
        RECT 108.640 144.625 109.585 144.825 ;
        RECT 109.595 144.625 113.070 145.535 ;
        RECT 114.205 144.665 114.635 145.450 ;
        RECT 115.345 144.855 119.245 145.535 ;
        RECT 118.315 144.625 119.245 144.855 ;
        RECT 119.265 144.625 120.615 145.535 ;
        RECT 121.095 144.755 122.465 145.535 ;
        RECT 122.475 144.725 126.145 145.535 ;
        RECT 126.155 144.725 127.525 145.535 ;
      LAYER nwell ;
        RECT 14.180 141.505 127.720 144.335 ;
      LAYER pwell ;
        RECT 14.375 140.305 15.745 141.115 ;
        RECT 15.755 140.305 18.505 141.115 ;
        RECT 18.515 140.305 24.025 141.115 ;
        RECT 24.045 140.390 24.475 141.175 ;
        RECT 24.955 140.305 28.625 141.115 ;
        RECT 28.635 140.305 34.145 141.115 ;
        RECT 34.155 141.015 35.100 141.215 ;
        RECT 34.155 140.335 36.905 141.015 ;
        RECT 34.155 140.305 35.100 140.335 ;
        RECT 14.515 140.095 14.685 140.305 ;
        RECT 18.195 140.115 18.365 140.305 ;
        RECT 23.715 140.115 23.885 140.305 ;
        RECT 24.690 140.145 24.810 140.255 ;
        RECT 25.095 140.095 25.265 140.285 ;
        RECT 27.855 140.095 28.025 140.285 ;
        RECT 28.315 140.115 28.485 140.305 ;
        RECT 33.375 140.095 33.545 140.285 ;
        RECT 33.835 140.115 34.005 140.305 ;
        RECT 36.590 140.115 36.760 140.335 ;
        RECT 37.835 140.305 41.505 141.115 ;
        RECT 41.515 140.305 47.025 141.115 ;
        RECT 47.035 141.015 47.980 141.215 ;
        RECT 47.035 140.335 49.785 141.015 ;
        RECT 49.805 140.390 50.235 141.175 ;
        RECT 47.035 140.305 47.980 140.335 ;
        RECT 37.515 140.150 37.675 140.260 ;
        RECT 37.975 140.140 38.135 140.250 ;
        RECT 33.855 140.095 34.005 140.115 ;
        RECT 14.375 139.285 15.745 140.095 ;
        RECT 16.125 139.415 25.405 140.095 ;
        RECT 16.125 139.295 18.460 139.415 ;
        RECT 16.125 139.185 17.045 139.295 ;
        RECT 23.125 139.195 24.045 139.415 ;
        RECT 25.415 139.285 28.165 140.095 ;
        RECT 28.175 139.285 33.685 140.095 ;
        RECT 33.855 139.275 35.785 140.095 ;
        RECT 38.295 140.065 39.240 140.095 ;
        RECT 40.730 140.065 40.900 140.285 ;
        RECT 41.195 140.255 41.365 140.305 ;
        RECT 41.195 140.145 41.370 140.255 ;
        RECT 41.195 140.115 41.365 140.145 ;
        RECT 43.955 140.095 44.125 140.285 ;
        RECT 46.715 140.115 46.885 140.305 ;
        RECT 49.470 140.285 49.640 140.335 ;
        RECT 50.255 140.305 52.085 141.115 ;
        RECT 52.095 140.305 55.570 141.215 ;
        RECT 58.430 140.985 59.350 141.215 ;
        RECT 55.885 140.305 59.350 140.985 ;
        RECT 59.455 140.985 60.375 141.215 ;
        RECT 63.205 140.985 64.135 141.205 ;
        RECT 59.455 140.305 68.645 140.985 ;
        RECT 68.655 140.305 70.025 141.085 ;
        RECT 70.035 140.305 71.405 141.115 ;
        RECT 71.425 140.305 72.775 141.215 ;
        RECT 72.795 140.305 75.545 141.115 ;
        RECT 75.565 140.390 75.995 141.175 ;
        RECT 76.475 140.305 79.225 141.115 ;
        RECT 79.235 140.305 84.745 141.115 ;
        RECT 84.755 140.305 90.265 141.115 ;
        RECT 90.275 140.305 95.785 141.115 ;
        RECT 95.795 140.305 101.305 141.115 ;
        RECT 101.325 140.390 101.755 141.175 ;
        RECT 101.775 140.305 104.525 141.115 ;
        RECT 104.535 140.305 110.045 141.115 ;
        RECT 110.055 140.305 115.565 141.115 ;
        RECT 118.775 140.985 119.705 141.215 ;
        RECT 115.805 140.305 119.705 140.985 ;
        RECT 119.725 140.305 121.075 141.215 ;
        RECT 121.095 140.305 122.465 141.115 ;
        RECT 122.475 140.305 126.145 141.115 ;
        RECT 126.155 140.305 127.525 141.115 ;
        RECT 49.470 140.115 49.645 140.285 ;
        RECT 51.775 140.115 51.945 140.305 ;
        RECT 52.240 140.115 52.410 140.305 ;
        RECT 49.475 140.095 49.645 140.115 ;
        RECT 54.995 140.095 55.165 140.285 ;
        RECT 55.455 140.095 55.625 140.285 ;
        RECT 55.915 140.115 56.085 140.305 ;
        RECT 56.890 140.145 57.010 140.255 ;
        RECT 58.675 140.095 58.845 140.285 ;
        RECT 59.140 140.095 59.310 140.285 ;
        RECT 63.330 140.145 63.450 140.255 ;
        RECT 63.740 140.095 63.910 140.285 ;
        RECT 68.335 140.115 68.505 140.305 ;
        RECT 69.715 140.115 69.885 140.305 ;
        RECT 71.095 140.115 71.265 140.305 ;
        RECT 72.475 140.115 72.645 140.305 ;
        RECT 75.235 140.115 75.405 140.305 ;
        RECT 76.210 140.145 76.330 140.255 ;
        RECT 76.615 140.095 76.785 140.285 ;
        RECT 77.130 140.145 77.250 140.255 ;
        RECT 78.915 140.095 79.085 140.305 ;
        RECT 79.380 140.095 79.550 140.285 ;
        RECT 83.975 140.095 84.145 140.285 ;
        RECT 84.435 140.115 84.605 140.305 ;
        RECT 87.840 140.095 88.010 140.285 ;
        RECT 89.035 140.095 89.205 140.285 ;
        RECT 89.955 140.115 90.125 140.305 ;
        RECT 91.795 140.095 91.965 140.285 ;
        RECT 95.475 140.115 95.645 140.305 ;
        RECT 97.315 140.095 97.485 140.285 ;
        RECT 100.995 140.115 101.165 140.305 ;
        RECT 104.215 140.115 104.385 140.305 ;
        RECT 106.975 140.095 107.145 140.285 ;
        RECT 107.490 140.145 107.610 140.255 ;
        RECT 109.275 140.095 109.445 140.285 ;
        RECT 109.735 140.115 109.905 140.305 ;
        RECT 112.950 140.095 113.120 140.285 ;
        RECT 113.875 140.140 114.035 140.250 ;
        RECT 114.850 140.145 114.970 140.255 ;
        RECT 115.255 140.095 115.425 140.305 ;
        RECT 119.120 140.115 119.290 140.305 ;
        RECT 119.855 140.115 120.025 140.305 ;
        RECT 122.155 140.115 122.325 140.305 ;
        RECT 125.835 140.095 126.005 140.305 ;
        RECT 127.215 140.095 127.385 140.305 ;
        RECT 34.835 139.185 35.785 139.275 ;
        RECT 36.925 139.225 37.355 140.010 ;
        RECT 38.295 139.385 41.045 140.065 ;
        RECT 38.295 139.185 39.240 139.385 ;
        RECT 41.515 139.285 44.265 140.095 ;
        RECT 44.275 139.285 49.785 140.095 ;
        RECT 49.795 139.285 55.305 140.095 ;
        RECT 55.325 139.185 56.675 140.095 ;
        RECT 57.155 139.285 58.985 140.095 ;
        RECT 58.995 139.185 62.470 140.095 ;
        RECT 62.685 139.225 63.115 140.010 ;
        RECT 63.595 139.185 67.070 140.095 ;
        RECT 67.645 139.415 76.925 140.095 ;
        RECT 67.645 139.295 69.980 139.415 ;
        RECT 67.645 139.185 68.565 139.295 ;
        RECT 74.645 139.195 75.565 139.415 ;
        RECT 77.395 139.285 79.225 140.095 ;
        RECT 79.235 139.185 82.710 140.095 ;
        RECT 82.915 139.285 84.285 140.095 ;
        RECT 84.525 139.415 88.425 140.095 ;
        RECT 87.495 139.185 88.425 139.415 ;
        RECT 88.445 139.225 88.875 140.010 ;
        RECT 88.895 139.315 90.265 140.095 ;
        RECT 90.275 139.285 92.105 140.095 ;
        RECT 92.115 139.285 97.625 140.095 ;
        RECT 98.005 139.415 107.285 140.095 ;
        RECT 98.005 139.295 100.340 139.415 ;
        RECT 98.005 139.185 98.925 139.295 ;
        RECT 105.005 139.195 105.925 139.415 ;
        RECT 107.755 139.285 109.585 140.095 ;
        RECT 109.790 139.185 113.265 140.095 ;
        RECT 114.205 139.225 114.635 140.010 ;
        RECT 115.125 139.185 116.475 140.095 ;
        RECT 116.865 139.415 126.145 140.095 ;
        RECT 116.865 139.295 119.200 139.415 ;
        RECT 116.865 139.185 117.785 139.295 ;
        RECT 123.865 139.195 124.785 139.415 ;
        RECT 126.155 139.285 127.525 140.095 ;
      LAYER nwell ;
        RECT 14.180 136.065 127.720 138.895 ;
      LAYER pwell ;
        RECT 14.375 134.865 15.745 135.675 ;
        RECT 16.215 134.865 19.885 135.675 ;
        RECT 19.895 135.545 20.825 135.775 ;
        RECT 19.895 134.865 23.795 135.545 ;
        RECT 24.045 134.950 24.475 135.735 ;
        RECT 24.495 134.865 28.165 135.675 ;
        RECT 28.175 135.545 29.105 135.775 ;
        RECT 33.455 135.685 34.405 135.775 ;
        RECT 28.175 134.865 32.075 135.545 ;
        RECT 32.475 134.865 34.405 135.685 ;
        RECT 34.615 135.575 35.560 135.775 ;
        RECT 37.375 135.575 38.320 135.775 ;
        RECT 34.615 134.895 37.365 135.575 ;
        RECT 37.375 134.895 40.125 135.575 ;
        RECT 34.615 134.865 35.560 134.895 ;
        RECT 14.515 134.655 14.685 134.865 ;
        RECT 15.950 134.705 16.070 134.815 ;
        RECT 17.275 134.655 17.445 134.845 ;
        RECT 17.735 134.655 17.905 134.845 ;
        RECT 19.115 134.655 19.285 134.845 ;
        RECT 19.575 134.675 19.745 134.865 ;
        RECT 20.310 134.675 20.480 134.865 ;
        RECT 27.855 134.675 28.025 134.865 ;
        RECT 28.590 134.675 28.760 134.865 ;
        RECT 32.475 134.845 32.625 134.865 ;
        RECT 29.695 134.655 29.865 134.845 ;
        RECT 30.210 134.705 30.330 134.815 ;
        RECT 30.615 134.675 30.785 134.845 ;
        RECT 32.455 134.675 32.625 134.845 ;
        RECT 30.635 134.655 30.785 134.675 ;
        RECT 36.320 134.655 36.490 134.845 ;
        RECT 37.050 134.675 37.220 134.895 ;
        RECT 37.375 134.865 38.320 134.895 ;
        RECT 38.895 134.655 39.065 134.845 ;
        RECT 14.375 133.845 15.745 134.655 ;
        RECT 16.225 133.745 17.575 134.655 ;
        RECT 17.595 133.875 18.965 134.655 ;
        RECT 18.985 133.745 20.335 134.655 ;
        RECT 20.725 133.975 30.005 134.655 ;
        RECT 20.725 133.855 23.060 133.975 ;
        RECT 20.725 133.745 21.645 133.855 ;
        RECT 27.725 133.755 28.645 133.975 ;
        RECT 30.635 133.835 32.565 134.655 ;
        RECT 33.005 133.975 36.905 134.655 ;
        RECT 31.615 133.745 32.565 133.835 ;
        RECT 35.975 133.745 36.905 133.975 ;
        RECT 36.925 133.785 37.355 134.570 ;
        RECT 37.375 133.845 39.205 134.655 ;
        RECT 39.360 134.625 39.530 134.845 ;
        RECT 39.810 134.675 39.980 134.895 ;
        RECT 40.595 134.865 43.345 135.675 ;
        RECT 43.355 135.575 44.300 135.775 ;
        RECT 43.355 134.895 46.105 135.575 ;
        RECT 43.355 134.865 44.300 134.895 ;
        RECT 40.330 134.705 40.450 134.815 ;
        RECT 41.020 134.625 41.965 134.655 ;
        RECT 42.120 134.625 42.290 134.845 ;
        RECT 43.035 134.675 43.205 134.865 ;
        RECT 44.880 134.655 45.050 134.845 ;
        RECT 45.790 134.675 45.960 134.895 ;
        RECT 46.115 134.865 49.590 135.775 ;
        RECT 49.805 134.950 50.235 135.735 ;
        RECT 50.255 134.865 53.005 135.675 ;
        RECT 56.215 135.545 57.145 135.775 ;
        RECT 53.245 134.865 57.145 135.545 ;
        RECT 57.615 134.865 58.985 135.645 ;
        RECT 58.995 134.865 60.825 135.675 ;
        RECT 60.835 134.865 64.310 135.775 ;
        RECT 67.170 135.545 68.090 135.775 ;
        RECT 64.625 134.865 68.090 135.545 ;
        RECT 68.195 134.865 71.405 135.775 ;
        RECT 71.875 134.865 75.545 135.675 ;
        RECT 75.565 134.950 75.995 135.735 ;
        RECT 76.935 135.575 77.880 135.775 ;
        RECT 76.935 134.895 79.685 135.575 ;
        RECT 76.935 134.865 77.880 134.895 ;
        RECT 46.260 134.675 46.430 134.865 ;
        RECT 48.560 134.655 48.730 134.845 ;
        RECT 52.695 134.675 52.865 134.865 ;
        RECT 56.560 134.675 56.730 134.865 ;
        RECT 57.350 134.705 57.470 134.815 ;
        RECT 57.755 134.675 57.925 134.865 ;
        RECT 60.515 134.675 60.685 134.865 ;
        RECT 60.980 134.675 61.150 134.865 ;
        RECT 61.435 134.655 61.605 134.845 ;
        RECT 62.355 134.700 62.515 134.810 ;
        RECT 63.280 134.655 63.450 134.845 ;
        RECT 64.655 134.675 64.825 134.865 ;
        RECT 67.415 134.700 67.575 134.810 ;
        RECT 68.335 134.675 68.505 134.865 ;
        RECT 71.610 134.705 71.730 134.815 ;
        RECT 72.935 134.655 73.105 134.845 ;
        RECT 75.235 134.675 75.405 134.865 ;
        RECT 76.615 134.710 76.775 134.820 ;
        RECT 78.455 134.655 78.625 134.845 ;
        RECT 43.780 134.625 44.725 134.655 ;
        RECT 39.215 133.945 41.965 134.625 ;
        RECT 41.975 133.945 44.725 134.625 ;
        RECT 41.020 133.745 41.965 133.945 ;
        RECT 43.780 133.745 44.725 133.945 ;
        RECT 44.735 133.745 48.210 134.655 ;
        RECT 48.415 133.745 51.890 134.655 ;
        RECT 52.465 133.975 61.745 134.655 ;
        RECT 52.465 133.855 54.800 133.975 ;
        RECT 52.465 133.745 53.385 133.855 ;
        RECT 59.465 133.755 60.385 133.975 ;
        RECT 62.685 133.785 63.115 134.570 ;
        RECT 63.135 133.745 66.610 134.655 ;
        RECT 67.735 133.845 73.245 134.655 ;
        RECT 73.255 133.845 78.765 134.655 ;
        RECT 78.920 134.625 79.090 134.845 ;
        RECT 79.370 134.675 79.540 134.895 ;
        RECT 79.695 134.865 83.170 135.775 ;
        RECT 83.745 135.665 84.665 135.775 ;
        RECT 83.745 135.545 86.080 135.665 ;
        RECT 90.745 135.545 91.665 135.765 ;
        RECT 93.035 135.545 93.965 135.775 ;
        RECT 83.745 134.865 93.025 135.545 ;
        RECT 93.035 134.865 96.935 135.545 ;
        RECT 97.830 134.865 101.305 135.775 ;
        RECT 101.325 134.950 101.755 135.735 ;
        RECT 105.895 135.545 106.825 135.775 ;
        RECT 102.925 134.865 106.825 135.545 ;
        RECT 106.835 134.865 108.205 135.645 ;
        RECT 112.335 135.545 113.265 135.775 ;
        RECT 109.365 134.865 113.265 135.545 ;
        RECT 113.645 135.665 114.565 135.775 ;
        RECT 113.645 135.545 115.980 135.665 ;
        RECT 120.645 135.545 121.565 135.765 ;
        RECT 113.645 134.865 122.925 135.545 ;
        RECT 122.935 134.865 124.305 135.645 ;
        RECT 124.315 134.865 126.145 135.675 ;
        RECT 126.155 134.865 127.525 135.675 ;
        RECT 79.840 134.675 80.010 134.865 ;
        RECT 86.735 134.655 86.905 134.845 ;
        RECT 88.115 134.655 88.285 134.845 ;
        RECT 92.715 134.675 92.885 134.865 ;
        RECT 93.450 134.675 93.620 134.865 ;
        RECT 97.370 134.705 97.490 134.815 ;
        RECT 98.235 134.655 98.405 134.845 ;
        RECT 80.580 134.625 81.525 134.655 ;
        RECT 78.775 133.945 81.525 134.625 ;
        RECT 80.580 133.745 81.525 133.945 ;
        RECT 81.535 133.845 87.045 134.655 ;
        RECT 87.065 133.745 88.415 134.655 ;
        RECT 88.445 133.785 88.875 134.570 ;
        RECT 89.265 133.975 98.545 134.655 ;
        RECT 98.555 134.625 99.500 134.655 ;
        RECT 100.990 134.625 101.160 134.865 ;
        RECT 102.375 134.655 102.545 134.845 ;
        RECT 102.890 134.705 103.010 134.815 ;
        RECT 89.265 133.855 91.600 133.975 ;
        RECT 89.265 133.745 90.185 133.855 ;
        RECT 96.265 133.755 97.185 133.975 ;
        RECT 98.555 133.945 101.305 134.625 ;
        RECT 98.555 133.745 99.500 133.945 ;
        RECT 101.325 133.745 102.675 134.655 ;
        RECT 103.155 134.625 104.100 134.655 ;
        RECT 105.590 134.625 105.760 134.845 ;
        RECT 106.060 134.655 106.230 134.845 ;
        RECT 106.240 134.675 106.410 134.865 ;
        RECT 107.895 134.675 108.065 134.865 ;
        RECT 108.815 134.710 108.975 134.820 ;
        RECT 103.155 133.945 105.905 134.625 ;
        RECT 103.155 133.745 104.100 133.945 ;
        RECT 105.915 133.745 109.390 134.655 ;
        RECT 109.595 134.625 110.540 134.655 ;
        RECT 112.030 134.625 112.200 134.845 ;
        RECT 112.680 134.675 112.850 134.865 ;
        RECT 113.875 134.655 114.045 134.845 ;
        RECT 114.850 134.705 114.970 134.815 ;
        RECT 118.475 134.655 118.645 134.845 ;
        RECT 118.935 134.655 119.105 134.845 ;
        RECT 120.370 134.705 120.490 134.815 ;
        RECT 122.615 134.675 122.785 134.865 ;
        RECT 123.075 134.675 123.245 134.865 ;
        RECT 125.835 134.655 126.005 134.865 ;
        RECT 127.215 134.655 127.385 134.865 ;
        RECT 109.595 133.945 112.345 134.625 ;
        RECT 109.595 133.745 110.540 133.945 ;
        RECT 112.355 133.845 114.185 134.655 ;
        RECT 114.205 133.785 114.635 134.570 ;
        RECT 115.115 133.845 118.785 134.655 ;
        RECT 118.795 133.875 120.165 134.655 ;
        RECT 120.635 133.845 126.145 134.655 ;
        RECT 126.155 133.845 127.525 134.655 ;
      LAYER nwell ;
        RECT 14.180 130.625 127.720 133.455 ;
      LAYER pwell ;
        RECT 14.375 129.425 15.745 130.235 ;
        RECT 16.215 129.425 19.885 130.235 ;
        RECT 23.095 130.105 24.025 130.335 ;
        RECT 20.125 129.425 24.025 130.105 ;
        RECT 24.045 129.510 24.475 130.295 ;
        RECT 24.955 129.425 28.625 130.235 ;
        RECT 30.385 130.225 31.305 130.335 ;
        RECT 28.635 129.425 30.005 130.205 ;
        RECT 30.385 130.105 32.720 130.225 ;
        RECT 37.385 130.105 38.305 130.325 ;
        RECT 30.385 129.425 39.665 130.105 ;
        RECT 39.760 129.425 48.865 130.105 ;
        RECT 49.805 129.510 50.235 130.295 ;
        RECT 50.715 129.425 54.385 130.235 ;
        RECT 54.395 129.425 59.905 130.235 ;
        RECT 59.915 129.425 65.425 130.235 ;
        RECT 68.635 130.105 69.565 130.335 ;
        RECT 71.615 130.245 72.565 130.335 ;
        RECT 65.665 129.425 69.565 130.105 ;
        RECT 69.575 129.425 71.405 130.105 ;
        RECT 71.615 129.425 73.545 130.245 ;
        RECT 73.715 129.425 75.545 130.105 ;
        RECT 75.565 129.510 75.995 130.295 ;
        RECT 78.515 130.245 79.465 130.335 ;
        RECT 76.475 129.425 78.305 130.235 ;
        RECT 78.515 129.425 80.445 130.245 ;
        RECT 80.615 129.425 83.365 130.235 ;
        RECT 83.375 129.425 88.885 130.235 ;
        RECT 88.905 129.425 90.255 130.335 ;
        RECT 90.295 129.425 101.305 130.335 ;
        RECT 101.325 129.510 101.755 130.295 ;
        RECT 109.795 130.245 110.745 130.335 ;
        RECT 102.235 129.425 104.065 130.235 ;
        RECT 104.075 129.425 109.585 130.235 ;
        RECT 109.795 129.425 111.725 130.245 ;
        RECT 112.355 129.425 115.105 130.235 ;
        RECT 115.115 129.425 120.625 130.235 ;
        RECT 120.635 129.425 126.145 130.235 ;
        RECT 126.155 129.425 127.525 130.235 ;
        RECT 14.515 129.215 14.685 129.425 ;
        RECT 15.950 129.265 16.070 129.375 ;
        RECT 16.815 129.215 16.985 129.405 ;
        RECT 19.575 129.235 19.745 129.425 ;
        RECT 23.440 129.235 23.610 129.425 ;
        RECT 24.690 129.265 24.810 129.375 ;
        RECT 26.475 129.215 26.645 129.405 ;
        RECT 27.395 129.260 27.555 129.370 ;
        RECT 28.315 129.235 28.485 129.425 ;
        RECT 29.695 129.235 29.865 129.425 ;
        RECT 32.915 129.215 33.085 129.405 ;
        RECT 33.375 129.215 33.545 129.405 ;
        RECT 34.810 129.265 34.930 129.375 ;
        RECT 36.595 129.215 36.765 129.405 ;
        RECT 37.975 129.260 38.135 129.370 ;
        RECT 39.355 129.215 39.525 129.425 ;
        RECT 39.815 129.235 39.985 129.405 ;
        RECT 42.115 129.235 42.285 129.405 ;
        RECT 39.835 129.215 39.985 129.235 ;
        RECT 42.135 129.215 42.285 129.235 ;
        RECT 46.715 129.215 46.885 129.405 ;
        RECT 47.175 129.235 47.345 129.405 ;
        RECT 48.555 129.235 48.725 129.425 ;
        RECT 49.475 129.270 49.635 129.380 ;
        RECT 50.395 129.375 50.565 129.405 ;
        RECT 50.395 129.265 50.570 129.375 ;
        RECT 47.195 129.215 47.345 129.235 ;
        RECT 50.395 129.215 50.565 129.265 ;
        RECT 54.075 129.215 54.245 129.425 ;
        RECT 57.940 129.215 58.110 129.405 ;
        RECT 58.730 129.265 58.850 129.375 ;
        RECT 59.595 129.235 59.765 129.425 ;
        RECT 62.355 129.215 62.525 129.405 ;
        RECT 64.195 129.215 64.365 129.405 ;
        RECT 65.115 129.235 65.285 129.425 ;
        RECT 68.980 129.235 69.150 129.425 ;
        RECT 71.095 129.235 71.265 129.425 ;
        RECT 73.395 129.405 73.545 129.425 ;
        RECT 73.395 129.235 73.565 129.405 ;
        RECT 73.855 129.215 74.025 129.425 ;
        RECT 74.315 129.235 74.485 129.405 ;
        RECT 76.210 129.265 76.330 129.375 ;
        RECT 76.615 129.235 76.785 129.405 ;
        RECT 77.995 129.235 78.165 129.425 ;
        RECT 80.295 129.405 80.445 129.425 ;
        RECT 80.295 129.235 80.465 129.405 ;
        RECT 74.335 129.215 74.485 129.235 ;
        RECT 76.635 129.215 76.785 129.235 ;
        RECT 82.320 129.215 82.490 129.405 ;
        RECT 83.055 129.235 83.225 129.425 ;
        RECT 84.895 129.235 85.065 129.405 ;
        RECT 84.895 129.215 85.045 129.235 ;
        RECT 86.735 129.215 86.905 129.405 ;
        RECT 87.195 129.215 87.365 129.405 ;
        RECT 88.575 129.235 88.745 129.425 ;
        RECT 89.035 129.375 89.205 129.425 ;
        RECT 89.035 129.265 89.210 129.375 ;
        RECT 89.035 129.235 89.205 129.265 ;
        RECT 89.770 129.215 89.940 129.405 ;
        RECT 93.690 129.265 93.810 129.375 ;
        RECT 94.095 129.215 94.265 129.405 ;
        RECT 95.475 129.215 95.645 129.405 ;
        RECT 100.990 129.235 101.160 129.425 ;
        RECT 101.970 129.265 102.090 129.375 ;
        RECT 103.755 129.235 103.925 129.425 ;
        RECT 106.515 129.235 106.685 129.405 ;
        RECT 108.815 129.235 108.985 129.405 ;
        RECT 109.275 129.235 109.445 129.425 ;
        RECT 111.575 129.405 111.725 129.425 ;
        RECT 111.575 129.235 111.745 129.405 ;
        RECT 112.090 129.265 112.210 129.375 ;
        RECT 113.415 129.235 113.585 129.405 ;
        RECT 114.795 129.375 114.965 129.425 ;
        RECT 113.930 129.265 114.050 129.375 ;
        RECT 114.795 129.265 114.970 129.375 ;
        RECT 114.795 129.235 114.965 129.265 ;
        RECT 106.515 129.215 106.665 129.235 ;
        RECT 108.815 129.215 108.965 129.235 ;
        RECT 14.375 128.405 15.745 129.215 ;
        RECT 15.755 128.405 17.125 129.215 ;
        RECT 17.505 128.535 26.785 129.215 ;
        RECT 17.505 128.415 19.840 128.535 ;
        RECT 17.505 128.305 18.425 128.415 ;
        RECT 24.505 128.315 25.425 128.535 ;
        RECT 27.715 128.405 33.225 129.215 ;
        RECT 33.245 128.305 34.595 129.215 ;
        RECT 35.075 128.405 36.905 129.215 ;
        RECT 36.925 128.345 37.355 129.130 ;
        RECT 38.295 128.435 39.665 129.215 ;
        RECT 39.835 128.395 41.765 129.215 ;
        RECT 42.135 128.395 44.065 129.215 ;
        RECT 44.935 128.405 47.025 129.215 ;
        RECT 47.195 128.395 49.125 129.215 ;
        RECT 49.335 128.405 50.705 129.215 ;
        RECT 50.715 128.405 54.385 129.215 ;
        RECT 54.625 128.535 58.525 129.215 ;
        RECT 40.815 128.305 41.765 128.395 ;
        RECT 43.115 128.305 44.065 128.395 ;
        RECT 48.175 128.305 49.125 128.395 ;
        RECT 57.595 128.305 58.525 128.535 ;
        RECT 58.995 128.405 62.665 129.215 ;
        RECT 62.685 128.345 63.115 129.130 ;
        RECT 63.135 128.405 64.505 129.215 ;
        RECT 64.885 128.535 74.165 129.215 ;
        RECT 64.885 128.415 67.220 128.535 ;
        RECT 64.885 128.305 65.805 128.415 ;
        RECT 71.885 128.315 72.805 128.535 ;
        RECT 74.335 128.395 76.265 129.215 ;
        RECT 76.635 128.395 78.565 129.215 ;
        RECT 79.005 128.535 82.905 129.215 ;
        RECT 75.315 128.305 76.265 128.395 ;
        RECT 77.615 128.305 78.565 128.395 ;
        RECT 81.975 128.305 82.905 128.535 ;
        RECT 83.115 128.395 85.045 129.215 ;
        RECT 85.215 128.405 87.045 129.215 ;
        RECT 87.055 128.435 88.425 129.215 ;
        RECT 83.115 128.305 84.065 128.395 ;
        RECT 88.445 128.345 88.875 129.130 ;
        RECT 89.355 128.535 93.255 129.215 ;
        RECT 89.355 128.305 90.285 128.535 ;
        RECT 93.955 128.435 95.325 129.215 ;
        RECT 95.335 128.535 104.440 129.215 ;
        RECT 104.735 128.395 106.665 129.215 ;
        RECT 107.035 128.395 108.965 129.215 ;
        RECT 109.295 129.215 109.445 129.235 ;
        RECT 113.415 129.215 113.565 129.235 ;
        RECT 117.555 129.215 117.725 129.405 ;
        RECT 118.015 129.215 118.185 129.405 ;
        RECT 119.395 129.215 119.565 129.405 ;
        RECT 120.315 129.235 120.485 129.425 ;
        RECT 125.835 129.215 126.005 129.425 ;
        RECT 127.215 129.215 127.385 129.425 ;
        RECT 109.295 128.395 111.225 129.215 ;
        RECT 104.735 128.305 105.685 128.395 ;
        RECT 107.035 128.305 107.985 128.395 ;
        RECT 110.275 128.305 111.225 128.395 ;
        RECT 111.635 128.395 113.565 129.215 ;
        RECT 111.635 128.305 112.585 128.395 ;
        RECT 114.205 128.345 114.635 129.130 ;
        RECT 115.115 128.405 117.865 129.215 ;
        RECT 117.885 128.305 119.235 129.215 ;
        RECT 119.255 128.435 120.625 129.215 ;
        RECT 120.635 128.405 126.145 129.215 ;
        RECT 126.155 128.405 127.525 129.215 ;
      LAYER nwell ;
        RECT 14.180 125.185 127.720 128.015 ;
      LAYER pwell ;
        RECT 14.375 123.985 15.745 124.795 ;
        RECT 15.755 123.985 17.125 124.795 ;
        RECT 17.135 123.985 20.805 124.795 ;
        RECT 20.825 123.985 22.175 124.895 ;
        RECT 22.655 123.985 24.025 124.765 ;
        RECT 24.045 124.070 24.475 124.855 ;
        RECT 37.595 124.805 38.545 124.895 ;
        RECT 25.415 123.985 30.925 124.795 ;
        RECT 30.935 123.985 36.445 124.795 ;
        RECT 36.615 123.985 38.545 124.805 ;
        RECT 40.335 124.805 41.285 124.895 ;
        RECT 43.575 124.805 44.525 124.895 ;
        RECT 38.755 123.985 40.125 124.795 ;
        RECT 40.335 123.985 42.265 124.805 ;
        RECT 14.515 123.775 14.685 123.985 ;
        RECT 16.815 123.775 16.985 123.985 ;
        RECT 20.495 123.795 20.665 123.985 ;
        RECT 21.875 123.795 22.045 123.985 ;
        RECT 22.335 123.935 22.505 123.965 ;
        RECT 22.335 123.825 22.510 123.935 ;
        RECT 22.335 123.775 22.505 123.825 ;
        RECT 22.795 123.795 22.965 123.985 ;
        RECT 25.095 123.830 25.255 123.940 ;
        RECT 26.200 123.775 26.370 123.965 ;
        RECT 26.990 123.825 27.110 123.935 ;
        RECT 30.615 123.795 30.785 123.985 ;
        RECT 32.455 123.775 32.625 123.965 ;
        RECT 36.135 123.795 36.305 123.985 ;
        RECT 36.615 123.965 36.765 123.985 ;
        RECT 36.320 123.775 36.490 123.965 ;
        RECT 36.595 123.795 36.765 123.965 ;
        RECT 37.570 123.825 37.690 123.935 ;
        RECT 39.815 123.795 39.985 123.985 ;
        RECT 42.115 123.965 42.265 123.985 ;
        RECT 42.595 123.985 44.525 124.805 ;
        RECT 44.935 124.805 45.885 124.895 ;
        RECT 44.935 123.985 46.865 124.805 ;
        RECT 47.045 123.985 49.785 124.665 ;
        RECT 49.805 124.070 50.235 124.855 ;
        RECT 50.255 123.985 52.085 124.795 ;
        RECT 52.095 123.985 57.605 124.795 ;
        RECT 57.615 123.985 58.985 124.765 ;
        RECT 62.195 124.665 63.125 124.895 ;
        RECT 59.225 123.985 63.125 124.665 ;
        RECT 63.135 123.985 64.505 124.795 ;
        RECT 64.515 123.985 68.185 124.795 ;
        RECT 68.205 123.985 69.555 124.895 ;
        RECT 70.035 123.985 71.405 124.765 ;
        RECT 72.335 123.985 75.075 124.665 ;
        RECT 75.565 124.070 75.995 124.855 ;
        RECT 76.015 123.985 77.845 124.795 ;
        RECT 78.225 124.785 79.145 124.895 ;
        RECT 78.225 124.665 80.560 124.785 ;
        RECT 85.225 124.665 86.145 124.885 ;
        RECT 78.225 123.985 87.505 124.665 ;
        RECT 87.515 123.985 89.345 124.795 ;
        RECT 90.715 124.665 91.635 124.885 ;
        RECT 97.715 124.785 98.635 124.895 ;
        RECT 100.155 124.805 101.105 124.895 ;
        RECT 96.300 124.665 98.635 124.785 ;
        RECT 89.355 123.985 98.635 124.665 ;
        RECT 99.175 123.985 101.105 124.805 ;
        RECT 101.325 124.070 101.755 124.855 ;
        RECT 101.775 123.985 105.445 124.795 ;
        RECT 105.455 123.985 110.965 124.795 ;
        RECT 114.175 124.665 115.105 124.895 ;
        RECT 111.205 123.985 115.105 124.665 ;
        RECT 115.485 124.785 116.405 124.895 ;
        RECT 115.485 124.665 117.820 124.785 ;
        RECT 122.485 124.665 123.405 124.885 ;
        RECT 115.485 123.985 124.765 124.665 ;
        RECT 124.775 123.985 126.145 124.795 ;
        RECT 126.155 123.985 127.525 124.795 ;
        RECT 42.595 123.965 42.745 123.985 ;
        RECT 41.195 123.775 41.365 123.965 ;
        RECT 42.115 123.795 42.285 123.965 ;
        RECT 42.575 123.795 42.745 123.965 ;
        RECT 46.715 123.965 46.865 123.985 ;
        RECT 46.715 123.775 46.885 123.965 ;
        RECT 49.475 123.795 49.645 123.985 ;
        RECT 51.775 123.795 51.945 123.985 ;
        RECT 52.235 123.775 52.405 123.965 ;
        RECT 57.295 123.795 57.465 123.985 ;
        RECT 57.755 123.795 57.925 123.985 ;
        RECT 61.895 123.775 62.065 123.965 ;
        RECT 62.410 123.825 62.530 123.935 ;
        RECT 62.540 123.795 62.710 123.985 ;
        RECT 63.330 123.825 63.450 123.935 ;
        RECT 64.195 123.795 64.365 123.985 ;
        RECT 67.140 123.775 67.310 123.965 ;
        RECT 67.875 123.795 68.045 123.985 ;
        RECT 69.255 123.795 69.425 123.985 ;
        RECT 69.770 123.825 69.890 123.935 ;
        RECT 70.175 123.775 70.345 123.985 ;
        RECT 72.015 123.830 72.175 123.940 ;
        RECT 72.475 123.795 72.645 123.985 ;
        RECT 75.290 123.825 75.410 123.935 ;
        RECT 75.695 123.775 75.865 123.965 ;
        RECT 77.535 123.795 77.705 123.985 ;
        RECT 81.215 123.775 81.385 123.965 ;
        RECT 82.595 123.775 82.765 123.965 ;
        RECT 83.110 123.825 83.230 123.935 ;
        RECT 83.515 123.775 83.685 123.965 ;
        RECT 87.195 123.795 87.365 123.985 ;
        RECT 88.115 123.775 88.285 123.965 ;
        RECT 89.035 123.795 89.205 123.985 ;
        RECT 89.495 123.795 89.665 123.985 ;
        RECT 99.175 123.965 99.325 123.985 ;
        RECT 92.255 123.775 92.425 123.965 ;
        RECT 92.715 123.775 92.885 123.965 ;
        RECT 95.015 123.775 95.185 123.965 ;
        RECT 98.695 123.775 98.865 123.965 ;
        RECT 99.155 123.795 99.325 123.965 ;
        RECT 104.215 123.775 104.385 123.965 ;
        RECT 105.135 123.795 105.305 123.985 ;
        RECT 109.735 123.775 109.905 123.965 ;
        RECT 110.655 123.795 110.825 123.985 ;
        RECT 113.600 123.775 113.770 123.965 ;
        RECT 114.520 123.795 114.690 123.985 ;
        RECT 114.850 123.825 114.970 123.935 ;
        RECT 124.455 123.775 124.625 123.985 ;
        RECT 125.835 123.775 126.005 123.985 ;
        RECT 127.215 123.775 127.385 123.985 ;
        RECT 14.375 122.965 15.745 123.775 ;
        RECT 15.755 122.965 17.125 123.775 ;
        RECT 17.135 122.965 22.645 123.775 ;
        RECT 22.885 123.095 26.785 123.775 ;
        RECT 25.855 122.865 26.785 123.095 ;
        RECT 27.255 122.965 32.765 123.775 ;
        RECT 33.005 123.095 36.905 123.775 ;
        RECT 35.975 122.865 36.905 123.095 ;
        RECT 36.925 122.905 37.355 123.690 ;
        RECT 37.835 122.965 41.505 123.775 ;
        RECT 41.515 122.965 47.025 123.775 ;
        RECT 47.035 122.965 52.545 123.775 ;
        RECT 52.925 123.095 62.205 123.775 ;
        RECT 52.925 122.975 55.260 123.095 ;
        RECT 52.925 122.865 53.845 122.975 ;
        RECT 59.925 122.875 60.845 123.095 ;
        RECT 62.685 122.905 63.115 123.690 ;
        RECT 63.825 123.095 67.725 123.775 ;
        RECT 66.795 122.865 67.725 123.095 ;
        RECT 67.735 122.965 70.485 123.775 ;
        RECT 70.495 122.965 76.005 123.775 ;
        RECT 76.015 122.965 81.525 123.775 ;
        RECT 81.545 122.865 82.895 123.775 ;
        RECT 83.375 122.995 84.745 123.775 ;
        RECT 84.755 122.965 88.425 123.775 ;
        RECT 88.445 122.905 88.875 123.690 ;
        RECT 88.895 122.965 92.565 123.775 ;
        RECT 92.585 122.865 93.935 123.775 ;
        RECT 93.955 122.965 95.325 123.775 ;
        RECT 95.335 122.965 99.005 123.775 ;
        RECT 99.015 122.965 104.525 123.775 ;
        RECT 104.535 122.965 110.045 123.775 ;
        RECT 110.285 123.095 114.185 123.775 ;
        RECT 113.255 122.865 114.185 123.095 ;
        RECT 114.205 122.905 114.635 123.690 ;
        RECT 115.485 123.095 124.765 123.775 ;
        RECT 115.485 122.975 117.820 123.095 ;
        RECT 115.485 122.865 116.405 122.975 ;
        RECT 122.485 122.875 123.405 123.095 ;
        RECT 124.775 122.965 126.145 123.775 ;
        RECT 126.155 122.965 127.525 123.775 ;
      LAYER nwell ;
        RECT 14.180 119.745 127.720 122.575 ;
      LAYER pwell ;
        RECT 14.375 118.545 15.745 119.355 ;
        RECT 16.215 118.545 19.885 119.355 ;
        RECT 19.895 119.225 20.825 119.455 ;
        RECT 19.895 118.545 23.795 119.225 ;
        RECT 24.045 118.630 24.475 119.415 ;
        RECT 24.495 118.545 25.865 119.355 ;
        RECT 25.875 118.545 27.245 119.325 ;
        RECT 27.255 118.545 30.005 119.355 ;
        RECT 30.385 119.345 31.305 119.455 ;
        RECT 30.385 119.225 32.720 119.345 ;
        RECT 37.385 119.225 38.305 119.445 ;
        RECT 39.675 119.225 40.605 119.455 ;
        RECT 30.385 118.545 39.665 119.225 ;
        RECT 39.675 118.545 43.575 119.225 ;
        RECT 44.275 118.545 45.645 119.325 ;
        RECT 48.855 119.225 49.785 119.455 ;
        RECT 45.885 118.545 49.785 119.225 ;
        RECT 49.805 118.630 50.235 119.415 ;
        RECT 50.265 118.545 51.615 119.455 ;
        RECT 51.635 118.545 53.005 119.355 ;
        RECT 53.155 118.545 55.765 119.455 ;
        RECT 56.705 118.545 58.055 119.455 ;
        RECT 59.365 119.345 60.285 119.455 ;
        RECT 59.365 119.225 61.700 119.345 ;
        RECT 66.365 119.225 67.285 119.445 ;
        RECT 59.365 118.545 68.645 119.225 ;
        RECT 68.655 118.545 70.025 119.325 ;
        RECT 70.495 118.545 74.165 119.355 ;
        RECT 74.185 118.545 75.535 119.455 ;
        RECT 75.565 118.630 75.995 119.415 ;
        RECT 79.675 119.225 80.605 119.455 ;
        RECT 76.705 118.545 80.605 119.225 ;
        RECT 80.615 118.545 81.985 119.325 ;
        RECT 82.005 118.545 83.355 119.455 ;
        RECT 83.835 118.545 85.205 119.325 ;
        RECT 85.215 118.545 90.725 119.355 ;
        RECT 90.735 119.225 91.665 119.455 ;
        RECT 90.735 118.545 94.635 119.225 ;
        RECT 95.335 118.545 97.165 119.355 ;
        RECT 100.375 119.225 101.305 119.455 ;
        RECT 97.405 118.545 101.305 119.225 ;
        RECT 101.325 118.630 101.755 119.415 ;
        RECT 101.775 118.545 103.145 119.355 ;
        RECT 103.165 118.545 104.515 119.455 ;
        RECT 107.735 119.225 108.665 119.455 ;
        RECT 104.765 118.545 108.665 119.225 ;
        RECT 109.045 119.345 109.965 119.455 ;
        RECT 109.045 119.225 111.380 119.345 ;
        RECT 116.045 119.225 116.965 119.445 ;
        RECT 109.045 118.545 118.325 119.225 ;
        RECT 118.345 118.545 119.695 119.455 ;
        RECT 120.175 118.545 121.545 119.325 ;
        RECT 122.475 118.545 126.145 119.355 ;
        RECT 126.155 118.545 127.525 119.355 ;
        RECT 14.515 118.335 14.685 118.545 ;
        RECT 15.950 118.385 16.070 118.495 ;
        RECT 17.275 118.335 17.445 118.525 ;
        RECT 19.575 118.355 19.745 118.545 ;
        RECT 20.310 118.355 20.480 118.545 ;
        RECT 25.555 118.355 25.725 118.545 ;
        RECT 26.935 118.335 27.105 118.545 ;
        RECT 27.395 118.335 27.565 118.525 ;
        RECT 29.695 118.355 29.865 118.545 ;
        RECT 39.355 118.355 39.525 118.545 ;
        RECT 40.090 118.355 40.260 118.545 ;
        RECT 44.010 118.385 44.130 118.495 ;
        RECT 45.335 118.355 45.505 118.545 ;
        RECT 46.715 118.335 46.885 118.525 ;
        RECT 49.200 118.355 49.370 118.545 ;
        RECT 50.395 118.355 50.565 118.545 ;
        RECT 52.695 118.355 52.865 118.545 ;
        RECT 55.450 118.355 55.620 118.545 ;
        RECT 56.375 118.335 56.545 118.525 ;
        RECT 57.295 118.380 57.455 118.490 ;
        RECT 57.755 118.355 57.925 118.545 ;
        RECT 58.675 118.390 58.835 118.500 ;
        RECT 60.975 118.335 61.145 118.525 ;
        RECT 61.435 118.335 61.605 118.525 ;
        RECT 68.335 118.355 68.505 118.545 ;
        RECT 69.715 118.355 69.885 118.545 ;
        RECT 70.230 118.385 70.350 118.495 ;
        RECT 72.475 118.335 72.645 118.525 ;
        RECT 73.855 118.355 74.025 118.545 ;
        RECT 74.315 118.355 74.485 118.545 ;
        RECT 76.210 118.385 76.330 118.495 ;
        RECT 80.020 118.355 80.190 118.545 ;
        RECT 81.675 118.355 81.845 118.545 ;
        RECT 82.135 118.335 82.305 118.525 ;
        RECT 82.870 118.335 83.040 118.525 ;
        RECT 83.055 118.355 83.225 118.545 ;
        RECT 83.570 118.385 83.690 118.495 ;
        RECT 83.975 118.355 84.145 118.545 ;
        RECT 86.790 118.385 86.910 118.495 ;
        RECT 87.195 118.335 87.365 118.525 ;
        RECT 89.035 118.335 89.205 118.525 ;
        RECT 90.415 118.335 90.585 118.545 ;
        RECT 91.150 118.355 91.320 118.545 ;
        RECT 92.255 118.380 92.415 118.490 ;
        RECT 95.070 118.385 95.190 118.495 ;
        RECT 96.855 118.355 97.025 118.545 ;
        RECT 100.720 118.355 100.890 118.545 ;
        RECT 101.915 118.335 102.085 118.525 ;
        RECT 102.835 118.355 103.005 118.545 ;
        RECT 103.295 118.355 103.465 118.545 ;
        RECT 108.080 118.355 108.250 118.545 ;
        RECT 111.575 118.335 111.745 118.525 ;
        RECT 112.495 118.380 112.655 118.490 ;
        RECT 113.875 118.335 114.045 118.525 ;
        RECT 114.850 118.385 114.970 118.495 ;
        RECT 115.255 118.335 115.425 118.525 ;
        RECT 116.690 118.385 116.810 118.495 ;
        RECT 118.015 118.355 118.185 118.545 ;
        RECT 118.475 118.355 118.645 118.545 ;
        RECT 119.910 118.385 120.030 118.495 ;
        RECT 120.315 118.335 120.485 118.545 ;
        RECT 122.155 118.390 122.315 118.500 ;
        RECT 125.835 118.335 126.005 118.545 ;
        RECT 127.215 118.335 127.385 118.545 ;
        RECT 14.375 117.525 15.745 118.335 ;
        RECT 16.225 117.425 17.575 118.335 ;
        RECT 17.965 117.655 27.245 118.335 ;
        RECT 27.255 117.655 36.535 118.335 ;
        RECT 17.965 117.535 20.300 117.655 ;
        RECT 17.965 117.425 18.885 117.535 ;
        RECT 24.965 117.435 25.885 117.655 ;
        RECT 28.615 117.435 29.535 117.655 ;
        RECT 34.200 117.535 36.535 117.655 ;
        RECT 35.615 117.425 36.535 117.535 ;
        RECT 36.925 117.465 37.355 118.250 ;
        RECT 37.745 117.655 47.025 118.335 ;
        RECT 47.405 117.655 56.685 118.335 ;
        RECT 37.745 117.535 40.080 117.655 ;
        RECT 37.745 117.425 38.665 117.535 ;
        RECT 44.745 117.435 45.665 117.655 ;
        RECT 47.405 117.535 49.740 117.655 ;
        RECT 47.405 117.425 48.325 117.535 ;
        RECT 54.405 117.435 55.325 117.655 ;
        RECT 57.615 117.525 61.285 118.335 ;
        RECT 61.305 117.425 62.655 118.335 ;
        RECT 62.685 117.465 63.115 118.250 ;
        RECT 63.505 117.655 72.785 118.335 ;
        RECT 73.165 117.655 82.445 118.335 ;
        RECT 82.455 117.655 86.355 118.335 ;
        RECT 63.505 117.535 65.840 117.655 ;
        RECT 63.505 117.425 64.425 117.535 ;
        RECT 70.505 117.435 71.425 117.655 ;
        RECT 73.165 117.535 75.500 117.655 ;
        RECT 73.165 117.425 74.085 117.535 ;
        RECT 80.165 117.435 81.085 117.655 ;
        RECT 82.455 117.425 83.385 117.655 ;
        RECT 87.055 117.555 88.425 118.335 ;
        RECT 88.445 117.465 88.875 118.250 ;
        RECT 88.905 117.425 90.255 118.335 ;
        RECT 90.285 117.425 91.635 118.335 ;
        RECT 92.945 117.655 102.225 118.335 ;
        RECT 102.605 117.655 111.885 118.335 ;
        RECT 92.945 117.535 95.280 117.655 ;
        RECT 92.945 117.425 93.865 117.535 ;
        RECT 99.945 117.435 100.865 117.655 ;
        RECT 102.605 117.535 104.940 117.655 ;
        RECT 102.605 117.425 103.525 117.535 ;
        RECT 109.605 117.435 110.525 117.655 ;
        RECT 112.825 117.425 114.175 118.335 ;
        RECT 114.205 117.465 114.635 118.250 ;
        RECT 115.115 117.555 116.485 118.335 ;
        RECT 116.955 117.525 120.625 118.335 ;
        RECT 120.635 117.525 126.145 118.335 ;
        RECT 126.155 117.525 127.525 118.335 ;
      LAYER nwell ;
        RECT 14.180 114.305 127.720 117.135 ;
      LAYER pwell ;
        RECT 14.375 113.105 15.745 113.915 ;
        RECT 15.755 113.105 17.125 113.915 ;
        RECT 17.135 113.105 20.805 113.915 ;
        RECT 20.815 113.105 22.185 113.885 ;
        RECT 22.205 113.105 23.555 114.015 ;
        RECT 24.045 113.190 24.475 113.975 ;
        RECT 25.855 113.785 26.775 114.005 ;
        RECT 32.855 113.905 33.775 114.015 ;
        RECT 31.440 113.785 33.775 113.905 ;
        RECT 24.495 113.105 33.775 113.785 ;
        RECT 34.625 113.105 35.975 114.015 ;
        RECT 36.455 113.105 37.825 113.885 ;
        RECT 38.755 113.105 40.125 113.885 ;
        RECT 40.135 113.105 43.805 113.915 ;
        RECT 43.825 113.105 45.175 114.015 ;
        RECT 45.195 113.785 46.125 114.015 ;
        RECT 45.195 113.105 49.095 113.785 ;
        RECT 49.805 113.190 50.235 113.975 ;
        RECT 50.255 113.105 52.085 113.915 ;
        RECT 52.095 113.105 53.465 113.885 ;
        RECT 53.475 113.105 54.845 113.915 ;
        RECT 54.855 113.105 60.365 113.915 ;
        RECT 60.375 113.105 65.885 113.915 ;
        RECT 65.905 113.105 67.255 114.015 ;
        RECT 67.735 113.105 69.105 113.885 ;
        RECT 70.035 113.105 75.545 113.915 ;
        RECT 75.565 113.190 75.995 113.975 ;
        RECT 77.305 113.905 78.225 114.015 ;
        RECT 77.305 113.785 79.640 113.905 ;
        RECT 84.305 113.785 85.225 114.005 ;
        RECT 88.415 113.785 89.335 114.005 ;
        RECT 95.415 113.905 96.335 114.015 ;
        RECT 94.000 113.785 96.335 113.905 ;
        RECT 77.305 113.105 86.585 113.785 ;
        RECT 87.055 113.105 96.335 113.785 ;
        RECT 97.175 113.105 99.925 113.915 ;
        RECT 99.935 113.105 101.305 113.885 ;
        RECT 101.325 113.190 101.755 113.975 ;
        RECT 102.235 113.105 107.745 113.915 ;
        RECT 107.755 113.105 109.125 113.885 ;
        RECT 109.135 113.105 110.965 113.915 ;
        RECT 114.175 113.785 115.105 114.015 ;
        RECT 111.205 113.105 115.105 113.785 ;
        RECT 115.115 113.105 120.625 113.915 ;
        RECT 120.635 113.105 126.145 113.915 ;
        RECT 126.155 113.105 127.525 113.915 ;
        RECT 14.515 112.895 14.685 113.105 ;
        RECT 16.815 112.915 16.985 113.105 ;
        RECT 20.495 112.915 20.665 113.105 ;
        RECT 20.955 112.915 21.125 113.105 ;
        RECT 23.255 112.915 23.425 113.105 ;
        RECT 23.770 112.945 23.890 113.055 ;
        RECT 24.635 112.915 24.805 113.105 ;
        RECT 26.015 112.895 26.185 113.085 ;
        RECT 27.855 112.895 28.025 113.085 ;
        RECT 33.375 112.895 33.545 113.085 ;
        RECT 34.350 112.945 34.470 113.055 ;
        RECT 34.755 112.895 34.925 113.085 ;
        RECT 35.675 112.915 35.845 113.105 ;
        RECT 36.190 112.945 36.310 113.055 ;
        RECT 36.595 112.895 36.765 113.105 ;
        RECT 37.570 112.945 37.690 113.055 ;
        RECT 38.435 112.950 38.595 113.060 ;
        RECT 39.815 112.915 39.985 113.105 ;
        RECT 43.495 112.915 43.665 113.105 ;
        RECT 44.875 112.915 45.045 113.105 ;
        RECT 45.610 112.915 45.780 113.105 ;
        RECT 46.715 112.895 46.885 113.085 ;
        RECT 47.635 112.940 47.795 113.050 ;
        RECT 49.530 112.945 49.650 113.055 ;
        RECT 51.315 112.895 51.485 113.085 ;
        RECT 51.775 112.915 51.945 113.105 ;
        RECT 52.235 112.915 52.405 113.105 ;
        RECT 54.535 112.915 54.705 113.105 ;
        RECT 56.835 112.895 57.005 113.085 ;
        RECT 60.055 112.915 60.225 113.105 ;
        RECT 62.355 112.895 62.525 113.085 ;
        RECT 63.330 112.945 63.450 113.055 ;
        RECT 65.575 112.915 65.745 113.105 ;
        RECT 66.035 112.915 66.205 113.105 ;
        RECT 67.470 112.945 67.590 113.055 ;
        RECT 67.875 112.915 68.045 113.105 ;
        RECT 68.795 112.895 68.965 113.085 ;
        RECT 69.715 112.950 69.875 113.060 ;
        RECT 74.315 112.895 74.485 113.085 ;
        RECT 75.235 112.915 75.405 113.105 ;
        RECT 76.615 112.950 76.775 113.060 ;
        RECT 79.835 112.895 80.005 113.085 ;
        RECT 81.215 112.895 81.385 113.085 ;
        RECT 82.595 112.895 82.765 113.085 ;
        RECT 86.275 112.915 86.445 113.105 ;
        RECT 86.790 112.945 86.910 113.055 ;
        RECT 87.195 112.915 87.365 113.105 ;
        RECT 88.115 112.895 88.285 113.085 ;
        RECT 92.255 112.895 92.425 113.085 ;
        RECT 92.715 112.895 92.885 113.085 ;
        RECT 96.910 112.945 97.030 113.055 ;
        RECT 99.615 112.915 99.785 113.105 ;
        RECT 100.995 112.915 101.165 113.105 ;
        RECT 101.970 112.945 102.090 113.055 ;
        RECT 102.835 112.915 103.005 113.085 ;
        RECT 107.435 112.915 107.605 113.105 ;
        RECT 107.895 112.915 108.065 113.105 ;
        RECT 108.355 112.895 108.525 113.085 ;
        RECT 110.655 112.915 110.825 113.105 ;
        RECT 113.875 112.895 114.045 113.085 ;
        RECT 114.520 112.915 114.690 113.105 ;
        RECT 115.255 112.940 115.415 113.050 ;
        RECT 118.935 112.895 119.105 113.085 ;
        RECT 119.395 112.895 119.565 113.085 ;
        RECT 120.315 112.915 120.485 113.105 ;
        RECT 121.695 112.895 121.865 113.085 ;
        RECT 123.075 112.895 123.245 113.085 ;
        RECT 125.835 112.895 126.005 113.105 ;
        RECT 127.215 112.895 127.385 113.105 ;
        RECT 14.375 112.085 15.745 112.895 ;
        RECT 15.955 112.215 26.325 112.895 ;
        RECT 15.955 111.985 18.165 112.215 ;
        RECT 20.885 111.995 21.815 112.215 ;
        RECT 26.335 112.085 28.165 112.895 ;
        RECT 28.175 112.085 33.685 112.895 ;
        RECT 33.705 111.985 35.055 112.895 ;
        RECT 35.075 112.085 36.905 112.895 ;
        RECT 36.925 112.025 37.355 112.810 ;
        RECT 37.920 112.215 47.025 112.895 ;
        RECT 47.955 112.085 51.625 112.895 ;
        RECT 51.635 112.085 57.145 112.895 ;
        RECT 57.155 112.085 62.665 112.895 ;
        RECT 62.685 112.025 63.115 112.810 ;
        RECT 63.595 112.085 69.105 112.895 ;
        RECT 69.115 112.085 74.625 112.895 ;
        RECT 74.635 112.085 80.145 112.895 ;
        RECT 80.165 111.985 81.515 112.895 ;
        RECT 81.535 112.085 82.905 112.895 ;
        RECT 82.915 112.085 88.425 112.895 ;
        RECT 88.445 112.025 88.875 112.810 ;
        RECT 88.895 112.085 92.565 112.895 ;
        RECT 92.575 112.215 101.680 112.895 ;
        RECT 101.775 112.215 102.730 112.895 ;
        RECT 103.155 112.085 108.665 112.895 ;
        RECT 108.675 112.085 114.185 112.895 ;
        RECT 114.205 112.025 114.635 112.810 ;
        RECT 115.575 112.085 119.245 112.895 ;
        RECT 119.265 111.985 120.615 112.895 ;
        RECT 120.635 112.115 122.005 112.895 ;
        RECT 122.015 112.115 123.385 112.895 ;
        RECT 123.395 112.085 126.145 112.895 ;
        RECT 126.155 112.085 127.525 112.895 ;
      LAYER nwell ;
        RECT 14.180 108.865 127.720 111.695 ;
      LAYER pwell ;
        RECT 14.375 107.665 15.745 108.475 ;
        RECT 16.675 107.665 20.345 108.475 ;
        RECT 20.365 107.665 21.715 108.575 ;
        RECT 22.665 107.665 24.015 108.575 ;
        RECT 24.045 107.750 24.475 108.535 ;
        RECT 24.495 107.665 27.245 108.475 ;
        RECT 27.255 107.665 28.625 108.445 ;
        RECT 28.635 107.665 30.465 108.475 ;
        RECT 30.485 107.665 31.835 108.575 ;
        RECT 31.855 107.665 33.225 108.445 ;
        RECT 34.155 107.665 35.525 108.445 ;
        RECT 35.995 107.665 38.745 108.475 ;
        RECT 38.755 107.665 44.265 108.475 ;
        RECT 44.275 107.665 49.785 108.475 ;
        RECT 49.805 107.750 50.235 108.535 ;
        RECT 50.715 107.665 52.085 108.445 ;
        RECT 53.015 107.665 56.685 108.475 ;
        RECT 56.695 107.665 58.065 108.445 ;
        RECT 58.075 107.665 59.445 108.475 ;
        RECT 59.455 107.665 62.065 108.575 ;
        RECT 62.675 107.665 64.505 108.475 ;
        RECT 64.525 107.665 65.875 108.575 ;
        RECT 66.355 107.665 68.185 108.475 ;
        RECT 68.195 107.665 69.565 108.445 ;
        RECT 70.035 107.665 75.545 108.475 ;
        RECT 75.565 107.750 75.995 108.535 ;
        RECT 76.025 107.665 77.375 108.575 ;
        RECT 77.405 107.665 78.755 108.575 ;
        RECT 79.695 107.665 82.305 108.575 ;
        RECT 82.455 107.665 83.825 108.445 ;
        RECT 84.295 107.665 87.045 108.475 ;
        RECT 87.065 107.665 88.415 108.575 ;
        RECT 88.435 107.665 92.105 108.475 ;
        RECT 92.125 107.665 93.475 108.575 ;
        RECT 93.495 107.665 94.865 108.445 ;
        RECT 94.875 107.665 96.245 108.475 ;
        RECT 96.255 107.665 99.925 108.475 ;
        RECT 99.935 107.665 101.305 108.445 ;
        RECT 101.325 107.750 101.755 108.535 ;
        RECT 102.235 107.665 105.905 108.475 ;
        RECT 105.915 107.665 107.285 108.445 ;
        RECT 107.295 107.665 108.665 108.475 ;
        RECT 108.685 107.665 110.035 108.575 ;
        RECT 110.055 107.665 111.425 108.445 ;
        RECT 111.435 107.665 112.805 108.445 ;
        RECT 112.815 107.665 114.185 108.475 ;
        RECT 114.205 107.665 115.555 108.575 ;
        RECT 120.085 108.345 121.015 108.565 ;
        RECT 123.735 108.345 125.945 108.575 ;
        RECT 115.575 107.665 125.945 108.345 ;
        RECT 126.155 107.665 127.525 108.475 ;
        RECT 14.515 107.455 14.685 107.665 ;
        RECT 16.355 107.510 16.515 107.620 ;
        RECT 20.035 107.475 20.205 107.665 ;
        RECT 21.415 107.475 21.585 107.665 ;
        RECT 22.335 107.510 22.495 107.620 ;
        RECT 23.715 107.475 23.885 107.665 ;
        RECT 26.015 107.455 26.185 107.645 ;
        RECT 26.935 107.475 27.105 107.665 ;
        RECT 28.315 107.475 28.485 107.665 ;
        RECT 30.155 107.475 30.325 107.665 ;
        RECT 31.535 107.475 31.705 107.665 ;
        RECT 32.915 107.475 33.085 107.665 ;
        RECT 33.835 107.510 33.995 107.620 ;
        RECT 35.215 107.475 35.385 107.665 ;
        RECT 35.730 107.505 35.850 107.615 ;
        RECT 36.595 107.455 36.765 107.645 ;
        RECT 38.435 107.455 38.605 107.665 ;
        RECT 38.950 107.505 39.070 107.615 ;
        RECT 40.275 107.455 40.445 107.645 ;
        RECT 41.655 107.455 41.825 107.645 ;
        RECT 43.035 107.455 43.205 107.645 ;
        RECT 43.550 107.505 43.670 107.615 ;
        RECT 43.955 107.475 44.125 107.665 ;
        RECT 44.875 107.455 45.045 107.645 ;
        RECT 45.335 107.455 45.505 107.645 ;
        RECT 49.475 107.475 49.645 107.665 ;
        RECT 50.450 107.505 50.570 107.615 ;
        RECT 50.855 107.475 51.025 107.665 ;
        RECT 52.695 107.510 52.855 107.620 ;
        RECT 56.375 107.475 56.545 107.665 ;
        RECT 56.835 107.455 57.005 107.665 ;
        RECT 58.215 107.455 58.385 107.645 ;
        RECT 59.135 107.475 59.305 107.665 ;
        RECT 59.600 107.645 59.770 107.665 ;
        RECT 59.595 107.475 59.770 107.645 ;
        RECT 59.595 107.455 59.765 107.475 ;
        RECT 60.055 107.455 60.225 107.645 ;
        RECT 61.435 107.455 61.605 107.645 ;
        RECT 62.410 107.505 62.530 107.615 ;
        RECT 64.195 107.475 64.365 107.665 ;
        RECT 64.655 107.475 64.825 107.665 ;
        RECT 66.090 107.505 66.210 107.615 ;
        RECT 67.875 107.475 68.045 107.665 ;
        RECT 68.335 107.475 68.505 107.665 ;
        RECT 69.770 107.505 69.890 107.615 ;
        RECT 73.395 107.455 73.565 107.645 ;
        RECT 74.315 107.500 74.475 107.610 ;
        RECT 74.775 107.455 74.945 107.645 ;
        RECT 75.235 107.475 75.405 107.665 ;
        RECT 77.075 107.475 77.245 107.665 ;
        RECT 78.455 107.475 78.625 107.665 ;
        RECT 79.375 107.510 79.535 107.620 ;
        RECT 79.840 107.475 80.010 107.665 ;
        RECT 82.595 107.475 82.765 107.665 ;
        RECT 84.030 107.505 84.150 107.615 ;
        RECT 86.275 107.455 86.445 107.645 ;
        RECT 86.735 107.615 86.905 107.665 ;
        RECT 86.735 107.505 86.910 107.615 ;
        RECT 86.735 107.475 86.905 107.505 ;
        RECT 87.195 107.455 87.365 107.665 ;
        RECT 91.795 107.475 91.965 107.665 ;
        RECT 92.255 107.475 92.425 107.665 ;
        RECT 93.635 107.475 93.805 107.665 ;
        RECT 95.935 107.475 96.105 107.665 ;
        RECT 99.155 107.455 99.325 107.645 ;
        RECT 99.615 107.475 99.785 107.665 ;
        RECT 100.535 107.455 100.705 107.645 ;
        RECT 100.995 107.475 101.165 107.665 ;
        RECT 101.915 107.615 102.085 107.645 ;
        RECT 101.915 107.505 102.090 107.615 ;
        RECT 101.915 107.455 102.085 107.505 ;
        RECT 102.375 107.455 102.545 107.645 ;
        RECT 105.595 107.475 105.765 107.665 ;
        RECT 106.055 107.475 106.225 107.665 ;
        RECT 108.355 107.475 108.525 107.665 ;
        RECT 109.735 107.475 109.905 107.665 ;
        RECT 110.195 107.475 110.365 107.665 ;
        RECT 111.575 107.475 111.745 107.665 ;
        RECT 113.875 107.455 114.045 107.665 ;
        RECT 114.335 107.475 114.505 107.665 ;
        RECT 115.255 107.500 115.415 107.610 ;
        RECT 115.715 107.455 115.885 107.665 ;
        RECT 127.215 107.455 127.385 107.665 ;
        RECT 14.375 106.645 15.745 107.455 ;
        RECT 15.955 106.775 26.325 107.455 ;
        RECT 26.535 106.775 36.905 107.455 ;
        RECT 15.955 106.545 18.165 106.775 ;
        RECT 20.885 106.555 21.815 106.775 ;
        RECT 26.535 106.545 28.745 106.775 ;
        RECT 31.465 106.555 32.395 106.775 ;
        RECT 36.925 106.585 37.355 107.370 ;
        RECT 37.375 106.675 38.745 107.455 ;
        RECT 39.225 106.545 40.575 107.455 ;
        RECT 40.595 106.645 41.965 107.455 ;
        RECT 41.975 106.675 43.345 107.455 ;
        RECT 43.825 106.545 45.175 107.455 ;
        RECT 45.195 106.675 46.565 107.455 ;
        RECT 46.775 106.775 57.145 107.455 ;
        RECT 46.775 106.545 48.985 106.775 ;
        RECT 51.705 106.555 52.635 106.775 ;
        RECT 57.165 106.545 58.515 107.455 ;
        RECT 58.535 106.645 59.905 107.455 ;
        RECT 59.925 106.545 61.275 107.455 ;
        RECT 61.295 106.675 62.665 107.455 ;
        RECT 62.685 106.585 63.115 107.370 ;
        RECT 63.335 106.775 73.705 107.455 ;
        RECT 63.335 106.545 65.545 106.775 ;
        RECT 68.265 106.555 69.195 106.775 ;
        RECT 74.635 106.675 76.005 107.455 ;
        RECT 76.215 106.775 86.585 107.455 ;
        RECT 76.215 106.545 78.425 106.775 ;
        RECT 81.145 106.555 82.075 106.775 ;
        RECT 87.055 106.675 88.425 107.455 ;
        RECT 88.445 106.585 88.875 107.370 ;
        RECT 89.095 106.775 99.465 107.455 ;
        RECT 89.095 106.545 91.305 106.775 ;
        RECT 94.025 106.555 94.955 106.775 ;
        RECT 99.485 106.545 100.835 107.455 ;
        RECT 100.855 106.645 102.225 107.455 ;
        RECT 102.245 106.545 103.595 107.455 ;
        RECT 103.815 106.775 114.185 107.455 ;
        RECT 103.815 106.545 106.025 106.775 ;
        RECT 108.745 106.555 109.675 106.775 ;
        RECT 114.205 106.585 114.635 107.370 ;
        RECT 115.575 106.775 125.945 107.455 ;
        RECT 120.085 106.555 121.015 106.775 ;
        RECT 123.735 106.545 125.945 106.775 ;
        RECT 126.155 106.645 127.525 107.455 ;
      LAYER nwell ;
        RECT 14.180 103.425 127.720 106.255 ;
      LAYER pwell ;
        RECT 14.375 102.225 15.745 103.035 ;
        RECT 15.755 102.225 18.505 103.035 ;
        RECT 18.515 102.225 24.025 103.035 ;
        RECT 24.045 102.310 24.475 103.095 ;
        RECT 24.495 102.225 27.245 103.035 ;
        RECT 27.265 102.225 28.615 103.135 ;
        RECT 33.145 102.905 34.075 103.125 ;
        RECT 36.795 102.905 39.005 103.135 ;
        RECT 28.635 102.225 39.005 102.905 ;
        RECT 39.415 102.905 41.625 103.135 ;
        RECT 44.345 102.905 45.275 103.125 ;
        RECT 39.415 102.225 49.785 102.905 ;
        RECT 49.805 102.310 50.235 103.095 ;
        RECT 51.185 102.225 52.535 103.135 ;
        RECT 52.755 102.905 54.965 103.135 ;
        RECT 57.685 102.905 58.615 103.125 ;
        RECT 63.335 102.905 65.545 103.135 ;
        RECT 68.265 102.905 69.195 103.125 ;
        RECT 52.755 102.225 63.125 102.905 ;
        RECT 63.335 102.225 73.705 102.905 ;
        RECT 73.715 102.225 75.545 103.035 ;
        RECT 75.565 102.310 75.995 103.095 ;
        RECT 76.215 102.905 78.425 103.135 ;
        RECT 81.145 102.905 82.075 103.125 ;
        RECT 86.795 102.905 89.005 103.135 ;
        RECT 91.725 102.905 92.655 103.125 ;
        RECT 76.215 102.225 86.585 102.905 ;
        RECT 86.795 102.225 97.165 102.905 ;
        RECT 97.635 102.225 101.305 103.035 ;
        RECT 101.325 102.310 101.755 103.095 ;
        RECT 101.975 102.905 104.185 103.135 ;
        RECT 106.905 102.905 107.835 103.125 ;
        RECT 116.865 102.905 117.795 103.125 ;
        RECT 120.515 102.905 122.725 103.135 ;
        RECT 101.975 102.225 112.345 102.905 ;
        RECT 112.355 102.225 122.725 102.905 ;
        RECT 122.935 102.225 124.765 103.035 ;
        RECT 124.775 102.225 126.145 103.005 ;
        RECT 126.155 102.225 127.525 103.035 ;
        RECT 14.515 102.015 14.685 102.225 ;
        RECT 18.195 102.015 18.365 102.225 ;
        RECT 23.715 102.015 23.885 102.225 ;
        RECT 26.935 102.035 27.105 102.225 ;
        RECT 27.395 102.035 27.565 102.225 ;
        RECT 28.775 102.035 28.945 102.225 ;
        RECT 34.755 102.015 34.925 102.205 ;
        RECT 36.595 102.015 36.765 102.205 ;
        RECT 38.435 102.015 38.605 102.205 ;
        RECT 43.955 102.015 44.125 102.205 ;
        RECT 49.475 102.015 49.645 102.225 ;
        RECT 50.855 102.070 51.015 102.180 ;
        RECT 51.315 102.015 51.485 102.205 ;
        RECT 52.235 102.035 52.405 102.225 ;
        RECT 56.835 102.015 57.005 102.205 ;
        RECT 62.355 102.015 62.525 102.205 ;
        RECT 62.815 102.035 62.985 102.225 ;
        RECT 64.195 102.015 64.365 102.205 ;
        RECT 69.715 102.015 69.885 102.205 ;
        RECT 73.395 102.035 73.565 102.225 ;
        RECT 75.235 102.015 75.405 102.225 ;
        RECT 77.075 102.015 77.245 102.205 ;
        RECT 82.595 102.015 82.765 102.205 ;
        RECT 86.275 102.035 86.445 102.225 ;
        RECT 88.115 102.015 88.285 102.205 ;
        RECT 90.415 102.015 90.585 102.205 ;
        RECT 96.855 102.035 97.025 102.225 ;
        RECT 97.370 102.065 97.490 102.175 ;
        RECT 100.995 102.015 101.165 102.225 ;
        RECT 102.835 102.015 103.005 102.205 ;
        RECT 108.355 102.015 108.525 102.205 ;
        RECT 112.035 102.035 112.205 102.225 ;
        RECT 112.495 102.035 112.665 102.225 ;
        RECT 113.875 102.015 114.045 102.205 ;
        RECT 115.255 102.060 115.415 102.170 ;
        RECT 118.935 102.015 119.105 102.205 ;
        RECT 119.395 102.015 119.565 102.205 ;
        RECT 124.455 102.035 124.625 102.225 ;
        RECT 125.825 102.205 125.995 102.225 ;
        RECT 125.825 102.035 126.005 102.205 ;
        RECT 125.835 102.015 126.005 102.035 ;
        RECT 127.215 102.015 127.385 102.225 ;
        RECT 14.375 101.205 15.745 102.015 ;
        RECT 15.755 101.205 18.505 102.015 ;
        RECT 18.515 101.205 24.025 102.015 ;
        RECT 24.045 101.145 24.475 101.930 ;
        RECT 24.695 101.335 35.065 102.015 ;
        RECT 24.695 101.105 26.905 101.335 ;
        RECT 29.625 101.115 30.555 101.335 ;
        RECT 35.075 101.205 36.905 102.015 ;
        RECT 36.925 101.145 37.355 101.930 ;
        RECT 37.375 101.205 38.745 102.015 ;
        RECT 38.755 101.205 44.265 102.015 ;
        RECT 44.275 101.205 49.785 102.015 ;
        RECT 49.805 101.145 50.235 101.930 ;
        RECT 50.255 101.205 51.625 102.015 ;
        RECT 51.635 101.205 57.145 102.015 ;
        RECT 57.155 101.205 62.665 102.015 ;
        RECT 62.685 101.145 63.115 101.930 ;
        RECT 63.135 101.205 64.505 102.015 ;
        RECT 64.515 101.205 70.025 102.015 ;
        RECT 70.035 101.205 75.545 102.015 ;
        RECT 75.565 101.145 75.995 101.930 ;
        RECT 76.015 101.205 77.385 102.015 ;
        RECT 77.395 101.205 82.905 102.015 ;
        RECT 82.915 101.205 88.425 102.015 ;
        RECT 88.445 101.145 88.875 101.930 ;
        RECT 88.895 101.205 90.725 102.015 ;
        RECT 90.935 101.335 101.305 102.015 ;
        RECT 90.935 101.105 93.145 101.335 ;
        RECT 95.865 101.115 96.795 101.335 ;
        RECT 101.325 101.145 101.755 101.930 ;
        RECT 101.775 101.205 103.145 102.015 ;
        RECT 103.155 101.205 108.665 102.015 ;
        RECT 108.675 101.205 114.185 102.015 ;
        RECT 114.205 101.145 114.635 101.930 ;
        RECT 115.575 101.205 119.245 102.015 ;
        RECT 119.265 101.105 120.615 102.015 ;
        RECT 120.635 101.205 126.145 102.015 ;
        RECT 126.155 101.205 127.525 102.015 ;
      LAYER nwell ;
        RECT 14.180 99.210 127.720 100.815 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 14.370 210.835 127.530 211.005 ;
        RECT 14.455 210.085 15.665 210.835 ;
        RECT 14.455 209.545 14.975 210.085 ;
        RECT 15.835 210.065 18.425 210.835 ;
        RECT 18.600 210.290 23.945 210.835 ;
        RECT 15.145 209.375 15.665 209.915 ;
        RECT 14.455 208.285 15.665 209.375 ;
        RECT 15.835 209.375 17.045 209.895 ;
        RECT 17.215 209.545 18.425 210.065 ;
        RECT 15.835 208.285 18.425 209.375 ;
        RECT 20.190 208.720 20.540 209.970 ;
        RECT 22.020 209.460 22.360 210.290 ;
        RECT 24.115 210.110 24.405 210.835 ;
        RECT 24.575 210.085 25.785 210.835 ;
        RECT 25.960 210.290 31.305 210.835 ;
        RECT 31.480 210.290 36.825 210.835 ;
        RECT 18.600 208.285 23.945 208.720 ;
        RECT 24.115 208.285 24.405 209.450 ;
        RECT 24.575 209.375 25.095 209.915 ;
        RECT 25.265 209.545 25.785 210.085 ;
        RECT 24.575 208.285 25.785 209.375 ;
        RECT 27.550 208.720 27.900 209.970 ;
        RECT 29.380 209.460 29.720 210.290 ;
        RECT 33.070 208.720 33.420 209.970 ;
        RECT 34.900 209.460 35.240 210.290 ;
        RECT 36.995 210.110 37.285 210.835 ;
        RECT 37.455 210.085 38.665 210.835 ;
        RECT 38.840 210.290 44.185 210.835 ;
        RECT 44.360 210.290 49.705 210.835 ;
        RECT 25.960 208.285 31.305 208.720 ;
        RECT 31.480 208.285 36.825 208.720 ;
        RECT 36.995 208.285 37.285 209.450 ;
        RECT 37.455 209.375 37.975 209.915 ;
        RECT 38.145 209.545 38.665 210.085 ;
        RECT 37.455 208.285 38.665 209.375 ;
        RECT 40.430 208.720 40.780 209.970 ;
        RECT 42.260 209.460 42.600 210.290 ;
        RECT 45.950 208.720 46.300 209.970 ;
        RECT 47.780 209.460 48.120 210.290 ;
        RECT 49.875 210.110 50.165 210.835 ;
        RECT 50.335 210.085 51.545 210.835 ;
        RECT 51.720 210.290 57.065 210.835 ;
        RECT 57.240 210.290 62.585 210.835 ;
        RECT 38.840 208.285 44.185 208.720 ;
        RECT 44.360 208.285 49.705 208.720 ;
        RECT 49.875 208.285 50.165 209.450 ;
        RECT 50.335 209.375 50.855 209.915 ;
        RECT 51.025 209.545 51.545 210.085 ;
        RECT 50.335 208.285 51.545 209.375 ;
        RECT 53.310 208.720 53.660 209.970 ;
        RECT 55.140 209.460 55.480 210.290 ;
        RECT 58.830 208.720 59.180 209.970 ;
        RECT 60.660 209.460 61.000 210.290 ;
        RECT 62.755 210.110 63.045 210.835 ;
        RECT 63.215 210.085 64.425 210.835 ;
        RECT 64.600 210.290 69.945 210.835 ;
        RECT 70.120 210.290 75.465 210.835 ;
        RECT 51.720 208.285 57.065 208.720 ;
        RECT 57.240 208.285 62.585 208.720 ;
        RECT 62.755 208.285 63.045 209.450 ;
        RECT 63.215 209.375 63.735 209.915 ;
        RECT 63.905 209.545 64.425 210.085 ;
        RECT 63.215 208.285 64.425 209.375 ;
        RECT 66.190 208.720 66.540 209.970 ;
        RECT 68.020 209.460 68.360 210.290 ;
        RECT 71.710 208.720 72.060 209.970 ;
        RECT 73.540 209.460 73.880 210.290 ;
        RECT 75.635 210.110 75.925 210.835 ;
        RECT 76.095 210.085 77.305 210.835 ;
        RECT 77.480 210.290 82.825 210.835 ;
        RECT 83.000 210.290 88.345 210.835 ;
        RECT 64.600 208.285 69.945 208.720 ;
        RECT 70.120 208.285 75.465 208.720 ;
        RECT 75.635 208.285 75.925 209.450 ;
        RECT 76.095 209.375 76.615 209.915 ;
        RECT 76.785 209.545 77.305 210.085 ;
        RECT 76.095 208.285 77.305 209.375 ;
        RECT 79.070 208.720 79.420 209.970 ;
        RECT 80.900 209.460 81.240 210.290 ;
        RECT 84.590 208.720 84.940 209.970 ;
        RECT 86.420 209.460 86.760 210.290 ;
        RECT 88.515 210.110 88.805 210.835 ;
        RECT 88.975 210.085 90.185 210.835 ;
        RECT 90.360 210.290 95.705 210.835 ;
        RECT 95.880 210.290 101.225 210.835 ;
        RECT 77.480 208.285 82.825 208.720 ;
        RECT 83.000 208.285 88.345 208.720 ;
        RECT 88.515 208.285 88.805 209.450 ;
        RECT 88.975 209.375 89.495 209.915 ;
        RECT 89.665 209.545 90.185 210.085 ;
        RECT 88.975 208.285 90.185 209.375 ;
        RECT 91.950 208.720 92.300 209.970 ;
        RECT 93.780 209.460 94.120 210.290 ;
        RECT 97.470 208.720 97.820 209.970 ;
        RECT 99.300 209.460 99.640 210.290 ;
        RECT 101.395 210.110 101.685 210.835 ;
        RECT 101.855 210.085 103.065 210.835 ;
        RECT 103.240 210.290 108.585 210.835 ;
        RECT 108.760 210.290 114.105 210.835 ;
        RECT 90.360 208.285 95.705 208.720 ;
        RECT 95.880 208.285 101.225 208.720 ;
        RECT 101.395 208.285 101.685 209.450 ;
        RECT 101.855 209.375 102.375 209.915 ;
        RECT 102.545 209.545 103.065 210.085 ;
        RECT 101.855 208.285 103.065 209.375 ;
        RECT 104.830 208.720 105.180 209.970 ;
        RECT 106.660 209.460 107.000 210.290 ;
        RECT 110.350 208.720 110.700 209.970 ;
        RECT 112.180 209.460 112.520 210.290 ;
        RECT 114.275 210.110 114.565 210.835 ;
        RECT 115.200 210.290 120.545 210.835 ;
        RECT 120.720 210.290 126.065 210.835 ;
        RECT 103.240 208.285 108.585 208.720 ;
        RECT 108.760 208.285 114.105 208.720 ;
        RECT 114.275 208.285 114.565 209.450 ;
        RECT 116.790 208.720 117.140 209.970 ;
        RECT 118.620 209.460 118.960 210.290 ;
        RECT 122.310 208.720 122.660 209.970 ;
        RECT 124.140 209.460 124.480 210.290 ;
        RECT 126.235 210.085 127.445 210.835 ;
        RECT 126.235 209.375 126.755 209.915 ;
        RECT 126.925 209.545 127.445 210.085 ;
        RECT 115.200 208.285 120.545 208.720 ;
        RECT 120.720 208.285 126.065 208.720 ;
        RECT 126.235 208.285 127.445 209.375 ;
        RECT 14.370 208.115 127.530 208.285 ;
        RECT 14.455 207.025 15.665 208.115 ;
        RECT 14.455 206.315 14.975 206.855 ;
        RECT 15.145 206.485 15.665 207.025 ;
        RECT 15.835 207.025 18.425 208.115 ;
        RECT 18.600 207.680 23.945 208.115 ;
        RECT 15.835 206.505 17.045 207.025 ;
        RECT 17.215 206.335 18.425 206.855 ;
        RECT 20.190 206.430 20.540 207.680 ;
        RECT 24.115 206.950 24.405 208.115 ;
        RECT 25.035 207.025 27.625 208.115 ;
        RECT 27.800 207.680 33.145 208.115 ;
        RECT 33.320 207.680 38.665 208.115 ;
        RECT 38.840 207.680 44.185 208.115 ;
        RECT 44.360 207.680 49.705 208.115 ;
        RECT 14.455 205.565 15.665 206.315 ;
        RECT 15.835 205.565 18.425 206.335 ;
        RECT 22.020 206.110 22.360 206.940 ;
        RECT 25.035 206.505 26.245 207.025 ;
        RECT 26.415 206.335 27.625 206.855 ;
        RECT 29.390 206.430 29.740 207.680 ;
        RECT 18.600 205.565 23.945 206.110 ;
        RECT 24.115 205.565 24.405 206.290 ;
        RECT 25.035 205.565 27.625 206.335 ;
        RECT 31.220 206.110 31.560 206.940 ;
        RECT 34.910 206.430 35.260 207.680 ;
        RECT 36.740 206.110 37.080 206.940 ;
        RECT 40.430 206.430 40.780 207.680 ;
        RECT 42.260 206.110 42.600 206.940 ;
        RECT 45.950 206.430 46.300 207.680 ;
        RECT 49.875 206.950 50.165 208.115 ;
        RECT 50.340 207.680 55.685 208.115 ;
        RECT 55.860 207.680 61.205 208.115 ;
        RECT 61.380 207.680 66.725 208.115 ;
        RECT 66.900 207.680 72.245 208.115 ;
        RECT 47.780 206.110 48.120 206.940 ;
        RECT 51.930 206.430 52.280 207.680 ;
        RECT 27.800 205.565 33.145 206.110 ;
        RECT 33.320 205.565 38.665 206.110 ;
        RECT 38.840 205.565 44.185 206.110 ;
        RECT 44.360 205.565 49.705 206.110 ;
        RECT 49.875 205.565 50.165 206.290 ;
        RECT 53.760 206.110 54.100 206.940 ;
        RECT 57.450 206.430 57.800 207.680 ;
        RECT 59.280 206.110 59.620 206.940 ;
        RECT 62.970 206.430 63.320 207.680 ;
        RECT 64.800 206.110 65.140 206.940 ;
        RECT 68.490 206.430 68.840 207.680 ;
        RECT 72.455 206.975 72.685 208.115 ;
        RECT 72.855 206.965 73.185 207.945 ;
        RECT 73.355 206.975 73.565 208.115 ;
        RECT 73.885 207.185 74.055 207.945 ;
        RECT 74.270 207.355 74.600 208.115 ;
        RECT 73.885 207.015 74.600 207.185 ;
        RECT 74.770 207.040 75.025 207.945 ;
        RECT 70.320 206.110 70.660 206.940 ;
        RECT 72.435 206.555 72.765 206.805 ;
        RECT 50.340 205.565 55.685 206.110 ;
        RECT 55.860 205.565 61.205 206.110 ;
        RECT 61.380 205.565 66.725 206.110 ;
        RECT 66.900 205.565 72.245 206.110 ;
        RECT 72.455 205.565 72.685 206.385 ;
        RECT 72.935 206.365 73.185 206.965 ;
        RECT 73.795 206.465 74.150 206.835 ;
        RECT 74.430 206.805 74.600 207.015 ;
        RECT 74.430 206.475 74.685 206.805 ;
        RECT 72.855 205.735 73.185 206.365 ;
        RECT 73.355 205.565 73.565 206.385 ;
        RECT 74.430 206.285 74.600 206.475 ;
        RECT 74.855 206.310 75.025 207.040 ;
        RECT 75.200 206.965 75.460 208.115 ;
        RECT 75.635 206.950 75.925 208.115 ;
        RECT 77.035 207.605 77.335 208.115 ;
        RECT 77.505 207.605 77.885 207.775 ;
        RECT 78.465 207.605 79.095 208.115 ;
        RECT 77.505 207.435 77.675 207.605 ;
        RECT 79.265 207.435 79.595 207.945 ;
        RECT 79.765 207.605 80.065 208.115 ;
        RECT 77.015 207.235 77.675 207.435 ;
        RECT 77.845 207.265 80.065 207.435 ;
        RECT 73.885 206.115 74.600 206.285 ;
        RECT 73.885 205.735 74.055 206.115 ;
        RECT 74.270 205.565 74.600 205.945 ;
        RECT 74.770 205.735 75.025 206.310 ;
        RECT 75.200 205.565 75.460 206.405 ;
        RECT 77.015 206.305 77.185 207.235 ;
        RECT 77.845 207.065 78.015 207.265 ;
        RECT 77.355 206.895 78.015 207.065 ;
        RECT 78.185 206.925 79.725 207.095 ;
        RECT 77.355 206.475 77.525 206.895 ;
        RECT 78.185 206.725 78.355 206.925 ;
        RECT 77.755 206.555 78.355 206.725 ;
        RECT 78.525 206.555 79.220 206.755 ;
        RECT 79.480 206.475 79.725 206.925 ;
        RECT 77.845 206.305 78.755 206.385 ;
        RECT 75.635 205.565 75.925 206.290 ;
        RECT 77.015 205.825 77.335 206.305 ;
        RECT 77.505 206.215 78.755 206.305 ;
        RECT 77.505 206.135 78.015 206.215 ;
        RECT 77.505 205.735 77.735 206.135 ;
        RECT 77.905 205.565 78.255 205.955 ;
        RECT 78.425 205.735 78.755 206.215 ;
        RECT 78.925 205.565 79.095 206.385 ;
        RECT 79.895 206.305 80.065 207.265 ;
        RECT 81.155 207.025 84.665 208.115 ;
        RECT 84.840 207.680 90.185 208.115 ;
        RECT 90.360 207.680 95.705 208.115 ;
        RECT 95.880 207.680 101.225 208.115 ;
        RECT 81.155 206.505 82.845 207.025 ;
        RECT 83.015 206.335 84.665 206.855 ;
        RECT 86.430 206.430 86.780 207.680 ;
        RECT 79.600 205.760 80.065 206.305 ;
        RECT 81.155 205.565 84.665 206.335 ;
        RECT 88.260 206.110 88.600 206.940 ;
        RECT 91.950 206.430 92.300 207.680 ;
        RECT 93.780 206.110 94.120 206.940 ;
        RECT 97.470 206.430 97.820 207.680 ;
        RECT 101.395 206.950 101.685 208.115 ;
        RECT 102.315 207.025 103.985 208.115 ;
        RECT 104.160 207.680 109.505 208.115 ;
        RECT 109.680 207.680 115.025 208.115 ;
        RECT 115.200 207.680 120.545 208.115 ;
        RECT 120.720 207.680 126.065 208.115 ;
        RECT 99.300 206.110 99.640 206.940 ;
        RECT 102.315 206.505 103.065 207.025 ;
        RECT 103.235 206.335 103.985 206.855 ;
        RECT 105.750 206.430 106.100 207.680 ;
        RECT 84.840 205.565 90.185 206.110 ;
        RECT 90.360 205.565 95.705 206.110 ;
        RECT 95.880 205.565 101.225 206.110 ;
        RECT 101.395 205.565 101.685 206.290 ;
        RECT 102.315 205.565 103.985 206.335 ;
        RECT 107.580 206.110 107.920 206.940 ;
        RECT 111.270 206.430 111.620 207.680 ;
        RECT 113.100 206.110 113.440 206.940 ;
        RECT 116.790 206.430 117.140 207.680 ;
        RECT 118.620 206.110 118.960 206.940 ;
        RECT 122.310 206.430 122.660 207.680 ;
        RECT 126.235 207.025 127.445 208.115 ;
        RECT 124.140 206.110 124.480 206.940 ;
        RECT 126.235 206.485 126.755 207.025 ;
        RECT 126.925 206.315 127.445 206.855 ;
        RECT 104.160 205.565 109.505 206.110 ;
        RECT 109.680 205.565 115.025 206.110 ;
        RECT 115.200 205.565 120.545 206.110 ;
        RECT 120.720 205.565 126.065 206.110 ;
        RECT 126.235 205.565 127.445 206.315 ;
        RECT 14.370 205.395 127.530 205.565 ;
        RECT 14.455 204.645 15.665 205.395 ;
        RECT 14.455 204.105 14.975 204.645 ;
        RECT 16.755 204.625 20.265 205.395 ;
        RECT 20.440 204.850 25.785 205.395 ;
        RECT 25.960 204.850 31.305 205.395 ;
        RECT 31.480 204.850 36.825 205.395 ;
        RECT 15.145 203.935 15.665 204.475 ;
        RECT 14.455 202.845 15.665 203.935 ;
        RECT 16.755 203.935 18.445 204.455 ;
        RECT 18.615 204.105 20.265 204.625 ;
        RECT 16.755 202.845 20.265 203.935 ;
        RECT 22.030 203.280 22.380 204.530 ;
        RECT 23.860 204.020 24.200 204.850 ;
        RECT 27.550 203.280 27.900 204.530 ;
        RECT 29.380 204.020 29.720 204.850 ;
        RECT 33.070 203.280 33.420 204.530 ;
        RECT 34.900 204.020 35.240 204.850 ;
        RECT 36.995 204.670 37.285 205.395 ;
        RECT 37.915 204.625 40.505 205.395 ;
        RECT 40.680 204.850 46.025 205.395 ;
        RECT 46.200 204.850 51.545 205.395 ;
        RECT 51.720 204.850 57.065 205.395 ;
        RECT 57.240 204.850 62.585 205.395 ;
        RECT 20.440 202.845 25.785 203.280 ;
        RECT 25.960 202.845 31.305 203.280 ;
        RECT 31.480 202.845 36.825 203.280 ;
        RECT 36.995 202.845 37.285 204.010 ;
        RECT 37.915 203.935 39.125 204.455 ;
        RECT 39.295 204.105 40.505 204.625 ;
        RECT 37.915 202.845 40.505 203.935 ;
        RECT 42.270 203.280 42.620 204.530 ;
        RECT 44.100 204.020 44.440 204.850 ;
        RECT 47.790 203.280 48.140 204.530 ;
        RECT 49.620 204.020 49.960 204.850 ;
        RECT 53.310 203.280 53.660 204.530 ;
        RECT 55.140 204.020 55.480 204.850 ;
        RECT 58.830 203.280 59.180 204.530 ;
        RECT 60.660 204.020 61.000 204.850 ;
        RECT 62.755 204.670 63.045 205.395 ;
        RECT 63.215 204.645 64.425 205.395 ;
        RECT 40.680 202.845 46.025 203.280 ;
        RECT 46.200 202.845 51.545 203.280 ;
        RECT 51.720 202.845 57.065 203.280 ;
        RECT 57.240 202.845 62.585 203.280 ;
        RECT 62.755 202.845 63.045 204.010 ;
        RECT 63.215 203.935 63.735 204.475 ;
        RECT 63.905 204.105 64.425 204.645 ;
        RECT 64.655 204.575 64.865 205.395 ;
        RECT 65.035 204.595 65.365 205.225 ;
        RECT 65.035 203.995 65.285 204.595 ;
        RECT 65.535 204.575 65.765 205.395 ;
        RECT 66.935 204.575 67.165 205.395 ;
        RECT 67.335 204.595 67.665 205.225 ;
        RECT 65.455 204.155 65.785 204.405 ;
        RECT 66.915 204.155 67.245 204.405 ;
        RECT 67.415 203.995 67.665 204.595 ;
        RECT 67.835 204.575 68.045 205.395 ;
        RECT 68.280 204.685 68.535 205.215 ;
        RECT 68.705 204.935 69.010 205.395 ;
        RECT 69.255 205.015 70.325 205.185 ;
        RECT 63.215 202.845 64.425 203.935 ;
        RECT 64.655 202.845 64.865 203.985 ;
        RECT 65.035 203.015 65.365 203.995 ;
        RECT 65.535 202.845 65.765 203.985 ;
        RECT 66.935 202.845 67.165 203.985 ;
        RECT 67.335 203.015 67.665 203.995 ;
        RECT 68.280 204.035 68.490 204.685 ;
        RECT 69.255 204.660 69.575 205.015 ;
        RECT 69.250 204.485 69.575 204.660 ;
        RECT 68.660 204.185 69.575 204.485 ;
        RECT 69.745 204.445 69.985 204.845 ;
        RECT 70.155 204.785 70.325 205.015 ;
        RECT 70.495 204.955 70.685 205.395 ;
        RECT 70.855 204.945 71.805 205.225 ;
        RECT 72.025 205.035 72.375 205.205 ;
        RECT 70.155 204.615 70.685 204.785 ;
        RECT 68.660 204.155 69.400 204.185 ;
        RECT 67.835 202.845 68.045 203.985 ;
        RECT 68.280 203.155 68.535 204.035 ;
        RECT 68.705 202.845 69.010 203.985 ;
        RECT 69.230 203.565 69.400 204.155 ;
        RECT 69.745 204.075 70.285 204.445 ;
        RECT 70.465 204.335 70.685 204.615 ;
        RECT 70.855 204.165 71.025 204.945 ;
        RECT 70.620 203.995 71.025 204.165 ;
        RECT 71.195 204.155 71.545 204.775 ;
        RECT 70.620 203.905 70.790 203.995 ;
        RECT 71.715 203.985 71.925 204.775 ;
        RECT 69.570 203.735 70.790 203.905 ;
        RECT 71.250 203.825 71.925 203.985 ;
        RECT 69.230 203.395 70.030 203.565 ;
        RECT 69.350 202.845 69.680 203.225 ;
        RECT 69.860 203.105 70.030 203.395 ;
        RECT 70.620 203.355 70.790 203.735 ;
        RECT 70.960 203.815 71.925 203.825 ;
        RECT 72.115 204.645 72.375 205.035 ;
        RECT 72.585 204.935 72.915 205.395 ;
        RECT 73.790 205.005 74.645 205.175 ;
        RECT 74.850 205.005 75.345 205.175 ;
        RECT 75.515 205.035 75.845 205.395 ;
        RECT 72.115 203.955 72.285 204.645 ;
        RECT 72.455 204.295 72.625 204.475 ;
        RECT 72.795 204.465 73.585 204.715 ;
        RECT 73.790 204.295 73.960 205.005 ;
        RECT 74.130 204.495 74.485 204.715 ;
        RECT 72.455 204.125 74.145 204.295 ;
        RECT 70.960 203.525 71.420 203.815 ;
        RECT 72.115 203.785 73.615 203.955 ;
        RECT 72.115 203.645 72.285 203.785 ;
        RECT 71.725 203.475 72.285 203.645 ;
        RECT 70.200 202.845 70.450 203.305 ;
        RECT 70.620 203.015 71.490 203.355 ;
        RECT 71.725 203.015 71.895 203.475 ;
        RECT 72.730 203.445 73.805 203.615 ;
        RECT 72.065 202.845 72.435 203.305 ;
        RECT 72.730 203.105 72.900 203.445 ;
        RECT 73.070 202.845 73.400 203.275 ;
        RECT 73.635 203.105 73.805 203.445 ;
        RECT 73.975 203.345 74.145 204.125 ;
        RECT 74.315 203.905 74.485 204.495 ;
        RECT 74.655 204.095 75.005 204.715 ;
        RECT 74.315 203.515 74.780 203.905 ;
        RECT 75.175 203.645 75.345 205.005 ;
        RECT 75.515 203.815 75.975 204.865 ;
        RECT 74.950 203.475 75.345 203.645 ;
        RECT 74.950 203.345 75.120 203.475 ;
        RECT 73.975 203.015 74.655 203.345 ;
        RECT 74.870 203.015 75.120 203.345 ;
        RECT 75.290 202.845 75.540 203.305 ;
        RECT 75.710 203.030 76.035 203.815 ;
        RECT 76.205 203.015 76.375 205.135 ;
        RECT 76.545 205.015 76.875 205.395 ;
        RECT 77.045 204.845 77.300 205.135 ;
        RECT 76.550 204.675 77.300 204.845 ;
        RECT 77.480 204.685 77.735 205.215 ;
        RECT 77.905 204.935 78.210 205.395 ;
        RECT 78.455 205.015 79.525 205.185 ;
        RECT 76.550 203.685 76.780 204.675 ;
        RECT 76.950 203.855 77.300 204.505 ;
        RECT 77.480 204.035 77.690 204.685 ;
        RECT 78.455 204.660 78.775 205.015 ;
        RECT 78.450 204.485 78.775 204.660 ;
        RECT 77.860 204.185 78.775 204.485 ;
        RECT 78.945 204.445 79.185 204.845 ;
        RECT 79.355 204.785 79.525 205.015 ;
        RECT 79.695 204.955 79.885 205.395 ;
        RECT 80.055 204.945 81.005 205.225 ;
        RECT 81.225 205.035 81.575 205.205 ;
        RECT 79.355 204.615 79.885 204.785 ;
        RECT 77.860 204.155 78.600 204.185 ;
        RECT 76.550 203.515 77.300 203.685 ;
        RECT 76.545 202.845 76.875 203.345 ;
        RECT 77.045 203.015 77.300 203.515 ;
        RECT 77.480 203.155 77.735 204.035 ;
        RECT 77.905 202.845 78.210 203.985 ;
        RECT 78.430 203.565 78.600 204.155 ;
        RECT 78.945 204.075 79.485 204.445 ;
        RECT 79.665 204.335 79.885 204.615 ;
        RECT 80.055 204.165 80.225 204.945 ;
        RECT 79.820 203.995 80.225 204.165 ;
        RECT 80.395 204.155 80.745 204.775 ;
        RECT 79.820 203.905 79.990 203.995 ;
        RECT 80.915 203.985 81.125 204.775 ;
        RECT 78.770 203.735 79.990 203.905 ;
        RECT 80.450 203.825 81.125 203.985 ;
        RECT 78.430 203.395 79.230 203.565 ;
        RECT 78.550 202.845 78.880 203.225 ;
        RECT 79.060 203.105 79.230 203.395 ;
        RECT 79.820 203.355 79.990 203.735 ;
        RECT 80.160 203.815 81.125 203.825 ;
        RECT 81.315 204.645 81.575 205.035 ;
        RECT 81.785 204.935 82.115 205.395 ;
        RECT 82.990 205.005 83.845 205.175 ;
        RECT 84.050 205.005 84.545 205.175 ;
        RECT 84.715 205.035 85.045 205.395 ;
        RECT 81.315 203.955 81.485 204.645 ;
        RECT 81.655 204.295 81.825 204.475 ;
        RECT 81.995 204.465 82.785 204.715 ;
        RECT 82.990 204.295 83.160 205.005 ;
        RECT 83.330 204.495 83.685 204.715 ;
        RECT 81.655 204.125 83.345 204.295 ;
        RECT 80.160 203.525 80.620 203.815 ;
        RECT 81.315 203.785 82.815 203.955 ;
        RECT 81.315 203.645 81.485 203.785 ;
        RECT 80.925 203.475 81.485 203.645 ;
        RECT 79.400 202.845 79.650 203.305 ;
        RECT 79.820 203.015 80.690 203.355 ;
        RECT 80.925 203.015 81.095 203.475 ;
        RECT 81.930 203.445 83.005 203.615 ;
        RECT 81.265 202.845 81.635 203.305 ;
        RECT 81.930 203.105 82.100 203.445 ;
        RECT 82.270 202.845 82.600 203.275 ;
        RECT 82.835 203.105 83.005 203.445 ;
        RECT 83.175 203.345 83.345 204.125 ;
        RECT 83.515 203.905 83.685 204.495 ;
        RECT 83.855 204.095 84.205 204.715 ;
        RECT 83.515 203.515 83.980 203.905 ;
        RECT 84.375 203.645 84.545 205.005 ;
        RECT 84.715 203.815 85.175 204.865 ;
        RECT 84.150 203.475 84.545 203.645 ;
        RECT 84.150 203.345 84.320 203.475 ;
        RECT 83.175 203.015 83.855 203.345 ;
        RECT 84.070 203.015 84.320 203.345 ;
        RECT 84.490 202.845 84.740 203.305 ;
        RECT 84.910 203.030 85.235 203.815 ;
        RECT 85.405 203.015 85.575 205.135 ;
        RECT 85.745 205.015 86.075 205.395 ;
        RECT 86.245 204.845 86.500 205.135 ;
        RECT 85.750 204.675 86.500 204.845 ;
        RECT 85.750 203.685 85.980 204.675 ;
        RECT 86.675 204.625 88.345 205.395 ;
        RECT 88.515 204.670 88.805 205.395 ;
        RECT 89.435 204.625 92.025 205.395 ;
        RECT 92.200 204.850 97.545 205.395 ;
        RECT 97.720 204.850 103.065 205.395 ;
        RECT 103.240 204.850 108.585 205.395 ;
        RECT 108.760 204.850 114.105 205.395 ;
        RECT 86.150 203.855 86.500 204.505 ;
        RECT 86.675 203.935 87.425 204.455 ;
        RECT 87.595 204.105 88.345 204.625 ;
        RECT 85.750 203.515 86.500 203.685 ;
        RECT 85.745 202.845 86.075 203.345 ;
        RECT 86.245 203.015 86.500 203.515 ;
        RECT 86.675 202.845 88.345 203.935 ;
        RECT 88.515 202.845 88.805 204.010 ;
        RECT 89.435 203.935 90.645 204.455 ;
        RECT 90.815 204.105 92.025 204.625 ;
        RECT 89.435 202.845 92.025 203.935 ;
        RECT 93.790 203.280 94.140 204.530 ;
        RECT 95.620 204.020 95.960 204.850 ;
        RECT 99.310 203.280 99.660 204.530 ;
        RECT 101.140 204.020 101.480 204.850 ;
        RECT 104.830 203.280 105.180 204.530 ;
        RECT 106.660 204.020 107.000 204.850 ;
        RECT 110.350 203.280 110.700 204.530 ;
        RECT 112.180 204.020 112.520 204.850 ;
        RECT 114.275 204.670 114.565 205.395 ;
        RECT 115.200 204.850 120.545 205.395 ;
        RECT 120.720 204.850 126.065 205.395 ;
        RECT 92.200 202.845 97.545 203.280 ;
        RECT 97.720 202.845 103.065 203.280 ;
        RECT 103.240 202.845 108.585 203.280 ;
        RECT 108.760 202.845 114.105 203.280 ;
        RECT 114.275 202.845 114.565 204.010 ;
        RECT 116.790 203.280 117.140 204.530 ;
        RECT 118.620 204.020 118.960 204.850 ;
        RECT 122.310 203.280 122.660 204.530 ;
        RECT 124.140 204.020 124.480 204.850 ;
        RECT 126.235 204.645 127.445 205.395 ;
        RECT 126.235 203.935 126.755 204.475 ;
        RECT 126.925 204.105 127.445 204.645 ;
        RECT 115.200 202.845 120.545 203.280 ;
        RECT 120.720 202.845 126.065 203.280 ;
        RECT 126.235 202.845 127.445 203.935 ;
        RECT 14.370 202.675 127.530 202.845 ;
        RECT 14.455 201.585 15.665 202.675 ;
        RECT 14.455 200.875 14.975 201.415 ;
        RECT 15.145 201.045 15.665 201.585 ;
        RECT 15.835 201.585 18.425 202.675 ;
        RECT 18.600 202.240 23.945 202.675 ;
        RECT 15.835 201.065 17.045 201.585 ;
        RECT 17.215 200.895 18.425 201.415 ;
        RECT 20.190 200.990 20.540 202.240 ;
        RECT 24.115 201.510 24.405 202.675 ;
        RECT 25.035 201.585 27.625 202.675 ;
        RECT 27.800 202.240 33.145 202.675 ;
        RECT 33.320 202.240 38.665 202.675 ;
        RECT 38.840 202.240 44.185 202.675 ;
        RECT 44.360 202.240 49.705 202.675 ;
        RECT 14.455 200.125 15.665 200.875 ;
        RECT 15.835 200.125 18.425 200.895 ;
        RECT 22.020 200.670 22.360 201.500 ;
        RECT 25.035 201.065 26.245 201.585 ;
        RECT 26.415 200.895 27.625 201.415 ;
        RECT 29.390 200.990 29.740 202.240 ;
        RECT 18.600 200.125 23.945 200.670 ;
        RECT 24.115 200.125 24.405 200.850 ;
        RECT 25.035 200.125 27.625 200.895 ;
        RECT 31.220 200.670 31.560 201.500 ;
        RECT 34.910 200.990 35.260 202.240 ;
        RECT 36.740 200.670 37.080 201.500 ;
        RECT 40.430 200.990 40.780 202.240 ;
        RECT 42.260 200.670 42.600 201.500 ;
        RECT 45.950 200.990 46.300 202.240 ;
        RECT 49.875 201.510 50.165 202.675 ;
        RECT 50.335 201.585 53.845 202.675 ;
        RECT 54.020 202.240 59.365 202.675 ;
        RECT 47.780 200.670 48.120 201.500 ;
        RECT 50.335 201.065 52.025 201.585 ;
        RECT 52.195 200.895 53.845 201.415 ;
        RECT 55.610 200.990 55.960 202.240 ;
        RECT 59.540 202.005 59.795 202.505 ;
        RECT 59.965 202.175 60.295 202.675 ;
        RECT 59.540 201.835 60.290 202.005 ;
        RECT 27.800 200.125 33.145 200.670 ;
        RECT 33.320 200.125 38.665 200.670 ;
        RECT 38.840 200.125 44.185 200.670 ;
        RECT 44.360 200.125 49.705 200.670 ;
        RECT 49.875 200.125 50.165 200.850 ;
        RECT 50.335 200.125 53.845 200.895 ;
        RECT 57.440 200.670 57.780 201.500 ;
        RECT 59.540 201.015 59.890 201.665 ;
        RECT 60.060 200.845 60.290 201.835 ;
        RECT 59.540 200.675 60.290 200.845 ;
        RECT 54.020 200.125 59.365 200.670 ;
        RECT 59.540 200.385 59.795 200.675 ;
        RECT 59.965 200.125 60.295 200.505 ;
        RECT 60.465 200.385 60.635 202.505 ;
        RECT 60.805 201.705 61.130 202.490 ;
        RECT 61.300 202.215 61.550 202.675 ;
        RECT 61.720 202.175 61.970 202.505 ;
        RECT 62.185 202.175 62.865 202.505 ;
        RECT 61.720 202.045 61.890 202.175 ;
        RECT 61.495 201.875 61.890 202.045 ;
        RECT 60.865 200.655 61.325 201.705 ;
        RECT 61.495 200.515 61.665 201.875 ;
        RECT 62.060 201.615 62.525 202.005 ;
        RECT 61.835 200.805 62.185 201.425 ;
        RECT 62.355 201.025 62.525 201.615 ;
        RECT 62.695 201.395 62.865 202.175 ;
        RECT 63.035 202.075 63.205 202.415 ;
        RECT 63.440 202.245 63.770 202.675 ;
        RECT 63.940 202.075 64.110 202.415 ;
        RECT 64.405 202.215 64.775 202.675 ;
        RECT 63.035 201.905 64.110 202.075 ;
        RECT 64.945 202.045 65.115 202.505 ;
        RECT 65.350 202.165 66.220 202.505 ;
        RECT 66.390 202.215 66.640 202.675 ;
        RECT 64.555 201.875 65.115 202.045 ;
        RECT 64.555 201.735 64.725 201.875 ;
        RECT 63.225 201.565 64.725 201.735 ;
        RECT 65.420 201.705 65.880 201.995 ;
        RECT 62.695 201.225 64.385 201.395 ;
        RECT 62.355 200.805 62.710 201.025 ;
        RECT 62.880 200.515 63.050 201.225 ;
        RECT 63.255 200.805 64.045 201.055 ;
        RECT 64.215 201.045 64.385 201.225 ;
        RECT 64.555 200.875 64.725 201.565 ;
        RECT 60.995 200.125 61.325 200.485 ;
        RECT 61.495 200.345 61.990 200.515 ;
        RECT 62.195 200.345 63.050 200.515 ;
        RECT 63.925 200.125 64.255 200.585 ;
        RECT 64.465 200.485 64.725 200.875 ;
        RECT 64.915 201.695 65.880 201.705 ;
        RECT 66.050 201.785 66.220 202.165 ;
        RECT 66.810 202.125 66.980 202.415 ;
        RECT 67.160 202.295 67.490 202.675 ;
        RECT 66.810 201.955 67.610 202.125 ;
        RECT 64.915 201.535 65.590 201.695 ;
        RECT 66.050 201.615 67.270 201.785 ;
        RECT 64.915 200.745 65.125 201.535 ;
        RECT 66.050 201.525 66.220 201.615 ;
        RECT 65.295 200.745 65.645 201.365 ;
        RECT 65.815 201.355 66.220 201.525 ;
        RECT 65.815 200.575 65.985 201.355 ;
        RECT 66.155 200.905 66.375 201.185 ;
        RECT 66.555 201.075 67.095 201.445 ;
        RECT 67.440 201.335 67.610 201.955 ;
        RECT 67.785 201.615 67.955 202.675 ;
        RECT 68.165 201.665 68.455 202.505 ;
        RECT 68.625 201.835 68.795 202.675 ;
        RECT 69.005 201.665 69.255 202.505 ;
        RECT 69.465 201.835 69.635 202.675 ;
        RECT 68.165 201.495 69.890 201.665 ;
        RECT 66.155 200.735 66.685 200.905 ;
        RECT 64.465 200.315 64.815 200.485 ;
        RECT 65.035 200.295 65.985 200.575 ;
        RECT 66.155 200.125 66.345 200.565 ;
        RECT 66.515 200.505 66.685 200.735 ;
        RECT 66.855 200.675 67.095 201.075 ;
        RECT 67.265 201.325 67.610 201.335 ;
        RECT 67.265 201.115 69.295 201.325 ;
        RECT 67.265 200.860 67.590 201.115 ;
        RECT 69.480 200.945 69.890 201.495 ;
        RECT 67.265 200.505 67.585 200.860 ;
        RECT 66.515 200.335 67.585 200.505 ;
        RECT 67.785 200.125 67.955 200.935 ;
        RECT 68.125 200.775 69.890 200.945 ;
        RECT 70.115 201.535 70.375 202.505 ;
        RECT 70.570 202.265 70.900 202.675 ;
        RECT 71.100 202.085 71.270 202.505 ;
        RECT 71.485 202.265 72.155 202.675 ;
        RECT 72.390 202.085 72.560 202.505 ;
        RECT 72.865 202.235 73.195 202.675 ;
        RECT 70.545 201.915 72.560 202.085 ;
        RECT 73.365 202.055 73.540 202.505 ;
        RECT 73.800 202.250 74.135 202.675 ;
        RECT 74.305 202.070 74.490 202.475 ;
        RECT 70.115 200.845 70.285 201.535 ;
        RECT 70.545 201.365 70.715 201.915 ;
        RECT 70.455 201.035 70.715 201.365 ;
        RECT 68.125 200.295 68.455 200.775 ;
        RECT 68.625 200.125 68.795 200.595 ;
        RECT 68.965 200.295 69.295 200.775 ;
        RECT 69.465 200.125 69.635 200.595 ;
        RECT 70.115 200.380 70.455 200.845 ;
        RECT 70.885 200.705 71.225 201.735 ;
        RECT 71.415 200.635 71.685 201.735 ;
        RECT 70.120 200.335 70.455 200.380 ;
        RECT 70.625 200.125 70.955 200.505 ;
        RECT 71.415 200.465 71.725 200.635 ;
        RECT 71.415 200.460 71.685 200.465 ;
        RECT 71.910 200.460 72.190 201.735 ;
        RECT 72.390 200.625 72.560 201.915 ;
        RECT 72.910 201.885 73.540 202.055 ;
        RECT 73.825 201.895 74.490 202.070 ;
        RECT 74.695 201.895 75.025 202.675 ;
        RECT 72.910 201.365 73.080 201.885 ;
        RECT 72.730 201.035 73.080 201.365 ;
        RECT 73.260 201.035 73.625 201.715 ;
        RECT 72.910 200.865 73.080 201.035 ;
        RECT 73.825 200.865 74.165 201.895 ;
        RECT 75.195 201.705 75.465 202.475 ;
        RECT 74.335 201.535 75.465 201.705 ;
        RECT 74.335 201.035 74.585 201.535 ;
        RECT 72.910 200.695 73.540 200.865 ;
        RECT 73.825 200.695 74.510 200.865 ;
        RECT 74.765 200.785 75.125 201.365 ;
        RECT 72.390 200.295 72.620 200.625 ;
        RECT 72.865 200.125 73.195 200.505 ;
        RECT 73.365 200.295 73.540 200.695 ;
        RECT 73.800 200.125 74.135 200.525 ;
        RECT 74.305 200.295 74.510 200.695 ;
        RECT 75.295 200.625 75.465 201.535 ;
        RECT 75.635 201.510 75.925 202.675 ;
        RECT 76.555 201.805 76.830 202.505 ;
        RECT 77.000 202.130 77.255 202.675 ;
        RECT 77.425 202.165 77.905 202.505 ;
        RECT 78.080 202.120 78.685 202.675 ;
        RECT 78.070 202.020 78.685 202.120 ;
        RECT 78.070 201.995 78.255 202.020 ;
        RECT 74.720 200.125 74.995 200.605 ;
        RECT 75.205 200.295 75.465 200.625 ;
        RECT 75.635 200.125 75.925 200.850 ;
        RECT 76.555 200.775 76.725 201.805 ;
        RECT 77.000 201.675 77.755 201.925 ;
        RECT 77.925 201.750 78.255 201.995 ;
        RECT 77.000 201.640 77.770 201.675 ;
        RECT 77.000 201.630 77.785 201.640 ;
        RECT 76.895 201.615 77.790 201.630 ;
        RECT 76.895 201.600 77.810 201.615 ;
        RECT 76.895 201.590 77.830 201.600 ;
        RECT 76.895 201.580 77.855 201.590 ;
        RECT 76.895 201.550 77.925 201.580 ;
        RECT 76.895 201.520 77.945 201.550 ;
        RECT 76.895 201.490 77.965 201.520 ;
        RECT 76.895 201.465 77.995 201.490 ;
        RECT 76.895 201.430 78.030 201.465 ;
        RECT 76.895 201.425 78.060 201.430 ;
        RECT 76.895 201.030 77.125 201.425 ;
        RECT 77.670 201.420 78.060 201.425 ;
        RECT 77.695 201.410 78.060 201.420 ;
        RECT 77.710 201.405 78.060 201.410 ;
        RECT 77.725 201.400 78.060 201.405 ;
        RECT 78.425 201.400 78.685 201.850 ;
        RECT 77.725 201.395 78.685 201.400 ;
        RECT 77.735 201.385 78.685 201.395 ;
        RECT 77.745 201.380 78.685 201.385 ;
        RECT 77.755 201.370 78.685 201.380 ;
        RECT 77.760 201.360 78.685 201.370 ;
        RECT 77.765 201.355 78.685 201.360 ;
        RECT 77.775 201.340 78.685 201.355 ;
        RECT 77.780 201.325 78.685 201.340 ;
        RECT 77.790 201.300 78.685 201.325 ;
        RECT 77.295 200.830 77.625 201.255 ;
        RECT 77.375 200.805 77.625 200.830 ;
        RECT 76.555 200.295 76.815 200.775 ;
        RECT 76.985 200.125 77.235 200.665 ;
        RECT 77.405 200.345 77.625 200.805 ;
        RECT 77.795 201.230 78.685 201.300 ;
        RECT 79.320 201.485 79.575 202.365 ;
        RECT 79.745 201.535 80.050 202.675 ;
        RECT 80.390 202.295 80.720 202.675 ;
        RECT 80.900 202.125 81.070 202.415 ;
        RECT 81.240 202.215 81.490 202.675 ;
        RECT 80.270 201.955 81.070 202.125 ;
        RECT 81.660 202.165 82.530 202.505 ;
        RECT 77.795 200.505 77.965 201.230 ;
        RECT 78.135 200.675 78.685 201.060 ;
        RECT 79.320 200.835 79.530 201.485 ;
        RECT 80.270 201.365 80.440 201.955 ;
        RECT 81.660 201.785 81.830 202.165 ;
        RECT 82.765 202.045 82.935 202.505 ;
        RECT 83.105 202.215 83.475 202.675 ;
        RECT 83.770 202.075 83.940 202.415 ;
        RECT 84.110 202.245 84.440 202.675 ;
        RECT 84.675 202.075 84.845 202.415 ;
        RECT 80.610 201.615 81.830 201.785 ;
        RECT 82.000 201.705 82.460 201.995 ;
        RECT 82.765 201.875 83.325 202.045 ;
        RECT 83.770 201.905 84.845 202.075 ;
        RECT 85.015 202.175 85.695 202.505 ;
        RECT 85.910 202.175 86.160 202.505 ;
        RECT 86.330 202.215 86.580 202.675 ;
        RECT 83.155 201.735 83.325 201.875 ;
        RECT 82.000 201.695 82.965 201.705 ;
        RECT 81.660 201.525 81.830 201.615 ;
        RECT 82.290 201.535 82.965 201.695 ;
        RECT 79.700 201.335 80.440 201.365 ;
        RECT 79.700 201.035 80.615 201.335 ;
        RECT 80.290 200.860 80.615 201.035 ;
        RECT 77.795 200.335 78.685 200.505 ;
        RECT 79.320 200.305 79.575 200.835 ;
        RECT 79.745 200.125 80.050 200.585 ;
        RECT 80.295 200.505 80.615 200.860 ;
        RECT 80.785 201.075 81.325 201.445 ;
        RECT 81.660 201.355 82.065 201.525 ;
        RECT 80.785 200.675 81.025 201.075 ;
        RECT 81.505 200.905 81.725 201.185 ;
        RECT 81.195 200.735 81.725 200.905 ;
        RECT 81.195 200.505 81.365 200.735 ;
        RECT 81.895 200.575 82.065 201.355 ;
        RECT 82.235 200.745 82.585 201.365 ;
        RECT 82.755 200.745 82.965 201.535 ;
        RECT 83.155 201.565 84.655 201.735 ;
        RECT 83.155 200.875 83.325 201.565 ;
        RECT 85.015 201.395 85.185 202.175 ;
        RECT 85.990 202.045 86.160 202.175 ;
        RECT 83.495 201.225 85.185 201.395 ;
        RECT 85.355 201.615 85.820 202.005 ;
        RECT 85.990 201.875 86.385 202.045 ;
        RECT 83.495 201.045 83.665 201.225 ;
        RECT 80.295 200.335 81.365 200.505 ;
        RECT 81.535 200.125 81.725 200.565 ;
        RECT 81.895 200.295 82.845 200.575 ;
        RECT 83.155 200.485 83.415 200.875 ;
        RECT 83.835 200.805 84.625 201.055 ;
        RECT 83.065 200.315 83.415 200.485 ;
        RECT 83.625 200.125 83.955 200.585 ;
        RECT 84.830 200.515 85.000 201.225 ;
        RECT 85.355 201.025 85.525 201.615 ;
        RECT 85.170 200.805 85.525 201.025 ;
        RECT 85.695 200.805 86.045 201.425 ;
        RECT 86.215 200.515 86.385 201.875 ;
        RECT 86.750 201.705 87.075 202.490 ;
        RECT 86.555 200.655 87.015 201.705 ;
        RECT 84.830 200.345 85.685 200.515 ;
        RECT 85.890 200.345 86.385 200.515 ;
        RECT 86.555 200.125 86.885 200.485 ;
        RECT 87.245 200.385 87.415 202.505 ;
        RECT 87.585 202.175 87.915 202.675 ;
        RECT 88.085 202.005 88.340 202.505 ;
        RECT 87.590 201.835 88.340 202.005 ;
        RECT 87.590 200.845 87.820 201.835 ;
        RECT 87.990 201.015 88.340 201.665 ;
        RECT 88.515 201.585 90.185 202.675 ;
        RECT 90.360 202.240 95.705 202.675 ;
        RECT 95.880 202.240 101.225 202.675 ;
        RECT 88.515 201.065 89.265 201.585 ;
        RECT 89.435 200.895 90.185 201.415 ;
        RECT 91.950 200.990 92.300 202.240 ;
        RECT 87.590 200.675 88.340 200.845 ;
        RECT 87.585 200.125 87.915 200.505 ;
        RECT 88.085 200.385 88.340 200.675 ;
        RECT 88.515 200.125 90.185 200.895 ;
        RECT 93.780 200.670 94.120 201.500 ;
        RECT 97.470 200.990 97.820 202.240 ;
        RECT 101.395 201.510 101.685 202.675 ;
        RECT 102.315 201.585 103.985 202.675 ;
        RECT 104.160 202.240 109.505 202.675 ;
        RECT 109.680 202.240 115.025 202.675 ;
        RECT 115.200 202.240 120.545 202.675 ;
        RECT 120.720 202.240 126.065 202.675 ;
        RECT 99.300 200.670 99.640 201.500 ;
        RECT 102.315 201.065 103.065 201.585 ;
        RECT 103.235 200.895 103.985 201.415 ;
        RECT 105.750 200.990 106.100 202.240 ;
        RECT 90.360 200.125 95.705 200.670 ;
        RECT 95.880 200.125 101.225 200.670 ;
        RECT 101.395 200.125 101.685 200.850 ;
        RECT 102.315 200.125 103.985 200.895 ;
        RECT 107.580 200.670 107.920 201.500 ;
        RECT 111.270 200.990 111.620 202.240 ;
        RECT 113.100 200.670 113.440 201.500 ;
        RECT 116.790 200.990 117.140 202.240 ;
        RECT 118.620 200.670 118.960 201.500 ;
        RECT 122.310 200.990 122.660 202.240 ;
        RECT 126.235 201.585 127.445 202.675 ;
        RECT 124.140 200.670 124.480 201.500 ;
        RECT 126.235 201.045 126.755 201.585 ;
        RECT 126.925 200.875 127.445 201.415 ;
        RECT 104.160 200.125 109.505 200.670 ;
        RECT 109.680 200.125 115.025 200.670 ;
        RECT 115.200 200.125 120.545 200.670 ;
        RECT 120.720 200.125 126.065 200.670 ;
        RECT 126.235 200.125 127.445 200.875 ;
        RECT 14.370 199.955 127.530 200.125 ;
        RECT 14.455 199.205 15.665 199.955 ;
        RECT 14.455 198.665 14.975 199.205 ;
        RECT 16.755 199.185 20.265 199.955 ;
        RECT 20.440 199.410 25.785 199.955 ;
        RECT 25.960 199.410 31.305 199.955 ;
        RECT 31.480 199.410 36.825 199.955 ;
        RECT 15.145 198.495 15.665 199.035 ;
        RECT 14.455 197.405 15.665 198.495 ;
        RECT 16.755 198.495 18.445 199.015 ;
        RECT 18.615 198.665 20.265 199.185 ;
        RECT 16.755 197.405 20.265 198.495 ;
        RECT 22.030 197.840 22.380 199.090 ;
        RECT 23.860 198.580 24.200 199.410 ;
        RECT 27.550 197.840 27.900 199.090 ;
        RECT 29.380 198.580 29.720 199.410 ;
        RECT 33.070 197.840 33.420 199.090 ;
        RECT 34.900 198.580 35.240 199.410 ;
        RECT 36.995 199.230 37.285 199.955 ;
        RECT 37.915 199.185 40.505 199.955 ;
        RECT 40.680 199.410 46.025 199.955 ;
        RECT 46.200 199.410 51.545 199.955 ;
        RECT 51.720 199.410 57.065 199.955 ;
        RECT 57.240 199.410 62.585 199.955 ;
        RECT 20.440 197.405 25.785 197.840 ;
        RECT 25.960 197.405 31.305 197.840 ;
        RECT 31.480 197.405 36.825 197.840 ;
        RECT 36.995 197.405 37.285 198.570 ;
        RECT 37.915 198.495 39.125 199.015 ;
        RECT 39.295 198.665 40.505 199.185 ;
        RECT 37.915 197.405 40.505 198.495 ;
        RECT 42.270 197.840 42.620 199.090 ;
        RECT 44.100 198.580 44.440 199.410 ;
        RECT 47.790 197.840 48.140 199.090 ;
        RECT 49.620 198.580 49.960 199.410 ;
        RECT 53.310 197.840 53.660 199.090 ;
        RECT 55.140 198.580 55.480 199.410 ;
        RECT 58.830 197.840 59.180 199.090 ;
        RECT 60.660 198.580 61.000 199.410 ;
        RECT 62.755 199.230 63.045 199.955 ;
        RECT 63.675 199.185 67.185 199.955 ;
        RECT 40.680 197.405 46.025 197.840 ;
        RECT 46.200 197.405 51.545 197.840 ;
        RECT 51.720 197.405 57.065 197.840 ;
        RECT 57.240 197.405 62.585 197.840 ;
        RECT 62.755 197.405 63.045 198.570 ;
        RECT 63.675 198.495 65.365 199.015 ;
        RECT 65.535 198.665 67.185 199.185 ;
        RECT 67.355 199.280 67.615 199.785 ;
        RECT 67.795 199.575 68.125 199.955 ;
        RECT 68.305 199.405 68.475 199.785 ;
        RECT 68.740 199.555 69.075 199.955 ;
        RECT 63.675 197.405 67.185 198.495 ;
        RECT 67.355 198.480 67.525 199.280 ;
        RECT 67.810 199.235 68.475 199.405 ;
        RECT 69.245 199.385 69.450 199.785 ;
        RECT 69.660 199.475 69.935 199.955 ;
        RECT 70.145 199.455 70.405 199.785 ;
        RECT 67.810 198.980 67.980 199.235 ;
        RECT 68.765 199.215 69.450 199.385 ;
        RECT 67.695 198.650 67.980 198.980 ;
        RECT 68.215 198.685 68.545 199.055 ;
        RECT 67.810 198.505 67.980 198.650 ;
        RECT 67.355 197.575 67.625 198.480 ;
        RECT 67.810 198.335 68.475 198.505 ;
        RECT 67.795 197.405 68.125 198.165 ;
        RECT 68.305 197.575 68.475 198.335 ;
        RECT 68.765 198.185 69.105 199.215 ;
        RECT 69.275 198.545 69.525 199.045 ;
        RECT 69.705 198.715 70.065 199.295 ;
        RECT 70.235 198.545 70.405 199.455 ;
        RECT 69.275 198.375 70.405 198.545 ;
        RECT 68.765 198.010 69.430 198.185 ;
        RECT 68.740 197.405 69.075 197.830 ;
        RECT 69.245 197.605 69.430 198.010 ;
        RECT 69.635 197.405 69.965 198.185 ;
        RECT 70.135 197.605 70.405 198.375 ;
        RECT 70.575 197.575 70.835 199.785 ;
        RECT 71.005 199.575 71.335 199.955 ;
        RECT 71.545 199.045 71.740 199.620 ;
        RECT 72.010 199.045 72.195 199.625 ;
        RECT 71.005 198.125 71.175 199.045 ;
        RECT 71.485 198.715 71.740 199.045 ;
        RECT 71.965 198.715 72.195 199.045 ;
        RECT 72.445 199.615 73.925 199.785 ;
        RECT 72.445 198.715 72.615 199.615 ;
        RECT 72.785 199.115 73.335 199.445 ;
        RECT 73.525 199.285 73.925 199.615 ;
        RECT 74.105 199.575 74.435 199.955 ;
        RECT 74.745 199.455 75.005 199.785 ;
        RECT 71.545 198.405 71.740 198.715 ;
        RECT 72.010 198.405 72.195 198.715 ;
        RECT 72.785 198.125 72.955 199.115 ;
        RECT 73.525 198.805 73.695 199.285 ;
        RECT 74.275 199.095 74.485 199.275 ;
        RECT 73.865 198.925 74.485 199.095 ;
        RECT 71.005 197.955 72.955 198.125 ;
        RECT 73.125 198.635 73.695 198.805 ;
        RECT 74.835 198.755 75.005 199.455 ;
        RECT 73.125 198.125 73.295 198.635 ;
        RECT 73.875 198.585 75.005 198.755 ;
        RECT 73.875 198.465 74.045 198.585 ;
        RECT 73.465 198.295 74.045 198.465 ;
        RECT 73.125 197.955 73.865 198.125 ;
        RECT 74.315 198.085 74.665 198.415 ;
        RECT 71.005 197.405 71.335 197.785 ;
        RECT 71.760 197.575 71.930 197.955 ;
        RECT 72.190 197.405 72.520 197.785 ;
        RECT 72.715 197.575 72.885 197.955 ;
        RECT 73.095 197.405 73.425 197.785 ;
        RECT 73.675 197.575 73.865 197.955 ;
        RECT 74.835 197.905 75.005 198.585 ;
        RECT 74.105 197.405 74.435 197.785 ;
        RECT 74.745 197.575 75.005 197.905 ;
        RECT 75.175 199.215 75.560 199.785 ;
        RECT 75.730 199.495 76.055 199.955 ;
        RECT 76.575 199.325 76.855 199.785 ;
        RECT 75.175 198.545 75.455 199.215 ;
        RECT 75.730 199.155 76.855 199.325 ;
        RECT 75.730 199.045 76.180 199.155 ;
        RECT 75.625 198.715 76.180 199.045 ;
        RECT 77.045 198.985 77.445 199.785 ;
        RECT 77.845 199.495 78.115 199.955 ;
        RECT 78.285 199.325 78.570 199.785 ;
        RECT 75.175 197.575 75.560 198.545 ;
        RECT 75.730 198.255 76.180 198.715 ;
        RECT 76.350 198.425 77.445 198.985 ;
        RECT 75.730 198.035 76.855 198.255 ;
        RECT 75.730 197.405 76.055 197.865 ;
        RECT 76.575 197.575 76.855 198.035 ;
        RECT 77.045 197.575 77.445 198.425 ;
        RECT 77.615 199.155 78.570 199.325 ;
        RECT 78.890 199.215 79.505 199.785 ;
        RECT 79.675 199.445 79.890 199.955 ;
        RECT 80.120 199.445 80.400 199.775 ;
        RECT 80.580 199.445 80.820 199.955 ;
        RECT 77.615 198.255 77.825 199.155 ;
        RECT 77.995 198.425 78.685 198.985 ;
        RECT 77.615 198.035 78.570 198.255 ;
        RECT 77.845 197.405 78.115 197.865 ;
        RECT 78.285 197.575 78.570 198.035 ;
        RECT 78.890 198.195 79.205 199.215 ;
        RECT 79.375 198.545 79.545 199.045 ;
        RECT 79.795 198.715 80.060 199.275 ;
        RECT 80.230 198.545 80.400 199.445 ;
        RECT 80.570 198.715 80.925 199.275 ;
        RECT 81.155 199.155 81.850 199.785 ;
        RECT 82.055 199.155 82.365 199.955 ;
        RECT 82.625 199.405 82.795 199.785 ;
        RECT 82.975 199.575 83.305 199.955 ;
        RECT 82.625 199.235 83.290 199.405 ;
        RECT 83.485 199.280 83.745 199.785 ;
        RECT 81.175 198.715 81.510 198.965 ;
        RECT 81.680 198.555 81.850 199.155 ;
        RECT 82.020 198.715 82.355 198.985 ;
        RECT 82.555 198.685 82.885 199.055 ;
        RECT 83.120 198.980 83.290 199.235 ;
        RECT 83.120 198.650 83.405 198.980 ;
        RECT 79.375 198.375 80.800 198.545 ;
        RECT 78.890 197.575 79.425 198.195 ;
        RECT 79.595 197.405 79.925 198.205 ;
        RECT 80.410 198.200 80.800 198.375 ;
        RECT 81.155 197.405 81.415 198.545 ;
        RECT 81.585 197.575 81.915 198.555 ;
        RECT 82.085 197.405 82.365 198.545 ;
        RECT 83.120 198.505 83.290 198.650 ;
        RECT 82.625 198.335 83.290 198.505 ;
        RECT 83.575 198.480 83.745 199.280 ;
        RECT 83.955 199.135 84.185 199.955 ;
        RECT 84.355 199.155 84.685 199.785 ;
        RECT 83.935 198.715 84.265 198.965 ;
        RECT 84.435 198.555 84.685 199.155 ;
        RECT 84.855 199.135 85.065 199.955 ;
        RECT 85.355 199.135 85.565 199.955 ;
        RECT 85.735 199.155 86.065 199.785 ;
        RECT 82.625 197.575 82.795 198.335 ;
        RECT 82.975 197.405 83.305 198.165 ;
        RECT 83.475 197.575 83.745 198.480 ;
        RECT 83.955 197.405 84.185 198.545 ;
        RECT 84.355 197.575 84.685 198.555 ;
        RECT 85.735 198.555 85.985 199.155 ;
        RECT 86.235 199.135 86.465 199.955 ;
        RECT 86.675 199.185 88.345 199.955 ;
        RECT 88.515 199.230 88.805 199.955 ;
        RECT 89.435 199.185 91.105 199.955 ;
        RECT 91.280 199.410 96.625 199.955 ;
        RECT 86.155 198.715 86.485 198.965 ;
        RECT 84.855 197.405 85.065 198.545 ;
        RECT 85.355 197.405 85.565 198.545 ;
        RECT 85.735 197.575 86.065 198.555 ;
        RECT 86.235 197.405 86.465 198.545 ;
        RECT 86.675 198.495 87.425 199.015 ;
        RECT 87.595 198.665 88.345 199.185 ;
        RECT 86.675 197.405 88.345 198.495 ;
        RECT 88.515 197.405 88.805 198.570 ;
        RECT 89.435 198.495 90.185 199.015 ;
        RECT 90.355 198.665 91.105 199.185 ;
        RECT 89.435 197.405 91.105 198.495 ;
        RECT 92.870 197.840 93.220 199.090 ;
        RECT 94.700 198.580 95.040 199.410 ;
        RECT 96.800 199.245 97.055 199.775 ;
        RECT 97.225 199.495 97.530 199.955 ;
        RECT 97.775 199.575 98.845 199.745 ;
        RECT 96.800 198.595 97.010 199.245 ;
        RECT 97.775 199.220 98.095 199.575 ;
        RECT 97.770 199.045 98.095 199.220 ;
        RECT 97.180 198.745 98.095 199.045 ;
        RECT 98.265 199.005 98.505 199.405 ;
        RECT 98.675 199.345 98.845 199.575 ;
        RECT 99.015 199.515 99.205 199.955 ;
        RECT 99.375 199.505 100.325 199.785 ;
        RECT 100.545 199.595 100.895 199.765 ;
        RECT 98.675 199.175 99.205 199.345 ;
        RECT 97.180 198.715 97.920 198.745 ;
        RECT 91.280 197.405 96.625 197.840 ;
        RECT 96.800 197.715 97.055 198.595 ;
        RECT 97.225 197.405 97.530 198.545 ;
        RECT 97.750 198.125 97.920 198.715 ;
        RECT 98.265 198.635 98.805 199.005 ;
        RECT 98.985 198.895 99.205 199.175 ;
        RECT 99.375 198.725 99.545 199.505 ;
        RECT 99.140 198.555 99.545 198.725 ;
        RECT 99.715 198.715 100.065 199.335 ;
        RECT 99.140 198.465 99.310 198.555 ;
        RECT 100.235 198.545 100.445 199.335 ;
        RECT 98.090 198.295 99.310 198.465 ;
        RECT 99.770 198.385 100.445 198.545 ;
        RECT 97.750 197.955 98.550 198.125 ;
        RECT 97.870 197.405 98.200 197.785 ;
        RECT 98.380 197.665 98.550 197.955 ;
        RECT 99.140 197.915 99.310 198.295 ;
        RECT 99.480 198.375 100.445 198.385 ;
        RECT 100.635 199.205 100.895 199.595 ;
        RECT 101.105 199.495 101.435 199.955 ;
        RECT 102.310 199.565 103.165 199.735 ;
        RECT 103.370 199.565 103.865 199.735 ;
        RECT 104.035 199.595 104.365 199.955 ;
        RECT 100.635 198.515 100.805 199.205 ;
        RECT 100.975 198.855 101.145 199.035 ;
        RECT 101.315 199.025 102.105 199.275 ;
        RECT 102.310 198.855 102.480 199.565 ;
        RECT 102.650 199.055 103.005 199.275 ;
        RECT 100.975 198.685 102.665 198.855 ;
        RECT 99.480 198.085 99.940 198.375 ;
        RECT 100.635 198.345 102.135 198.515 ;
        RECT 100.635 198.205 100.805 198.345 ;
        RECT 100.245 198.035 100.805 198.205 ;
        RECT 98.720 197.405 98.970 197.865 ;
        RECT 99.140 197.575 100.010 197.915 ;
        RECT 100.245 197.575 100.415 198.035 ;
        RECT 101.250 198.005 102.325 198.175 ;
        RECT 100.585 197.405 100.955 197.865 ;
        RECT 101.250 197.665 101.420 198.005 ;
        RECT 101.590 197.405 101.920 197.835 ;
        RECT 102.155 197.665 102.325 198.005 ;
        RECT 102.495 197.905 102.665 198.685 ;
        RECT 102.835 198.465 103.005 199.055 ;
        RECT 103.175 198.655 103.525 199.275 ;
        RECT 102.835 198.075 103.300 198.465 ;
        RECT 103.695 198.205 103.865 199.565 ;
        RECT 104.035 198.375 104.495 199.425 ;
        RECT 103.470 198.035 103.865 198.205 ;
        RECT 103.470 197.905 103.640 198.035 ;
        RECT 102.495 197.575 103.175 197.905 ;
        RECT 103.390 197.575 103.640 197.905 ;
        RECT 103.810 197.405 104.060 197.865 ;
        RECT 104.230 197.590 104.555 198.375 ;
        RECT 104.725 197.575 104.895 199.695 ;
        RECT 105.065 199.575 105.395 199.955 ;
        RECT 105.565 199.405 105.820 199.695 ;
        RECT 105.070 199.235 105.820 199.405 ;
        RECT 105.070 198.245 105.300 199.235 ;
        RECT 105.995 199.185 108.585 199.955 ;
        RECT 108.760 199.410 114.105 199.955 ;
        RECT 105.470 198.415 105.820 199.065 ;
        RECT 105.995 198.495 107.205 199.015 ;
        RECT 107.375 198.665 108.585 199.185 ;
        RECT 105.070 198.075 105.820 198.245 ;
        RECT 105.065 197.405 105.395 197.905 ;
        RECT 105.565 197.575 105.820 198.075 ;
        RECT 105.995 197.405 108.585 198.495 ;
        RECT 110.350 197.840 110.700 199.090 ;
        RECT 112.180 198.580 112.520 199.410 ;
        RECT 114.275 199.230 114.565 199.955 ;
        RECT 115.200 199.410 120.545 199.955 ;
        RECT 120.720 199.410 126.065 199.955 ;
        RECT 108.760 197.405 114.105 197.840 ;
        RECT 114.275 197.405 114.565 198.570 ;
        RECT 116.790 197.840 117.140 199.090 ;
        RECT 118.620 198.580 118.960 199.410 ;
        RECT 122.310 197.840 122.660 199.090 ;
        RECT 124.140 198.580 124.480 199.410 ;
        RECT 126.235 199.205 127.445 199.955 ;
        RECT 126.235 198.495 126.755 199.035 ;
        RECT 126.925 198.665 127.445 199.205 ;
        RECT 115.200 197.405 120.545 197.840 ;
        RECT 120.720 197.405 126.065 197.840 ;
        RECT 126.235 197.405 127.445 198.495 ;
        RECT 14.370 197.235 127.530 197.405 ;
        RECT 14.455 196.145 15.665 197.235 ;
        RECT 14.455 195.435 14.975 195.975 ;
        RECT 15.145 195.605 15.665 196.145 ;
        RECT 15.835 196.145 18.425 197.235 ;
        RECT 18.600 196.800 23.945 197.235 ;
        RECT 15.835 195.625 17.045 196.145 ;
        RECT 17.215 195.455 18.425 195.975 ;
        RECT 20.190 195.550 20.540 196.800 ;
        RECT 24.115 196.070 24.405 197.235 ;
        RECT 25.035 196.145 27.625 197.235 ;
        RECT 27.800 196.800 33.145 197.235 ;
        RECT 33.320 196.800 38.665 197.235 ;
        RECT 38.840 196.800 44.185 197.235 ;
        RECT 44.360 196.800 49.705 197.235 ;
        RECT 14.455 194.685 15.665 195.435 ;
        RECT 15.835 194.685 18.425 195.455 ;
        RECT 22.020 195.230 22.360 196.060 ;
        RECT 25.035 195.625 26.245 196.145 ;
        RECT 26.415 195.455 27.625 195.975 ;
        RECT 29.390 195.550 29.740 196.800 ;
        RECT 18.600 194.685 23.945 195.230 ;
        RECT 24.115 194.685 24.405 195.410 ;
        RECT 25.035 194.685 27.625 195.455 ;
        RECT 31.220 195.230 31.560 196.060 ;
        RECT 34.910 195.550 35.260 196.800 ;
        RECT 36.740 195.230 37.080 196.060 ;
        RECT 40.430 195.550 40.780 196.800 ;
        RECT 42.260 195.230 42.600 196.060 ;
        RECT 45.950 195.550 46.300 196.800 ;
        RECT 49.875 196.070 50.165 197.235 ;
        RECT 50.795 196.145 52.465 197.235 ;
        RECT 47.780 195.230 48.120 196.060 ;
        RECT 50.795 195.625 51.545 196.145 ;
        RECT 52.695 196.095 52.905 197.235 ;
        RECT 53.075 196.085 53.405 197.065 ;
        RECT 53.575 196.095 53.805 197.235 ;
        RECT 54.130 196.605 54.415 197.065 ;
        RECT 54.585 196.775 54.855 197.235 ;
        RECT 54.130 196.385 55.085 196.605 ;
        RECT 51.715 195.455 52.465 195.975 ;
        RECT 27.800 194.685 33.145 195.230 ;
        RECT 33.320 194.685 38.665 195.230 ;
        RECT 38.840 194.685 44.185 195.230 ;
        RECT 44.360 194.685 49.705 195.230 ;
        RECT 49.875 194.685 50.165 195.410 ;
        RECT 50.795 194.685 52.465 195.455 ;
        RECT 52.695 194.685 52.905 195.505 ;
        RECT 53.075 195.485 53.325 196.085 ;
        RECT 53.495 195.675 53.825 195.925 ;
        RECT 54.015 195.655 54.705 196.215 ;
        RECT 53.075 194.855 53.405 195.485 ;
        RECT 53.575 194.685 53.805 195.505 ;
        RECT 54.875 195.485 55.085 196.385 ;
        RECT 54.130 195.315 55.085 195.485 ;
        RECT 55.255 196.215 55.655 197.065 ;
        RECT 55.845 196.605 56.125 197.065 ;
        RECT 56.645 196.775 56.970 197.235 ;
        RECT 55.845 196.385 56.970 196.605 ;
        RECT 55.255 195.655 56.350 196.215 ;
        RECT 56.520 195.925 56.970 196.385 ;
        RECT 57.140 196.095 57.525 197.065 ;
        RECT 57.700 196.800 63.045 197.235 ;
        RECT 63.220 196.800 68.565 197.235 ;
        RECT 54.130 194.855 54.415 195.315 ;
        RECT 54.585 194.685 54.855 195.145 ;
        RECT 55.255 194.855 55.655 195.655 ;
        RECT 56.520 195.595 57.075 195.925 ;
        RECT 56.520 195.485 56.970 195.595 ;
        RECT 55.845 195.315 56.970 195.485 ;
        RECT 57.245 195.425 57.525 196.095 ;
        RECT 59.290 195.550 59.640 196.800 ;
        RECT 55.845 194.855 56.125 195.315 ;
        RECT 56.645 194.685 56.970 195.145 ;
        RECT 57.140 194.855 57.525 195.425 ;
        RECT 61.120 195.230 61.460 196.060 ;
        RECT 64.810 195.550 65.160 196.800 ;
        RECT 68.735 196.365 69.010 197.065 ;
        RECT 69.180 196.690 69.435 197.235 ;
        RECT 69.605 196.725 70.085 197.065 ;
        RECT 70.260 196.680 70.865 197.235 ;
        RECT 70.250 196.580 70.865 196.680 ;
        RECT 70.250 196.555 70.435 196.580 ;
        RECT 66.640 195.230 66.980 196.060 ;
        RECT 68.735 195.335 68.905 196.365 ;
        RECT 69.180 196.235 69.935 196.485 ;
        RECT 70.105 196.310 70.435 196.555 ;
        RECT 69.180 196.200 69.950 196.235 ;
        RECT 69.180 196.190 69.965 196.200 ;
        RECT 69.075 196.175 69.970 196.190 ;
        RECT 69.075 196.160 69.990 196.175 ;
        RECT 69.075 196.150 70.010 196.160 ;
        RECT 69.075 196.140 70.035 196.150 ;
        RECT 69.075 196.110 70.105 196.140 ;
        RECT 69.075 196.080 70.125 196.110 ;
        RECT 69.075 196.050 70.145 196.080 ;
        RECT 69.075 196.025 70.175 196.050 ;
        RECT 69.075 195.990 70.210 196.025 ;
        RECT 69.075 195.985 70.240 195.990 ;
        RECT 69.075 195.590 69.305 195.985 ;
        RECT 69.850 195.980 70.240 195.985 ;
        RECT 69.875 195.970 70.240 195.980 ;
        RECT 69.890 195.965 70.240 195.970 ;
        RECT 69.905 195.960 70.240 195.965 ;
        RECT 70.605 195.960 70.865 196.410 ;
        RECT 69.905 195.955 70.865 195.960 ;
        RECT 69.915 195.945 70.865 195.955 ;
        RECT 69.925 195.940 70.865 195.945 ;
        RECT 69.935 195.930 70.865 195.940 ;
        RECT 69.940 195.920 70.865 195.930 ;
        RECT 69.945 195.915 70.865 195.920 ;
        RECT 69.955 195.900 70.865 195.915 ;
        RECT 69.960 195.885 70.865 195.900 ;
        RECT 69.970 195.860 70.865 195.885 ;
        RECT 69.475 195.390 69.805 195.815 ;
        RECT 57.700 194.685 63.045 195.230 ;
        RECT 63.220 194.685 68.565 195.230 ;
        RECT 68.735 194.855 68.995 195.335 ;
        RECT 69.165 194.685 69.415 195.225 ;
        RECT 69.585 194.905 69.805 195.390 ;
        RECT 69.975 195.790 70.865 195.860 ;
        RECT 71.045 196.175 71.375 197.025 ;
        RECT 69.975 195.065 70.145 195.790 ;
        RECT 70.315 195.235 70.865 195.620 ;
        RECT 71.045 195.410 71.235 196.175 ;
        RECT 71.545 196.095 71.795 197.235 ;
        RECT 71.985 196.595 72.235 197.015 ;
        RECT 72.465 196.765 72.795 197.235 ;
        RECT 73.025 196.595 73.275 197.015 ;
        RECT 71.985 196.425 73.275 196.595 ;
        RECT 73.455 196.595 73.785 197.025 ;
        RECT 73.455 196.425 73.910 196.595 ;
        RECT 71.975 195.925 72.190 196.255 ;
        RECT 71.405 195.595 71.715 195.925 ;
        RECT 71.885 195.595 72.190 195.925 ;
        RECT 72.365 195.595 72.650 196.255 ;
        RECT 72.845 195.595 73.110 196.255 ;
        RECT 73.325 195.595 73.570 196.255 ;
        RECT 71.545 195.425 71.715 195.595 ;
        RECT 73.740 195.425 73.910 196.425 ;
        RECT 74.255 196.145 75.465 197.235 ;
        RECT 74.255 195.605 74.775 196.145 ;
        RECT 75.635 196.070 75.925 197.235 ;
        RECT 76.095 196.145 79.605 197.235 ;
        RECT 79.780 196.800 85.125 197.235 ;
        RECT 74.945 195.435 75.465 195.975 ;
        RECT 76.095 195.625 77.785 196.145 ;
        RECT 77.955 195.455 79.605 195.975 ;
        RECT 81.370 195.550 81.720 196.800 ;
        RECT 85.670 196.255 85.925 196.925 ;
        RECT 86.105 196.435 86.390 197.235 ;
        RECT 86.570 196.515 86.900 197.025 ;
        RECT 69.975 194.895 70.865 195.065 ;
        RECT 71.045 194.900 71.375 195.410 ;
        RECT 71.545 195.255 73.910 195.425 ;
        RECT 71.545 194.685 71.875 195.085 ;
        RECT 72.925 194.915 73.255 195.255 ;
        RECT 73.425 194.685 73.755 195.085 ;
        RECT 74.255 194.685 75.465 195.435 ;
        RECT 75.635 194.685 75.925 195.410 ;
        RECT 76.095 194.685 79.605 195.455 ;
        RECT 83.200 195.230 83.540 196.060 ;
        RECT 85.670 195.395 85.850 196.255 ;
        RECT 86.570 195.925 86.820 196.515 ;
        RECT 87.170 196.365 87.340 196.975 ;
        RECT 87.510 196.545 87.840 197.235 ;
        RECT 88.070 196.685 88.310 196.975 ;
        RECT 88.510 196.855 88.930 197.235 ;
        RECT 89.110 196.765 89.740 197.015 ;
        RECT 90.210 196.855 90.540 197.235 ;
        RECT 89.110 196.685 89.280 196.765 ;
        RECT 90.710 196.685 90.880 196.975 ;
        RECT 91.060 196.855 91.440 197.235 ;
        RECT 91.680 196.850 92.510 197.020 ;
        RECT 88.070 196.515 89.280 196.685 ;
        RECT 86.020 195.595 86.820 195.925 ;
        RECT 79.780 194.685 85.125 195.230 ;
        RECT 85.670 195.195 85.925 195.395 ;
        RECT 85.585 195.025 85.925 195.195 ;
        RECT 85.670 194.865 85.925 195.025 ;
        RECT 86.105 194.685 86.390 195.145 ;
        RECT 86.570 194.945 86.820 195.595 ;
        RECT 87.020 196.345 87.340 196.365 ;
        RECT 87.020 196.175 88.940 196.345 ;
        RECT 87.020 195.280 87.210 196.175 ;
        RECT 89.110 196.005 89.280 196.515 ;
        RECT 89.450 196.255 89.970 196.565 ;
        RECT 87.380 195.835 89.280 196.005 ;
        RECT 87.380 195.775 87.710 195.835 ;
        RECT 87.860 195.605 88.190 195.665 ;
        RECT 87.530 195.335 88.190 195.605 ;
        RECT 87.020 194.950 87.340 195.280 ;
        RECT 87.520 194.685 88.180 195.165 ;
        RECT 88.380 195.075 88.550 195.835 ;
        RECT 89.450 195.665 89.630 196.075 ;
        RECT 88.720 195.495 89.050 195.615 ;
        RECT 89.800 195.495 89.970 196.255 ;
        RECT 88.720 195.325 89.970 195.495 ;
        RECT 90.140 196.435 91.510 196.685 ;
        RECT 90.140 195.665 90.330 196.435 ;
        RECT 91.260 196.175 91.510 196.435 ;
        RECT 90.500 196.005 90.750 196.165 ;
        RECT 91.680 196.005 91.850 196.850 ;
        RECT 92.745 196.565 92.915 197.065 ;
        RECT 93.085 196.735 93.415 197.235 ;
        RECT 92.020 196.175 92.520 196.555 ;
        RECT 92.745 196.395 93.440 196.565 ;
        RECT 90.500 195.835 91.850 196.005 ;
        RECT 91.430 195.795 91.850 195.835 ;
        RECT 90.140 195.325 90.560 195.665 ;
        RECT 90.850 195.335 91.260 195.665 ;
        RECT 88.380 194.905 89.230 195.075 ;
        RECT 89.790 194.685 90.110 195.145 ;
        RECT 90.310 194.895 90.560 195.325 ;
        RECT 90.850 194.685 91.260 195.125 ;
        RECT 91.430 195.065 91.600 195.795 ;
        RECT 91.770 195.245 92.120 195.615 ;
        RECT 92.300 195.305 92.520 196.175 ;
        RECT 92.690 195.605 93.100 196.225 ;
        RECT 93.270 195.425 93.440 196.395 ;
        RECT 92.745 195.235 93.440 195.425 ;
        RECT 91.430 194.865 92.445 195.065 ;
        RECT 92.745 194.905 92.915 195.235 ;
        RECT 93.085 194.685 93.415 195.065 ;
        RECT 93.630 194.945 93.855 197.065 ;
        RECT 94.025 196.735 94.355 197.235 ;
        RECT 94.525 196.565 94.695 197.065 ;
        RECT 94.030 196.395 94.695 196.565 ;
        RECT 94.030 195.405 94.260 196.395 ;
        RECT 94.430 195.575 94.780 196.225 ;
        RECT 94.955 196.145 97.545 197.235 ;
        RECT 97.830 196.605 98.115 197.065 ;
        RECT 98.285 196.775 98.555 197.235 ;
        RECT 97.830 196.385 98.785 196.605 ;
        RECT 94.955 195.625 96.165 196.145 ;
        RECT 96.335 195.455 97.545 195.975 ;
        RECT 97.715 195.655 98.405 196.215 ;
        RECT 98.575 195.485 98.785 196.385 ;
        RECT 94.030 195.235 94.695 195.405 ;
        RECT 94.025 194.685 94.355 195.065 ;
        RECT 94.525 194.945 94.695 195.235 ;
        RECT 94.955 194.685 97.545 195.455 ;
        RECT 97.830 195.315 98.785 195.485 ;
        RECT 98.955 196.215 99.355 197.065 ;
        RECT 99.545 196.605 99.825 197.065 ;
        RECT 100.345 196.775 100.670 197.235 ;
        RECT 99.545 196.385 100.670 196.605 ;
        RECT 98.955 195.655 100.050 196.215 ;
        RECT 100.220 195.925 100.670 196.385 ;
        RECT 100.840 196.095 101.225 197.065 ;
        RECT 97.830 194.855 98.115 195.315 ;
        RECT 98.285 194.685 98.555 195.145 ;
        RECT 98.955 194.855 99.355 195.655 ;
        RECT 100.220 195.595 100.775 195.925 ;
        RECT 100.220 195.485 100.670 195.595 ;
        RECT 99.545 195.315 100.670 195.485 ;
        RECT 100.945 195.425 101.225 196.095 ;
        RECT 101.395 196.070 101.685 197.235 ;
        RECT 101.855 196.145 104.445 197.235 ;
        RECT 104.620 196.800 109.965 197.235 ;
        RECT 101.855 195.625 103.065 196.145 ;
        RECT 103.235 195.455 104.445 195.975 ;
        RECT 106.210 195.550 106.560 196.800 ;
        RECT 99.545 194.855 99.825 195.315 ;
        RECT 100.345 194.685 100.670 195.145 ;
        RECT 100.840 194.855 101.225 195.425 ;
        RECT 101.395 194.685 101.685 195.410 ;
        RECT 101.855 194.685 104.445 195.455 ;
        RECT 108.040 195.230 108.380 196.060 ;
        RECT 110.140 196.045 110.395 196.925 ;
        RECT 110.565 196.095 110.870 197.235 ;
        RECT 111.210 196.855 111.540 197.235 ;
        RECT 111.720 196.685 111.890 196.975 ;
        RECT 112.060 196.775 112.310 197.235 ;
        RECT 111.090 196.515 111.890 196.685 ;
        RECT 112.480 196.725 113.350 197.065 ;
        RECT 110.140 195.395 110.350 196.045 ;
        RECT 111.090 195.925 111.260 196.515 ;
        RECT 112.480 196.345 112.650 196.725 ;
        RECT 113.585 196.605 113.755 197.065 ;
        RECT 113.925 196.775 114.295 197.235 ;
        RECT 114.590 196.635 114.760 196.975 ;
        RECT 114.930 196.805 115.260 197.235 ;
        RECT 115.495 196.635 115.665 196.975 ;
        RECT 111.430 196.175 112.650 196.345 ;
        RECT 112.820 196.265 113.280 196.555 ;
        RECT 113.585 196.435 114.145 196.605 ;
        RECT 114.590 196.465 115.665 196.635 ;
        RECT 115.835 196.735 116.515 197.065 ;
        RECT 116.730 196.735 116.980 197.065 ;
        RECT 117.150 196.775 117.400 197.235 ;
        RECT 113.975 196.295 114.145 196.435 ;
        RECT 112.820 196.255 113.785 196.265 ;
        RECT 112.480 196.085 112.650 196.175 ;
        RECT 113.110 196.095 113.785 196.255 ;
        RECT 110.520 195.895 111.260 195.925 ;
        RECT 110.520 195.595 111.435 195.895 ;
        RECT 111.110 195.420 111.435 195.595 ;
        RECT 104.620 194.685 109.965 195.230 ;
        RECT 110.140 194.865 110.395 195.395 ;
        RECT 110.565 194.685 110.870 195.145 ;
        RECT 111.115 195.065 111.435 195.420 ;
        RECT 111.605 195.635 112.145 196.005 ;
        RECT 112.480 195.915 112.885 196.085 ;
        RECT 111.605 195.235 111.845 195.635 ;
        RECT 112.325 195.465 112.545 195.745 ;
        RECT 112.015 195.295 112.545 195.465 ;
        RECT 112.015 195.065 112.185 195.295 ;
        RECT 112.715 195.135 112.885 195.915 ;
        RECT 113.055 195.305 113.405 195.925 ;
        RECT 113.575 195.305 113.785 196.095 ;
        RECT 113.975 196.125 115.475 196.295 ;
        RECT 113.975 195.435 114.145 196.125 ;
        RECT 115.835 195.955 116.005 196.735 ;
        RECT 116.810 196.605 116.980 196.735 ;
        RECT 114.315 195.785 116.005 195.955 ;
        RECT 116.175 196.175 116.640 196.565 ;
        RECT 116.810 196.435 117.205 196.605 ;
        RECT 114.315 195.605 114.485 195.785 ;
        RECT 111.115 194.895 112.185 195.065 ;
        RECT 112.355 194.685 112.545 195.125 ;
        RECT 112.715 194.855 113.665 195.135 ;
        RECT 113.975 195.045 114.235 195.435 ;
        RECT 114.655 195.365 115.445 195.615 ;
        RECT 113.885 194.875 114.235 195.045 ;
        RECT 114.445 194.685 114.775 195.145 ;
        RECT 115.650 195.075 115.820 195.785 ;
        RECT 116.175 195.585 116.345 196.175 ;
        RECT 115.990 195.365 116.345 195.585 ;
        RECT 116.515 195.365 116.865 195.985 ;
        RECT 117.035 195.075 117.205 196.435 ;
        RECT 117.570 196.265 117.895 197.050 ;
        RECT 117.375 195.215 117.835 196.265 ;
        RECT 115.650 194.905 116.505 195.075 ;
        RECT 116.710 194.905 117.205 195.075 ;
        RECT 117.375 194.685 117.705 195.045 ;
        RECT 118.065 194.945 118.235 197.065 ;
        RECT 118.405 196.735 118.735 197.235 ;
        RECT 118.905 196.565 119.160 197.065 ;
        RECT 118.410 196.395 119.160 196.565 ;
        RECT 118.410 195.405 118.640 196.395 ;
        RECT 118.810 195.575 119.160 196.225 ;
        RECT 119.335 196.145 120.545 197.235 ;
        RECT 120.720 196.800 126.065 197.235 ;
        RECT 119.335 195.605 119.855 196.145 ;
        RECT 120.025 195.435 120.545 195.975 ;
        RECT 122.310 195.550 122.660 196.800 ;
        RECT 126.235 196.145 127.445 197.235 ;
        RECT 118.410 195.235 119.160 195.405 ;
        RECT 118.405 194.685 118.735 195.065 ;
        RECT 118.905 194.945 119.160 195.235 ;
        RECT 119.335 194.685 120.545 195.435 ;
        RECT 124.140 195.230 124.480 196.060 ;
        RECT 126.235 195.605 126.755 196.145 ;
        RECT 126.925 195.435 127.445 195.975 ;
        RECT 120.720 194.685 126.065 195.230 ;
        RECT 126.235 194.685 127.445 195.435 ;
        RECT 14.370 194.515 127.530 194.685 ;
        RECT 14.455 193.765 15.665 194.515 ;
        RECT 14.455 193.225 14.975 193.765 ;
        RECT 16.755 193.745 20.265 194.515 ;
        RECT 20.440 193.970 25.785 194.515 ;
        RECT 25.960 193.970 31.305 194.515 ;
        RECT 31.480 193.970 36.825 194.515 ;
        RECT 15.145 193.055 15.665 193.595 ;
        RECT 14.455 191.965 15.665 193.055 ;
        RECT 16.755 193.055 18.445 193.575 ;
        RECT 18.615 193.225 20.265 193.745 ;
        RECT 16.755 191.965 20.265 193.055 ;
        RECT 22.030 192.400 22.380 193.650 ;
        RECT 23.860 193.140 24.200 193.970 ;
        RECT 27.550 192.400 27.900 193.650 ;
        RECT 29.380 193.140 29.720 193.970 ;
        RECT 33.070 192.400 33.420 193.650 ;
        RECT 34.900 193.140 35.240 193.970 ;
        RECT 36.995 193.790 37.285 194.515 ;
        RECT 38.375 193.745 41.885 194.515 ;
        RECT 42.060 193.970 47.405 194.515 ;
        RECT 20.440 191.965 25.785 192.400 ;
        RECT 25.960 191.965 31.305 192.400 ;
        RECT 31.480 191.965 36.825 192.400 ;
        RECT 36.995 191.965 37.285 193.130 ;
        RECT 38.375 193.055 40.065 193.575 ;
        RECT 40.235 193.225 41.885 193.745 ;
        RECT 38.375 191.965 41.885 193.055 ;
        RECT 43.650 192.400 44.000 193.650 ;
        RECT 45.480 193.140 45.820 193.970 ;
        RECT 47.635 193.695 47.845 194.515 ;
        RECT 48.015 193.715 48.345 194.345 ;
        RECT 48.015 193.115 48.265 193.715 ;
        RECT 48.515 193.695 48.745 194.515 ;
        RECT 48.960 193.965 49.215 194.255 ;
        RECT 49.385 194.135 49.715 194.515 ;
        RECT 48.960 193.795 49.710 193.965 ;
        RECT 48.435 193.275 48.765 193.525 ;
        RECT 42.060 191.965 47.405 192.400 ;
        RECT 47.635 191.965 47.845 193.105 ;
        RECT 48.015 192.135 48.345 193.115 ;
        RECT 48.515 191.965 48.745 193.105 ;
        RECT 48.960 192.975 49.310 193.625 ;
        RECT 49.480 192.805 49.710 193.795 ;
        RECT 48.960 192.635 49.710 192.805 ;
        RECT 48.960 192.135 49.215 192.635 ;
        RECT 49.385 191.965 49.715 192.465 ;
        RECT 49.885 192.135 50.055 194.255 ;
        RECT 50.415 194.155 50.745 194.515 ;
        RECT 50.915 194.125 51.410 194.295 ;
        RECT 51.615 194.125 52.470 194.295 ;
        RECT 50.285 192.935 50.745 193.985 ;
        RECT 50.225 192.150 50.550 192.935 ;
        RECT 50.915 192.765 51.085 194.125 ;
        RECT 51.255 193.215 51.605 193.835 ;
        RECT 51.775 193.615 52.130 193.835 ;
        RECT 51.775 193.025 51.945 193.615 ;
        RECT 52.300 193.415 52.470 194.125 ;
        RECT 53.345 194.055 53.675 194.515 ;
        RECT 53.885 194.155 54.235 194.325 ;
        RECT 52.675 193.585 53.465 193.835 ;
        RECT 53.885 193.765 54.145 194.155 ;
        RECT 54.455 194.065 55.405 194.345 ;
        RECT 55.575 194.075 55.765 194.515 ;
        RECT 55.935 194.135 57.005 194.305 ;
        RECT 53.635 193.415 53.805 193.595 ;
        RECT 50.915 192.595 51.310 192.765 ;
        RECT 51.480 192.635 51.945 193.025 ;
        RECT 52.115 193.245 53.805 193.415 ;
        RECT 51.140 192.465 51.310 192.595 ;
        RECT 52.115 192.465 52.285 193.245 ;
        RECT 53.975 193.075 54.145 193.765 ;
        RECT 52.645 192.905 54.145 193.075 ;
        RECT 54.335 193.105 54.545 193.895 ;
        RECT 54.715 193.275 55.065 193.895 ;
        RECT 55.235 193.285 55.405 194.065 ;
        RECT 55.935 193.905 56.105 194.135 ;
        RECT 55.575 193.735 56.105 193.905 ;
        RECT 55.575 193.455 55.795 193.735 ;
        RECT 56.275 193.565 56.515 193.965 ;
        RECT 55.235 193.115 55.640 193.285 ;
        RECT 55.975 193.195 56.515 193.565 ;
        RECT 56.685 193.780 57.005 194.135 ;
        RECT 57.250 194.055 57.555 194.515 ;
        RECT 57.725 193.805 57.980 194.335 ;
        RECT 56.685 193.605 57.010 193.780 ;
        RECT 56.685 193.305 57.600 193.605 ;
        RECT 56.860 193.275 57.600 193.305 ;
        RECT 54.335 192.945 55.010 193.105 ;
        RECT 55.470 193.025 55.640 193.115 ;
        RECT 54.335 192.935 55.300 192.945 ;
        RECT 53.975 192.765 54.145 192.905 ;
        RECT 50.720 191.965 50.970 192.425 ;
        RECT 51.140 192.135 51.390 192.465 ;
        RECT 51.605 192.135 52.285 192.465 ;
        RECT 52.455 192.565 53.530 192.735 ;
        RECT 53.975 192.595 54.535 192.765 ;
        RECT 54.840 192.645 55.300 192.935 ;
        RECT 55.470 192.855 56.690 193.025 ;
        RECT 52.455 192.225 52.625 192.565 ;
        RECT 52.860 191.965 53.190 192.395 ;
        RECT 53.360 192.225 53.530 192.565 ;
        RECT 53.825 191.965 54.195 192.425 ;
        RECT 54.365 192.135 54.535 192.595 ;
        RECT 55.470 192.475 55.640 192.855 ;
        RECT 56.860 192.685 57.030 193.275 ;
        RECT 57.770 193.155 57.980 193.805 ;
        RECT 59.075 193.745 62.585 194.515 ;
        RECT 62.755 193.790 63.045 194.515 ;
        RECT 63.215 193.745 64.885 194.515 ;
        RECT 54.770 192.135 55.640 192.475 ;
        RECT 56.230 192.515 57.030 192.685 ;
        RECT 55.810 191.965 56.060 192.425 ;
        RECT 56.230 192.225 56.400 192.515 ;
        RECT 56.580 191.965 56.910 192.345 ;
        RECT 57.250 191.965 57.555 193.105 ;
        RECT 57.725 192.275 57.980 193.155 ;
        RECT 59.075 193.055 60.765 193.575 ;
        RECT 60.935 193.225 62.585 193.745 ;
        RECT 59.075 191.965 62.585 193.055 ;
        RECT 62.755 191.965 63.045 193.130 ;
        RECT 63.215 193.055 63.965 193.575 ;
        RECT 64.135 193.225 64.885 193.745 ;
        RECT 65.115 193.695 65.325 194.515 ;
        RECT 65.495 193.715 65.825 194.345 ;
        RECT 65.495 193.115 65.745 193.715 ;
        RECT 65.995 193.695 66.225 194.515 ;
        RECT 66.895 193.745 68.565 194.515 ;
        RECT 65.915 193.275 66.245 193.525 ;
        RECT 63.215 191.965 64.885 193.055 ;
        RECT 65.115 191.965 65.325 193.105 ;
        RECT 65.495 192.135 65.825 193.115 ;
        RECT 65.995 191.965 66.225 193.105 ;
        RECT 66.895 193.055 67.645 193.575 ;
        RECT 67.815 193.225 68.565 193.745 ;
        RECT 68.735 193.695 68.995 194.515 ;
        RECT 69.165 193.695 69.495 194.115 ;
        RECT 69.675 193.945 69.935 194.345 ;
        RECT 70.105 194.115 70.435 194.515 ;
        RECT 70.605 193.945 70.775 194.295 ;
        RECT 70.945 194.115 71.320 194.515 ;
        RECT 69.675 193.775 71.340 193.945 ;
        RECT 71.510 193.840 71.785 194.185 ;
        RECT 69.245 193.605 69.495 193.695 ;
        RECT 71.170 193.605 71.340 193.775 ;
        RECT 68.740 193.275 69.075 193.525 ;
        RECT 69.245 193.275 69.960 193.605 ;
        RECT 70.175 193.275 71.000 193.605 ;
        RECT 71.170 193.275 71.445 193.605 ;
        RECT 66.895 191.965 68.565 193.055 ;
        RECT 68.735 191.965 68.995 193.105 ;
        RECT 69.245 192.715 69.415 193.275 ;
        RECT 69.675 192.815 70.005 193.105 ;
        RECT 70.175 192.985 70.420 193.275 ;
        RECT 71.170 193.105 71.340 193.275 ;
        RECT 71.615 193.105 71.785 193.840 ;
        RECT 70.680 192.935 71.340 193.105 ;
        RECT 70.680 192.815 70.850 192.935 ;
        RECT 69.675 192.645 70.850 192.815 ;
        RECT 69.235 192.145 70.850 192.475 ;
        RECT 71.020 191.965 71.300 192.765 ;
        RECT 71.510 192.135 71.785 193.105 ;
        RECT 71.955 193.840 72.230 194.185 ;
        RECT 72.420 194.115 72.795 194.515 ;
        RECT 72.965 193.945 73.135 194.295 ;
        RECT 73.305 194.115 73.635 194.515 ;
        RECT 73.805 193.945 74.065 194.345 ;
        RECT 71.955 193.105 72.125 193.840 ;
        RECT 72.400 193.775 74.065 193.945 ;
        RECT 72.400 193.605 72.570 193.775 ;
        RECT 74.245 193.695 74.575 194.115 ;
        RECT 74.745 193.695 75.005 194.515 ;
        RECT 75.175 193.745 78.685 194.515 ;
        RECT 78.860 193.970 84.205 194.515 ;
        RECT 74.245 193.605 74.495 193.695 ;
        RECT 72.295 193.275 72.570 193.605 ;
        RECT 72.740 193.275 73.565 193.605 ;
        RECT 73.780 193.275 74.495 193.605 ;
        RECT 74.665 193.275 75.000 193.525 ;
        RECT 72.400 193.105 72.570 193.275 ;
        RECT 71.955 192.135 72.230 193.105 ;
        RECT 72.400 192.935 73.060 193.105 ;
        RECT 73.320 192.985 73.565 193.275 ;
        RECT 72.890 192.815 73.060 192.935 ;
        RECT 73.735 192.815 74.065 193.105 ;
        RECT 72.440 191.965 72.720 192.765 ;
        RECT 72.890 192.645 74.065 192.815 ;
        RECT 74.325 192.715 74.495 193.275 ;
        RECT 72.890 192.145 74.505 192.475 ;
        RECT 74.745 191.965 75.005 193.105 ;
        RECT 75.175 193.055 76.865 193.575 ;
        RECT 77.035 193.225 78.685 193.745 ;
        RECT 75.175 191.965 78.685 193.055 ;
        RECT 80.450 192.400 80.800 193.650 ;
        RECT 82.280 193.140 82.620 193.970 ;
        RECT 84.650 193.705 84.895 194.310 ;
        RECT 85.115 193.980 85.625 194.515 ;
        RECT 84.375 193.535 85.605 193.705 ;
        RECT 84.375 192.725 84.715 193.535 ;
        RECT 84.885 192.970 85.635 193.160 ;
        RECT 78.860 191.965 84.205 192.400 ;
        RECT 84.375 192.315 84.890 192.725 ;
        RECT 85.125 191.965 85.295 192.725 ;
        RECT 85.465 192.305 85.635 192.970 ;
        RECT 85.805 192.985 85.995 194.345 ;
        RECT 86.165 193.495 86.440 194.345 ;
        RECT 86.630 193.980 87.160 194.345 ;
        RECT 87.585 194.115 87.915 194.515 ;
        RECT 86.985 193.945 87.160 193.980 ;
        RECT 86.165 193.325 86.445 193.495 ;
        RECT 86.165 193.185 86.440 193.325 ;
        RECT 86.645 192.985 86.815 193.785 ;
        RECT 85.805 192.815 86.815 192.985 ;
        RECT 86.985 193.775 87.915 193.945 ;
        RECT 88.085 193.775 88.340 194.345 ;
        RECT 88.515 193.790 88.805 194.515 ;
        RECT 86.985 192.645 87.155 193.775 ;
        RECT 87.745 193.605 87.915 193.775 ;
        RECT 86.030 192.475 87.155 192.645 ;
        RECT 87.325 193.275 87.520 193.605 ;
        RECT 87.745 193.275 88.000 193.605 ;
        RECT 87.325 192.305 87.495 193.275 ;
        RECT 88.170 193.105 88.340 193.775 ;
        RECT 89.035 193.695 89.245 194.515 ;
        RECT 89.415 193.715 89.745 194.345 ;
        RECT 85.465 192.135 87.495 192.305 ;
        RECT 87.665 191.965 87.835 193.105 ;
        RECT 88.005 192.135 88.340 193.105 ;
        RECT 88.515 191.965 88.805 193.130 ;
        RECT 89.415 193.115 89.665 193.715 ;
        RECT 89.915 193.695 90.145 194.515 ;
        RECT 90.355 193.745 92.945 194.515 ;
        RECT 89.835 193.275 90.165 193.525 ;
        RECT 89.035 191.965 89.245 193.105 ;
        RECT 89.415 192.135 89.745 193.115 ;
        RECT 89.915 191.965 90.145 193.105 ;
        RECT 90.355 193.055 91.565 193.575 ;
        RECT 91.735 193.225 92.945 193.745 ;
        RECT 93.155 193.695 93.385 194.515 ;
        RECT 93.555 193.715 93.885 194.345 ;
        RECT 93.135 193.275 93.465 193.525 ;
        RECT 93.635 193.115 93.885 193.715 ;
        RECT 94.055 193.695 94.265 194.515 ;
        RECT 94.495 194.005 94.800 194.515 ;
        RECT 94.495 193.275 94.810 193.835 ;
        RECT 94.980 193.525 95.230 194.335 ;
        RECT 95.400 193.990 95.660 194.515 ;
        RECT 95.840 193.525 96.090 194.335 ;
        RECT 96.260 193.955 96.520 194.515 ;
        RECT 96.690 193.865 96.950 194.320 ;
        RECT 97.120 194.035 97.380 194.515 ;
        RECT 97.550 193.865 97.810 194.320 ;
        RECT 97.980 194.035 98.240 194.515 ;
        RECT 98.410 193.865 98.670 194.320 ;
        RECT 98.840 194.035 99.085 194.515 ;
        RECT 99.255 193.865 99.530 194.320 ;
        RECT 99.700 194.035 99.945 194.515 ;
        RECT 100.115 193.865 100.375 194.320 ;
        RECT 100.555 194.035 100.805 194.515 ;
        RECT 100.975 193.865 101.235 194.320 ;
        RECT 101.415 194.035 101.665 194.515 ;
        RECT 101.835 193.865 102.095 194.320 ;
        RECT 102.275 194.035 102.535 194.515 ;
        RECT 102.705 193.865 102.965 194.320 ;
        RECT 103.135 194.035 103.435 194.515 ;
        RECT 96.690 193.835 103.435 193.865 ;
        RECT 96.690 193.695 103.465 193.835 ;
        RECT 103.695 193.765 104.905 194.515 ;
        RECT 102.270 193.665 103.465 193.695 ;
        RECT 94.980 193.275 102.100 193.525 ;
        RECT 90.355 191.965 92.945 193.055 ;
        RECT 93.155 191.965 93.385 193.105 ;
        RECT 93.555 192.135 93.885 193.115 ;
        RECT 94.055 191.965 94.265 193.105 ;
        RECT 94.505 191.965 94.800 192.775 ;
        RECT 94.980 192.135 95.225 193.275 ;
        RECT 95.400 191.965 95.660 192.775 ;
        RECT 95.840 192.140 96.090 193.275 ;
        RECT 102.270 193.105 103.435 193.665 ;
        RECT 96.690 192.880 103.435 193.105 ;
        RECT 103.695 193.055 104.215 193.595 ;
        RECT 104.385 193.225 104.905 193.765 ;
        RECT 105.075 193.745 108.585 194.515 ;
        RECT 105.075 193.055 106.765 193.575 ;
        RECT 106.935 193.225 108.585 193.745 ;
        RECT 108.795 193.695 109.025 194.515 ;
        RECT 109.195 193.715 109.525 194.345 ;
        RECT 108.775 193.275 109.105 193.525 ;
        RECT 109.275 193.115 109.525 193.715 ;
        RECT 109.695 193.695 109.905 194.515 ;
        RECT 110.410 193.705 110.655 194.310 ;
        RECT 110.875 193.980 111.385 194.515 ;
        RECT 96.690 192.865 102.095 192.880 ;
        RECT 96.260 191.970 96.520 192.765 ;
        RECT 96.690 192.140 96.950 192.865 ;
        RECT 97.120 191.970 97.380 192.695 ;
        RECT 97.550 192.140 97.810 192.865 ;
        RECT 97.980 191.970 98.240 192.695 ;
        RECT 98.410 192.140 98.670 192.865 ;
        RECT 98.840 191.970 99.100 192.695 ;
        RECT 99.270 192.140 99.530 192.865 ;
        RECT 99.700 191.970 99.945 192.695 ;
        RECT 100.115 192.140 100.375 192.865 ;
        RECT 100.560 191.970 100.805 192.695 ;
        RECT 100.975 192.140 101.235 192.865 ;
        RECT 101.420 191.970 101.665 192.695 ;
        RECT 101.835 192.140 102.095 192.865 ;
        RECT 102.280 191.970 102.535 192.695 ;
        RECT 102.705 192.140 102.995 192.880 ;
        RECT 96.260 191.965 102.535 191.970 ;
        RECT 103.165 191.965 103.435 192.710 ;
        RECT 103.695 191.965 104.905 193.055 ;
        RECT 105.075 191.965 108.585 193.055 ;
        RECT 108.795 191.965 109.025 193.105 ;
        RECT 109.195 192.135 109.525 193.115 ;
        RECT 110.135 193.535 111.365 193.705 ;
        RECT 109.695 191.965 109.905 193.105 ;
        RECT 110.135 192.725 110.475 193.535 ;
        RECT 110.645 192.970 111.395 193.160 ;
        RECT 110.135 192.315 110.650 192.725 ;
        RECT 110.885 191.965 111.055 192.725 ;
        RECT 111.225 192.305 111.395 192.970 ;
        RECT 111.565 192.985 111.755 194.345 ;
        RECT 111.925 194.175 112.200 194.345 ;
        RECT 111.925 194.005 112.205 194.175 ;
        RECT 111.925 193.185 112.200 194.005 ;
        RECT 112.390 193.980 112.920 194.345 ;
        RECT 113.345 194.115 113.675 194.515 ;
        RECT 112.745 193.945 112.920 193.980 ;
        RECT 112.405 192.985 112.575 193.785 ;
        RECT 111.565 192.815 112.575 192.985 ;
        RECT 112.745 193.775 113.675 193.945 ;
        RECT 113.845 193.775 114.100 194.345 ;
        RECT 114.275 193.790 114.565 194.515 ;
        RECT 112.745 192.645 112.915 193.775 ;
        RECT 113.505 193.605 113.675 193.775 ;
        RECT 111.790 192.475 112.915 192.645 ;
        RECT 113.085 193.275 113.280 193.605 ;
        RECT 113.505 193.275 113.760 193.605 ;
        RECT 113.085 192.305 113.255 193.275 ;
        RECT 113.930 193.105 114.100 193.775 ;
        RECT 114.795 193.695 115.005 194.515 ;
        RECT 115.175 193.715 115.505 194.345 ;
        RECT 111.225 192.135 113.255 192.305 ;
        RECT 113.425 191.965 113.595 193.105 ;
        RECT 113.765 192.135 114.100 193.105 ;
        RECT 114.275 191.965 114.565 193.130 ;
        RECT 115.175 193.115 115.425 193.715 ;
        RECT 115.675 193.695 115.905 194.515 ;
        RECT 117.035 193.745 120.545 194.515 ;
        RECT 120.720 193.970 126.065 194.515 ;
        RECT 115.595 193.275 115.925 193.525 ;
        RECT 114.795 191.965 115.005 193.105 ;
        RECT 115.175 192.135 115.505 193.115 ;
        RECT 115.675 191.965 115.905 193.105 ;
        RECT 117.035 193.055 118.725 193.575 ;
        RECT 118.895 193.225 120.545 193.745 ;
        RECT 117.035 191.965 120.545 193.055 ;
        RECT 122.310 192.400 122.660 193.650 ;
        RECT 124.140 193.140 124.480 193.970 ;
        RECT 126.235 193.765 127.445 194.515 ;
        RECT 126.235 193.055 126.755 193.595 ;
        RECT 126.925 193.225 127.445 193.765 ;
        RECT 120.720 191.965 126.065 192.400 ;
        RECT 126.235 191.965 127.445 193.055 ;
        RECT 14.370 191.795 127.530 191.965 ;
        RECT 14.455 190.705 15.665 191.795 ;
        RECT 14.455 189.995 14.975 190.535 ;
        RECT 15.145 190.165 15.665 190.705 ;
        RECT 15.835 190.705 18.425 191.795 ;
        RECT 18.600 191.360 23.945 191.795 ;
        RECT 15.835 190.185 17.045 190.705 ;
        RECT 17.215 190.015 18.425 190.535 ;
        RECT 20.190 190.110 20.540 191.360 ;
        RECT 24.115 190.630 24.405 191.795 ;
        RECT 25.040 191.360 30.385 191.795 ;
        RECT 30.560 191.360 35.905 191.795 ;
        RECT 14.455 189.245 15.665 189.995 ;
        RECT 15.835 189.245 18.425 190.015 ;
        RECT 22.020 189.790 22.360 190.620 ;
        RECT 26.630 190.110 26.980 191.360 ;
        RECT 18.600 189.245 23.945 189.790 ;
        RECT 24.115 189.245 24.405 189.970 ;
        RECT 28.460 189.790 28.800 190.620 ;
        RECT 32.150 190.110 32.500 191.360 ;
        RECT 36.450 190.815 36.705 191.485 ;
        RECT 36.885 190.995 37.170 191.795 ;
        RECT 37.350 191.075 37.680 191.585 ;
        RECT 36.450 190.775 36.630 190.815 ;
        RECT 33.980 189.790 34.320 190.620 ;
        RECT 36.365 190.605 36.630 190.775 ;
        RECT 36.450 189.955 36.630 190.605 ;
        RECT 37.350 190.485 37.600 191.075 ;
        RECT 37.950 190.925 38.120 191.535 ;
        RECT 38.290 191.105 38.620 191.795 ;
        RECT 38.850 191.245 39.090 191.535 ;
        RECT 39.290 191.415 39.710 191.795 ;
        RECT 39.890 191.325 40.520 191.575 ;
        RECT 40.990 191.415 41.320 191.795 ;
        RECT 39.890 191.245 40.060 191.325 ;
        RECT 41.490 191.245 41.660 191.535 ;
        RECT 41.840 191.415 42.220 191.795 ;
        RECT 42.460 191.410 43.290 191.580 ;
        RECT 38.850 191.075 40.060 191.245 ;
        RECT 36.800 190.155 37.600 190.485 ;
        RECT 25.040 189.245 30.385 189.790 ;
        RECT 30.560 189.245 35.905 189.790 ;
        RECT 36.450 189.425 36.705 189.955 ;
        RECT 36.885 189.245 37.170 189.705 ;
        RECT 37.350 189.505 37.600 190.155 ;
        RECT 37.800 190.905 38.120 190.925 ;
        RECT 37.800 190.735 39.720 190.905 ;
        RECT 37.800 189.840 37.990 190.735 ;
        RECT 39.890 190.565 40.060 191.075 ;
        RECT 40.230 190.815 40.750 191.125 ;
        RECT 38.160 190.395 40.060 190.565 ;
        RECT 38.160 190.335 38.490 190.395 ;
        RECT 38.640 190.165 38.970 190.225 ;
        RECT 38.310 189.895 38.970 190.165 ;
        RECT 37.800 189.510 38.120 189.840 ;
        RECT 38.300 189.245 38.960 189.725 ;
        RECT 39.160 189.635 39.330 190.395 ;
        RECT 40.230 190.225 40.410 190.635 ;
        RECT 39.500 190.055 39.830 190.175 ;
        RECT 40.580 190.055 40.750 190.815 ;
        RECT 39.500 189.885 40.750 190.055 ;
        RECT 40.920 190.995 42.290 191.245 ;
        RECT 40.920 190.225 41.110 190.995 ;
        RECT 42.040 190.735 42.290 190.995 ;
        RECT 41.280 190.565 41.530 190.725 ;
        RECT 42.460 190.565 42.630 191.410 ;
        RECT 43.525 191.125 43.695 191.625 ;
        RECT 43.865 191.295 44.195 191.795 ;
        RECT 42.800 190.735 43.300 191.115 ;
        RECT 43.525 190.955 44.220 191.125 ;
        RECT 41.280 190.395 42.630 190.565 ;
        RECT 42.210 190.355 42.630 190.395 ;
        RECT 40.920 189.885 41.340 190.225 ;
        RECT 41.630 189.895 42.040 190.225 ;
        RECT 39.160 189.465 40.010 189.635 ;
        RECT 40.570 189.245 40.890 189.705 ;
        RECT 41.090 189.455 41.340 189.885 ;
        RECT 41.630 189.245 42.040 189.685 ;
        RECT 42.210 189.625 42.380 190.355 ;
        RECT 42.550 189.805 42.900 190.175 ;
        RECT 43.080 189.865 43.300 190.735 ;
        RECT 43.470 190.165 43.880 190.785 ;
        RECT 44.050 189.985 44.220 190.955 ;
        RECT 43.525 189.795 44.220 189.985 ;
        RECT 42.210 189.425 43.225 189.625 ;
        RECT 43.525 189.465 43.695 189.795 ;
        RECT 43.865 189.245 44.195 189.625 ;
        RECT 44.410 189.505 44.635 191.625 ;
        RECT 44.805 191.295 45.135 191.795 ;
        RECT 45.305 191.125 45.475 191.625 ;
        RECT 44.810 190.955 45.475 191.125 ;
        RECT 45.735 191.035 46.250 191.445 ;
        RECT 46.485 191.035 46.655 191.795 ;
        RECT 46.825 191.455 48.855 191.625 ;
        RECT 44.810 189.965 45.040 190.955 ;
        RECT 45.210 190.135 45.560 190.785 ;
        RECT 45.735 190.225 46.075 191.035 ;
        RECT 46.825 190.790 46.995 191.455 ;
        RECT 47.390 191.115 48.515 191.285 ;
        RECT 46.245 190.600 46.995 190.790 ;
        RECT 47.165 190.775 48.175 190.945 ;
        RECT 45.735 190.055 46.965 190.225 ;
        RECT 44.810 189.795 45.475 189.965 ;
        RECT 44.805 189.245 45.135 189.625 ;
        RECT 45.305 189.505 45.475 189.795 ;
        RECT 46.010 189.450 46.255 190.055 ;
        RECT 46.475 189.245 46.985 189.780 ;
        RECT 47.165 189.415 47.355 190.775 ;
        RECT 47.525 190.435 47.800 190.575 ;
        RECT 47.525 190.265 47.805 190.435 ;
        RECT 47.525 189.415 47.800 190.265 ;
        RECT 48.005 189.975 48.175 190.775 ;
        RECT 48.345 189.985 48.515 191.115 ;
        RECT 48.685 190.485 48.855 191.455 ;
        RECT 49.025 190.655 49.195 191.795 ;
        RECT 49.365 190.655 49.700 191.625 ;
        RECT 48.685 190.155 48.880 190.485 ;
        RECT 49.105 190.155 49.360 190.485 ;
        RECT 49.105 189.985 49.275 190.155 ;
        RECT 49.530 189.985 49.700 190.655 ;
        RECT 49.875 190.630 50.165 191.795 ;
        RECT 50.795 190.720 51.065 191.625 ;
        RECT 51.235 191.035 51.565 191.795 ;
        RECT 51.745 190.865 51.915 191.625 ;
        RECT 48.345 189.815 49.275 189.985 ;
        RECT 48.345 189.780 48.520 189.815 ;
        RECT 47.990 189.415 48.520 189.780 ;
        RECT 48.945 189.245 49.275 189.645 ;
        RECT 49.445 189.415 49.700 189.985 ;
        RECT 49.875 189.245 50.165 189.970 ;
        RECT 50.795 189.920 50.965 190.720 ;
        RECT 51.250 190.695 51.915 190.865 ;
        RECT 51.250 190.550 51.420 190.695 ;
        RECT 51.135 190.220 51.420 190.550 ;
        RECT 52.180 190.605 52.435 191.485 ;
        RECT 52.605 190.655 52.910 191.795 ;
        RECT 53.250 191.415 53.580 191.795 ;
        RECT 53.760 191.245 53.930 191.535 ;
        RECT 54.100 191.335 54.350 191.795 ;
        RECT 53.130 191.075 53.930 191.245 ;
        RECT 54.520 191.285 55.390 191.625 ;
        RECT 51.250 189.965 51.420 190.220 ;
        RECT 51.655 190.145 51.985 190.515 ;
        RECT 50.795 189.415 51.055 189.920 ;
        RECT 51.250 189.795 51.915 189.965 ;
        RECT 51.235 189.245 51.565 189.625 ;
        RECT 51.745 189.415 51.915 189.795 ;
        RECT 52.180 189.955 52.390 190.605 ;
        RECT 53.130 190.485 53.300 191.075 ;
        RECT 54.520 190.905 54.690 191.285 ;
        RECT 55.625 191.165 55.795 191.625 ;
        RECT 55.965 191.335 56.335 191.795 ;
        RECT 56.630 191.195 56.800 191.535 ;
        RECT 56.970 191.365 57.300 191.795 ;
        RECT 57.535 191.195 57.705 191.535 ;
        RECT 53.470 190.735 54.690 190.905 ;
        RECT 54.860 190.825 55.320 191.115 ;
        RECT 55.625 190.995 56.185 191.165 ;
        RECT 56.630 191.025 57.705 191.195 ;
        RECT 57.875 191.295 58.555 191.625 ;
        RECT 58.770 191.295 59.020 191.625 ;
        RECT 59.190 191.335 59.440 191.795 ;
        RECT 56.015 190.855 56.185 190.995 ;
        RECT 54.860 190.815 55.825 190.825 ;
        RECT 54.520 190.645 54.690 190.735 ;
        RECT 55.150 190.655 55.825 190.815 ;
        RECT 52.560 190.455 53.300 190.485 ;
        RECT 52.560 190.155 53.475 190.455 ;
        RECT 53.150 189.980 53.475 190.155 ;
        RECT 52.180 189.425 52.435 189.955 ;
        RECT 52.605 189.245 52.910 189.705 ;
        RECT 53.155 189.625 53.475 189.980 ;
        RECT 53.645 190.195 54.185 190.565 ;
        RECT 54.520 190.475 54.925 190.645 ;
        RECT 53.645 189.795 53.885 190.195 ;
        RECT 54.365 190.025 54.585 190.305 ;
        RECT 54.055 189.855 54.585 190.025 ;
        RECT 54.055 189.625 54.225 189.855 ;
        RECT 54.755 189.695 54.925 190.475 ;
        RECT 55.095 189.865 55.445 190.485 ;
        RECT 55.615 189.865 55.825 190.655 ;
        RECT 56.015 190.685 57.515 190.855 ;
        RECT 56.015 189.995 56.185 190.685 ;
        RECT 57.875 190.515 58.045 191.295 ;
        RECT 58.850 191.165 59.020 191.295 ;
        RECT 56.355 190.345 58.045 190.515 ;
        RECT 58.215 190.735 58.680 191.125 ;
        RECT 58.850 190.995 59.245 191.165 ;
        RECT 56.355 190.165 56.525 190.345 ;
        RECT 53.155 189.455 54.225 189.625 ;
        RECT 54.395 189.245 54.585 189.685 ;
        RECT 54.755 189.415 55.705 189.695 ;
        RECT 56.015 189.605 56.275 189.995 ;
        RECT 56.695 189.925 57.485 190.175 ;
        RECT 55.925 189.435 56.275 189.605 ;
        RECT 56.485 189.245 56.815 189.705 ;
        RECT 57.690 189.635 57.860 190.345 ;
        RECT 58.215 190.145 58.385 190.735 ;
        RECT 58.030 189.925 58.385 190.145 ;
        RECT 58.555 189.925 58.905 190.545 ;
        RECT 59.075 189.635 59.245 190.995 ;
        RECT 59.610 190.825 59.935 191.610 ;
        RECT 59.415 189.775 59.875 190.825 ;
        RECT 57.690 189.465 58.545 189.635 ;
        RECT 58.750 189.465 59.245 189.635 ;
        RECT 59.415 189.245 59.745 189.605 ;
        RECT 60.105 189.505 60.275 191.625 ;
        RECT 60.445 191.295 60.775 191.795 ;
        RECT 60.945 191.125 61.200 191.625 ;
        RECT 60.450 190.955 61.200 191.125 ;
        RECT 60.450 189.965 60.680 190.955 ;
        RECT 60.850 190.135 61.200 190.785 ;
        RECT 61.425 190.655 61.675 191.795 ;
        RECT 61.845 190.605 62.095 191.485 ;
        RECT 62.265 190.655 62.570 191.795 ;
        RECT 62.910 191.415 63.240 191.795 ;
        RECT 63.420 191.245 63.590 191.535 ;
        RECT 63.760 191.335 64.010 191.795 ;
        RECT 62.790 191.075 63.590 191.245 ;
        RECT 64.180 191.285 65.050 191.625 ;
        RECT 60.450 189.795 61.200 189.965 ;
        RECT 60.445 189.245 60.775 189.625 ;
        RECT 60.945 189.505 61.200 189.795 ;
        RECT 61.425 189.245 61.675 190.000 ;
        RECT 61.845 189.955 62.050 190.605 ;
        RECT 62.790 190.485 62.960 191.075 ;
        RECT 64.180 190.905 64.350 191.285 ;
        RECT 65.285 191.165 65.455 191.625 ;
        RECT 65.625 191.335 65.995 191.795 ;
        RECT 66.290 191.195 66.460 191.535 ;
        RECT 66.630 191.365 66.960 191.795 ;
        RECT 67.195 191.195 67.365 191.535 ;
        RECT 63.130 190.735 64.350 190.905 ;
        RECT 64.520 190.825 64.980 191.115 ;
        RECT 65.285 190.995 65.845 191.165 ;
        RECT 66.290 191.025 67.365 191.195 ;
        RECT 67.535 191.295 68.215 191.625 ;
        RECT 68.430 191.295 68.680 191.625 ;
        RECT 68.850 191.335 69.100 191.795 ;
        RECT 65.675 190.855 65.845 190.995 ;
        RECT 64.520 190.815 65.485 190.825 ;
        RECT 64.180 190.645 64.350 190.735 ;
        RECT 64.810 190.655 65.485 190.815 ;
        RECT 62.220 190.455 62.960 190.485 ;
        RECT 62.220 190.155 63.135 190.455 ;
        RECT 62.810 189.980 63.135 190.155 ;
        RECT 61.845 189.425 62.095 189.955 ;
        RECT 62.265 189.245 62.570 189.705 ;
        RECT 62.815 189.625 63.135 189.980 ;
        RECT 63.305 190.195 63.845 190.565 ;
        RECT 64.180 190.475 64.585 190.645 ;
        RECT 63.305 189.795 63.545 190.195 ;
        RECT 64.025 190.025 64.245 190.305 ;
        RECT 63.715 189.855 64.245 190.025 ;
        RECT 63.715 189.625 63.885 189.855 ;
        RECT 64.415 189.695 64.585 190.475 ;
        RECT 64.755 189.865 65.105 190.485 ;
        RECT 65.275 189.865 65.485 190.655 ;
        RECT 65.675 190.685 67.175 190.855 ;
        RECT 65.675 189.995 65.845 190.685 ;
        RECT 67.535 190.515 67.705 191.295 ;
        RECT 68.510 191.165 68.680 191.295 ;
        RECT 66.015 190.345 67.705 190.515 ;
        RECT 67.875 190.735 68.340 191.125 ;
        RECT 68.510 190.995 68.905 191.165 ;
        RECT 66.015 190.165 66.185 190.345 ;
        RECT 62.815 189.455 63.885 189.625 ;
        RECT 64.055 189.245 64.245 189.685 ;
        RECT 64.415 189.415 65.365 189.695 ;
        RECT 65.675 189.605 65.935 189.995 ;
        RECT 66.355 189.925 67.145 190.175 ;
        RECT 65.585 189.435 65.935 189.605 ;
        RECT 66.145 189.245 66.475 189.705 ;
        RECT 67.350 189.635 67.520 190.345 ;
        RECT 67.875 190.145 68.045 190.735 ;
        RECT 67.690 189.925 68.045 190.145 ;
        RECT 68.215 189.925 68.565 190.545 ;
        RECT 68.735 189.635 68.905 190.995 ;
        RECT 69.270 190.825 69.595 191.610 ;
        RECT 69.075 189.775 69.535 190.825 ;
        RECT 67.350 189.465 68.205 189.635 ;
        RECT 68.410 189.465 68.905 189.635 ;
        RECT 69.075 189.245 69.405 189.605 ;
        RECT 69.765 189.505 69.935 191.625 ;
        RECT 70.105 191.295 70.435 191.795 ;
        RECT 70.605 191.125 70.860 191.625 ;
        RECT 71.055 191.285 71.355 191.795 ;
        RECT 71.525 191.285 71.905 191.455 ;
        RECT 72.485 191.285 73.115 191.795 ;
        RECT 70.110 190.955 70.860 191.125 ;
        RECT 71.525 191.115 71.695 191.285 ;
        RECT 73.285 191.115 73.615 191.625 ;
        RECT 73.785 191.285 74.085 191.795 ;
        RECT 70.110 189.965 70.340 190.955 ;
        RECT 71.035 190.915 71.695 191.115 ;
        RECT 71.865 190.945 74.085 191.115 ;
        RECT 70.510 190.135 70.860 190.785 ;
        RECT 71.035 189.985 71.205 190.915 ;
        RECT 71.865 190.745 72.035 190.945 ;
        RECT 71.375 190.575 72.035 190.745 ;
        RECT 72.205 190.605 73.745 190.775 ;
        RECT 71.375 190.155 71.545 190.575 ;
        RECT 72.205 190.405 72.375 190.605 ;
        RECT 71.775 190.235 72.375 190.405 ;
        RECT 72.545 190.235 73.240 190.435 ;
        RECT 73.500 190.155 73.745 190.605 ;
        RECT 71.865 189.985 72.775 190.065 ;
        RECT 70.110 189.795 70.860 189.965 ;
        RECT 70.105 189.245 70.435 189.625 ;
        RECT 70.605 189.505 70.860 189.795 ;
        RECT 71.035 189.505 71.355 189.985 ;
        RECT 71.525 189.895 72.775 189.985 ;
        RECT 71.525 189.815 72.035 189.895 ;
        RECT 71.525 189.415 71.755 189.815 ;
        RECT 71.925 189.245 72.275 189.635 ;
        RECT 72.445 189.415 72.775 189.895 ;
        RECT 72.945 189.245 73.115 190.065 ;
        RECT 73.915 189.985 74.085 190.945 ;
        RECT 74.255 190.705 75.465 191.795 ;
        RECT 74.255 190.165 74.775 190.705 ;
        RECT 75.635 190.630 75.925 191.795 ;
        RECT 76.095 190.655 76.355 191.795 ;
        RECT 76.525 190.825 76.855 191.625 ;
        RECT 77.025 190.995 77.195 191.795 ;
        RECT 77.395 190.825 77.725 191.625 ;
        RECT 77.925 190.995 78.205 191.795 ;
        RECT 76.525 190.655 77.805 190.825 ;
        RECT 74.945 189.995 75.465 190.535 ;
        RECT 76.120 190.155 76.405 190.485 ;
        RECT 76.605 190.155 76.985 190.485 ;
        RECT 77.155 190.155 77.465 190.485 ;
        RECT 73.620 189.440 74.085 189.985 ;
        RECT 74.255 189.245 75.465 189.995 ;
        RECT 75.635 189.245 75.925 189.970 ;
        RECT 76.100 189.245 76.435 189.985 ;
        RECT 76.605 189.460 76.820 190.155 ;
        RECT 77.155 189.985 77.360 190.155 ;
        RECT 77.635 189.985 77.805 190.655 ;
        RECT 77.985 190.155 78.225 190.825 ;
        RECT 79.315 190.705 82.825 191.795 ;
        RECT 83.370 190.815 83.625 191.485 ;
        RECT 83.805 190.995 84.090 191.795 ;
        RECT 84.270 191.075 84.600 191.585 ;
        RECT 79.315 190.185 81.005 190.705 ;
        RECT 81.175 190.015 82.825 190.535 ;
        RECT 77.010 189.460 77.360 189.985 ;
        RECT 77.530 189.415 78.225 189.985 ;
        RECT 79.315 189.245 82.825 190.015 ;
        RECT 83.370 189.955 83.550 190.815 ;
        RECT 84.270 190.485 84.520 191.075 ;
        RECT 84.870 190.925 85.040 191.535 ;
        RECT 85.210 191.105 85.540 191.795 ;
        RECT 85.770 191.245 86.010 191.535 ;
        RECT 86.210 191.415 86.630 191.795 ;
        RECT 86.810 191.325 87.440 191.575 ;
        RECT 87.910 191.415 88.240 191.795 ;
        RECT 86.810 191.245 86.980 191.325 ;
        RECT 88.410 191.245 88.580 191.535 ;
        RECT 88.760 191.415 89.140 191.795 ;
        RECT 89.380 191.410 90.210 191.580 ;
        RECT 85.770 191.075 86.980 191.245 ;
        RECT 83.720 190.155 84.520 190.485 ;
        RECT 83.370 189.755 83.625 189.955 ;
        RECT 83.285 189.585 83.625 189.755 ;
        RECT 83.370 189.425 83.625 189.585 ;
        RECT 83.805 189.245 84.090 189.705 ;
        RECT 84.270 189.505 84.520 190.155 ;
        RECT 84.720 190.905 85.040 190.925 ;
        RECT 84.720 190.735 86.640 190.905 ;
        RECT 84.720 189.840 84.910 190.735 ;
        RECT 86.810 190.565 86.980 191.075 ;
        RECT 87.150 190.815 87.670 191.125 ;
        RECT 85.080 190.395 86.980 190.565 ;
        RECT 85.080 190.335 85.410 190.395 ;
        RECT 85.560 190.165 85.890 190.225 ;
        RECT 85.230 189.895 85.890 190.165 ;
        RECT 84.720 189.510 85.040 189.840 ;
        RECT 85.220 189.245 85.880 189.725 ;
        RECT 86.080 189.635 86.250 190.395 ;
        RECT 87.150 190.225 87.330 190.635 ;
        RECT 86.420 190.055 86.750 190.175 ;
        RECT 87.500 190.055 87.670 190.815 ;
        RECT 86.420 189.885 87.670 190.055 ;
        RECT 87.840 190.995 89.210 191.245 ;
        RECT 87.840 190.225 88.030 190.995 ;
        RECT 88.960 190.735 89.210 190.995 ;
        RECT 88.200 190.565 88.450 190.725 ;
        RECT 89.380 190.565 89.550 191.410 ;
        RECT 90.445 191.125 90.615 191.625 ;
        RECT 90.785 191.295 91.115 191.795 ;
        RECT 89.720 190.735 90.220 191.115 ;
        RECT 90.445 190.955 91.140 191.125 ;
        RECT 88.200 190.395 89.550 190.565 ;
        RECT 89.130 190.355 89.550 190.395 ;
        RECT 87.840 189.885 88.260 190.225 ;
        RECT 88.550 189.895 88.960 190.225 ;
        RECT 86.080 189.465 86.930 189.635 ;
        RECT 87.490 189.245 87.810 189.705 ;
        RECT 88.010 189.455 88.260 189.885 ;
        RECT 88.550 189.245 88.960 189.685 ;
        RECT 89.130 189.625 89.300 190.355 ;
        RECT 89.470 189.805 89.820 190.175 ;
        RECT 90.000 189.865 90.220 190.735 ;
        RECT 90.390 190.165 90.800 190.785 ;
        RECT 90.970 189.985 91.140 190.955 ;
        RECT 90.445 189.795 91.140 189.985 ;
        RECT 89.130 189.425 90.145 189.625 ;
        RECT 90.445 189.465 90.615 189.795 ;
        RECT 90.785 189.245 91.115 189.625 ;
        RECT 91.330 189.505 91.555 191.625 ;
        RECT 91.725 191.295 92.055 191.795 ;
        RECT 92.225 191.125 92.395 191.625 ;
        RECT 91.730 190.955 92.395 191.125 ;
        RECT 91.730 189.965 91.960 190.955 ;
        RECT 92.745 190.865 92.915 191.625 ;
        RECT 93.095 191.035 93.425 191.795 ;
        RECT 92.130 190.135 92.480 190.785 ;
        RECT 92.745 190.695 93.410 190.865 ;
        RECT 93.595 190.720 93.865 191.625 ;
        RECT 94.035 190.960 94.420 191.795 ;
        RECT 94.590 190.790 94.850 191.595 ;
        RECT 95.020 190.960 95.280 191.795 ;
        RECT 95.450 190.790 95.705 191.595 ;
        RECT 95.880 190.960 96.140 191.795 ;
        RECT 96.310 190.790 96.565 191.595 ;
        RECT 96.740 190.960 97.085 191.795 ;
        RECT 97.255 191.035 97.770 191.445 ;
        RECT 98.005 191.035 98.175 191.795 ;
        RECT 98.345 191.455 100.375 191.625 ;
        RECT 93.240 190.550 93.410 190.695 ;
        RECT 92.675 190.145 93.005 190.515 ;
        RECT 93.240 190.220 93.525 190.550 ;
        RECT 93.240 189.965 93.410 190.220 ;
        RECT 91.730 189.795 92.395 189.965 ;
        RECT 91.725 189.245 92.055 189.625 ;
        RECT 92.225 189.505 92.395 189.795 ;
        RECT 92.745 189.795 93.410 189.965 ;
        RECT 93.695 189.920 93.865 190.720 ;
        RECT 92.745 189.415 92.915 189.795 ;
        RECT 93.095 189.245 93.425 189.625 ;
        RECT 93.605 189.415 93.865 189.920 ;
        RECT 94.035 190.620 97.065 190.790 ;
        RECT 94.035 190.055 94.335 190.620 ;
        RECT 94.510 190.225 96.725 190.450 ;
        RECT 96.895 190.055 97.065 190.620 ;
        RECT 97.255 190.225 97.595 191.035 ;
        RECT 98.345 190.790 98.515 191.455 ;
        RECT 98.910 191.115 100.035 191.285 ;
        RECT 97.765 190.600 98.515 190.790 ;
        RECT 98.685 190.775 99.695 190.945 ;
        RECT 97.255 190.055 98.485 190.225 ;
        RECT 94.035 189.885 97.065 190.055 ;
        RECT 94.555 189.245 94.855 189.715 ;
        RECT 95.025 189.440 95.280 189.885 ;
        RECT 95.450 189.245 95.710 189.715 ;
        RECT 95.880 189.440 96.140 189.885 ;
        RECT 96.310 189.245 96.605 189.715 ;
        RECT 97.530 189.450 97.775 190.055 ;
        RECT 97.995 189.245 98.505 189.780 ;
        RECT 98.685 189.415 98.875 190.775 ;
        RECT 99.045 190.435 99.320 190.575 ;
        RECT 99.045 190.265 99.325 190.435 ;
        RECT 99.045 189.415 99.320 190.265 ;
        RECT 99.525 189.975 99.695 190.775 ;
        RECT 99.865 189.985 100.035 191.115 ;
        RECT 100.205 190.485 100.375 191.455 ;
        RECT 100.545 190.655 100.715 191.795 ;
        RECT 100.885 190.655 101.220 191.625 ;
        RECT 100.205 190.155 100.400 190.485 ;
        RECT 100.625 190.155 100.880 190.485 ;
        RECT 100.625 189.985 100.795 190.155 ;
        RECT 101.050 189.985 101.220 190.655 ;
        RECT 101.395 190.630 101.685 191.795 ;
        RECT 101.945 190.865 102.115 191.625 ;
        RECT 102.295 191.035 102.625 191.795 ;
        RECT 101.945 190.695 102.610 190.865 ;
        RECT 102.795 190.720 103.065 191.625 ;
        RECT 102.440 190.550 102.610 190.695 ;
        RECT 101.875 190.145 102.205 190.515 ;
        RECT 102.440 190.220 102.725 190.550 ;
        RECT 99.865 189.815 100.795 189.985 ;
        RECT 99.865 189.780 100.040 189.815 ;
        RECT 99.510 189.415 100.040 189.780 ;
        RECT 100.465 189.245 100.795 189.645 ;
        RECT 100.965 189.415 101.220 189.985 ;
        RECT 101.395 189.245 101.685 189.970 ;
        RECT 102.440 189.965 102.610 190.220 ;
        RECT 101.945 189.795 102.610 189.965 ;
        RECT 102.895 189.920 103.065 190.720 ;
        RECT 103.235 190.705 104.445 191.795 ;
        RECT 104.615 191.035 105.130 191.445 ;
        RECT 105.365 191.035 105.535 191.795 ;
        RECT 105.705 191.455 107.735 191.625 ;
        RECT 103.235 190.165 103.755 190.705 ;
        RECT 103.925 189.995 104.445 190.535 ;
        RECT 104.615 190.225 104.955 191.035 ;
        RECT 105.705 190.790 105.875 191.455 ;
        RECT 106.270 191.115 107.395 191.285 ;
        RECT 105.125 190.600 105.875 190.790 ;
        RECT 106.045 190.775 107.055 190.945 ;
        RECT 104.615 190.055 105.845 190.225 ;
        RECT 101.945 189.415 102.115 189.795 ;
        RECT 102.295 189.245 102.625 189.625 ;
        RECT 102.805 189.415 103.065 189.920 ;
        RECT 103.235 189.245 104.445 189.995 ;
        RECT 104.890 189.450 105.135 190.055 ;
        RECT 105.355 189.245 105.865 189.780 ;
        RECT 106.045 189.415 106.235 190.775 ;
        RECT 106.405 190.435 106.680 190.575 ;
        RECT 106.405 190.265 106.685 190.435 ;
        RECT 106.405 189.415 106.680 190.265 ;
        RECT 106.885 189.975 107.055 190.775 ;
        RECT 107.225 189.985 107.395 191.115 ;
        RECT 107.565 190.485 107.735 191.455 ;
        RECT 107.905 190.655 108.075 191.795 ;
        RECT 108.245 190.655 108.580 191.625 ;
        RECT 107.565 190.155 107.760 190.485 ;
        RECT 107.985 190.155 108.240 190.485 ;
        RECT 107.985 189.985 108.155 190.155 ;
        RECT 108.410 189.985 108.580 190.655 ;
        RECT 107.225 189.815 108.155 189.985 ;
        RECT 107.225 189.780 107.400 189.815 ;
        RECT 106.870 189.415 107.400 189.780 ;
        RECT 107.825 189.245 108.155 189.645 ;
        RECT 108.325 189.415 108.580 189.985 ;
        RECT 108.760 190.605 109.015 191.485 ;
        RECT 109.185 190.655 109.490 191.795 ;
        RECT 109.830 191.415 110.160 191.795 ;
        RECT 110.340 191.245 110.510 191.535 ;
        RECT 110.680 191.335 110.930 191.795 ;
        RECT 109.710 191.075 110.510 191.245 ;
        RECT 111.100 191.285 111.970 191.625 ;
        RECT 108.760 189.955 108.970 190.605 ;
        RECT 109.710 190.485 109.880 191.075 ;
        RECT 111.100 190.905 111.270 191.285 ;
        RECT 112.205 191.165 112.375 191.625 ;
        RECT 112.545 191.335 112.915 191.795 ;
        RECT 113.210 191.195 113.380 191.535 ;
        RECT 113.550 191.365 113.880 191.795 ;
        RECT 114.115 191.195 114.285 191.535 ;
        RECT 110.050 190.735 111.270 190.905 ;
        RECT 111.440 190.825 111.900 191.115 ;
        RECT 112.205 190.995 112.765 191.165 ;
        RECT 113.210 191.025 114.285 191.195 ;
        RECT 114.455 191.295 115.135 191.625 ;
        RECT 115.350 191.295 115.600 191.625 ;
        RECT 115.770 191.335 116.020 191.795 ;
        RECT 112.595 190.855 112.765 190.995 ;
        RECT 111.440 190.815 112.405 190.825 ;
        RECT 111.100 190.645 111.270 190.735 ;
        RECT 111.730 190.655 112.405 190.815 ;
        RECT 109.140 190.455 109.880 190.485 ;
        RECT 109.140 190.155 110.055 190.455 ;
        RECT 109.730 189.980 110.055 190.155 ;
        RECT 108.760 189.425 109.015 189.955 ;
        RECT 109.185 189.245 109.490 189.705 ;
        RECT 109.735 189.625 110.055 189.980 ;
        RECT 110.225 190.195 110.765 190.565 ;
        RECT 111.100 190.475 111.505 190.645 ;
        RECT 110.225 189.795 110.465 190.195 ;
        RECT 110.945 190.025 111.165 190.305 ;
        RECT 110.635 189.855 111.165 190.025 ;
        RECT 110.635 189.625 110.805 189.855 ;
        RECT 111.335 189.695 111.505 190.475 ;
        RECT 111.675 189.865 112.025 190.485 ;
        RECT 112.195 189.865 112.405 190.655 ;
        RECT 112.595 190.685 114.095 190.855 ;
        RECT 112.595 189.995 112.765 190.685 ;
        RECT 114.455 190.515 114.625 191.295 ;
        RECT 115.430 191.165 115.600 191.295 ;
        RECT 112.935 190.345 114.625 190.515 ;
        RECT 114.795 190.735 115.260 191.125 ;
        RECT 115.430 190.995 115.825 191.165 ;
        RECT 112.935 190.165 113.105 190.345 ;
        RECT 109.735 189.455 110.805 189.625 ;
        RECT 110.975 189.245 111.165 189.685 ;
        RECT 111.335 189.415 112.285 189.695 ;
        RECT 112.595 189.605 112.855 189.995 ;
        RECT 113.275 189.925 114.065 190.175 ;
        RECT 112.505 189.435 112.855 189.605 ;
        RECT 113.065 189.245 113.395 189.705 ;
        RECT 114.270 189.635 114.440 190.345 ;
        RECT 114.795 190.145 114.965 190.735 ;
        RECT 114.610 189.925 114.965 190.145 ;
        RECT 115.135 189.925 115.485 190.545 ;
        RECT 115.655 189.635 115.825 190.995 ;
        RECT 116.190 190.825 116.515 191.610 ;
        RECT 115.995 189.775 116.455 190.825 ;
        RECT 114.270 189.465 115.125 189.635 ;
        RECT 115.330 189.465 115.825 189.635 ;
        RECT 115.995 189.245 116.325 189.605 ;
        RECT 116.685 189.505 116.855 191.625 ;
        RECT 117.025 191.295 117.355 191.795 ;
        RECT 117.525 191.125 117.780 191.625 ;
        RECT 117.030 190.955 117.780 191.125 ;
        RECT 117.030 189.965 117.260 190.955 ;
        RECT 117.430 190.135 117.780 190.785 ;
        RECT 117.955 190.720 118.225 191.625 ;
        RECT 118.395 191.035 118.725 191.795 ;
        RECT 118.905 190.865 119.075 191.625 ;
        RECT 117.030 189.795 117.780 189.965 ;
        RECT 117.025 189.245 117.355 189.625 ;
        RECT 117.525 189.505 117.780 189.795 ;
        RECT 117.955 189.920 118.125 190.720 ;
        RECT 118.410 190.695 119.075 190.865 ;
        RECT 119.335 190.705 120.545 191.795 ;
        RECT 120.720 191.360 126.065 191.795 ;
        RECT 118.410 190.550 118.580 190.695 ;
        RECT 118.295 190.220 118.580 190.550 ;
        RECT 118.410 189.965 118.580 190.220 ;
        RECT 118.815 190.145 119.145 190.515 ;
        RECT 119.335 190.165 119.855 190.705 ;
        RECT 120.025 189.995 120.545 190.535 ;
        RECT 122.310 190.110 122.660 191.360 ;
        RECT 126.235 190.705 127.445 191.795 ;
        RECT 117.955 189.415 118.215 189.920 ;
        RECT 118.410 189.795 119.075 189.965 ;
        RECT 118.395 189.245 118.725 189.625 ;
        RECT 118.905 189.415 119.075 189.795 ;
        RECT 119.335 189.245 120.545 189.995 ;
        RECT 124.140 189.790 124.480 190.620 ;
        RECT 126.235 190.165 126.755 190.705 ;
        RECT 126.925 189.995 127.445 190.535 ;
        RECT 120.720 189.245 126.065 189.790 ;
        RECT 126.235 189.245 127.445 189.995 ;
        RECT 14.370 189.075 127.530 189.245 ;
        RECT 14.455 188.325 15.665 189.075 ;
        RECT 14.455 187.785 14.975 188.325 ;
        RECT 16.295 188.305 17.965 189.075 ;
        RECT 18.140 188.530 23.485 189.075 ;
        RECT 23.660 188.530 29.005 189.075 ;
        RECT 15.145 187.615 15.665 188.155 ;
        RECT 14.455 186.525 15.665 187.615 ;
        RECT 16.295 187.615 17.045 188.135 ;
        RECT 17.215 187.785 17.965 188.305 ;
        RECT 16.295 186.525 17.965 187.615 ;
        RECT 19.730 186.960 20.080 188.210 ;
        RECT 21.560 187.700 21.900 188.530 ;
        RECT 25.250 186.960 25.600 188.210 ;
        RECT 27.080 187.700 27.420 188.530 ;
        RECT 29.235 188.255 29.445 189.075 ;
        RECT 29.615 188.275 29.945 188.905 ;
        RECT 29.615 187.675 29.865 188.275 ;
        RECT 30.115 188.255 30.345 189.075 ;
        RECT 30.555 188.325 31.765 189.075 ;
        RECT 30.035 187.835 30.365 188.085 ;
        RECT 18.140 186.525 23.485 186.960 ;
        RECT 23.660 186.525 29.005 186.960 ;
        RECT 29.235 186.525 29.445 187.665 ;
        RECT 29.615 186.695 29.945 187.675 ;
        RECT 30.115 186.525 30.345 187.665 ;
        RECT 30.555 187.615 31.075 188.155 ;
        RECT 31.245 187.785 31.765 188.325 ;
        RECT 31.935 188.305 35.445 189.075 ;
        RECT 31.935 187.615 33.625 188.135 ;
        RECT 33.795 187.785 35.445 188.305 ;
        RECT 35.655 188.255 35.885 189.075 ;
        RECT 36.055 188.275 36.385 188.905 ;
        RECT 35.635 187.835 35.965 188.085 ;
        RECT 36.135 187.675 36.385 188.275 ;
        RECT 36.555 188.255 36.765 189.075 ;
        RECT 36.995 188.350 37.285 189.075 ;
        RECT 37.460 188.365 37.715 188.895 ;
        RECT 37.885 188.615 38.190 189.075 ;
        RECT 38.435 188.695 39.505 188.865 ;
        RECT 37.460 187.715 37.670 188.365 ;
        RECT 38.435 188.340 38.755 188.695 ;
        RECT 38.430 188.165 38.755 188.340 ;
        RECT 37.840 187.865 38.755 188.165 ;
        RECT 38.925 188.125 39.165 188.525 ;
        RECT 39.335 188.465 39.505 188.695 ;
        RECT 39.675 188.635 39.865 189.075 ;
        RECT 40.035 188.625 40.985 188.905 ;
        RECT 41.205 188.715 41.555 188.885 ;
        RECT 39.335 188.295 39.865 188.465 ;
        RECT 37.840 187.835 38.580 187.865 ;
        RECT 30.555 186.525 31.765 187.615 ;
        RECT 31.935 186.525 35.445 187.615 ;
        RECT 35.655 186.525 35.885 187.665 ;
        RECT 36.055 186.695 36.385 187.675 ;
        RECT 36.555 186.525 36.765 187.665 ;
        RECT 36.995 186.525 37.285 187.690 ;
        RECT 37.460 186.835 37.715 187.715 ;
        RECT 37.885 186.525 38.190 187.665 ;
        RECT 38.410 187.245 38.580 187.835 ;
        RECT 38.925 187.755 39.465 188.125 ;
        RECT 39.645 188.015 39.865 188.295 ;
        RECT 40.035 187.845 40.205 188.625 ;
        RECT 39.800 187.675 40.205 187.845 ;
        RECT 40.375 187.835 40.725 188.455 ;
        RECT 39.800 187.585 39.970 187.675 ;
        RECT 40.895 187.665 41.105 188.455 ;
        RECT 38.750 187.415 39.970 187.585 ;
        RECT 40.430 187.505 41.105 187.665 ;
        RECT 38.410 187.075 39.210 187.245 ;
        RECT 38.530 186.525 38.860 186.905 ;
        RECT 39.040 186.785 39.210 187.075 ;
        RECT 39.800 187.035 39.970 187.415 ;
        RECT 40.140 187.495 41.105 187.505 ;
        RECT 41.295 188.325 41.555 188.715 ;
        RECT 41.765 188.615 42.095 189.075 ;
        RECT 42.970 188.685 43.825 188.855 ;
        RECT 44.030 188.685 44.525 188.855 ;
        RECT 44.695 188.715 45.025 189.075 ;
        RECT 41.295 187.635 41.465 188.325 ;
        RECT 41.635 187.975 41.805 188.155 ;
        RECT 41.975 188.145 42.765 188.395 ;
        RECT 42.970 187.975 43.140 188.685 ;
        RECT 43.310 188.175 43.665 188.395 ;
        RECT 41.635 187.805 43.325 187.975 ;
        RECT 40.140 187.205 40.600 187.495 ;
        RECT 41.295 187.465 42.795 187.635 ;
        RECT 41.295 187.325 41.465 187.465 ;
        RECT 40.905 187.155 41.465 187.325 ;
        RECT 39.380 186.525 39.630 186.985 ;
        RECT 39.800 186.695 40.670 187.035 ;
        RECT 40.905 186.695 41.075 187.155 ;
        RECT 41.910 187.125 42.985 187.295 ;
        RECT 41.245 186.525 41.615 186.985 ;
        RECT 41.910 186.785 42.080 187.125 ;
        RECT 42.250 186.525 42.580 186.955 ;
        RECT 42.815 186.785 42.985 187.125 ;
        RECT 43.155 187.025 43.325 187.805 ;
        RECT 43.495 187.585 43.665 188.175 ;
        RECT 43.835 187.775 44.185 188.395 ;
        RECT 43.495 187.195 43.960 187.585 ;
        RECT 44.355 187.325 44.525 188.685 ;
        RECT 44.695 187.495 45.155 188.545 ;
        RECT 44.130 187.155 44.525 187.325 ;
        RECT 44.130 187.025 44.300 187.155 ;
        RECT 43.155 186.695 43.835 187.025 ;
        RECT 44.050 186.695 44.300 187.025 ;
        RECT 44.470 186.525 44.720 186.985 ;
        RECT 44.890 186.710 45.215 187.495 ;
        RECT 45.385 186.695 45.555 188.815 ;
        RECT 45.725 188.695 46.055 189.075 ;
        RECT 46.225 188.525 46.480 188.815 ;
        RECT 46.745 188.595 47.045 189.075 ;
        RECT 45.730 188.355 46.480 188.525 ;
        RECT 47.215 188.425 47.475 188.880 ;
        RECT 47.645 188.595 47.905 189.075 ;
        RECT 48.085 188.425 48.345 188.880 ;
        RECT 48.515 188.595 48.765 189.075 ;
        RECT 48.945 188.425 49.205 188.880 ;
        RECT 49.375 188.595 49.625 189.075 ;
        RECT 49.805 188.425 50.065 188.880 ;
        RECT 50.235 188.595 50.480 189.075 ;
        RECT 50.650 188.425 50.925 188.880 ;
        RECT 51.095 188.595 51.340 189.075 ;
        RECT 51.510 188.425 51.770 188.880 ;
        RECT 51.940 188.595 52.200 189.075 ;
        RECT 52.370 188.425 52.630 188.880 ;
        RECT 52.800 188.595 53.060 189.075 ;
        RECT 53.230 188.425 53.490 188.880 ;
        RECT 53.660 188.515 53.920 189.075 ;
        RECT 45.730 187.365 45.960 188.355 ;
        RECT 46.745 188.255 53.490 188.425 ;
        RECT 46.130 187.535 46.480 188.185 ;
        RECT 46.745 187.665 47.910 188.255 ;
        RECT 54.090 188.085 54.340 188.895 ;
        RECT 54.520 188.550 54.780 189.075 ;
        RECT 54.950 188.085 55.200 188.895 ;
        RECT 55.380 188.565 55.685 189.075 ;
        RECT 48.080 187.835 55.200 188.085 ;
        RECT 55.370 187.835 55.685 188.395 ;
        RECT 56.130 188.265 56.375 188.870 ;
        RECT 56.595 188.540 57.105 189.075 ;
        RECT 55.855 188.095 57.085 188.265 ;
        RECT 46.745 187.440 53.490 187.665 ;
        RECT 45.730 187.195 46.480 187.365 ;
        RECT 45.725 186.525 46.055 187.025 ;
        RECT 46.225 186.695 46.480 187.195 ;
        RECT 46.745 186.525 47.015 187.270 ;
        RECT 47.185 186.700 47.475 187.440 ;
        RECT 48.085 187.425 53.490 187.440 ;
        RECT 47.645 186.530 47.900 187.255 ;
        RECT 48.085 186.700 48.345 187.425 ;
        RECT 48.515 186.530 48.760 187.255 ;
        RECT 48.945 186.700 49.205 187.425 ;
        RECT 49.375 186.530 49.620 187.255 ;
        RECT 49.805 186.700 50.065 187.425 ;
        RECT 50.235 186.530 50.480 187.255 ;
        RECT 50.650 186.700 50.910 187.425 ;
        RECT 51.080 186.530 51.340 187.255 ;
        RECT 51.510 186.700 51.770 187.425 ;
        RECT 51.940 186.530 52.200 187.255 ;
        RECT 52.370 186.700 52.630 187.425 ;
        RECT 52.800 186.530 53.060 187.255 ;
        RECT 53.230 186.700 53.490 187.425 ;
        RECT 53.660 186.530 53.920 187.325 ;
        RECT 54.090 186.700 54.340 187.835 ;
        RECT 47.645 186.525 53.920 186.530 ;
        RECT 54.520 186.525 54.780 187.335 ;
        RECT 54.955 186.695 55.200 187.835 ;
        RECT 55.380 186.525 55.675 187.335 ;
        RECT 55.855 187.285 56.195 188.095 ;
        RECT 56.365 187.530 57.115 187.720 ;
        RECT 55.855 186.875 56.370 187.285 ;
        RECT 56.605 186.525 56.775 187.285 ;
        RECT 56.945 186.865 57.115 187.530 ;
        RECT 57.285 187.545 57.475 188.905 ;
        RECT 57.645 188.735 57.920 188.905 ;
        RECT 57.645 188.565 57.925 188.735 ;
        RECT 57.645 187.745 57.920 188.565 ;
        RECT 58.110 188.540 58.640 188.905 ;
        RECT 59.065 188.675 59.395 189.075 ;
        RECT 58.465 188.505 58.640 188.540 ;
        RECT 58.125 187.545 58.295 188.345 ;
        RECT 57.285 187.375 58.295 187.545 ;
        RECT 58.465 188.335 59.395 188.505 ;
        RECT 59.565 188.335 59.820 188.905 ;
        RECT 58.465 187.205 58.635 188.335 ;
        RECT 59.225 188.165 59.395 188.335 ;
        RECT 57.510 187.035 58.635 187.205 ;
        RECT 58.805 187.835 59.000 188.165 ;
        RECT 59.225 187.835 59.480 188.165 ;
        RECT 58.805 186.865 58.975 187.835 ;
        RECT 59.650 187.665 59.820 188.335 ;
        RECT 56.945 186.695 58.975 186.865 ;
        RECT 59.145 186.525 59.315 187.665 ;
        RECT 59.485 186.695 59.820 187.665 ;
        RECT 59.995 188.400 60.255 188.905 ;
        RECT 60.435 188.695 60.765 189.075 ;
        RECT 60.945 188.525 61.115 188.905 ;
        RECT 59.995 187.600 60.165 188.400 ;
        RECT 60.450 188.355 61.115 188.525 ;
        RECT 60.450 188.100 60.620 188.355 ;
        RECT 61.375 188.325 62.585 189.075 ;
        RECT 62.755 188.350 63.045 189.075 ;
        RECT 63.790 188.445 64.075 188.905 ;
        RECT 64.245 188.615 64.515 189.075 ;
        RECT 60.335 187.770 60.620 188.100 ;
        RECT 60.855 187.805 61.185 188.175 ;
        RECT 60.450 187.625 60.620 187.770 ;
        RECT 59.995 186.695 60.265 187.600 ;
        RECT 60.450 187.455 61.115 187.625 ;
        RECT 60.435 186.525 60.765 187.285 ;
        RECT 60.945 186.695 61.115 187.455 ;
        RECT 61.375 187.615 61.895 188.155 ;
        RECT 62.065 187.785 62.585 188.325 ;
        RECT 63.790 188.275 64.745 188.445 ;
        RECT 61.375 186.525 62.585 187.615 ;
        RECT 62.755 186.525 63.045 187.690 ;
        RECT 63.675 187.545 64.365 188.105 ;
        RECT 64.535 187.375 64.745 188.275 ;
        RECT 63.790 187.155 64.745 187.375 ;
        RECT 64.915 188.105 65.315 188.905 ;
        RECT 65.505 188.445 65.785 188.905 ;
        RECT 66.305 188.615 66.630 189.075 ;
        RECT 65.505 188.275 66.630 188.445 ;
        RECT 66.800 188.335 67.185 188.905 ;
        RECT 66.180 188.165 66.630 188.275 ;
        RECT 64.915 187.545 66.010 188.105 ;
        RECT 66.180 187.835 66.735 188.165 ;
        RECT 63.790 186.695 64.075 187.155 ;
        RECT 64.245 186.525 64.515 186.985 ;
        RECT 64.915 186.695 65.315 187.545 ;
        RECT 66.180 187.375 66.630 187.835 ;
        RECT 66.905 187.665 67.185 188.335 ;
        RECT 67.355 188.305 69.945 189.075 ;
        RECT 70.120 188.530 75.465 189.075 ;
        RECT 75.640 188.530 80.985 189.075 ;
        RECT 81.160 188.530 86.505 189.075 ;
        RECT 65.505 187.155 66.630 187.375 ;
        RECT 65.505 186.695 65.785 187.155 ;
        RECT 66.305 186.525 66.630 186.985 ;
        RECT 66.800 186.695 67.185 187.665 ;
        RECT 67.355 187.615 68.565 188.135 ;
        RECT 68.735 187.785 69.945 188.305 ;
        RECT 67.355 186.525 69.945 187.615 ;
        RECT 71.710 186.960 72.060 188.210 ;
        RECT 73.540 187.700 73.880 188.530 ;
        RECT 77.230 186.960 77.580 188.210 ;
        RECT 79.060 187.700 79.400 188.530 ;
        RECT 82.750 186.960 83.100 188.210 ;
        RECT 84.580 187.700 84.920 188.530 ;
        RECT 86.735 188.255 86.945 189.075 ;
        RECT 87.115 188.275 87.445 188.905 ;
        RECT 87.115 187.675 87.365 188.275 ;
        RECT 87.615 188.255 87.845 189.075 ;
        RECT 88.515 188.350 88.805 189.075 ;
        RECT 89.065 188.525 89.235 188.905 ;
        RECT 89.415 188.695 89.745 189.075 ;
        RECT 89.065 188.355 89.730 188.525 ;
        RECT 89.925 188.400 90.185 188.905 ;
        RECT 87.535 187.835 87.865 188.085 ;
        RECT 88.995 187.805 89.325 188.175 ;
        RECT 89.560 188.100 89.730 188.355 ;
        RECT 89.560 187.770 89.845 188.100 ;
        RECT 70.120 186.525 75.465 186.960 ;
        RECT 75.640 186.525 80.985 186.960 ;
        RECT 81.160 186.525 86.505 186.960 ;
        RECT 86.735 186.525 86.945 187.665 ;
        RECT 87.115 186.695 87.445 187.675 ;
        RECT 87.615 186.525 87.845 187.665 ;
        RECT 88.515 186.525 88.805 187.690 ;
        RECT 89.560 187.625 89.730 187.770 ;
        RECT 89.065 187.455 89.730 187.625 ;
        RECT 90.015 187.600 90.185 188.400 ;
        RECT 90.355 188.305 92.025 189.075 ;
        RECT 92.200 188.530 97.545 189.075 ;
        RECT 89.065 186.695 89.235 187.455 ;
        RECT 89.415 186.525 89.745 187.285 ;
        RECT 89.915 186.695 90.185 187.600 ;
        RECT 90.355 187.615 91.105 188.135 ;
        RECT 91.275 187.785 92.025 188.305 ;
        RECT 90.355 186.525 92.025 187.615 ;
        RECT 93.790 186.960 94.140 188.210 ;
        RECT 95.620 187.700 95.960 188.530 ;
        RECT 97.720 188.365 97.975 188.895 ;
        RECT 98.145 188.615 98.450 189.075 ;
        RECT 98.695 188.695 99.765 188.865 ;
        RECT 97.720 187.715 97.930 188.365 ;
        RECT 98.695 188.340 99.015 188.695 ;
        RECT 98.690 188.165 99.015 188.340 ;
        RECT 98.100 187.865 99.015 188.165 ;
        RECT 99.185 188.125 99.425 188.525 ;
        RECT 99.595 188.465 99.765 188.695 ;
        RECT 99.935 188.635 100.125 189.075 ;
        RECT 100.295 188.625 101.245 188.905 ;
        RECT 101.465 188.715 101.815 188.885 ;
        RECT 99.595 188.295 100.125 188.465 ;
        RECT 98.100 187.835 98.840 187.865 ;
        RECT 92.200 186.525 97.545 186.960 ;
        RECT 97.720 186.835 97.975 187.715 ;
        RECT 98.145 186.525 98.450 187.665 ;
        RECT 98.670 187.245 98.840 187.835 ;
        RECT 99.185 187.755 99.725 188.125 ;
        RECT 99.905 188.015 100.125 188.295 ;
        RECT 100.295 187.845 100.465 188.625 ;
        RECT 100.060 187.675 100.465 187.845 ;
        RECT 100.635 187.835 100.985 188.455 ;
        RECT 100.060 187.585 100.230 187.675 ;
        RECT 101.155 187.665 101.365 188.455 ;
        RECT 99.010 187.415 100.230 187.585 ;
        RECT 100.690 187.505 101.365 187.665 ;
        RECT 98.670 187.075 99.470 187.245 ;
        RECT 98.790 186.525 99.120 186.905 ;
        RECT 99.300 186.785 99.470 187.075 ;
        RECT 100.060 187.035 100.230 187.415 ;
        RECT 100.400 187.495 101.365 187.505 ;
        RECT 101.555 188.325 101.815 188.715 ;
        RECT 102.025 188.615 102.355 189.075 ;
        RECT 103.230 188.685 104.085 188.855 ;
        RECT 104.290 188.685 104.785 188.855 ;
        RECT 104.955 188.715 105.285 189.075 ;
        RECT 101.555 187.635 101.725 188.325 ;
        RECT 101.895 187.975 102.065 188.155 ;
        RECT 102.235 188.145 103.025 188.395 ;
        RECT 103.230 187.975 103.400 188.685 ;
        RECT 103.570 188.175 103.925 188.395 ;
        RECT 101.895 187.805 103.585 187.975 ;
        RECT 100.400 187.205 100.860 187.495 ;
        RECT 101.555 187.465 103.055 187.635 ;
        RECT 101.555 187.325 101.725 187.465 ;
        RECT 101.165 187.155 101.725 187.325 ;
        RECT 99.640 186.525 99.890 186.985 ;
        RECT 100.060 186.695 100.930 187.035 ;
        RECT 101.165 186.695 101.335 187.155 ;
        RECT 102.170 187.125 103.245 187.295 ;
        RECT 101.505 186.525 101.875 186.985 ;
        RECT 102.170 186.785 102.340 187.125 ;
        RECT 102.510 186.525 102.840 186.955 ;
        RECT 103.075 186.785 103.245 187.125 ;
        RECT 103.415 187.025 103.585 187.805 ;
        RECT 103.755 187.585 103.925 188.175 ;
        RECT 104.095 187.775 104.445 188.395 ;
        RECT 103.755 187.195 104.220 187.585 ;
        RECT 104.615 187.325 104.785 188.685 ;
        RECT 104.955 187.495 105.415 188.545 ;
        RECT 104.390 187.155 104.785 187.325 ;
        RECT 104.390 187.025 104.560 187.155 ;
        RECT 103.415 186.695 104.095 187.025 ;
        RECT 104.310 186.695 104.560 187.025 ;
        RECT 104.730 186.525 104.980 186.985 ;
        RECT 105.150 186.710 105.475 187.495 ;
        RECT 105.645 186.695 105.815 188.815 ;
        RECT 105.985 188.695 106.315 189.075 ;
        RECT 106.485 188.525 106.740 188.815 ;
        RECT 105.990 188.355 106.740 188.525 ;
        RECT 105.990 187.365 106.220 188.355 ;
        RECT 106.915 188.335 107.300 188.905 ;
        RECT 107.470 188.615 107.795 189.075 ;
        RECT 108.315 188.445 108.595 188.905 ;
        RECT 106.390 187.535 106.740 188.185 ;
        RECT 106.915 187.665 107.195 188.335 ;
        RECT 107.470 188.275 108.595 188.445 ;
        RECT 107.470 188.165 107.920 188.275 ;
        RECT 107.365 187.835 107.920 188.165 ;
        RECT 108.785 188.105 109.185 188.905 ;
        RECT 109.585 188.615 109.855 189.075 ;
        RECT 110.025 188.445 110.310 188.905 ;
        RECT 105.990 187.195 106.740 187.365 ;
        RECT 105.985 186.525 106.315 187.025 ;
        RECT 106.485 186.695 106.740 187.195 ;
        RECT 106.915 186.695 107.300 187.665 ;
        RECT 107.470 187.375 107.920 187.835 ;
        RECT 108.090 187.545 109.185 188.105 ;
        RECT 107.470 187.155 108.595 187.375 ;
        RECT 107.470 186.525 107.795 186.985 ;
        RECT 108.315 186.695 108.595 187.155 ;
        RECT 108.785 186.695 109.185 187.545 ;
        RECT 109.355 188.275 110.310 188.445 ;
        RECT 111.055 188.305 112.725 189.075 ;
        RECT 112.985 188.525 113.155 188.905 ;
        RECT 113.335 188.695 113.665 189.075 ;
        RECT 112.985 188.355 113.650 188.525 ;
        RECT 113.845 188.400 114.105 188.905 ;
        RECT 109.355 187.375 109.565 188.275 ;
        RECT 109.735 187.545 110.425 188.105 ;
        RECT 111.055 187.615 111.805 188.135 ;
        RECT 111.975 187.785 112.725 188.305 ;
        RECT 112.915 187.805 113.245 188.175 ;
        RECT 113.480 188.100 113.650 188.355 ;
        RECT 113.480 187.770 113.765 188.100 ;
        RECT 113.480 187.625 113.650 187.770 ;
        RECT 109.355 187.155 110.310 187.375 ;
        RECT 109.585 186.525 109.855 186.985 ;
        RECT 110.025 186.695 110.310 187.155 ;
        RECT 111.055 186.525 112.725 187.615 ;
        RECT 112.985 187.455 113.650 187.625 ;
        RECT 113.935 187.600 114.105 188.400 ;
        RECT 114.275 188.350 114.565 189.075 ;
        RECT 115.200 188.530 120.545 189.075 ;
        RECT 120.720 188.530 126.065 189.075 ;
        RECT 112.985 186.695 113.155 187.455 ;
        RECT 113.335 186.525 113.665 187.285 ;
        RECT 113.835 186.695 114.105 187.600 ;
        RECT 114.275 186.525 114.565 187.690 ;
        RECT 116.790 186.960 117.140 188.210 ;
        RECT 118.620 187.700 118.960 188.530 ;
        RECT 122.310 186.960 122.660 188.210 ;
        RECT 124.140 187.700 124.480 188.530 ;
        RECT 126.235 188.325 127.445 189.075 ;
        RECT 126.235 187.615 126.755 188.155 ;
        RECT 126.925 187.785 127.445 188.325 ;
        RECT 115.200 186.525 120.545 186.960 ;
        RECT 120.720 186.525 126.065 186.960 ;
        RECT 126.235 186.525 127.445 187.615 ;
        RECT 14.370 186.355 127.530 186.525 ;
        RECT 14.455 185.265 15.665 186.355 ;
        RECT 14.455 184.555 14.975 185.095 ;
        RECT 15.145 184.725 15.665 185.265 ;
        RECT 15.835 185.265 18.425 186.355 ;
        RECT 18.600 185.920 23.945 186.355 ;
        RECT 15.835 184.745 17.045 185.265 ;
        RECT 17.215 184.575 18.425 185.095 ;
        RECT 20.190 184.670 20.540 185.920 ;
        RECT 24.115 185.190 24.405 186.355 ;
        RECT 24.575 185.265 25.785 186.355 ;
        RECT 14.455 183.805 15.665 184.555 ;
        RECT 15.835 183.805 18.425 184.575 ;
        RECT 22.020 184.350 22.360 185.180 ;
        RECT 24.575 184.725 25.095 185.265 ;
        RECT 25.960 185.165 26.215 186.045 ;
        RECT 26.385 185.215 26.690 186.355 ;
        RECT 27.030 185.975 27.360 186.355 ;
        RECT 27.540 185.805 27.710 186.095 ;
        RECT 27.880 185.895 28.130 186.355 ;
        RECT 26.910 185.635 27.710 185.805 ;
        RECT 28.300 185.845 29.170 186.185 ;
        RECT 25.265 184.555 25.785 185.095 ;
        RECT 18.600 183.805 23.945 184.350 ;
        RECT 24.115 183.805 24.405 184.530 ;
        RECT 24.575 183.805 25.785 184.555 ;
        RECT 25.960 184.515 26.170 185.165 ;
        RECT 26.910 185.045 27.080 185.635 ;
        RECT 28.300 185.465 28.470 185.845 ;
        RECT 29.405 185.725 29.575 186.185 ;
        RECT 29.745 185.895 30.115 186.355 ;
        RECT 30.410 185.755 30.580 186.095 ;
        RECT 30.750 185.925 31.080 186.355 ;
        RECT 31.315 185.755 31.485 186.095 ;
        RECT 27.250 185.295 28.470 185.465 ;
        RECT 28.640 185.385 29.100 185.675 ;
        RECT 29.405 185.555 29.965 185.725 ;
        RECT 30.410 185.585 31.485 185.755 ;
        RECT 31.655 185.855 32.335 186.185 ;
        RECT 32.550 185.855 32.800 186.185 ;
        RECT 32.970 185.895 33.220 186.355 ;
        RECT 29.795 185.415 29.965 185.555 ;
        RECT 28.640 185.375 29.605 185.385 ;
        RECT 28.300 185.205 28.470 185.295 ;
        RECT 28.930 185.215 29.605 185.375 ;
        RECT 26.340 185.015 27.080 185.045 ;
        RECT 26.340 184.715 27.255 185.015 ;
        RECT 26.930 184.540 27.255 184.715 ;
        RECT 25.960 183.985 26.215 184.515 ;
        RECT 26.385 183.805 26.690 184.265 ;
        RECT 26.935 184.185 27.255 184.540 ;
        RECT 27.425 184.755 27.965 185.125 ;
        RECT 28.300 185.035 28.705 185.205 ;
        RECT 27.425 184.355 27.665 184.755 ;
        RECT 28.145 184.585 28.365 184.865 ;
        RECT 27.835 184.415 28.365 184.585 ;
        RECT 27.835 184.185 28.005 184.415 ;
        RECT 28.535 184.255 28.705 185.035 ;
        RECT 28.875 184.425 29.225 185.045 ;
        RECT 29.395 184.425 29.605 185.215 ;
        RECT 29.795 185.245 31.295 185.415 ;
        RECT 29.795 184.555 29.965 185.245 ;
        RECT 31.655 185.075 31.825 185.855 ;
        RECT 32.630 185.725 32.800 185.855 ;
        RECT 30.135 184.905 31.825 185.075 ;
        RECT 31.995 185.295 32.460 185.685 ;
        RECT 32.630 185.555 33.025 185.725 ;
        RECT 30.135 184.725 30.305 184.905 ;
        RECT 26.935 184.015 28.005 184.185 ;
        RECT 28.175 183.805 28.365 184.245 ;
        RECT 28.535 183.975 29.485 184.255 ;
        RECT 29.795 184.165 30.055 184.555 ;
        RECT 30.475 184.485 31.265 184.735 ;
        RECT 29.705 183.995 30.055 184.165 ;
        RECT 30.265 183.805 30.595 184.265 ;
        RECT 31.470 184.195 31.640 184.905 ;
        RECT 31.995 184.705 32.165 185.295 ;
        RECT 31.810 184.485 32.165 184.705 ;
        RECT 32.335 184.485 32.685 185.105 ;
        RECT 32.855 184.195 33.025 185.555 ;
        RECT 33.390 185.385 33.715 186.170 ;
        RECT 33.195 184.335 33.655 185.385 ;
        RECT 31.470 184.025 32.325 184.195 ;
        RECT 32.530 184.025 33.025 184.195 ;
        RECT 33.195 183.805 33.525 184.165 ;
        RECT 33.885 184.065 34.055 186.185 ;
        RECT 34.225 185.855 34.555 186.355 ;
        RECT 34.725 185.685 34.980 186.185 ;
        RECT 34.230 185.515 34.980 185.685 ;
        RECT 34.230 184.525 34.460 185.515 ;
        RECT 34.630 184.695 34.980 185.345 ;
        RECT 35.615 185.265 38.205 186.355 ;
        RECT 35.615 184.745 36.825 185.265 ;
        RECT 38.415 185.215 38.645 186.355 ;
        RECT 38.815 185.205 39.145 186.185 ;
        RECT 39.315 185.215 39.525 186.355 ;
        RECT 39.755 185.595 40.270 186.005 ;
        RECT 40.505 185.595 40.675 186.355 ;
        RECT 40.845 186.015 42.875 186.185 ;
        RECT 36.995 184.575 38.205 185.095 ;
        RECT 38.395 184.795 38.725 185.045 ;
        RECT 34.230 184.355 34.980 184.525 ;
        RECT 34.225 183.805 34.555 184.185 ;
        RECT 34.725 184.065 34.980 184.355 ;
        RECT 35.615 183.805 38.205 184.575 ;
        RECT 38.415 183.805 38.645 184.625 ;
        RECT 38.895 184.605 39.145 185.205 ;
        RECT 39.755 184.785 40.095 185.595 ;
        RECT 40.845 185.350 41.015 186.015 ;
        RECT 41.410 185.675 42.535 185.845 ;
        RECT 40.265 185.160 41.015 185.350 ;
        RECT 41.185 185.335 42.195 185.505 ;
        RECT 38.815 183.975 39.145 184.605 ;
        RECT 39.315 183.805 39.525 184.625 ;
        RECT 39.755 184.615 40.985 184.785 ;
        RECT 40.030 184.010 40.275 184.615 ;
        RECT 40.495 183.805 41.005 184.340 ;
        RECT 41.185 183.975 41.375 185.335 ;
        RECT 41.545 184.315 41.820 185.135 ;
        RECT 42.025 184.535 42.195 185.335 ;
        RECT 42.365 184.545 42.535 185.675 ;
        RECT 42.705 185.045 42.875 186.015 ;
        RECT 43.045 185.215 43.215 186.355 ;
        RECT 43.385 185.215 43.720 186.185 ;
        RECT 42.705 184.715 42.900 185.045 ;
        RECT 43.125 184.715 43.380 185.045 ;
        RECT 43.125 184.545 43.295 184.715 ;
        RECT 43.550 184.545 43.720 185.215 ;
        RECT 42.365 184.375 43.295 184.545 ;
        RECT 42.365 184.340 42.540 184.375 ;
        RECT 41.545 184.145 41.825 184.315 ;
        RECT 41.545 183.975 41.820 184.145 ;
        RECT 42.010 183.975 42.540 184.340 ;
        RECT 42.965 183.805 43.295 184.205 ;
        RECT 43.465 183.975 43.720 184.545 ;
        RECT 43.900 185.215 44.235 186.185 ;
        RECT 44.405 185.215 44.575 186.355 ;
        RECT 44.745 186.015 46.775 186.185 ;
        RECT 43.900 184.545 44.070 185.215 ;
        RECT 44.745 185.045 44.915 186.015 ;
        RECT 44.240 184.715 44.495 185.045 ;
        RECT 44.720 184.715 44.915 185.045 ;
        RECT 45.085 185.675 46.210 185.845 ;
        RECT 44.325 184.545 44.495 184.715 ;
        RECT 45.085 184.545 45.255 185.675 ;
        RECT 43.900 183.975 44.155 184.545 ;
        RECT 44.325 184.375 45.255 184.545 ;
        RECT 45.425 185.335 46.435 185.505 ;
        RECT 45.425 184.535 45.595 185.335 ;
        RECT 45.080 184.340 45.255 184.375 ;
        RECT 44.325 183.805 44.655 184.205 ;
        RECT 45.080 183.975 45.610 184.340 ;
        RECT 45.800 184.315 46.075 185.135 ;
        RECT 45.795 184.145 46.075 184.315 ;
        RECT 45.800 183.975 46.075 184.145 ;
        RECT 46.245 183.975 46.435 185.335 ;
        RECT 46.605 185.350 46.775 186.015 ;
        RECT 46.945 185.595 47.115 186.355 ;
        RECT 47.350 185.595 47.865 186.005 ;
        RECT 46.605 185.160 47.355 185.350 ;
        RECT 47.525 184.785 47.865 185.595 ;
        RECT 48.535 185.215 48.765 186.355 ;
        RECT 48.935 185.205 49.265 186.185 ;
        RECT 49.435 185.215 49.645 186.355 ;
        RECT 48.515 184.795 48.845 185.045 ;
        RECT 46.635 184.615 47.865 184.785 ;
        RECT 46.615 183.805 47.125 184.340 ;
        RECT 47.345 184.010 47.590 184.615 ;
        RECT 48.535 183.805 48.765 184.625 ;
        RECT 49.015 184.605 49.265 185.205 ;
        RECT 49.875 185.190 50.165 186.355 ;
        RECT 50.340 185.165 50.595 186.045 ;
        RECT 50.765 185.215 51.070 186.355 ;
        RECT 51.410 185.975 51.740 186.355 ;
        RECT 51.920 185.805 52.090 186.095 ;
        RECT 52.260 185.895 52.510 186.355 ;
        RECT 51.290 185.635 52.090 185.805 ;
        RECT 52.680 185.845 53.550 186.185 ;
        RECT 48.935 183.975 49.265 184.605 ;
        RECT 49.435 183.805 49.645 184.625 ;
        RECT 49.875 183.805 50.165 184.530 ;
        RECT 50.340 184.515 50.550 185.165 ;
        RECT 51.290 185.045 51.460 185.635 ;
        RECT 52.680 185.465 52.850 185.845 ;
        RECT 53.785 185.725 53.955 186.185 ;
        RECT 54.125 185.895 54.495 186.355 ;
        RECT 54.790 185.755 54.960 186.095 ;
        RECT 55.130 185.925 55.460 186.355 ;
        RECT 55.695 185.755 55.865 186.095 ;
        RECT 51.630 185.295 52.850 185.465 ;
        RECT 53.020 185.385 53.480 185.675 ;
        RECT 53.785 185.555 54.345 185.725 ;
        RECT 54.790 185.585 55.865 185.755 ;
        RECT 56.035 185.855 56.715 186.185 ;
        RECT 56.930 185.855 57.180 186.185 ;
        RECT 57.350 185.895 57.600 186.355 ;
        RECT 54.175 185.415 54.345 185.555 ;
        RECT 53.020 185.375 53.985 185.385 ;
        RECT 52.680 185.205 52.850 185.295 ;
        RECT 53.310 185.215 53.985 185.375 ;
        RECT 50.720 185.015 51.460 185.045 ;
        RECT 50.720 184.715 51.635 185.015 ;
        RECT 51.310 184.540 51.635 184.715 ;
        RECT 50.340 183.985 50.595 184.515 ;
        RECT 50.765 183.805 51.070 184.265 ;
        RECT 51.315 184.185 51.635 184.540 ;
        RECT 51.805 184.755 52.345 185.125 ;
        RECT 52.680 185.035 53.085 185.205 ;
        RECT 51.805 184.355 52.045 184.755 ;
        RECT 52.525 184.585 52.745 184.865 ;
        RECT 52.215 184.415 52.745 184.585 ;
        RECT 52.215 184.185 52.385 184.415 ;
        RECT 52.915 184.255 53.085 185.035 ;
        RECT 53.255 184.425 53.605 185.045 ;
        RECT 53.775 184.425 53.985 185.215 ;
        RECT 54.175 185.245 55.675 185.415 ;
        RECT 54.175 184.555 54.345 185.245 ;
        RECT 56.035 185.075 56.205 185.855 ;
        RECT 57.010 185.725 57.180 185.855 ;
        RECT 54.515 184.905 56.205 185.075 ;
        RECT 56.375 185.295 56.840 185.685 ;
        RECT 57.010 185.555 57.405 185.725 ;
        RECT 54.515 184.725 54.685 184.905 ;
        RECT 51.315 184.015 52.385 184.185 ;
        RECT 52.555 183.805 52.745 184.245 ;
        RECT 52.915 183.975 53.865 184.255 ;
        RECT 54.175 184.165 54.435 184.555 ;
        RECT 54.855 184.485 55.645 184.735 ;
        RECT 54.085 183.995 54.435 184.165 ;
        RECT 54.645 183.805 54.975 184.265 ;
        RECT 55.850 184.195 56.020 184.905 ;
        RECT 56.375 184.705 56.545 185.295 ;
        RECT 56.190 184.485 56.545 184.705 ;
        RECT 56.715 184.485 57.065 185.105 ;
        RECT 57.235 184.195 57.405 185.555 ;
        RECT 57.770 185.385 58.095 186.170 ;
        RECT 57.575 184.335 58.035 185.385 ;
        RECT 55.850 184.025 56.705 184.195 ;
        RECT 56.910 184.025 57.405 184.195 ;
        RECT 57.575 183.805 57.905 184.165 ;
        RECT 58.265 184.065 58.435 186.185 ;
        RECT 58.605 185.855 58.935 186.355 ;
        RECT 59.105 185.685 59.360 186.185 ;
        RECT 60.000 185.920 65.345 186.355 ;
        RECT 65.520 185.920 70.865 186.355 ;
        RECT 58.610 185.515 59.360 185.685 ;
        RECT 58.610 184.525 58.840 185.515 ;
        RECT 59.010 184.695 59.360 185.345 ;
        RECT 61.590 184.670 61.940 185.920 ;
        RECT 58.610 184.355 59.360 184.525 ;
        RECT 58.605 183.805 58.935 184.185 ;
        RECT 59.105 184.065 59.360 184.355 ;
        RECT 63.420 184.350 63.760 185.180 ;
        RECT 67.110 184.670 67.460 185.920 ;
        RECT 68.940 184.350 69.280 185.180 ;
        RECT 60.000 183.805 65.345 184.350 ;
        RECT 65.520 183.805 70.865 184.350 ;
        RECT 71.035 183.975 71.295 186.185 ;
        RECT 71.465 185.975 71.795 186.355 ;
        RECT 72.220 185.805 72.390 186.185 ;
        RECT 72.650 185.975 72.980 186.355 ;
        RECT 73.175 185.805 73.345 186.185 ;
        RECT 73.555 185.975 73.885 186.355 ;
        RECT 74.135 185.805 74.325 186.185 ;
        RECT 74.565 185.975 74.895 186.355 ;
        RECT 75.205 185.855 75.465 186.185 ;
        RECT 71.465 185.635 73.415 185.805 ;
        RECT 71.465 184.715 71.635 185.635 ;
        RECT 72.005 185.045 72.200 185.355 ;
        RECT 72.470 185.045 72.655 185.355 ;
        RECT 71.945 184.715 72.200 185.045 ;
        RECT 72.425 184.715 72.655 185.045 ;
        RECT 71.465 183.805 71.795 184.185 ;
        RECT 72.005 184.140 72.200 184.715 ;
        RECT 72.470 184.135 72.655 184.715 ;
        RECT 72.905 184.145 73.075 185.045 ;
        RECT 73.245 184.645 73.415 185.635 ;
        RECT 73.585 185.635 74.325 185.805 ;
        RECT 73.585 185.125 73.755 185.635 ;
        RECT 73.925 185.295 74.505 185.465 ;
        RECT 74.775 185.345 75.125 185.675 ;
        RECT 74.335 185.175 74.505 185.295 ;
        RECT 75.295 185.175 75.465 185.855 ;
        RECT 75.635 185.190 75.925 186.355 ;
        RECT 76.095 185.265 78.685 186.355 ;
        RECT 78.860 185.920 84.205 186.355 ;
        RECT 73.585 184.955 74.155 185.125 ;
        RECT 74.335 185.005 75.465 185.175 ;
        RECT 73.245 184.315 73.795 184.645 ;
        RECT 73.985 184.475 74.155 184.955 ;
        RECT 74.325 184.665 74.945 184.835 ;
        RECT 74.735 184.485 74.945 184.665 ;
        RECT 73.985 184.145 74.385 184.475 ;
        RECT 75.295 184.305 75.465 185.005 ;
        RECT 76.095 184.745 77.305 185.265 ;
        RECT 77.475 184.575 78.685 185.095 ;
        RECT 80.450 184.670 80.800 185.920 ;
        RECT 84.375 185.595 84.890 186.005 ;
        RECT 85.125 185.595 85.295 186.355 ;
        RECT 85.465 186.015 87.495 186.185 ;
        RECT 72.905 183.975 74.385 184.145 ;
        RECT 74.565 183.805 74.895 184.185 ;
        RECT 75.205 183.975 75.465 184.305 ;
        RECT 75.635 183.805 75.925 184.530 ;
        RECT 76.095 183.805 78.685 184.575 ;
        RECT 82.280 184.350 82.620 185.180 ;
        RECT 84.375 184.785 84.715 185.595 ;
        RECT 85.465 185.350 85.635 186.015 ;
        RECT 86.030 185.675 87.155 185.845 ;
        RECT 84.885 185.160 85.635 185.350 ;
        RECT 85.805 185.335 86.815 185.505 ;
        RECT 84.375 184.615 85.605 184.785 ;
        RECT 78.860 183.805 84.205 184.350 ;
        RECT 84.650 184.010 84.895 184.615 ;
        RECT 85.115 183.805 85.625 184.340 ;
        RECT 85.805 183.975 85.995 185.335 ;
        RECT 86.165 184.315 86.440 185.135 ;
        RECT 86.645 184.535 86.815 185.335 ;
        RECT 86.985 184.545 87.155 185.675 ;
        RECT 87.325 185.045 87.495 186.015 ;
        RECT 87.665 185.215 87.835 186.355 ;
        RECT 88.005 185.215 88.340 186.185 ;
        RECT 88.520 185.920 93.865 186.355 ;
        RECT 87.325 184.715 87.520 185.045 ;
        RECT 87.745 184.715 88.000 185.045 ;
        RECT 87.745 184.545 87.915 184.715 ;
        RECT 88.170 184.545 88.340 185.215 ;
        RECT 90.110 184.670 90.460 185.920 ;
        RECT 94.150 185.725 94.435 186.185 ;
        RECT 94.605 185.895 94.875 186.355 ;
        RECT 94.150 185.505 95.105 185.725 ;
        RECT 86.985 184.375 87.915 184.545 ;
        RECT 86.985 184.340 87.160 184.375 ;
        RECT 86.165 184.145 86.445 184.315 ;
        RECT 86.165 183.975 86.440 184.145 ;
        RECT 86.630 183.975 87.160 184.340 ;
        RECT 87.585 183.805 87.915 184.205 ;
        RECT 88.085 183.975 88.340 184.545 ;
        RECT 91.940 184.350 92.280 185.180 ;
        RECT 94.035 184.775 94.725 185.335 ;
        RECT 94.895 184.605 95.105 185.505 ;
        RECT 94.150 184.435 95.105 184.605 ;
        RECT 95.275 185.335 95.675 186.185 ;
        RECT 95.865 185.725 96.145 186.185 ;
        RECT 96.665 185.895 96.990 186.355 ;
        RECT 95.865 185.505 96.990 185.725 ;
        RECT 95.275 184.775 96.370 185.335 ;
        RECT 96.540 185.045 96.990 185.505 ;
        RECT 97.160 185.215 97.545 186.185 ;
        RECT 98.725 185.425 98.895 186.185 ;
        RECT 99.075 185.595 99.405 186.355 ;
        RECT 98.725 185.255 99.390 185.425 ;
        RECT 99.575 185.280 99.845 186.185 ;
        RECT 88.520 183.805 93.865 184.350 ;
        RECT 94.150 183.975 94.435 184.435 ;
        RECT 94.605 183.805 94.875 184.265 ;
        RECT 95.275 183.975 95.675 184.775 ;
        RECT 96.540 184.715 97.095 185.045 ;
        RECT 96.540 184.605 96.990 184.715 ;
        RECT 95.865 184.435 96.990 184.605 ;
        RECT 97.265 184.545 97.545 185.215 ;
        RECT 99.220 185.110 99.390 185.255 ;
        RECT 98.655 184.705 98.985 185.075 ;
        RECT 99.220 184.780 99.505 185.110 ;
        RECT 95.865 183.975 96.145 184.435 ;
        RECT 96.665 183.805 96.990 184.265 ;
        RECT 97.160 183.975 97.545 184.545 ;
        RECT 99.220 184.525 99.390 184.780 ;
        RECT 98.725 184.355 99.390 184.525 ;
        RECT 99.675 184.480 99.845 185.280 ;
        RECT 100.055 185.215 100.285 186.355 ;
        RECT 100.455 185.205 100.785 186.185 ;
        RECT 100.955 185.215 101.165 186.355 ;
        RECT 100.035 184.795 100.365 185.045 ;
        RECT 98.725 183.975 98.895 184.355 ;
        RECT 99.075 183.805 99.405 184.185 ;
        RECT 99.585 183.975 99.845 184.480 ;
        RECT 100.055 183.805 100.285 184.625 ;
        RECT 100.535 184.605 100.785 185.205 ;
        RECT 101.395 185.190 101.685 186.355 ;
        RECT 102.315 185.215 102.700 186.185 ;
        RECT 102.870 185.895 103.195 186.355 ;
        RECT 103.715 185.725 103.995 186.185 ;
        RECT 102.870 185.505 103.995 185.725 ;
        RECT 100.455 183.975 100.785 184.605 ;
        RECT 100.955 183.805 101.165 184.625 ;
        RECT 102.315 184.545 102.595 185.215 ;
        RECT 102.870 185.045 103.320 185.505 ;
        RECT 104.185 185.335 104.585 186.185 ;
        RECT 104.985 185.895 105.255 186.355 ;
        RECT 105.425 185.725 105.710 186.185 ;
        RECT 102.765 184.715 103.320 185.045 ;
        RECT 103.490 184.775 104.585 185.335 ;
        RECT 102.870 184.605 103.320 184.715 ;
        RECT 101.395 183.805 101.685 184.530 ;
        RECT 102.315 183.975 102.700 184.545 ;
        RECT 102.870 184.435 103.995 184.605 ;
        RECT 102.870 183.805 103.195 184.265 ;
        RECT 103.715 183.975 103.995 184.435 ;
        RECT 104.185 183.975 104.585 184.775 ;
        RECT 104.755 185.505 105.710 185.725 ;
        RECT 106.570 185.725 106.855 186.185 ;
        RECT 107.025 185.895 107.295 186.355 ;
        RECT 106.570 185.505 107.525 185.725 ;
        RECT 104.755 184.605 104.965 185.505 ;
        RECT 105.135 184.775 105.825 185.335 ;
        RECT 106.455 184.775 107.145 185.335 ;
        RECT 107.315 184.605 107.525 185.505 ;
        RECT 104.755 184.435 105.710 184.605 ;
        RECT 104.985 183.805 105.255 184.265 ;
        RECT 105.425 183.975 105.710 184.435 ;
        RECT 106.570 184.435 107.525 184.605 ;
        RECT 107.695 185.335 108.095 186.185 ;
        RECT 108.285 185.725 108.565 186.185 ;
        RECT 109.085 185.895 109.410 186.355 ;
        RECT 108.285 185.505 109.410 185.725 ;
        RECT 107.695 184.775 108.790 185.335 ;
        RECT 108.960 185.045 109.410 185.505 ;
        RECT 109.580 185.215 109.965 186.185 ;
        RECT 110.250 185.725 110.535 186.185 ;
        RECT 110.705 185.895 110.975 186.355 ;
        RECT 110.250 185.505 111.205 185.725 ;
        RECT 106.570 183.975 106.855 184.435 ;
        RECT 107.025 183.805 107.295 184.265 ;
        RECT 107.695 183.975 108.095 184.775 ;
        RECT 108.960 184.715 109.515 185.045 ;
        RECT 108.960 184.605 109.410 184.715 ;
        RECT 108.285 184.435 109.410 184.605 ;
        RECT 109.685 184.545 109.965 185.215 ;
        RECT 110.135 184.775 110.825 185.335 ;
        RECT 110.995 184.605 111.205 185.505 ;
        RECT 108.285 183.975 108.565 184.435 ;
        RECT 109.085 183.805 109.410 184.265 ;
        RECT 109.580 183.975 109.965 184.545 ;
        RECT 110.250 184.435 111.205 184.605 ;
        RECT 111.375 185.335 111.775 186.185 ;
        RECT 111.965 185.725 112.245 186.185 ;
        RECT 112.765 185.895 113.090 186.355 ;
        RECT 111.965 185.505 113.090 185.725 ;
        RECT 111.375 184.775 112.470 185.335 ;
        RECT 112.640 185.045 113.090 185.505 ;
        RECT 113.260 185.215 113.645 186.185 ;
        RECT 110.250 183.975 110.535 184.435 ;
        RECT 110.705 183.805 110.975 184.265 ;
        RECT 111.375 183.975 111.775 184.775 ;
        RECT 112.640 184.715 113.195 185.045 ;
        RECT 112.640 184.605 113.090 184.715 ;
        RECT 111.965 184.435 113.090 184.605 ;
        RECT 113.365 184.545 113.645 185.215 ;
        RECT 113.815 185.265 115.025 186.355 ;
        RECT 115.200 185.920 120.545 186.355 ;
        RECT 120.720 185.920 126.065 186.355 ;
        RECT 113.815 184.725 114.335 185.265 ;
        RECT 114.505 184.555 115.025 185.095 ;
        RECT 116.790 184.670 117.140 185.920 ;
        RECT 111.965 183.975 112.245 184.435 ;
        RECT 112.765 183.805 113.090 184.265 ;
        RECT 113.260 183.975 113.645 184.545 ;
        RECT 113.815 183.805 115.025 184.555 ;
        RECT 118.620 184.350 118.960 185.180 ;
        RECT 122.310 184.670 122.660 185.920 ;
        RECT 126.235 185.265 127.445 186.355 ;
        RECT 124.140 184.350 124.480 185.180 ;
        RECT 126.235 184.725 126.755 185.265 ;
        RECT 126.925 184.555 127.445 185.095 ;
        RECT 115.200 183.805 120.545 184.350 ;
        RECT 120.720 183.805 126.065 184.350 ;
        RECT 126.235 183.805 127.445 184.555 ;
        RECT 14.370 183.635 127.530 183.805 ;
        RECT 14.455 182.885 15.665 183.635 ;
        RECT 16.300 183.090 21.645 183.635 ;
        RECT 14.455 182.345 14.975 182.885 ;
        RECT 15.145 182.175 15.665 182.715 ;
        RECT 14.455 181.085 15.665 182.175 ;
        RECT 17.890 181.520 18.240 182.770 ;
        RECT 19.720 182.260 20.060 183.090 ;
        RECT 21.905 183.085 22.075 183.465 ;
        RECT 22.255 183.255 22.585 183.635 ;
        RECT 21.905 182.915 22.570 183.085 ;
        RECT 22.765 182.960 23.025 183.465 ;
        RECT 21.835 182.365 22.165 182.735 ;
        RECT 22.400 182.660 22.570 182.915 ;
        RECT 22.400 182.330 22.685 182.660 ;
        RECT 22.400 182.185 22.570 182.330 ;
        RECT 21.905 182.015 22.570 182.185 ;
        RECT 22.855 182.160 23.025 182.960 ;
        RECT 16.300 181.085 21.645 181.520 ;
        RECT 21.905 181.255 22.075 182.015 ;
        RECT 22.255 181.085 22.585 181.845 ;
        RECT 22.755 181.255 23.025 182.160 ;
        RECT 23.195 182.895 23.580 183.465 ;
        RECT 23.750 183.175 24.075 183.635 ;
        RECT 24.595 183.005 24.875 183.465 ;
        RECT 23.195 182.225 23.475 182.895 ;
        RECT 23.750 182.835 24.875 183.005 ;
        RECT 23.750 182.725 24.200 182.835 ;
        RECT 23.645 182.395 24.200 182.725 ;
        RECT 25.065 182.665 25.465 183.465 ;
        RECT 25.865 183.175 26.135 183.635 ;
        RECT 26.305 183.005 26.590 183.465 ;
        RECT 23.195 181.255 23.580 182.225 ;
        RECT 23.750 181.935 24.200 182.395 ;
        RECT 24.370 182.105 25.465 182.665 ;
        RECT 23.750 181.715 24.875 181.935 ;
        RECT 23.750 181.085 24.075 181.545 ;
        RECT 24.595 181.255 24.875 181.715 ;
        RECT 25.065 181.255 25.465 182.105 ;
        RECT 25.635 182.835 26.590 183.005 ;
        RECT 26.990 183.005 27.275 183.465 ;
        RECT 27.445 183.175 27.715 183.635 ;
        RECT 26.990 182.835 27.945 183.005 ;
        RECT 25.635 181.935 25.845 182.835 ;
        RECT 26.015 182.105 26.705 182.665 ;
        RECT 26.875 182.105 27.565 182.665 ;
        RECT 27.735 181.935 27.945 182.835 ;
        RECT 25.635 181.715 26.590 181.935 ;
        RECT 25.865 181.085 26.135 181.545 ;
        RECT 26.305 181.255 26.590 181.715 ;
        RECT 26.990 181.715 27.945 181.935 ;
        RECT 28.115 182.665 28.515 183.465 ;
        RECT 28.705 183.005 28.985 183.465 ;
        RECT 29.505 183.175 29.830 183.635 ;
        RECT 28.705 182.835 29.830 183.005 ;
        RECT 30.000 182.895 30.385 183.465 ;
        RECT 29.380 182.725 29.830 182.835 ;
        RECT 28.115 182.105 29.210 182.665 ;
        RECT 29.380 182.395 29.935 182.725 ;
        RECT 26.990 181.255 27.275 181.715 ;
        RECT 27.445 181.085 27.715 181.545 ;
        RECT 28.115 181.255 28.515 182.105 ;
        RECT 29.380 181.935 29.830 182.395 ;
        RECT 30.105 182.225 30.385 182.895 ;
        RECT 28.705 181.715 29.830 181.935 ;
        RECT 28.705 181.255 28.985 181.715 ;
        RECT 29.505 181.085 29.830 181.545 ;
        RECT 30.000 181.255 30.385 182.225 ;
        RECT 30.560 182.895 30.815 183.465 ;
        RECT 30.985 183.235 31.315 183.635 ;
        RECT 31.740 183.100 32.270 183.465 ;
        RECT 31.740 183.065 31.915 183.100 ;
        RECT 30.985 182.895 31.915 183.065 ;
        RECT 32.460 182.955 32.735 183.465 ;
        RECT 30.560 182.225 30.730 182.895 ;
        RECT 30.985 182.725 31.155 182.895 ;
        RECT 30.900 182.395 31.155 182.725 ;
        RECT 31.380 182.395 31.575 182.725 ;
        RECT 30.560 181.255 30.895 182.225 ;
        RECT 31.065 181.085 31.235 182.225 ;
        RECT 31.405 181.425 31.575 182.395 ;
        RECT 31.745 181.765 31.915 182.895 ;
        RECT 32.085 182.105 32.255 182.905 ;
        RECT 32.455 182.785 32.735 182.955 ;
        RECT 32.460 182.305 32.735 182.785 ;
        RECT 32.905 182.105 33.095 183.465 ;
        RECT 33.275 183.100 33.785 183.635 ;
        RECT 34.005 182.825 34.250 183.430 ;
        RECT 35.155 182.865 36.825 183.635 ;
        RECT 36.995 182.910 37.285 183.635 ;
        RECT 37.570 183.005 37.855 183.465 ;
        RECT 38.025 183.175 38.295 183.635 ;
        RECT 33.295 182.655 34.525 182.825 ;
        RECT 32.085 181.935 33.095 182.105 ;
        RECT 33.265 182.090 34.015 182.280 ;
        RECT 31.745 181.595 32.870 181.765 ;
        RECT 33.265 181.425 33.435 182.090 ;
        RECT 34.185 181.845 34.525 182.655 ;
        RECT 31.405 181.255 33.435 181.425 ;
        RECT 33.605 181.085 33.775 181.845 ;
        RECT 34.010 181.435 34.525 181.845 ;
        RECT 35.155 182.175 35.905 182.695 ;
        RECT 36.075 182.345 36.825 182.865 ;
        RECT 37.570 182.835 38.525 183.005 ;
        RECT 35.155 181.085 36.825 182.175 ;
        RECT 36.995 181.085 37.285 182.250 ;
        RECT 37.455 182.105 38.145 182.665 ;
        RECT 38.315 181.935 38.525 182.835 ;
        RECT 37.570 181.715 38.525 181.935 ;
        RECT 38.695 182.665 39.095 183.465 ;
        RECT 39.285 183.005 39.565 183.465 ;
        RECT 40.085 183.175 40.410 183.635 ;
        RECT 39.285 182.835 40.410 183.005 ;
        RECT 40.580 182.895 40.965 183.465 ;
        RECT 39.960 182.725 40.410 182.835 ;
        RECT 38.695 182.105 39.790 182.665 ;
        RECT 39.960 182.395 40.515 182.725 ;
        RECT 37.570 181.255 37.855 181.715 ;
        RECT 38.025 181.085 38.295 181.545 ;
        RECT 38.695 181.255 39.095 182.105 ;
        RECT 39.960 181.935 40.410 182.395 ;
        RECT 40.685 182.225 40.965 182.895 ;
        RECT 41.250 183.005 41.535 183.465 ;
        RECT 41.705 183.175 41.975 183.635 ;
        RECT 41.250 182.835 42.205 183.005 ;
        RECT 39.285 181.715 40.410 181.935 ;
        RECT 39.285 181.255 39.565 181.715 ;
        RECT 40.085 181.085 40.410 181.545 ;
        RECT 40.580 181.255 40.965 182.225 ;
        RECT 41.135 182.105 41.825 182.665 ;
        RECT 41.995 181.935 42.205 182.835 ;
        RECT 41.250 181.715 42.205 181.935 ;
        RECT 42.375 182.665 42.775 183.465 ;
        RECT 42.965 183.005 43.245 183.465 ;
        RECT 43.765 183.175 44.090 183.635 ;
        RECT 42.965 182.835 44.090 183.005 ;
        RECT 44.260 182.895 44.645 183.465 ;
        RECT 43.640 182.725 44.090 182.835 ;
        RECT 42.375 182.105 43.470 182.665 ;
        RECT 43.640 182.395 44.195 182.725 ;
        RECT 41.250 181.255 41.535 181.715 ;
        RECT 41.705 181.085 41.975 181.545 ;
        RECT 42.375 181.255 42.775 182.105 ;
        RECT 43.640 181.935 44.090 182.395 ;
        RECT 44.365 182.225 44.645 182.895 ;
        RECT 44.930 183.005 45.215 183.465 ;
        RECT 45.385 183.175 45.655 183.635 ;
        RECT 44.930 182.835 45.885 183.005 ;
        RECT 42.965 181.715 44.090 181.935 ;
        RECT 42.965 181.255 43.245 181.715 ;
        RECT 43.765 181.085 44.090 181.545 ;
        RECT 44.260 181.255 44.645 182.225 ;
        RECT 44.815 182.105 45.505 182.665 ;
        RECT 45.675 181.935 45.885 182.835 ;
        RECT 44.930 181.715 45.885 181.935 ;
        RECT 46.055 182.665 46.455 183.465 ;
        RECT 46.645 183.005 46.925 183.465 ;
        RECT 47.445 183.175 47.770 183.635 ;
        RECT 46.645 182.835 47.770 183.005 ;
        RECT 47.940 182.895 48.325 183.465 ;
        RECT 47.320 182.725 47.770 182.835 ;
        RECT 46.055 182.105 47.150 182.665 ;
        RECT 47.320 182.395 47.875 182.725 ;
        RECT 44.930 181.255 45.215 181.715 ;
        RECT 45.385 181.085 45.655 181.545 ;
        RECT 46.055 181.255 46.455 182.105 ;
        RECT 47.320 181.935 47.770 182.395 ;
        RECT 48.045 182.225 48.325 182.895 ;
        RECT 46.645 181.715 47.770 181.935 ;
        RECT 46.645 181.255 46.925 181.715 ;
        RECT 47.445 181.085 47.770 181.545 ;
        RECT 47.940 181.255 48.325 182.225 ;
        RECT 48.495 182.960 48.755 183.465 ;
        RECT 48.935 183.255 49.265 183.635 ;
        RECT 49.445 183.085 49.615 183.465 ;
        RECT 48.495 182.160 48.665 182.960 ;
        RECT 48.950 182.915 49.615 183.085 ;
        RECT 49.875 182.960 50.135 183.465 ;
        RECT 50.315 183.255 50.645 183.635 ;
        RECT 50.825 183.085 50.995 183.465 ;
        RECT 48.950 182.660 49.120 182.915 ;
        RECT 48.835 182.330 49.120 182.660 ;
        RECT 49.355 182.365 49.685 182.735 ;
        RECT 48.950 182.185 49.120 182.330 ;
        RECT 48.495 181.255 48.765 182.160 ;
        RECT 48.950 182.015 49.615 182.185 ;
        RECT 48.935 181.085 49.265 181.845 ;
        RECT 49.445 181.255 49.615 182.015 ;
        RECT 49.875 182.160 50.045 182.960 ;
        RECT 50.330 182.915 50.995 183.085 ;
        RECT 51.345 183.085 51.515 183.465 ;
        RECT 51.695 183.255 52.025 183.635 ;
        RECT 51.345 182.915 52.010 183.085 ;
        RECT 52.205 182.960 52.465 183.465 ;
        RECT 52.735 183.170 52.985 183.635 ;
        RECT 53.155 182.995 53.325 183.465 ;
        RECT 53.575 183.175 53.745 183.635 ;
        RECT 53.995 182.995 54.165 183.465 ;
        RECT 54.415 183.175 54.585 183.635 ;
        RECT 54.835 182.995 55.005 183.465 ;
        RECT 55.375 183.175 55.640 183.635 ;
        RECT 50.330 182.660 50.500 182.915 ;
        RECT 50.215 182.330 50.500 182.660 ;
        RECT 50.735 182.365 51.065 182.735 ;
        RECT 51.275 182.365 51.605 182.735 ;
        RECT 51.840 182.660 52.010 182.915 ;
        RECT 50.330 182.185 50.500 182.330 ;
        RECT 51.840 182.330 52.125 182.660 ;
        RECT 51.840 182.185 52.010 182.330 ;
        RECT 49.875 181.255 50.145 182.160 ;
        RECT 50.330 182.015 50.995 182.185 ;
        RECT 50.315 181.085 50.645 181.845 ;
        RECT 50.825 181.255 50.995 182.015 ;
        RECT 51.345 182.015 52.010 182.185 ;
        RECT 52.295 182.160 52.465 182.960 ;
        RECT 51.345 181.255 51.515 182.015 ;
        RECT 51.695 181.085 52.025 181.845 ;
        RECT 52.195 181.255 52.465 182.160 ;
        RECT 52.635 182.815 55.005 182.995 ;
        RECT 56.315 182.865 58.905 183.635 ;
        RECT 52.635 182.225 52.985 182.815 ;
        RECT 53.155 182.395 55.665 182.645 ;
        RECT 52.635 182.055 55.085 182.225 ;
        RECT 52.635 182.035 53.405 182.055 ;
        RECT 52.735 181.085 52.905 181.545 ;
        RECT 53.075 181.255 53.405 182.035 ;
        RECT 53.575 181.085 53.745 181.885 ;
        RECT 53.915 181.255 54.245 182.055 ;
        RECT 54.415 181.085 54.585 181.885 ;
        RECT 54.755 181.255 55.085 182.055 ;
        RECT 55.345 181.085 55.640 182.225 ;
        RECT 56.315 182.175 57.525 182.695 ;
        RECT 57.695 182.345 58.905 182.865 ;
        RECT 59.135 182.815 59.345 183.635 ;
        RECT 59.515 182.835 59.845 183.465 ;
        RECT 59.515 182.235 59.765 182.835 ;
        RECT 60.015 182.815 60.245 183.635 ;
        RECT 60.915 182.865 62.585 183.635 ;
        RECT 62.755 182.910 63.045 183.635 ;
        RECT 63.675 182.865 66.265 183.635 ;
        RECT 66.705 183.240 67.035 183.635 ;
        RECT 67.205 183.065 67.405 183.420 ;
        RECT 67.575 183.235 67.905 183.635 ;
        RECT 68.075 183.065 68.275 183.410 ;
        RECT 59.935 182.395 60.265 182.645 ;
        RECT 56.315 181.085 58.905 182.175 ;
        RECT 59.135 181.085 59.345 182.225 ;
        RECT 59.515 181.255 59.845 182.235 ;
        RECT 60.015 181.085 60.245 182.225 ;
        RECT 60.915 182.175 61.665 182.695 ;
        RECT 61.835 182.345 62.585 182.865 ;
        RECT 60.915 181.085 62.585 182.175 ;
        RECT 62.755 181.085 63.045 182.250 ;
        RECT 63.675 182.175 64.885 182.695 ;
        RECT 65.055 182.345 66.265 182.865 ;
        RECT 66.435 182.895 68.275 183.065 ;
        RECT 68.445 182.895 68.775 183.635 ;
        RECT 69.010 183.065 69.180 183.315 ;
        RECT 69.010 182.895 69.485 183.065 ;
        RECT 63.675 181.085 66.265 182.175 ;
        RECT 66.435 181.270 66.695 182.895 ;
        RECT 66.875 181.925 67.095 182.725 ;
        RECT 67.335 182.105 67.635 182.725 ;
        RECT 67.805 182.105 68.135 182.725 ;
        RECT 68.305 182.105 68.625 182.725 ;
        RECT 68.795 182.105 69.145 182.725 ;
        RECT 69.315 181.925 69.485 182.895 ;
        RECT 69.655 182.815 69.915 183.635 ;
        RECT 70.085 182.995 70.415 183.465 ;
        RECT 70.585 183.165 70.755 183.635 ;
        RECT 70.925 182.995 71.255 183.465 ;
        RECT 71.425 183.165 72.150 183.635 ;
        RECT 72.320 182.995 72.650 183.465 ;
        RECT 72.820 183.165 72.990 183.635 ;
        RECT 73.160 182.995 73.490 183.465 ;
        RECT 70.085 182.815 73.490 182.995 ;
        RECT 73.660 182.825 73.865 183.635 ;
        RECT 73.285 182.645 73.490 182.815 ;
        RECT 74.035 182.815 74.390 183.340 ;
        RECT 74.560 182.895 74.810 183.635 ;
        RECT 75.480 183.065 75.650 183.315 ;
        RECT 75.175 182.895 75.650 183.065 ;
        RECT 75.885 182.895 76.215 183.635 ;
        RECT 76.385 183.065 76.585 183.410 ;
        RECT 76.755 183.235 77.085 183.635 ;
        RECT 77.255 183.065 77.455 183.420 ;
        RECT 77.625 183.240 77.955 183.635 ;
        RECT 76.385 182.895 78.225 183.065 ;
        RECT 74.035 182.645 74.205 182.815 ;
        RECT 69.670 182.435 70.810 182.645 ;
        RECT 70.990 182.435 72.205 182.645 ;
        RECT 72.385 182.435 73.105 182.645 ;
        RECT 73.285 182.265 73.605 182.645 ;
        RECT 73.890 182.475 74.205 182.645 ;
        RECT 66.875 181.715 69.485 181.925 ;
        RECT 69.655 182.095 71.675 182.265 ;
        RECT 68.445 181.085 68.775 181.535 ;
        RECT 69.655 181.255 69.995 182.095 ;
        RECT 70.165 181.085 70.375 181.925 ;
        RECT 70.545 181.255 70.795 182.095 ;
        RECT 70.965 181.425 71.175 181.925 ;
        RECT 71.345 181.595 71.675 182.095 ;
        RECT 71.845 182.095 73.030 182.265 ;
        RECT 71.845 181.595 72.230 182.095 ;
        RECT 72.400 181.425 72.610 181.925 ;
        RECT 70.965 181.255 72.610 181.425 ;
        RECT 72.780 181.425 73.030 182.095 ;
        RECT 73.200 182.095 73.605 182.265 ;
        RECT 73.200 181.595 73.450 182.095 ;
        RECT 73.620 181.425 73.865 181.925 ;
        RECT 72.780 181.255 73.865 181.425 ;
        RECT 74.035 181.685 74.205 182.475 ;
        RECT 74.375 182.435 75.005 182.645 ;
        RECT 74.755 181.765 75.005 182.435 ;
        RECT 75.175 181.925 75.345 182.895 ;
        RECT 75.515 182.105 75.865 182.725 ;
        RECT 76.035 182.105 76.355 182.725 ;
        RECT 76.525 182.105 76.855 182.725 ;
        RECT 77.025 182.105 77.325 182.725 ;
        RECT 77.565 181.925 77.785 182.725 ;
        RECT 75.175 181.715 77.785 181.925 ;
        RECT 74.035 181.270 74.390 181.685 ;
        RECT 74.560 181.085 74.810 181.585 ;
        RECT 75.885 181.085 76.215 181.535 ;
        RECT 77.965 181.270 78.225 182.895 ;
        RECT 79.320 182.925 79.575 183.455 ;
        RECT 79.745 183.175 80.050 183.635 ;
        RECT 80.295 183.255 81.365 183.425 ;
        RECT 79.320 182.275 79.530 182.925 ;
        RECT 80.295 182.900 80.615 183.255 ;
        RECT 80.290 182.725 80.615 182.900 ;
        RECT 79.700 182.425 80.615 182.725 ;
        RECT 80.785 182.685 81.025 183.085 ;
        RECT 81.195 183.025 81.365 183.255 ;
        RECT 81.535 183.195 81.725 183.635 ;
        RECT 81.895 183.185 82.845 183.465 ;
        RECT 83.065 183.275 83.415 183.445 ;
        RECT 81.195 182.855 81.725 183.025 ;
        RECT 79.700 182.395 80.440 182.425 ;
        RECT 79.320 181.395 79.575 182.275 ;
        RECT 79.745 181.085 80.050 182.225 ;
        RECT 80.270 181.805 80.440 182.395 ;
        RECT 80.785 182.315 81.325 182.685 ;
        RECT 81.505 182.575 81.725 182.855 ;
        RECT 81.895 182.405 82.065 183.185 ;
        RECT 81.660 182.235 82.065 182.405 ;
        RECT 82.235 182.395 82.585 183.015 ;
        RECT 81.660 182.145 81.830 182.235 ;
        RECT 82.755 182.225 82.965 183.015 ;
        RECT 80.610 181.975 81.830 182.145 ;
        RECT 82.290 182.065 82.965 182.225 ;
        RECT 80.270 181.635 81.070 181.805 ;
        RECT 80.390 181.085 80.720 181.465 ;
        RECT 80.900 181.345 81.070 181.635 ;
        RECT 81.660 181.595 81.830 181.975 ;
        RECT 82.000 182.055 82.965 182.065 ;
        RECT 83.155 182.885 83.415 183.275 ;
        RECT 83.625 183.175 83.955 183.635 ;
        RECT 84.830 183.245 85.685 183.415 ;
        RECT 85.890 183.245 86.385 183.415 ;
        RECT 86.555 183.275 86.885 183.635 ;
        RECT 83.155 182.195 83.325 182.885 ;
        RECT 83.495 182.535 83.665 182.715 ;
        RECT 83.835 182.705 84.625 182.955 ;
        RECT 84.830 182.535 85.000 183.245 ;
        RECT 85.170 182.735 85.525 182.955 ;
        RECT 83.495 182.365 85.185 182.535 ;
        RECT 82.000 181.765 82.460 182.055 ;
        RECT 83.155 182.025 84.655 182.195 ;
        RECT 83.155 181.885 83.325 182.025 ;
        RECT 82.765 181.715 83.325 181.885 ;
        RECT 81.240 181.085 81.490 181.545 ;
        RECT 81.660 181.255 82.530 181.595 ;
        RECT 82.765 181.255 82.935 181.715 ;
        RECT 83.770 181.685 84.845 181.855 ;
        RECT 83.105 181.085 83.475 181.545 ;
        RECT 83.770 181.345 83.940 181.685 ;
        RECT 84.110 181.085 84.440 181.515 ;
        RECT 84.675 181.345 84.845 181.685 ;
        RECT 85.015 181.585 85.185 182.365 ;
        RECT 85.355 182.145 85.525 182.735 ;
        RECT 85.695 182.335 86.045 182.955 ;
        RECT 85.355 181.755 85.820 182.145 ;
        RECT 86.215 181.885 86.385 183.245 ;
        RECT 86.555 182.055 87.015 183.105 ;
        RECT 85.990 181.715 86.385 181.885 ;
        RECT 85.990 181.585 86.160 181.715 ;
        RECT 85.015 181.255 85.695 181.585 ;
        RECT 85.910 181.255 86.160 181.585 ;
        RECT 86.330 181.085 86.580 181.545 ;
        RECT 86.750 181.270 87.075 182.055 ;
        RECT 87.245 181.255 87.415 183.375 ;
        RECT 87.585 183.255 87.915 183.635 ;
        RECT 88.085 183.085 88.340 183.375 ;
        RECT 87.590 182.915 88.340 183.085 ;
        RECT 87.590 181.925 87.820 182.915 ;
        RECT 88.515 182.910 88.805 183.635 ;
        RECT 89.035 182.815 89.245 183.635 ;
        RECT 89.415 182.835 89.745 183.465 ;
        RECT 87.990 182.095 88.340 182.745 ;
        RECT 87.590 181.755 88.340 181.925 ;
        RECT 87.585 181.085 87.915 181.585 ;
        RECT 88.085 181.255 88.340 181.755 ;
        RECT 88.515 181.085 88.805 182.250 ;
        RECT 89.415 182.235 89.665 182.835 ;
        RECT 89.915 182.815 90.145 183.635 ;
        RECT 90.355 182.885 91.565 183.635 ;
        RECT 89.835 182.395 90.165 182.645 ;
        RECT 89.035 181.085 89.245 182.225 ;
        RECT 89.415 181.255 89.745 182.235 ;
        RECT 89.915 181.085 90.145 182.225 ;
        RECT 90.355 182.175 90.875 182.715 ;
        RECT 91.045 182.345 91.565 182.885 ;
        RECT 91.735 182.865 95.245 183.635 ;
        RECT 91.735 182.175 93.425 182.695 ;
        RECT 93.595 182.345 95.245 182.865 ;
        RECT 95.690 182.825 95.935 183.430 ;
        RECT 96.155 183.100 96.665 183.635 ;
        RECT 95.415 182.655 96.645 182.825 ;
        RECT 90.355 181.085 91.565 182.175 ;
        RECT 91.735 181.085 95.245 182.175 ;
        RECT 95.415 181.845 95.755 182.655 ;
        RECT 95.925 182.090 96.675 182.280 ;
        RECT 95.415 181.435 95.930 181.845 ;
        RECT 96.165 181.085 96.335 181.845 ;
        RECT 96.505 181.425 96.675 182.090 ;
        RECT 96.845 182.105 97.035 183.465 ;
        RECT 97.205 183.295 97.480 183.465 ;
        RECT 97.205 183.125 97.485 183.295 ;
        RECT 97.205 182.305 97.480 183.125 ;
        RECT 97.670 183.100 98.200 183.465 ;
        RECT 98.625 183.235 98.955 183.635 ;
        RECT 98.025 183.065 98.200 183.100 ;
        RECT 97.685 182.105 97.855 182.905 ;
        RECT 96.845 181.935 97.855 182.105 ;
        RECT 98.025 182.895 98.955 183.065 ;
        RECT 99.125 182.895 99.380 183.465 ;
        RECT 98.025 181.765 98.195 182.895 ;
        RECT 98.785 182.725 98.955 182.895 ;
        RECT 97.070 181.595 98.195 181.765 ;
        RECT 98.365 182.395 98.560 182.725 ;
        RECT 98.785 182.395 99.040 182.725 ;
        RECT 98.365 181.425 98.535 182.395 ;
        RECT 99.210 182.225 99.380 182.895 ;
        RECT 99.555 182.865 102.145 183.635 ;
        RECT 96.505 181.255 98.535 181.425 ;
        RECT 98.705 181.085 98.875 182.225 ;
        RECT 99.045 181.255 99.380 182.225 ;
        RECT 99.555 182.175 100.765 182.695 ;
        RECT 100.935 182.345 102.145 182.865 ;
        RECT 102.590 182.825 102.835 183.430 ;
        RECT 103.055 183.100 103.565 183.635 ;
        RECT 102.315 182.655 103.545 182.825 ;
        RECT 99.555 181.085 102.145 182.175 ;
        RECT 102.315 181.845 102.655 182.655 ;
        RECT 102.825 182.090 103.575 182.280 ;
        RECT 102.315 181.435 102.830 181.845 ;
        RECT 103.065 181.085 103.235 181.845 ;
        RECT 103.405 181.425 103.575 182.090 ;
        RECT 103.745 182.105 103.935 183.465 ;
        RECT 104.105 182.955 104.380 183.465 ;
        RECT 104.570 183.100 105.100 183.465 ;
        RECT 105.525 183.235 105.855 183.635 ;
        RECT 104.925 183.065 105.100 183.100 ;
        RECT 104.105 182.785 104.385 182.955 ;
        RECT 104.105 182.305 104.380 182.785 ;
        RECT 104.585 182.105 104.755 182.905 ;
        RECT 103.745 181.935 104.755 182.105 ;
        RECT 104.925 182.895 105.855 183.065 ;
        RECT 106.025 182.895 106.280 183.465 ;
        RECT 104.925 181.765 105.095 182.895 ;
        RECT 105.685 182.725 105.855 182.895 ;
        RECT 103.970 181.595 105.095 181.765 ;
        RECT 105.265 182.395 105.460 182.725 ;
        RECT 105.685 182.395 105.940 182.725 ;
        RECT 105.265 181.425 105.435 182.395 ;
        RECT 106.110 182.225 106.280 182.895 ;
        RECT 103.405 181.255 105.435 181.425 ;
        RECT 105.605 181.085 105.775 182.225 ;
        RECT 105.945 181.255 106.280 182.225 ;
        RECT 106.455 182.835 106.795 183.465 ;
        RECT 106.965 182.835 107.215 183.635 ;
        RECT 107.405 182.985 107.735 183.465 ;
        RECT 107.905 183.175 108.130 183.635 ;
        RECT 108.300 182.985 108.630 183.465 ;
        RECT 106.455 182.275 106.630 182.835 ;
        RECT 107.405 182.815 108.630 182.985 ;
        RECT 109.260 182.855 109.760 183.465 ;
        RECT 106.800 182.475 107.495 182.645 ;
        RECT 106.455 182.225 106.685 182.275 ;
        RECT 107.325 182.225 107.495 182.475 ;
        RECT 107.670 182.445 108.090 182.645 ;
        RECT 108.260 182.445 108.590 182.645 ;
        RECT 108.760 182.445 109.090 182.645 ;
        RECT 109.260 182.225 109.430 182.855 ;
        RECT 110.410 182.825 110.655 183.430 ;
        RECT 110.875 183.100 111.385 183.635 ;
        RECT 110.135 182.655 111.365 182.825 ;
        RECT 109.615 182.395 109.965 182.645 ;
        RECT 106.455 181.255 106.795 182.225 ;
        RECT 106.965 181.085 107.135 182.225 ;
        RECT 107.325 182.055 109.760 182.225 ;
        RECT 107.405 181.085 107.655 181.885 ;
        RECT 108.300 181.255 108.630 182.055 ;
        RECT 108.930 181.085 109.260 181.885 ;
        RECT 109.430 181.255 109.760 182.055 ;
        RECT 110.135 181.845 110.475 182.655 ;
        RECT 110.645 182.090 111.395 182.280 ;
        RECT 110.135 181.435 110.650 181.845 ;
        RECT 110.885 181.085 111.055 181.845 ;
        RECT 111.225 181.425 111.395 182.090 ;
        RECT 111.565 182.105 111.755 183.465 ;
        RECT 111.925 182.615 112.200 183.465 ;
        RECT 112.390 183.100 112.920 183.465 ;
        RECT 113.345 183.235 113.675 183.635 ;
        RECT 112.745 183.065 112.920 183.100 ;
        RECT 111.925 182.445 112.205 182.615 ;
        RECT 111.925 182.305 112.200 182.445 ;
        RECT 112.405 182.105 112.575 182.905 ;
        RECT 111.565 181.935 112.575 182.105 ;
        RECT 112.745 182.895 113.675 183.065 ;
        RECT 113.845 182.895 114.100 183.465 ;
        RECT 114.275 182.910 114.565 183.635 ;
        RECT 115.660 182.925 115.915 183.455 ;
        RECT 116.085 183.175 116.390 183.635 ;
        RECT 116.635 183.255 117.705 183.425 ;
        RECT 112.745 181.765 112.915 182.895 ;
        RECT 113.505 182.725 113.675 182.895 ;
        RECT 111.790 181.595 112.915 181.765 ;
        RECT 113.085 182.395 113.280 182.725 ;
        RECT 113.505 182.395 113.760 182.725 ;
        RECT 113.085 181.425 113.255 182.395 ;
        RECT 113.930 182.225 114.100 182.895 ;
        RECT 115.660 182.275 115.870 182.925 ;
        RECT 116.635 182.900 116.955 183.255 ;
        RECT 116.630 182.725 116.955 182.900 ;
        RECT 116.040 182.425 116.955 182.725 ;
        RECT 117.125 182.685 117.365 183.085 ;
        RECT 117.535 183.025 117.705 183.255 ;
        RECT 117.875 183.195 118.065 183.635 ;
        RECT 118.235 183.185 119.185 183.465 ;
        RECT 119.405 183.275 119.755 183.445 ;
        RECT 117.535 182.855 118.065 183.025 ;
        RECT 116.040 182.395 116.780 182.425 ;
        RECT 111.225 181.255 113.255 181.425 ;
        RECT 113.425 181.085 113.595 182.225 ;
        RECT 113.765 181.255 114.100 182.225 ;
        RECT 114.275 181.085 114.565 182.250 ;
        RECT 115.660 181.395 115.915 182.275 ;
        RECT 116.085 181.085 116.390 182.225 ;
        RECT 116.610 181.805 116.780 182.395 ;
        RECT 117.125 182.315 117.665 182.685 ;
        RECT 117.845 182.575 118.065 182.855 ;
        RECT 118.235 182.405 118.405 183.185 ;
        RECT 118.000 182.235 118.405 182.405 ;
        RECT 118.575 182.395 118.925 183.015 ;
        RECT 118.000 182.145 118.170 182.235 ;
        RECT 119.095 182.225 119.305 183.015 ;
        RECT 116.950 181.975 118.170 182.145 ;
        RECT 118.630 182.065 119.305 182.225 ;
        RECT 116.610 181.635 117.410 181.805 ;
        RECT 116.730 181.085 117.060 181.465 ;
        RECT 117.240 181.345 117.410 181.635 ;
        RECT 118.000 181.595 118.170 181.975 ;
        RECT 118.340 182.055 119.305 182.065 ;
        RECT 119.495 182.885 119.755 183.275 ;
        RECT 119.965 183.175 120.295 183.635 ;
        RECT 121.170 183.245 122.025 183.415 ;
        RECT 122.230 183.245 122.725 183.415 ;
        RECT 122.895 183.275 123.225 183.635 ;
        RECT 119.495 182.195 119.665 182.885 ;
        RECT 119.835 182.535 120.005 182.715 ;
        RECT 120.175 182.705 120.965 182.955 ;
        RECT 121.170 182.535 121.340 183.245 ;
        RECT 121.510 182.735 121.865 182.955 ;
        RECT 119.835 182.365 121.525 182.535 ;
        RECT 118.340 181.765 118.800 182.055 ;
        RECT 119.495 182.025 120.995 182.195 ;
        RECT 119.495 181.885 119.665 182.025 ;
        RECT 119.105 181.715 119.665 181.885 ;
        RECT 117.580 181.085 117.830 181.545 ;
        RECT 118.000 181.255 118.870 181.595 ;
        RECT 119.105 181.255 119.275 181.715 ;
        RECT 120.110 181.685 121.185 181.855 ;
        RECT 119.445 181.085 119.815 181.545 ;
        RECT 120.110 181.345 120.280 181.685 ;
        RECT 120.450 181.085 120.780 181.515 ;
        RECT 121.015 181.345 121.185 181.685 ;
        RECT 121.355 181.585 121.525 182.365 ;
        RECT 121.695 182.145 121.865 182.735 ;
        RECT 122.035 182.335 122.385 182.955 ;
        RECT 121.695 181.755 122.160 182.145 ;
        RECT 122.555 181.885 122.725 183.245 ;
        RECT 122.895 182.055 123.355 183.105 ;
        RECT 122.330 181.715 122.725 181.885 ;
        RECT 122.330 181.585 122.500 181.715 ;
        RECT 121.355 181.255 122.035 181.585 ;
        RECT 122.250 181.255 122.500 181.585 ;
        RECT 122.670 181.085 122.920 181.545 ;
        RECT 123.090 181.270 123.415 182.055 ;
        RECT 123.585 181.255 123.755 183.375 ;
        RECT 123.925 183.255 124.255 183.635 ;
        RECT 124.425 183.085 124.680 183.375 ;
        RECT 123.930 182.915 124.680 183.085 ;
        RECT 123.930 181.925 124.160 182.915 ;
        RECT 124.855 182.885 126.065 183.635 ;
        RECT 126.235 182.885 127.445 183.635 ;
        RECT 124.330 182.095 124.680 182.745 ;
        RECT 124.855 182.175 125.375 182.715 ;
        RECT 125.545 182.345 126.065 182.885 ;
        RECT 126.235 182.175 126.755 182.715 ;
        RECT 126.925 182.345 127.445 182.885 ;
        RECT 123.930 181.755 124.680 181.925 ;
        RECT 123.925 181.085 124.255 181.585 ;
        RECT 124.425 181.255 124.680 181.755 ;
        RECT 124.855 181.085 126.065 182.175 ;
        RECT 126.235 181.085 127.445 182.175 ;
        RECT 14.370 180.915 127.530 181.085 ;
        RECT 14.455 179.825 15.665 180.915 ;
        RECT 14.455 179.115 14.975 179.655 ;
        RECT 15.145 179.285 15.665 179.825 ;
        RECT 15.835 179.825 18.425 180.915 ;
        RECT 18.600 180.480 23.945 180.915 ;
        RECT 15.835 179.305 17.045 179.825 ;
        RECT 17.215 179.135 18.425 179.655 ;
        RECT 20.190 179.230 20.540 180.480 ;
        RECT 24.115 179.750 24.405 180.915 ;
        RECT 24.580 180.245 24.835 180.745 ;
        RECT 25.005 180.415 25.335 180.915 ;
        RECT 24.580 180.075 25.330 180.245 ;
        RECT 14.455 178.365 15.665 179.115 ;
        RECT 15.835 178.365 18.425 179.135 ;
        RECT 22.020 178.910 22.360 179.740 ;
        RECT 24.580 179.255 24.930 179.905 ;
        RECT 18.600 178.365 23.945 178.910 ;
        RECT 24.115 178.365 24.405 179.090 ;
        RECT 25.100 179.085 25.330 180.075 ;
        RECT 24.580 178.915 25.330 179.085 ;
        RECT 24.580 178.625 24.835 178.915 ;
        RECT 25.005 178.365 25.335 178.745 ;
        RECT 25.505 178.625 25.675 180.745 ;
        RECT 25.845 179.945 26.170 180.730 ;
        RECT 26.340 180.455 26.590 180.915 ;
        RECT 26.760 180.415 27.010 180.745 ;
        RECT 27.225 180.415 27.905 180.745 ;
        RECT 26.760 180.285 26.930 180.415 ;
        RECT 26.535 180.115 26.930 180.285 ;
        RECT 25.905 178.895 26.365 179.945 ;
        RECT 26.535 178.755 26.705 180.115 ;
        RECT 27.100 179.855 27.565 180.245 ;
        RECT 26.875 179.045 27.225 179.665 ;
        RECT 27.395 179.265 27.565 179.855 ;
        RECT 27.735 179.635 27.905 180.415 ;
        RECT 28.075 180.315 28.245 180.655 ;
        RECT 28.480 180.485 28.810 180.915 ;
        RECT 28.980 180.315 29.150 180.655 ;
        RECT 29.445 180.455 29.815 180.915 ;
        RECT 28.075 180.145 29.150 180.315 ;
        RECT 29.985 180.285 30.155 180.745 ;
        RECT 30.390 180.405 31.260 180.745 ;
        RECT 31.430 180.455 31.680 180.915 ;
        RECT 29.595 180.115 30.155 180.285 ;
        RECT 29.595 179.975 29.765 180.115 ;
        RECT 28.265 179.805 29.765 179.975 ;
        RECT 30.460 179.945 30.920 180.235 ;
        RECT 27.735 179.465 29.425 179.635 ;
        RECT 27.395 179.045 27.750 179.265 ;
        RECT 27.920 178.755 28.090 179.465 ;
        RECT 28.295 179.045 29.085 179.295 ;
        RECT 29.255 179.285 29.425 179.465 ;
        RECT 29.595 179.115 29.765 179.805 ;
        RECT 26.035 178.365 26.365 178.725 ;
        RECT 26.535 178.585 27.030 178.755 ;
        RECT 27.235 178.585 28.090 178.755 ;
        RECT 28.965 178.365 29.295 178.825 ;
        RECT 29.505 178.725 29.765 179.115 ;
        RECT 29.955 179.935 30.920 179.945 ;
        RECT 31.090 180.025 31.260 180.405 ;
        RECT 31.850 180.365 32.020 180.655 ;
        RECT 32.200 180.535 32.530 180.915 ;
        RECT 31.850 180.195 32.650 180.365 ;
        RECT 29.955 179.775 30.630 179.935 ;
        RECT 31.090 179.855 32.310 180.025 ;
        RECT 29.955 178.985 30.165 179.775 ;
        RECT 31.090 179.765 31.260 179.855 ;
        RECT 30.335 178.985 30.685 179.605 ;
        RECT 30.855 179.595 31.260 179.765 ;
        RECT 30.855 178.815 31.025 179.595 ;
        RECT 31.195 179.145 31.415 179.425 ;
        RECT 31.595 179.315 32.135 179.685 ;
        RECT 32.480 179.605 32.650 180.195 ;
        RECT 32.870 179.775 33.175 180.915 ;
        RECT 33.345 179.725 33.600 180.605 ;
        RECT 32.480 179.575 33.220 179.605 ;
        RECT 31.195 178.975 31.725 179.145 ;
        RECT 29.505 178.555 29.855 178.725 ;
        RECT 30.075 178.535 31.025 178.815 ;
        RECT 31.195 178.365 31.385 178.805 ;
        RECT 31.555 178.745 31.725 178.975 ;
        RECT 31.895 178.915 32.135 179.315 ;
        RECT 32.305 179.275 33.220 179.575 ;
        RECT 32.305 179.100 32.630 179.275 ;
        RECT 32.305 178.745 32.625 179.100 ;
        RECT 33.390 179.075 33.600 179.725 ;
        RECT 31.555 178.575 32.625 178.745 ;
        RECT 32.870 178.365 33.175 178.825 ;
        RECT 33.345 178.545 33.600 179.075 ;
        RECT 33.775 179.775 34.160 180.745 ;
        RECT 34.330 180.455 34.655 180.915 ;
        RECT 35.175 180.285 35.455 180.745 ;
        RECT 34.330 180.065 35.455 180.285 ;
        RECT 33.775 179.105 34.055 179.775 ;
        RECT 34.330 179.605 34.780 180.065 ;
        RECT 35.645 179.895 36.045 180.745 ;
        RECT 36.445 180.455 36.715 180.915 ;
        RECT 36.885 180.285 37.170 180.745 ;
        RECT 34.225 179.275 34.780 179.605 ;
        RECT 34.950 179.335 36.045 179.895 ;
        RECT 34.330 179.165 34.780 179.275 ;
        RECT 33.775 178.535 34.160 179.105 ;
        RECT 34.330 178.995 35.455 179.165 ;
        RECT 34.330 178.365 34.655 178.825 ;
        RECT 35.175 178.535 35.455 178.995 ;
        RECT 35.645 178.535 36.045 179.335 ;
        RECT 36.215 180.065 37.170 180.285 ;
        RECT 36.215 179.165 36.425 180.065 ;
        RECT 36.595 179.335 37.285 179.895 ;
        RECT 37.915 179.775 38.255 180.745 ;
        RECT 38.425 179.775 38.595 180.915 ;
        RECT 38.865 180.115 39.115 180.915 ;
        RECT 39.760 179.945 40.090 180.745 ;
        RECT 40.390 180.115 40.720 180.915 ;
        RECT 40.890 179.945 41.220 180.745 ;
        RECT 38.785 179.775 41.220 179.945 ;
        RECT 42.055 179.775 42.395 180.745 ;
        RECT 42.565 179.775 42.735 180.915 ;
        RECT 43.005 180.115 43.255 180.915 ;
        RECT 43.900 179.945 44.230 180.745 ;
        RECT 44.530 180.115 44.860 180.915 ;
        RECT 45.030 179.945 45.360 180.745 ;
        RECT 42.925 179.775 45.360 179.945 ;
        RECT 45.735 180.155 46.250 180.565 ;
        RECT 46.485 180.155 46.655 180.915 ;
        RECT 46.825 180.575 48.855 180.745 ;
        RECT 37.915 179.215 38.090 179.775 ;
        RECT 38.785 179.525 38.955 179.775 ;
        RECT 38.260 179.355 38.955 179.525 ;
        RECT 39.130 179.355 39.550 179.555 ;
        RECT 39.720 179.355 40.050 179.555 ;
        RECT 40.220 179.355 40.550 179.555 ;
        RECT 37.915 179.165 38.145 179.215 ;
        RECT 36.215 178.995 37.170 179.165 ;
        RECT 36.445 178.365 36.715 178.825 ;
        RECT 36.885 178.535 37.170 178.995 ;
        RECT 37.915 178.535 38.255 179.165 ;
        RECT 38.425 178.365 38.675 179.165 ;
        RECT 38.865 179.015 40.090 179.185 ;
        RECT 38.865 178.535 39.195 179.015 ;
        RECT 39.365 178.365 39.590 178.825 ;
        RECT 39.760 178.535 40.090 179.015 ;
        RECT 40.720 179.145 40.890 179.775 ;
        RECT 41.075 179.355 41.425 179.605 ;
        RECT 42.055 179.165 42.230 179.775 ;
        RECT 42.925 179.525 43.095 179.775 ;
        RECT 42.400 179.355 43.095 179.525 ;
        RECT 43.270 179.355 43.690 179.555 ;
        RECT 43.860 179.355 44.190 179.555 ;
        RECT 44.360 179.355 44.690 179.555 ;
        RECT 40.720 178.535 41.220 179.145 ;
        RECT 42.055 178.535 42.395 179.165 ;
        RECT 42.565 178.365 42.815 179.165 ;
        RECT 43.005 179.015 44.230 179.185 ;
        RECT 43.005 178.535 43.335 179.015 ;
        RECT 43.505 178.365 43.730 178.825 ;
        RECT 43.900 178.535 44.230 179.015 ;
        RECT 44.860 179.145 45.030 179.775 ;
        RECT 45.215 179.355 45.565 179.605 ;
        RECT 45.735 179.345 46.075 180.155 ;
        RECT 46.825 179.910 46.995 180.575 ;
        RECT 47.390 180.235 48.515 180.405 ;
        RECT 46.245 179.720 46.995 179.910 ;
        RECT 47.165 179.895 48.175 180.065 ;
        RECT 45.735 179.175 46.965 179.345 ;
        RECT 44.860 178.535 45.360 179.145 ;
        RECT 46.010 178.570 46.255 179.175 ;
        RECT 46.475 178.365 46.985 178.900 ;
        RECT 47.165 178.535 47.355 179.895 ;
        RECT 47.525 178.875 47.800 179.695 ;
        RECT 48.005 179.095 48.175 179.895 ;
        RECT 48.345 179.105 48.515 180.235 ;
        RECT 48.685 179.605 48.855 180.575 ;
        RECT 49.025 179.775 49.195 180.915 ;
        RECT 49.365 179.775 49.700 180.745 ;
        RECT 48.685 179.275 48.880 179.605 ;
        RECT 49.105 179.275 49.360 179.605 ;
        RECT 49.105 179.105 49.275 179.275 ;
        RECT 49.530 179.105 49.700 179.775 ;
        RECT 49.875 179.750 50.165 180.915 ;
        RECT 50.450 180.285 50.735 180.745 ;
        RECT 50.905 180.455 51.175 180.915 ;
        RECT 50.450 180.065 51.405 180.285 ;
        RECT 50.335 179.335 51.025 179.895 ;
        RECT 51.195 179.165 51.405 180.065 ;
        RECT 48.345 178.935 49.275 179.105 ;
        RECT 48.345 178.900 48.520 178.935 ;
        RECT 47.525 178.705 47.805 178.875 ;
        RECT 47.525 178.535 47.800 178.705 ;
        RECT 47.990 178.535 48.520 178.900 ;
        RECT 48.945 178.365 49.275 178.765 ;
        RECT 49.445 178.535 49.700 179.105 ;
        RECT 49.875 178.365 50.165 179.090 ;
        RECT 50.450 178.995 51.405 179.165 ;
        RECT 51.575 179.895 51.975 180.745 ;
        RECT 52.165 180.285 52.445 180.745 ;
        RECT 52.965 180.455 53.290 180.915 ;
        RECT 52.165 180.065 53.290 180.285 ;
        RECT 51.575 179.335 52.670 179.895 ;
        RECT 52.840 179.605 53.290 180.065 ;
        RECT 53.460 179.775 53.845 180.745 ;
        RECT 50.450 178.535 50.735 178.995 ;
        RECT 50.905 178.365 51.175 178.825 ;
        RECT 51.575 178.535 51.975 179.335 ;
        RECT 52.840 179.275 53.395 179.605 ;
        RECT 52.840 179.165 53.290 179.275 ;
        RECT 52.165 178.995 53.290 179.165 ;
        RECT 53.565 179.105 53.845 179.775 ;
        RECT 54.015 179.825 55.685 180.915 ;
        RECT 54.015 179.305 54.765 179.825 ;
        RECT 55.860 179.775 56.195 180.745 ;
        RECT 56.365 179.775 56.535 180.915 ;
        RECT 56.705 180.575 58.735 180.745 ;
        RECT 54.935 179.135 55.685 179.655 ;
        RECT 52.165 178.535 52.445 178.995 ;
        RECT 52.965 178.365 53.290 178.825 ;
        RECT 53.460 178.535 53.845 179.105 ;
        RECT 54.015 178.365 55.685 179.135 ;
        RECT 55.860 179.105 56.030 179.775 ;
        RECT 56.705 179.605 56.875 180.575 ;
        RECT 56.200 179.275 56.455 179.605 ;
        RECT 56.680 179.275 56.875 179.605 ;
        RECT 57.045 180.235 58.170 180.405 ;
        RECT 56.285 179.105 56.455 179.275 ;
        RECT 57.045 179.105 57.215 180.235 ;
        RECT 55.860 178.535 56.115 179.105 ;
        RECT 56.285 178.935 57.215 179.105 ;
        RECT 57.385 179.895 58.395 180.065 ;
        RECT 57.385 179.095 57.555 179.895 ;
        RECT 57.040 178.900 57.215 178.935 ;
        RECT 56.285 178.365 56.615 178.765 ;
        RECT 57.040 178.535 57.570 178.900 ;
        RECT 57.760 178.875 58.035 179.695 ;
        RECT 57.755 178.705 58.035 178.875 ;
        RECT 57.760 178.535 58.035 178.705 ;
        RECT 58.205 178.535 58.395 179.895 ;
        RECT 58.565 179.910 58.735 180.575 ;
        RECT 58.905 180.155 59.075 180.915 ;
        RECT 59.310 180.155 59.825 180.565 ;
        RECT 58.565 179.720 59.315 179.910 ;
        RECT 59.485 179.345 59.825 180.155 ;
        RECT 60.050 180.045 60.335 180.915 ;
        RECT 60.505 180.285 60.765 180.745 ;
        RECT 60.940 180.455 61.195 180.915 ;
        RECT 61.365 180.285 61.625 180.745 ;
        RECT 60.505 180.115 61.625 180.285 ;
        RECT 61.795 180.115 62.105 180.915 ;
        RECT 60.505 179.865 60.765 180.115 ;
        RECT 62.275 179.945 62.585 180.745 ;
        RECT 58.595 179.175 59.825 179.345 ;
        RECT 60.010 179.695 60.765 179.865 ;
        RECT 61.555 179.775 62.585 179.945 ;
        RECT 60.010 179.185 60.415 179.695 ;
        RECT 61.555 179.525 61.725 179.775 ;
        RECT 60.585 179.355 61.725 179.525 ;
        RECT 58.575 178.365 59.085 178.900 ;
        RECT 59.305 178.570 59.550 179.175 ;
        RECT 60.010 179.015 61.660 179.185 ;
        RECT 61.895 179.035 62.245 179.605 ;
        RECT 60.055 178.365 60.335 178.845 ;
        RECT 60.505 178.625 60.765 179.015 ;
        RECT 60.940 178.365 61.195 178.845 ;
        RECT 61.365 178.625 61.660 179.015 ;
        RECT 62.415 178.865 62.585 179.775 ;
        RECT 62.755 179.825 65.345 180.915 ;
        RECT 62.755 179.305 63.965 179.825 ;
        RECT 65.555 179.775 65.785 180.915 ;
        RECT 65.955 179.765 66.285 180.745 ;
        RECT 66.455 179.775 66.665 180.915 ;
        RECT 66.900 179.765 67.160 180.915 ;
        RECT 67.335 179.840 67.590 180.745 ;
        RECT 67.760 180.155 68.090 180.915 ;
        RECT 68.305 179.985 68.475 180.745 ;
        RECT 64.135 179.135 65.345 179.655 ;
        RECT 65.535 179.355 65.865 179.605 ;
        RECT 61.840 178.365 62.115 178.845 ;
        RECT 62.285 178.535 62.585 178.865 ;
        RECT 62.755 178.365 65.345 179.135 ;
        RECT 65.555 178.365 65.785 179.185 ;
        RECT 66.035 179.165 66.285 179.765 ;
        RECT 65.955 178.535 66.285 179.165 ;
        RECT 66.455 178.365 66.665 179.185 ;
        RECT 66.900 178.365 67.160 179.205 ;
        RECT 67.335 179.110 67.505 179.840 ;
        RECT 67.760 179.815 68.475 179.985 ;
        RECT 68.735 179.945 69.045 180.745 ;
        RECT 69.215 180.115 69.525 180.915 ;
        RECT 69.695 180.285 69.955 180.745 ;
        RECT 70.125 180.455 70.380 180.915 ;
        RECT 70.555 180.285 70.815 180.745 ;
        RECT 69.695 180.115 70.815 180.285 ;
        RECT 67.760 179.605 67.930 179.815 ;
        RECT 68.735 179.775 69.765 179.945 ;
        RECT 67.675 179.275 67.930 179.605 ;
        RECT 67.335 178.535 67.590 179.110 ;
        RECT 67.760 179.085 67.930 179.275 ;
        RECT 68.210 179.265 68.565 179.635 ;
        RECT 67.760 178.915 68.475 179.085 ;
        RECT 67.760 178.365 68.090 178.745 ;
        RECT 68.305 178.535 68.475 178.915 ;
        RECT 68.735 178.865 68.905 179.775 ;
        RECT 69.075 179.035 69.425 179.605 ;
        RECT 69.595 179.525 69.765 179.775 ;
        RECT 70.555 179.865 70.815 180.115 ;
        RECT 70.985 180.045 71.270 180.915 ;
        RECT 70.555 179.695 71.310 179.865 ;
        RECT 69.595 179.355 70.735 179.525 ;
        RECT 70.905 179.185 71.310 179.695 ;
        RECT 69.660 179.015 71.310 179.185 ;
        RECT 71.495 179.105 71.755 180.730 ;
        RECT 73.505 180.465 73.835 180.915 ;
        RECT 71.935 180.075 74.545 180.285 ;
        RECT 71.935 179.275 72.155 180.075 ;
        RECT 72.395 179.275 72.695 179.895 ;
        RECT 72.865 179.275 73.195 179.895 ;
        RECT 73.365 179.275 73.685 179.895 ;
        RECT 73.855 179.275 74.205 179.895 ;
        RECT 74.375 179.105 74.545 180.075 ;
        RECT 75.635 179.750 75.925 180.915 ;
        RECT 76.210 180.285 76.495 180.745 ;
        RECT 76.665 180.455 76.935 180.915 ;
        RECT 76.210 180.065 77.165 180.285 ;
        RECT 76.095 179.335 76.785 179.895 ;
        RECT 76.955 179.165 77.165 180.065 ;
        RECT 68.735 178.535 69.035 178.865 ;
        RECT 69.205 178.365 69.480 178.845 ;
        RECT 69.660 178.625 69.955 179.015 ;
        RECT 70.125 178.365 70.380 178.845 ;
        RECT 70.555 178.625 70.815 179.015 ;
        RECT 71.495 178.935 73.335 179.105 ;
        RECT 70.985 178.365 71.265 178.845 ;
        RECT 71.765 178.365 72.095 178.760 ;
        RECT 72.265 178.580 72.465 178.935 ;
        RECT 72.635 178.365 72.965 178.765 ;
        RECT 73.135 178.590 73.335 178.935 ;
        RECT 73.505 178.365 73.835 179.105 ;
        RECT 74.070 178.935 74.545 179.105 ;
        RECT 74.070 178.685 74.240 178.935 ;
        RECT 75.635 178.365 75.925 179.090 ;
        RECT 76.210 178.995 77.165 179.165 ;
        RECT 77.335 179.895 77.735 180.745 ;
        RECT 77.925 180.285 78.205 180.745 ;
        RECT 78.725 180.455 79.050 180.915 ;
        RECT 77.925 180.065 79.050 180.285 ;
        RECT 77.335 179.335 78.430 179.895 ;
        RECT 78.600 179.605 79.050 180.065 ;
        RECT 79.220 179.775 79.605 180.745 ;
        RECT 79.980 179.945 80.310 180.745 ;
        RECT 80.480 180.115 80.810 180.915 ;
        RECT 81.110 179.945 81.440 180.745 ;
        RECT 82.085 180.115 82.335 180.915 ;
        RECT 79.980 179.775 82.415 179.945 ;
        RECT 82.605 179.775 82.775 180.915 ;
        RECT 82.945 179.775 83.285 180.745 ;
        RECT 76.210 178.535 76.495 178.995 ;
        RECT 76.665 178.365 76.935 178.825 ;
        RECT 77.335 178.535 77.735 179.335 ;
        RECT 78.600 179.275 79.155 179.605 ;
        RECT 78.600 179.165 79.050 179.275 ;
        RECT 77.925 178.995 79.050 179.165 ;
        RECT 79.325 179.105 79.605 179.775 ;
        RECT 79.775 179.355 80.125 179.605 ;
        RECT 80.310 179.145 80.480 179.775 ;
        RECT 80.650 179.355 80.980 179.555 ;
        RECT 81.150 179.355 81.480 179.555 ;
        RECT 81.650 179.355 82.070 179.555 ;
        RECT 82.245 179.525 82.415 179.775 ;
        RECT 82.245 179.355 82.940 179.525 ;
        RECT 77.925 178.535 78.205 178.995 ;
        RECT 78.725 178.365 79.050 178.825 ;
        RECT 79.220 178.535 79.605 179.105 ;
        RECT 79.980 178.535 80.480 179.145 ;
        RECT 81.110 179.015 82.335 179.185 ;
        RECT 83.110 179.165 83.285 179.775 ;
        RECT 83.455 179.825 85.125 180.915 ;
        RECT 85.295 180.155 85.810 180.565 ;
        RECT 86.045 180.155 86.215 180.915 ;
        RECT 86.385 180.575 88.415 180.745 ;
        RECT 83.455 179.305 84.205 179.825 ;
        RECT 81.110 178.535 81.440 179.015 ;
        RECT 81.610 178.365 81.835 178.825 ;
        RECT 82.005 178.535 82.335 179.015 ;
        RECT 82.525 178.365 82.775 179.165 ;
        RECT 82.945 178.535 83.285 179.165 ;
        RECT 84.375 179.135 85.125 179.655 ;
        RECT 85.295 179.345 85.635 180.155 ;
        RECT 86.385 179.910 86.555 180.575 ;
        RECT 86.950 180.235 88.075 180.405 ;
        RECT 85.805 179.720 86.555 179.910 ;
        RECT 86.725 179.895 87.735 180.065 ;
        RECT 85.295 179.175 86.525 179.345 ;
        RECT 83.455 178.365 85.125 179.135 ;
        RECT 85.570 178.570 85.815 179.175 ;
        RECT 86.035 178.365 86.545 178.900 ;
        RECT 86.725 178.535 86.915 179.895 ;
        RECT 87.085 178.875 87.360 179.695 ;
        RECT 87.565 179.095 87.735 179.895 ;
        RECT 87.905 179.105 88.075 180.235 ;
        RECT 88.245 179.605 88.415 180.575 ;
        RECT 88.585 179.775 88.755 180.915 ;
        RECT 88.925 179.775 89.260 180.745 ;
        RECT 88.245 179.275 88.440 179.605 ;
        RECT 88.665 179.275 88.920 179.605 ;
        RECT 88.665 179.105 88.835 179.275 ;
        RECT 89.090 179.105 89.260 179.775 ;
        RECT 87.905 178.935 88.835 179.105 ;
        RECT 87.905 178.900 88.080 178.935 ;
        RECT 87.085 178.705 87.365 178.875 ;
        RECT 87.085 178.535 87.360 178.705 ;
        RECT 87.550 178.535 88.080 178.900 ;
        RECT 88.505 178.365 88.835 178.765 ;
        RECT 89.005 178.535 89.260 179.105 ;
        RECT 89.435 179.840 89.705 180.745 ;
        RECT 89.875 180.155 90.205 180.915 ;
        RECT 90.385 179.985 90.555 180.745 ;
        RECT 89.435 179.040 89.605 179.840 ;
        RECT 89.890 179.815 90.555 179.985 ;
        RECT 89.890 179.670 90.060 179.815 ;
        RECT 90.855 179.775 91.085 180.915 ;
        RECT 91.255 179.765 91.585 180.745 ;
        RECT 91.755 179.775 91.965 180.915 ;
        RECT 89.775 179.340 90.060 179.670 ;
        RECT 89.890 179.085 90.060 179.340 ;
        RECT 90.295 179.265 90.625 179.635 ;
        RECT 90.835 179.355 91.165 179.605 ;
        RECT 89.435 178.535 89.695 179.040 ;
        RECT 89.890 178.915 90.555 179.085 ;
        RECT 89.875 178.365 90.205 178.745 ;
        RECT 90.385 178.535 90.555 178.915 ;
        RECT 90.855 178.365 91.085 179.185 ;
        RECT 91.335 179.165 91.585 179.765 ;
        RECT 92.200 179.725 92.455 180.605 ;
        RECT 92.625 179.775 92.930 180.915 ;
        RECT 93.270 180.535 93.600 180.915 ;
        RECT 93.780 180.365 93.950 180.655 ;
        RECT 94.120 180.455 94.370 180.915 ;
        RECT 93.150 180.195 93.950 180.365 ;
        RECT 94.540 180.405 95.410 180.745 ;
        RECT 91.255 178.535 91.585 179.165 ;
        RECT 91.755 178.365 91.965 179.185 ;
        RECT 92.200 179.075 92.410 179.725 ;
        RECT 93.150 179.605 93.320 180.195 ;
        RECT 94.540 180.025 94.710 180.405 ;
        RECT 95.645 180.285 95.815 180.745 ;
        RECT 95.985 180.455 96.355 180.915 ;
        RECT 96.650 180.315 96.820 180.655 ;
        RECT 96.990 180.485 97.320 180.915 ;
        RECT 97.555 180.315 97.725 180.655 ;
        RECT 93.490 179.855 94.710 180.025 ;
        RECT 94.880 179.945 95.340 180.235 ;
        RECT 95.645 180.115 96.205 180.285 ;
        RECT 96.650 180.145 97.725 180.315 ;
        RECT 97.895 180.415 98.575 180.745 ;
        RECT 98.790 180.415 99.040 180.745 ;
        RECT 99.210 180.455 99.460 180.915 ;
        RECT 96.035 179.975 96.205 180.115 ;
        RECT 94.880 179.935 95.845 179.945 ;
        RECT 94.540 179.765 94.710 179.855 ;
        RECT 95.170 179.775 95.845 179.935 ;
        RECT 92.580 179.575 93.320 179.605 ;
        RECT 92.580 179.275 93.495 179.575 ;
        RECT 93.170 179.100 93.495 179.275 ;
        RECT 92.200 178.545 92.455 179.075 ;
        RECT 92.625 178.365 92.930 178.825 ;
        RECT 93.175 178.745 93.495 179.100 ;
        RECT 93.665 179.315 94.205 179.685 ;
        RECT 94.540 179.595 94.945 179.765 ;
        RECT 93.665 178.915 93.905 179.315 ;
        RECT 94.385 179.145 94.605 179.425 ;
        RECT 94.075 178.975 94.605 179.145 ;
        RECT 94.075 178.745 94.245 178.975 ;
        RECT 94.775 178.815 94.945 179.595 ;
        RECT 95.115 178.985 95.465 179.605 ;
        RECT 95.635 178.985 95.845 179.775 ;
        RECT 96.035 179.805 97.535 179.975 ;
        RECT 96.035 179.115 96.205 179.805 ;
        RECT 97.895 179.635 98.065 180.415 ;
        RECT 98.870 180.285 99.040 180.415 ;
        RECT 96.375 179.465 98.065 179.635 ;
        RECT 98.235 179.855 98.700 180.245 ;
        RECT 98.870 180.115 99.265 180.285 ;
        RECT 96.375 179.285 96.545 179.465 ;
        RECT 93.175 178.575 94.245 178.745 ;
        RECT 94.415 178.365 94.605 178.805 ;
        RECT 94.775 178.535 95.725 178.815 ;
        RECT 96.035 178.725 96.295 179.115 ;
        RECT 96.715 179.045 97.505 179.295 ;
        RECT 95.945 178.555 96.295 178.725 ;
        RECT 96.505 178.365 96.835 178.825 ;
        RECT 97.710 178.755 97.880 179.465 ;
        RECT 98.235 179.265 98.405 179.855 ;
        RECT 98.050 179.045 98.405 179.265 ;
        RECT 98.575 179.045 98.925 179.665 ;
        RECT 99.095 178.755 99.265 180.115 ;
        RECT 99.630 179.945 99.955 180.730 ;
        RECT 99.435 178.895 99.895 179.945 ;
        RECT 97.710 178.585 98.565 178.755 ;
        RECT 98.770 178.585 99.265 178.755 ;
        RECT 99.435 178.365 99.765 178.725 ;
        RECT 100.125 178.625 100.295 180.745 ;
        RECT 100.465 180.415 100.795 180.915 ;
        RECT 100.965 180.245 101.220 180.745 ;
        RECT 100.470 180.075 101.220 180.245 ;
        RECT 100.470 179.085 100.700 180.075 ;
        RECT 100.870 179.255 101.220 179.905 ;
        RECT 101.395 179.750 101.685 180.915 ;
        RECT 101.855 179.775 102.240 180.745 ;
        RECT 102.410 180.455 102.735 180.915 ;
        RECT 103.255 180.285 103.535 180.745 ;
        RECT 102.410 180.065 103.535 180.285 ;
        RECT 101.855 179.105 102.135 179.775 ;
        RECT 102.410 179.605 102.860 180.065 ;
        RECT 103.725 179.895 104.125 180.745 ;
        RECT 104.525 180.455 104.795 180.915 ;
        RECT 104.965 180.285 105.250 180.745 ;
        RECT 102.305 179.275 102.860 179.605 ;
        RECT 103.030 179.335 104.125 179.895 ;
        RECT 102.410 179.165 102.860 179.275 ;
        RECT 100.470 178.915 101.220 179.085 ;
        RECT 100.465 178.365 100.795 178.745 ;
        RECT 100.965 178.625 101.220 178.915 ;
        RECT 101.395 178.365 101.685 179.090 ;
        RECT 101.855 178.535 102.240 179.105 ;
        RECT 102.410 178.995 103.535 179.165 ;
        RECT 102.410 178.365 102.735 178.825 ;
        RECT 103.255 178.535 103.535 178.995 ;
        RECT 103.725 178.535 104.125 179.335 ;
        RECT 104.295 180.065 105.250 180.285 ;
        RECT 104.295 179.165 104.505 180.065 ;
        RECT 104.675 179.335 105.365 179.895 ;
        RECT 105.535 179.775 105.920 180.745 ;
        RECT 106.090 180.455 106.415 180.915 ;
        RECT 106.935 180.285 107.215 180.745 ;
        RECT 106.090 180.065 107.215 180.285 ;
        RECT 104.295 178.995 105.250 179.165 ;
        RECT 104.525 178.365 104.795 178.825 ;
        RECT 104.965 178.535 105.250 178.995 ;
        RECT 105.535 179.105 105.815 179.775 ;
        RECT 106.090 179.605 106.540 180.065 ;
        RECT 107.405 179.895 107.805 180.745 ;
        RECT 108.205 180.455 108.475 180.915 ;
        RECT 108.645 180.285 108.930 180.745 ;
        RECT 105.985 179.275 106.540 179.605 ;
        RECT 106.710 179.335 107.805 179.895 ;
        RECT 106.090 179.165 106.540 179.275 ;
        RECT 105.535 178.535 105.920 179.105 ;
        RECT 106.090 178.995 107.215 179.165 ;
        RECT 106.090 178.365 106.415 178.825 ;
        RECT 106.935 178.535 107.215 178.995 ;
        RECT 107.405 178.535 107.805 179.335 ;
        RECT 107.975 180.065 108.930 180.285 ;
        RECT 107.975 179.165 108.185 180.065 ;
        RECT 108.355 179.335 109.045 179.895 ;
        RECT 109.715 179.775 109.945 180.915 ;
        RECT 110.115 179.765 110.445 180.745 ;
        RECT 110.615 179.775 110.825 180.915 ;
        RECT 109.695 179.355 110.025 179.605 ;
        RECT 107.975 178.995 108.930 179.165 ;
        RECT 108.205 178.365 108.475 178.825 ;
        RECT 108.645 178.535 108.930 178.995 ;
        RECT 109.715 178.365 109.945 179.185 ;
        RECT 110.195 179.165 110.445 179.765 ;
        RECT 111.060 179.725 111.315 180.605 ;
        RECT 111.485 179.775 111.790 180.915 ;
        RECT 112.130 180.535 112.460 180.915 ;
        RECT 112.640 180.365 112.810 180.655 ;
        RECT 112.980 180.455 113.230 180.915 ;
        RECT 112.010 180.195 112.810 180.365 ;
        RECT 113.400 180.405 114.270 180.745 ;
        RECT 110.115 178.535 110.445 179.165 ;
        RECT 110.615 178.365 110.825 179.185 ;
        RECT 111.060 179.075 111.270 179.725 ;
        RECT 112.010 179.605 112.180 180.195 ;
        RECT 113.400 180.025 113.570 180.405 ;
        RECT 114.505 180.285 114.675 180.745 ;
        RECT 114.845 180.455 115.215 180.915 ;
        RECT 115.510 180.315 115.680 180.655 ;
        RECT 115.850 180.485 116.180 180.915 ;
        RECT 116.415 180.315 116.585 180.655 ;
        RECT 112.350 179.855 113.570 180.025 ;
        RECT 113.740 179.945 114.200 180.235 ;
        RECT 114.505 180.115 115.065 180.285 ;
        RECT 115.510 180.145 116.585 180.315 ;
        RECT 116.755 180.415 117.435 180.745 ;
        RECT 117.650 180.415 117.900 180.745 ;
        RECT 118.070 180.455 118.320 180.915 ;
        RECT 114.895 179.975 115.065 180.115 ;
        RECT 113.740 179.935 114.705 179.945 ;
        RECT 113.400 179.765 113.570 179.855 ;
        RECT 114.030 179.775 114.705 179.935 ;
        RECT 111.440 179.575 112.180 179.605 ;
        RECT 111.440 179.275 112.355 179.575 ;
        RECT 112.030 179.100 112.355 179.275 ;
        RECT 111.060 178.545 111.315 179.075 ;
        RECT 111.485 178.365 111.790 178.825 ;
        RECT 112.035 178.745 112.355 179.100 ;
        RECT 112.525 179.315 113.065 179.685 ;
        RECT 113.400 179.595 113.805 179.765 ;
        RECT 112.525 178.915 112.765 179.315 ;
        RECT 113.245 179.145 113.465 179.425 ;
        RECT 112.935 178.975 113.465 179.145 ;
        RECT 112.935 178.745 113.105 178.975 ;
        RECT 113.635 178.815 113.805 179.595 ;
        RECT 113.975 178.985 114.325 179.605 ;
        RECT 114.495 178.985 114.705 179.775 ;
        RECT 114.895 179.805 116.395 179.975 ;
        RECT 114.895 179.115 115.065 179.805 ;
        RECT 116.755 179.635 116.925 180.415 ;
        RECT 117.730 180.285 117.900 180.415 ;
        RECT 115.235 179.465 116.925 179.635 ;
        RECT 117.095 179.855 117.560 180.245 ;
        RECT 117.730 180.115 118.125 180.285 ;
        RECT 115.235 179.285 115.405 179.465 ;
        RECT 112.035 178.575 113.105 178.745 ;
        RECT 113.275 178.365 113.465 178.805 ;
        RECT 113.635 178.535 114.585 178.815 ;
        RECT 114.895 178.725 115.155 179.115 ;
        RECT 115.575 179.045 116.365 179.295 ;
        RECT 114.805 178.555 115.155 178.725 ;
        RECT 115.365 178.365 115.695 178.825 ;
        RECT 116.570 178.755 116.740 179.465 ;
        RECT 117.095 179.265 117.265 179.855 ;
        RECT 116.910 179.045 117.265 179.265 ;
        RECT 117.435 179.045 117.785 179.665 ;
        RECT 117.955 178.755 118.125 180.115 ;
        RECT 118.490 179.945 118.815 180.730 ;
        RECT 118.295 178.895 118.755 179.945 ;
        RECT 116.570 178.585 117.425 178.755 ;
        RECT 117.630 178.585 118.125 178.755 ;
        RECT 118.295 178.365 118.625 178.725 ;
        RECT 118.985 178.625 119.155 180.745 ;
        RECT 119.325 180.415 119.655 180.915 ;
        RECT 119.825 180.245 120.080 180.745 ;
        RECT 119.330 180.075 120.080 180.245 ;
        RECT 119.330 179.085 119.560 180.075 ;
        RECT 119.730 179.255 120.080 179.905 ;
        RECT 120.295 179.775 120.525 180.915 ;
        RECT 120.695 179.765 121.025 180.745 ;
        RECT 121.195 179.775 121.405 180.915 ;
        RECT 121.725 179.985 121.895 180.745 ;
        RECT 122.075 180.155 122.405 180.915 ;
        RECT 121.725 179.815 122.390 179.985 ;
        RECT 122.575 179.840 122.845 180.745 ;
        RECT 120.275 179.355 120.605 179.605 ;
        RECT 119.330 178.915 120.080 179.085 ;
        RECT 119.325 178.365 119.655 178.745 ;
        RECT 119.825 178.625 120.080 178.915 ;
        RECT 120.295 178.365 120.525 179.185 ;
        RECT 120.775 179.165 121.025 179.765 ;
        RECT 122.220 179.670 122.390 179.815 ;
        RECT 121.655 179.265 121.985 179.635 ;
        RECT 122.220 179.340 122.505 179.670 ;
        RECT 120.695 178.535 121.025 179.165 ;
        RECT 121.195 178.365 121.405 179.185 ;
        RECT 122.220 179.085 122.390 179.340 ;
        RECT 121.725 178.915 122.390 179.085 ;
        RECT 122.675 179.040 122.845 179.840 ;
        RECT 123.475 179.825 126.065 180.915 ;
        RECT 126.235 179.825 127.445 180.915 ;
        RECT 123.475 179.305 124.685 179.825 ;
        RECT 124.855 179.135 126.065 179.655 ;
        RECT 126.235 179.285 126.755 179.825 ;
        RECT 121.725 178.535 121.895 178.915 ;
        RECT 122.075 178.365 122.405 178.745 ;
        RECT 122.585 178.535 122.845 179.040 ;
        RECT 123.475 178.365 126.065 179.135 ;
        RECT 126.925 179.115 127.445 179.655 ;
        RECT 126.235 178.365 127.445 179.115 ;
        RECT 14.370 178.195 127.530 178.365 ;
        RECT 14.455 177.445 15.665 178.195 ;
        RECT 14.455 176.905 14.975 177.445 ;
        RECT 15.835 177.425 19.345 178.195 ;
        RECT 19.520 177.650 24.865 178.195 ;
        RECT 15.145 176.735 15.665 177.275 ;
        RECT 14.455 175.645 15.665 176.735 ;
        RECT 15.835 176.735 17.525 177.255 ;
        RECT 17.695 176.905 19.345 177.425 ;
        RECT 15.835 175.645 19.345 176.735 ;
        RECT 21.110 176.080 21.460 177.330 ;
        RECT 22.940 176.820 23.280 177.650 ;
        RECT 25.095 177.375 25.305 178.195 ;
        RECT 25.475 177.395 25.805 178.025 ;
        RECT 25.475 176.795 25.725 177.395 ;
        RECT 25.975 177.375 26.205 178.195 ;
        RECT 26.455 177.375 26.685 178.195 ;
        RECT 26.855 177.395 27.185 178.025 ;
        RECT 25.895 176.955 26.225 177.205 ;
        RECT 26.435 176.955 26.765 177.205 ;
        RECT 26.935 176.795 27.185 177.395 ;
        RECT 27.355 177.375 27.565 178.195 ;
        RECT 27.800 177.485 28.055 178.015 ;
        RECT 28.225 177.735 28.530 178.195 ;
        RECT 28.775 177.815 29.845 177.985 ;
        RECT 19.520 175.645 24.865 176.080 ;
        RECT 25.095 175.645 25.305 176.785 ;
        RECT 25.475 175.815 25.805 176.795 ;
        RECT 25.975 175.645 26.205 176.785 ;
        RECT 26.455 175.645 26.685 176.785 ;
        RECT 26.855 175.815 27.185 176.795 ;
        RECT 27.800 176.835 28.010 177.485 ;
        RECT 28.775 177.460 29.095 177.815 ;
        RECT 28.770 177.285 29.095 177.460 ;
        RECT 28.180 176.985 29.095 177.285 ;
        RECT 29.265 177.245 29.505 177.645 ;
        RECT 29.675 177.585 29.845 177.815 ;
        RECT 30.015 177.755 30.205 178.195 ;
        RECT 30.375 177.745 31.325 178.025 ;
        RECT 31.545 177.835 31.895 178.005 ;
        RECT 29.675 177.415 30.205 177.585 ;
        RECT 28.180 176.955 28.920 176.985 ;
        RECT 27.355 175.645 27.565 176.785 ;
        RECT 27.800 175.955 28.055 176.835 ;
        RECT 28.225 175.645 28.530 176.785 ;
        RECT 28.750 176.365 28.920 176.955 ;
        RECT 29.265 176.875 29.805 177.245 ;
        RECT 29.985 177.135 30.205 177.415 ;
        RECT 30.375 176.965 30.545 177.745 ;
        RECT 30.140 176.795 30.545 176.965 ;
        RECT 30.715 176.955 31.065 177.575 ;
        RECT 30.140 176.705 30.310 176.795 ;
        RECT 31.235 176.785 31.445 177.575 ;
        RECT 29.090 176.535 30.310 176.705 ;
        RECT 30.770 176.625 31.445 176.785 ;
        RECT 28.750 176.195 29.550 176.365 ;
        RECT 28.870 175.645 29.200 176.025 ;
        RECT 29.380 175.905 29.550 176.195 ;
        RECT 30.140 176.155 30.310 176.535 ;
        RECT 30.480 176.615 31.445 176.625 ;
        RECT 31.635 177.445 31.895 177.835 ;
        RECT 32.105 177.735 32.435 178.195 ;
        RECT 33.310 177.805 34.165 177.975 ;
        RECT 34.370 177.805 34.865 177.975 ;
        RECT 35.035 177.835 35.365 178.195 ;
        RECT 31.635 176.755 31.805 177.445 ;
        RECT 31.975 177.095 32.145 177.275 ;
        RECT 32.315 177.265 33.105 177.515 ;
        RECT 33.310 177.095 33.480 177.805 ;
        RECT 33.650 177.295 34.005 177.515 ;
        RECT 31.975 176.925 33.665 177.095 ;
        RECT 30.480 176.325 30.940 176.615 ;
        RECT 31.635 176.585 33.135 176.755 ;
        RECT 31.635 176.445 31.805 176.585 ;
        RECT 31.245 176.275 31.805 176.445 ;
        RECT 29.720 175.645 29.970 176.105 ;
        RECT 30.140 175.815 31.010 176.155 ;
        RECT 31.245 175.815 31.415 176.275 ;
        RECT 32.250 176.245 33.325 176.415 ;
        RECT 31.585 175.645 31.955 176.105 ;
        RECT 32.250 175.905 32.420 176.245 ;
        RECT 32.590 175.645 32.920 176.075 ;
        RECT 33.155 175.905 33.325 176.245 ;
        RECT 33.495 176.145 33.665 176.925 ;
        RECT 33.835 176.705 34.005 177.295 ;
        RECT 34.175 176.895 34.525 177.515 ;
        RECT 33.835 176.315 34.300 176.705 ;
        RECT 34.695 176.445 34.865 177.805 ;
        RECT 35.035 176.615 35.495 177.665 ;
        RECT 34.470 176.275 34.865 176.445 ;
        RECT 34.470 176.145 34.640 176.275 ;
        RECT 33.495 175.815 34.175 176.145 ;
        RECT 34.390 175.815 34.640 176.145 ;
        RECT 34.810 175.645 35.060 176.105 ;
        RECT 35.230 175.830 35.555 176.615 ;
        RECT 35.725 175.815 35.895 177.935 ;
        RECT 36.065 177.815 36.395 178.195 ;
        RECT 36.565 177.645 36.820 177.935 ;
        RECT 36.070 177.475 36.820 177.645 ;
        RECT 36.070 176.485 36.300 177.475 ;
        RECT 36.995 177.470 37.285 178.195 ;
        RECT 37.730 177.385 37.975 177.990 ;
        RECT 38.195 177.660 38.705 178.195 ;
        RECT 36.470 176.655 36.820 177.305 ;
        RECT 37.455 177.215 38.685 177.385 ;
        RECT 36.070 176.315 36.820 176.485 ;
        RECT 36.065 175.645 36.395 176.145 ;
        RECT 36.565 175.815 36.820 176.315 ;
        RECT 36.995 175.645 37.285 176.810 ;
        RECT 37.455 176.405 37.795 177.215 ;
        RECT 37.965 176.650 38.715 176.840 ;
        RECT 37.455 175.995 37.970 176.405 ;
        RECT 38.205 175.645 38.375 176.405 ;
        RECT 38.545 175.985 38.715 176.650 ;
        RECT 38.885 176.665 39.075 178.025 ;
        RECT 39.245 177.855 39.520 178.025 ;
        RECT 39.245 177.685 39.525 177.855 ;
        RECT 39.245 176.865 39.520 177.685 ;
        RECT 39.710 177.660 40.240 178.025 ;
        RECT 40.665 177.795 40.995 178.195 ;
        RECT 40.065 177.625 40.240 177.660 ;
        RECT 39.725 176.665 39.895 177.465 ;
        RECT 38.885 176.495 39.895 176.665 ;
        RECT 40.065 177.455 40.995 177.625 ;
        RECT 41.165 177.455 41.420 178.025 ;
        RECT 40.065 176.325 40.235 177.455 ;
        RECT 40.825 177.285 40.995 177.455 ;
        RECT 39.110 176.155 40.235 176.325 ;
        RECT 40.405 176.955 40.600 177.285 ;
        RECT 40.825 176.955 41.080 177.285 ;
        RECT 40.405 175.985 40.575 176.955 ;
        RECT 41.250 176.785 41.420 177.455 ;
        RECT 42.630 177.565 42.915 178.025 ;
        RECT 43.085 177.735 43.355 178.195 ;
        RECT 42.630 177.395 43.585 177.565 ;
        RECT 38.545 175.815 40.575 175.985 ;
        RECT 40.745 175.645 40.915 176.785 ;
        RECT 41.085 175.815 41.420 176.785 ;
        RECT 42.515 176.665 43.205 177.225 ;
        RECT 43.375 176.495 43.585 177.395 ;
        RECT 42.630 176.275 43.585 176.495 ;
        RECT 43.755 177.225 44.155 178.025 ;
        RECT 44.345 177.565 44.625 178.025 ;
        RECT 45.145 177.735 45.470 178.195 ;
        RECT 44.345 177.395 45.470 177.565 ;
        RECT 45.640 177.455 46.025 178.025 ;
        RECT 45.020 177.285 45.470 177.395 ;
        RECT 43.755 176.665 44.850 177.225 ;
        RECT 45.020 176.955 45.575 177.285 ;
        RECT 42.630 175.815 42.915 176.275 ;
        RECT 43.085 175.645 43.355 176.105 ;
        RECT 43.755 175.815 44.155 176.665 ;
        RECT 45.020 176.495 45.470 176.955 ;
        RECT 45.745 176.785 46.025 177.455 ;
        RECT 46.400 177.415 46.900 178.025 ;
        RECT 46.195 176.955 46.545 177.205 ;
        RECT 46.730 176.785 46.900 177.415 ;
        RECT 47.530 177.545 47.860 178.025 ;
        RECT 48.030 177.735 48.255 178.195 ;
        RECT 48.425 177.545 48.755 178.025 ;
        RECT 47.530 177.375 48.755 177.545 ;
        RECT 48.945 177.395 49.195 178.195 ;
        RECT 49.365 177.395 49.705 178.025 ;
        RECT 49.990 177.565 50.275 178.025 ;
        RECT 50.445 177.735 50.715 178.195 ;
        RECT 49.990 177.395 50.945 177.565 ;
        RECT 47.070 177.005 47.400 177.205 ;
        RECT 47.570 177.005 47.900 177.205 ;
        RECT 48.070 177.005 48.490 177.205 ;
        RECT 48.665 177.035 49.360 177.205 ;
        RECT 48.665 176.785 48.835 177.035 ;
        RECT 49.530 176.785 49.705 177.395 ;
        RECT 44.345 176.275 45.470 176.495 ;
        RECT 44.345 175.815 44.625 176.275 ;
        RECT 45.145 175.645 45.470 176.105 ;
        RECT 45.640 175.815 46.025 176.785 ;
        RECT 46.400 176.615 48.835 176.785 ;
        RECT 46.400 175.815 46.730 176.615 ;
        RECT 46.900 175.645 47.230 176.445 ;
        RECT 47.530 175.815 47.860 176.615 ;
        RECT 48.505 175.645 48.755 176.445 ;
        RECT 49.025 175.645 49.195 176.785 ;
        RECT 49.365 175.815 49.705 176.785 ;
        RECT 49.875 176.665 50.565 177.225 ;
        RECT 50.735 176.495 50.945 177.395 ;
        RECT 49.990 176.275 50.945 176.495 ;
        RECT 51.115 177.225 51.515 178.025 ;
        RECT 51.705 177.565 51.985 178.025 ;
        RECT 52.505 177.735 52.830 178.195 ;
        RECT 51.705 177.395 52.830 177.565 ;
        RECT 53.000 177.455 53.385 178.025 ;
        RECT 52.380 177.285 52.830 177.395 ;
        RECT 51.115 176.665 52.210 177.225 ;
        RECT 52.380 176.955 52.935 177.285 ;
        RECT 49.990 175.815 50.275 176.275 ;
        RECT 50.445 175.645 50.715 176.105 ;
        RECT 51.115 175.815 51.515 176.665 ;
        RECT 52.380 176.495 52.830 176.955 ;
        RECT 53.105 176.785 53.385 177.455 ;
        RECT 51.705 176.275 52.830 176.495 ;
        RECT 51.705 175.815 51.985 176.275 ;
        RECT 52.505 175.645 52.830 176.105 ;
        RECT 53.000 175.815 53.385 176.785 ;
        RECT 53.560 177.485 53.815 178.015 ;
        RECT 53.985 177.735 54.290 178.195 ;
        RECT 54.535 177.815 55.605 177.985 ;
        RECT 53.560 176.835 53.770 177.485 ;
        RECT 54.535 177.460 54.855 177.815 ;
        RECT 54.530 177.285 54.855 177.460 ;
        RECT 53.940 176.985 54.855 177.285 ;
        RECT 55.025 177.245 55.265 177.645 ;
        RECT 55.435 177.585 55.605 177.815 ;
        RECT 55.775 177.755 55.965 178.195 ;
        RECT 56.135 177.745 57.085 178.025 ;
        RECT 57.305 177.835 57.655 178.005 ;
        RECT 55.435 177.415 55.965 177.585 ;
        RECT 53.940 176.955 54.680 176.985 ;
        RECT 53.560 175.955 53.815 176.835 ;
        RECT 53.985 175.645 54.290 176.785 ;
        RECT 54.510 176.365 54.680 176.955 ;
        RECT 55.025 176.875 55.565 177.245 ;
        RECT 55.745 177.135 55.965 177.415 ;
        RECT 56.135 176.965 56.305 177.745 ;
        RECT 55.900 176.795 56.305 176.965 ;
        RECT 56.475 176.955 56.825 177.575 ;
        RECT 55.900 176.705 56.070 176.795 ;
        RECT 56.995 176.785 57.205 177.575 ;
        RECT 54.850 176.535 56.070 176.705 ;
        RECT 56.530 176.625 57.205 176.785 ;
        RECT 54.510 176.195 55.310 176.365 ;
        RECT 54.630 175.645 54.960 176.025 ;
        RECT 55.140 175.905 55.310 176.195 ;
        RECT 55.900 176.155 56.070 176.535 ;
        RECT 56.240 176.615 57.205 176.625 ;
        RECT 57.395 177.445 57.655 177.835 ;
        RECT 57.865 177.735 58.195 178.195 ;
        RECT 59.070 177.805 59.925 177.975 ;
        RECT 60.130 177.805 60.625 177.975 ;
        RECT 60.795 177.835 61.125 178.195 ;
        RECT 57.395 176.755 57.565 177.445 ;
        RECT 57.735 177.095 57.905 177.275 ;
        RECT 58.075 177.265 58.865 177.515 ;
        RECT 59.070 177.095 59.240 177.805 ;
        RECT 59.410 177.295 59.765 177.515 ;
        RECT 57.735 176.925 59.425 177.095 ;
        RECT 56.240 176.325 56.700 176.615 ;
        RECT 57.395 176.585 58.895 176.755 ;
        RECT 57.395 176.445 57.565 176.585 ;
        RECT 57.005 176.275 57.565 176.445 ;
        RECT 55.480 175.645 55.730 176.105 ;
        RECT 55.900 175.815 56.770 176.155 ;
        RECT 57.005 175.815 57.175 176.275 ;
        RECT 58.010 176.245 59.085 176.415 ;
        RECT 57.345 175.645 57.715 176.105 ;
        RECT 58.010 175.905 58.180 176.245 ;
        RECT 58.350 175.645 58.680 176.075 ;
        RECT 58.915 175.905 59.085 176.245 ;
        RECT 59.255 176.145 59.425 176.925 ;
        RECT 59.595 176.705 59.765 177.295 ;
        RECT 59.935 176.895 60.285 177.515 ;
        RECT 59.595 176.315 60.060 176.705 ;
        RECT 60.455 176.445 60.625 177.805 ;
        RECT 60.795 176.615 61.255 177.665 ;
        RECT 60.230 176.275 60.625 176.445 ;
        RECT 60.230 176.145 60.400 176.275 ;
        RECT 59.255 175.815 59.935 176.145 ;
        RECT 60.150 175.815 60.400 176.145 ;
        RECT 60.570 175.645 60.820 176.105 ;
        RECT 60.990 175.830 61.315 176.615 ;
        RECT 61.485 175.815 61.655 177.935 ;
        RECT 61.825 177.815 62.155 178.195 ;
        RECT 62.325 177.645 62.580 177.935 ;
        RECT 61.830 177.475 62.580 177.645 ;
        RECT 61.830 176.485 62.060 177.475 ;
        RECT 62.755 177.470 63.045 178.195 ;
        RECT 63.215 177.520 63.475 178.025 ;
        RECT 63.655 177.815 63.985 178.195 ;
        RECT 64.165 177.645 64.335 178.025 ;
        RECT 62.230 176.655 62.580 177.305 ;
        RECT 61.830 176.315 62.580 176.485 ;
        RECT 61.825 175.645 62.155 176.145 ;
        RECT 62.325 175.815 62.580 176.315 ;
        RECT 62.755 175.645 63.045 176.810 ;
        RECT 63.215 176.720 63.385 177.520 ;
        RECT 63.670 177.475 64.335 177.645 ;
        RECT 63.670 177.220 63.840 177.475 ;
        RECT 64.595 177.425 67.185 178.195 ;
        RECT 63.555 176.890 63.840 177.220 ;
        RECT 64.075 176.925 64.405 177.295 ;
        RECT 63.670 176.745 63.840 176.890 ;
        RECT 63.215 175.815 63.485 176.720 ;
        RECT 63.670 176.575 64.335 176.745 ;
        RECT 63.655 175.645 63.985 176.405 ;
        RECT 64.165 175.815 64.335 176.575 ;
        RECT 64.595 176.735 65.805 177.255 ;
        RECT 65.975 176.905 67.185 177.425 ;
        RECT 67.360 177.355 67.620 178.195 ;
        RECT 67.795 177.450 68.050 178.025 ;
        RECT 68.220 177.815 68.550 178.195 ;
        RECT 68.765 177.645 68.935 178.025 ;
        RECT 68.220 177.475 68.935 177.645 ;
        RECT 69.285 177.645 69.455 178.025 ;
        RECT 69.670 177.815 70.000 178.195 ;
        RECT 69.285 177.475 70.000 177.645 ;
        RECT 64.595 175.645 67.185 176.735 ;
        RECT 67.360 175.645 67.620 176.795 ;
        RECT 67.795 176.720 67.965 177.450 ;
        RECT 68.220 177.285 68.390 177.475 ;
        RECT 68.135 176.955 68.390 177.285 ;
        RECT 68.220 176.745 68.390 176.955 ;
        RECT 68.670 176.925 69.025 177.295 ;
        RECT 69.195 176.925 69.550 177.295 ;
        RECT 69.830 177.285 70.000 177.475 ;
        RECT 70.170 177.450 70.425 178.025 ;
        RECT 69.830 176.955 70.085 177.285 ;
        RECT 69.830 176.745 70.000 176.955 ;
        RECT 67.795 175.815 68.050 176.720 ;
        RECT 68.220 176.575 68.935 176.745 ;
        RECT 68.220 175.645 68.550 176.405 ;
        RECT 68.765 175.815 68.935 176.575 ;
        RECT 69.285 176.575 70.000 176.745 ;
        RECT 70.255 176.720 70.425 177.450 ;
        RECT 70.600 177.355 70.860 178.195 ;
        RECT 71.125 177.645 71.295 178.025 ;
        RECT 71.510 177.815 71.840 178.195 ;
        RECT 71.125 177.475 71.840 177.645 ;
        RECT 71.035 176.925 71.390 177.295 ;
        RECT 71.670 177.285 71.840 177.475 ;
        RECT 72.010 177.450 72.265 178.025 ;
        RECT 71.670 176.955 71.925 177.285 ;
        RECT 69.285 175.815 69.455 176.575 ;
        RECT 69.670 175.645 70.000 176.405 ;
        RECT 70.170 175.815 70.425 176.720 ;
        RECT 70.600 175.645 70.860 176.795 ;
        RECT 71.670 176.745 71.840 176.955 ;
        RECT 71.125 176.575 71.840 176.745 ;
        RECT 72.095 176.720 72.265 177.450 ;
        RECT 72.440 177.355 72.700 178.195 ;
        RECT 72.875 177.435 73.585 178.025 ;
        RECT 74.095 177.665 74.425 178.025 ;
        RECT 74.625 177.835 74.955 178.195 ;
        RECT 75.125 177.665 75.455 178.025 ;
        RECT 74.095 177.455 75.455 177.665 ;
        RECT 71.125 175.815 71.295 176.575 ;
        RECT 71.510 175.645 71.840 176.405 ;
        RECT 72.010 175.815 72.265 176.720 ;
        RECT 72.440 175.645 72.700 176.795 ;
        RECT 72.875 176.465 73.080 177.435 ;
        RECT 76.300 177.415 76.800 178.025 ;
        RECT 73.250 176.665 73.580 177.205 ;
        RECT 73.755 176.955 74.250 177.285 ;
        RECT 74.570 176.955 74.945 177.285 ;
        RECT 75.155 176.955 75.465 177.285 ;
        RECT 76.095 176.955 76.445 177.205 ;
        RECT 73.755 176.665 74.080 176.955 ;
        RECT 74.275 176.465 74.605 176.685 ;
        RECT 72.875 176.235 74.605 176.465 ;
        RECT 72.875 175.815 73.575 176.235 ;
        RECT 73.775 175.645 74.105 176.005 ;
        RECT 74.275 175.835 74.605 176.235 ;
        RECT 74.775 176.030 74.945 176.955 ;
        RECT 76.630 176.785 76.800 177.415 ;
        RECT 77.430 177.545 77.760 178.025 ;
        RECT 77.930 177.735 78.155 178.195 ;
        RECT 78.325 177.545 78.655 178.025 ;
        RECT 77.430 177.375 78.655 177.545 ;
        RECT 78.845 177.395 79.095 178.195 ;
        RECT 79.265 177.395 79.605 178.025 ;
        RECT 76.970 177.005 77.300 177.205 ;
        RECT 77.470 177.005 77.800 177.205 ;
        RECT 77.970 177.005 78.390 177.205 ;
        RECT 78.565 177.035 79.260 177.205 ;
        RECT 78.565 176.785 78.735 177.035 ;
        RECT 79.430 176.835 79.605 177.395 ;
        RECT 79.375 176.785 79.605 176.835 ;
        RECT 75.125 175.645 75.455 176.705 ;
        RECT 76.300 176.615 78.735 176.785 ;
        RECT 76.300 175.815 76.630 176.615 ;
        RECT 76.800 175.645 77.130 176.445 ;
        RECT 77.430 175.815 77.760 176.615 ;
        RECT 78.405 175.645 78.655 176.445 ;
        RECT 78.925 175.645 79.095 176.785 ;
        RECT 79.265 175.815 79.605 176.785 ;
        RECT 79.775 177.395 80.115 178.025 ;
        RECT 80.285 177.395 80.535 178.195 ;
        RECT 80.725 177.545 81.055 178.025 ;
        RECT 81.225 177.735 81.450 178.195 ;
        RECT 81.620 177.545 81.950 178.025 ;
        RECT 79.775 177.345 80.005 177.395 ;
        RECT 80.725 177.375 81.950 177.545 ;
        RECT 82.580 177.415 83.080 178.025 ;
        RECT 83.455 177.445 84.665 178.195 ;
        RECT 79.775 176.785 79.950 177.345 ;
        RECT 80.120 177.035 80.815 177.205 ;
        RECT 80.645 176.785 80.815 177.035 ;
        RECT 80.990 177.005 81.410 177.205 ;
        RECT 81.580 177.005 81.910 177.205 ;
        RECT 82.080 177.005 82.410 177.205 ;
        RECT 82.580 176.785 82.750 177.415 ;
        RECT 82.935 176.955 83.285 177.205 ;
        RECT 79.775 175.815 80.115 176.785 ;
        RECT 80.285 175.645 80.455 176.785 ;
        RECT 80.645 176.615 83.080 176.785 ;
        RECT 80.725 175.645 80.975 176.445 ;
        RECT 81.620 175.815 81.950 176.615 ;
        RECT 82.250 175.645 82.580 176.445 ;
        RECT 82.750 175.815 83.080 176.615 ;
        RECT 83.455 176.735 83.975 177.275 ;
        RECT 84.145 176.905 84.665 177.445 ;
        RECT 84.950 177.565 85.235 178.025 ;
        RECT 85.405 177.735 85.675 178.195 ;
        RECT 84.950 177.395 85.905 177.565 ;
        RECT 83.455 175.645 84.665 176.735 ;
        RECT 84.835 176.665 85.525 177.225 ;
        RECT 85.695 176.495 85.905 177.395 ;
        RECT 84.950 176.275 85.905 176.495 ;
        RECT 86.075 177.225 86.475 178.025 ;
        RECT 86.665 177.565 86.945 178.025 ;
        RECT 87.465 177.735 87.790 178.195 ;
        RECT 86.665 177.395 87.790 177.565 ;
        RECT 87.960 177.455 88.345 178.025 ;
        RECT 88.515 177.470 88.805 178.195 ;
        RECT 87.340 177.285 87.790 177.395 ;
        RECT 86.075 176.665 87.170 177.225 ;
        RECT 87.340 176.955 87.895 177.285 ;
        RECT 84.950 175.815 85.235 176.275 ;
        RECT 85.405 175.645 85.675 176.105 ;
        RECT 86.075 175.815 86.475 176.665 ;
        RECT 87.340 176.495 87.790 176.955 ;
        RECT 88.065 176.785 88.345 177.455 ;
        RECT 88.975 177.425 92.485 178.195 ;
        RECT 92.660 177.650 98.005 178.195 ;
        RECT 86.665 176.275 87.790 176.495 ;
        RECT 86.665 175.815 86.945 176.275 ;
        RECT 87.465 175.645 87.790 176.105 ;
        RECT 87.960 175.815 88.345 176.785 ;
        RECT 88.515 175.645 88.805 176.810 ;
        RECT 88.975 176.735 90.665 177.255 ;
        RECT 90.835 176.905 92.485 177.425 ;
        RECT 88.975 175.645 92.485 176.735 ;
        RECT 94.250 176.080 94.600 177.330 ;
        RECT 96.080 176.820 96.420 177.650 ;
        RECT 98.380 177.415 98.880 178.025 ;
        RECT 98.175 176.955 98.525 177.205 ;
        RECT 98.710 176.785 98.880 177.415 ;
        RECT 99.510 177.545 99.840 178.025 ;
        RECT 100.010 177.735 100.235 178.195 ;
        RECT 100.405 177.545 100.735 178.025 ;
        RECT 99.510 177.375 100.735 177.545 ;
        RECT 100.925 177.395 101.175 178.195 ;
        RECT 101.345 177.395 101.685 178.025 ;
        RECT 99.050 177.005 99.380 177.205 ;
        RECT 99.550 177.005 99.880 177.205 ;
        RECT 100.050 177.005 100.470 177.205 ;
        RECT 100.645 177.035 101.340 177.205 ;
        RECT 100.645 176.785 100.815 177.035 ;
        RECT 101.510 176.785 101.685 177.395 ;
        RECT 98.380 176.615 100.815 176.785 ;
        RECT 92.660 175.645 98.005 176.080 ;
        RECT 98.380 175.815 98.710 176.615 ;
        RECT 98.880 175.645 99.210 176.445 ;
        RECT 99.510 175.815 99.840 176.615 ;
        RECT 100.485 175.645 100.735 176.445 ;
        RECT 101.005 175.645 101.175 176.785 ;
        RECT 101.345 175.815 101.685 176.785 ;
        RECT 101.855 177.520 102.115 178.025 ;
        RECT 102.295 177.815 102.625 178.195 ;
        RECT 102.805 177.645 102.975 178.025 ;
        RECT 101.855 176.720 102.025 177.520 ;
        RECT 102.310 177.475 102.975 177.645 ;
        RECT 102.310 177.220 102.480 177.475 ;
        RECT 103.235 177.445 104.445 178.195 ;
        RECT 102.195 176.890 102.480 177.220 ;
        RECT 102.715 176.925 103.045 177.295 ;
        RECT 102.310 176.745 102.480 176.890 ;
        RECT 101.855 175.815 102.125 176.720 ;
        RECT 102.310 176.575 102.975 176.745 ;
        RECT 102.295 175.645 102.625 176.405 ;
        RECT 102.805 175.815 102.975 176.575 ;
        RECT 103.235 176.735 103.755 177.275 ;
        RECT 103.925 176.905 104.445 177.445 ;
        RECT 104.615 177.395 104.955 178.025 ;
        RECT 105.125 177.395 105.375 178.195 ;
        RECT 105.565 177.545 105.895 178.025 ;
        RECT 106.065 177.735 106.290 178.195 ;
        RECT 106.460 177.545 106.790 178.025 ;
        RECT 104.615 176.785 104.790 177.395 ;
        RECT 105.565 177.375 106.790 177.545 ;
        RECT 107.420 177.415 107.920 178.025 ;
        RECT 108.295 177.425 109.965 178.195 ;
        RECT 104.960 177.035 105.655 177.205 ;
        RECT 105.485 176.785 105.655 177.035 ;
        RECT 105.830 177.005 106.250 177.205 ;
        RECT 106.420 177.005 106.750 177.205 ;
        RECT 106.920 177.005 107.250 177.205 ;
        RECT 107.420 176.785 107.590 177.415 ;
        RECT 107.775 176.955 108.125 177.205 ;
        RECT 103.235 175.645 104.445 176.735 ;
        RECT 104.615 175.815 104.955 176.785 ;
        RECT 105.125 175.645 105.295 176.785 ;
        RECT 105.485 176.615 107.920 176.785 ;
        RECT 105.565 175.645 105.815 176.445 ;
        RECT 106.460 175.815 106.790 176.615 ;
        RECT 107.090 175.645 107.420 176.445 ;
        RECT 107.590 175.815 107.920 176.615 ;
        RECT 108.295 176.735 109.045 177.255 ;
        RECT 109.215 176.905 109.965 177.425 ;
        RECT 110.410 177.385 110.655 177.990 ;
        RECT 110.875 177.660 111.385 178.195 ;
        RECT 110.135 177.215 111.365 177.385 ;
        RECT 108.295 175.645 109.965 176.735 ;
        RECT 110.135 176.405 110.475 177.215 ;
        RECT 110.645 176.650 111.395 176.840 ;
        RECT 110.135 175.995 110.650 176.405 ;
        RECT 110.885 175.645 111.055 176.405 ;
        RECT 111.225 175.985 111.395 176.650 ;
        RECT 111.565 176.665 111.755 178.025 ;
        RECT 111.925 177.855 112.200 178.025 ;
        RECT 111.925 177.685 112.205 177.855 ;
        RECT 111.925 176.865 112.200 177.685 ;
        RECT 112.390 177.660 112.920 178.025 ;
        RECT 113.345 177.795 113.675 178.195 ;
        RECT 112.745 177.625 112.920 177.660 ;
        RECT 112.405 176.665 112.575 177.465 ;
        RECT 111.565 176.495 112.575 176.665 ;
        RECT 112.745 177.455 113.675 177.625 ;
        RECT 113.845 177.455 114.100 178.025 ;
        RECT 114.275 177.470 114.565 178.195 ;
        RECT 112.745 176.325 112.915 177.455 ;
        RECT 113.505 177.285 113.675 177.455 ;
        RECT 111.790 176.155 112.915 176.325 ;
        RECT 113.085 176.955 113.280 177.285 ;
        RECT 113.505 176.955 113.760 177.285 ;
        RECT 113.085 175.985 113.255 176.955 ;
        RECT 113.930 176.785 114.100 177.455 ;
        RECT 114.735 177.425 116.405 178.195 ;
        RECT 116.665 177.645 116.835 178.025 ;
        RECT 117.015 177.815 117.345 178.195 ;
        RECT 116.665 177.475 117.330 177.645 ;
        RECT 117.525 177.520 117.785 178.025 ;
        RECT 111.225 175.815 113.255 175.985 ;
        RECT 113.425 175.645 113.595 176.785 ;
        RECT 113.765 175.815 114.100 176.785 ;
        RECT 114.275 175.645 114.565 176.810 ;
        RECT 114.735 176.735 115.485 177.255 ;
        RECT 115.655 176.905 116.405 177.425 ;
        RECT 116.595 176.925 116.925 177.295 ;
        RECT 117.160 177.220 117.330 177.475 ;
        RECT 117.160 176.890 117.445 177.220 ;
        RECT 117.160 176.745 117.330 176.890 ;
        RECT 114.735 175.645 116.405 176.735 ;
        RECT 116.665 176.575 117.330 176.745 ;
        RECT 117.615 176.720 117.785 177.520 ;
        RECT 117.955 177.425 120.545 178.195 ;
        RECT 120.720 177.650 126.065 178.195 ;
        RECT 116.665 175.815 116.835 176.575 ;
        RECT 117.015 175.645 117.345 176.405 ;
        RECT 117.515 175.815 117.785 176.720 ;
        RECT 117.955 176.735 119.165 177.255 ;
        RECT 119.335 176.905 120.545 177.425 ;
        RECT 117.955 175.645 120.545 176.735 ;
        RECT 122.310 176.080 122.660 177.330 ;
        RECT 124.140 176.820 124.480 177.650 ;
        RECT 126.235 177.445 127.445 178.195 ;
        RECT 126.235 176.735 126.755 177.275 ;
        RECT 126.925 176.905 127.445 177.445 ;
        RECT 120.720 175.645 126.065 176.080 ;
        RECT 126.235 175.645 127.445 176.735 ;
        RECT 14.370 175.475 127.530 175.645 ;
        RECT 14.455 174.385 15.665 175.475 ;
        RECT 14.455 173.675 14.975 174.215 ;
        RECT 15.145 173.845 15.665 174.385 ;
        RECT 15.835 174.385 18.425 175.475 ;
        RECT 18.600 175.040 23.945 175.475 ;
        RECT 15.835 173.865 17.045 174.385 ;
        RECT 17.215 173.695 18.425 174.215 ;
        RECT 20.190 173.790 20.540 175.040 ;
        RECT 24.115 174.310 24.405 175.475 ;
        RECT 25.495 174.400 25.765 175.305 ;
        RECT 25.935 174.715 26.265 175.475 ;
        RECT 26.445 174.545 26.615 175.305 ;
        RECT 26.990 174.845 27.275 175.305 ;
        RECT 27.445 175.015 27.715 175.475 ;
        RECT 26.990 174.625 27.945 174.845 ;
        RECT 14.455 172.925 15.665 173.675 ;
        RECT 15.835 172.925 18.425 173.695 ;
        RECT 22.020 173.470 22.360 174.300 ;
        RECT 18.600 172.925 23.945 173.470 ;
        RECT 24.115 172.925 24.405 173.650 ;
        RECT 25.495 173.600 25.665 174.400 ;
        RECT 25.950 174.375 26.615 174.545 ;
        RECT 25.950 174.230 26.120 174.375 ;
        RECT 25.835 173.900 26.120 174.230 ;
        RECT 25.950 173.645 26.120 173.900 ;
        RECT 26.355 173.825 26.685 174.195 ;
        RECT 26.875 173.895 27.565 174.455 ;
        RECT 27.735 173.725 27.945 174.625 ;
        RECT 25.495 173.095 25.755 173.600 ;
        RECT 25.950 173.475 26.615 173.645 ;
        RECT 25.935 172.925 26.265 173.305 ;
        RECT 26.445 173.095 26.615 173.475 ;
        RECT 26.990 173.555 27.945 173.725 ;
        RECT 28.115 174.455 28.515 175.305 ;
        RECT 28.705 174.845 28.985 175.305 ;
        RECT 29.505 175.015 29.830 175.475 ;
        RECT 28.705 174.625 29.830 174.845 ;
        RECT 28.115 173.895 29.210 174.455 ;
        RECT 29.380 174.165 29.830 174.625 ;
        RECT 30.000 174.335 30.385 175.305 ;
        RECT 26.990 173.095 27.275 173.555 ;
        RECT 27.445 172.925 27.715 173.385 ;
        RECT 28.115 173.095 28.515 173.895 ;
        RECT 29.380 173.835 29.935 174.165 ;
        RECT 29.380 173.725 29.830 173.835 ;
        RECT 28.705 173.555 29.830 173.725 ;
        RECT 30.105 173.665 30.385 174.335 ;
        RECT 28.705 173.095 28.985 173.555 ;
        RECT 29.505 172.925 29.830 173.385 ;
        RECT 30.000 173.095 30.385 173.665 ;
        RECT 30.560 174.335 30.895 175.305 ;
        RECT 31.065 174.335 31.235 175.475 ;
        RECT 31.405 175.135 33.435 175.305 ;
        RECT 30.560 173.665 30.730 174.335 ;
        RECT 31.405 174.165 31.575 175.135 ;
        RECT 30.900 173.835 31.155 174.165 ;
        RECT 31.380 173.835 31.575 174.165 ;
        RECT 31.745 174.795 32.870 174.965 ;
        RECT 30.985 173.665 31.155 173.835 ;
        RECT 31.745 173.665 31.915 174.795 ;
        RECT 30.560 173.095 30.815 173.665 ;
        RECT 30.985 173.495 31.915 173.665 ;
        RECT 32.085 174.455 33.095 174.625 ;
        RECT 32.085 173.655 32.255 174.455 ;
        RECT 32.460 174.115 32.735 174.255 ;
        RECT 32.455 173.945 32.735 174.115 ;
        RECT 31.740 173.460 31.915 173.495 ;
        RECT 30.985 172.925 31.315 173.325 ;
        RECT 31.740 173.095 32.270 173.460 ;
        RECT 32.460 173.095 32.735 173.945 ;
        RECT 32.905 173.095 33.095 174.455 ;
        RECT 33.265 174.470 33.435 175.135 ;
        RECT 33.605 174.715 33.775 175.475 ;
        RECT 34.010 174.715 34.525 175.125 ;
        RECT 33.265 174.280 34.015 174.470 ;
        RECT 34.185 173.905 34.525 174.715 ;
        RECT 35.360 174.505 35.690 175.305 ;
        RECT 35.860 174.675 36.190 175.475 ;
        RECT 36.490 174.505 36.820 175.305 ;
        RECT 37.465 174.675 37.715 175.475 ;
        RECT 35.360 174.335 37.795 174.505 ;
        RECT 37.985 174.335 38.155 175.475 ;
        RECT 38.325 174.335 38.665 175.305 ;
        RECT 35.155 173.915 35.505 174.165 ;
        RECT 33.295 173.735 34.525 173.905 ;
        RECT 33.275 172.925 33.785 173.460 ;
        RECT 34.005 173.130 34.250 173.735 ;
        RECT 35.690 173.705 35.860 174.335 ;
        RECT 36.030 173.915 36.360 174.115 ;
        RECT 36.530 173.915 36.860 174.115 ;
        RECT 37.030 173.915 37.450 174.115 ;
        RECT 37.625 174.085 37.795 174.335 ;
        RECT 37.625 173.915 38.320 174.085 ;
        RECT 38.490 173.775 38.665 174.335 ;
        RECT 35.360 173.095 35.860 173.705 ;
        RECT 36.490 173.575 37.715 173.745 ;
        RECT 38.435 173.725 38.665 173.775 ;
        RECT 36.490 173.095 36.820 173.575 ;
        RECT 36.990 172.925 37.215 173.385 ;
        RECT 37.385 173.095 37.715 173.575 ;
        RECT 37.905 172.925 38.155 173.725 ;
        RECT 38.325 173.095 38.665 173.725 ;
        RECT 38.835 174.335 39.175 175.305 ;
        RECT 39.345 174.335 39.515 175.475 ;
        RECT 39.785 174.675 40.035 175.475 ;
        RECT 40.680 174.505 41.010 175.305 ;
        RECT 41.310 174.675 41.640 175.475 ;
        RECT 41.810 174.505 42.140 175.305 ;
        RECT 39.705 174.335 42.140 174.505 ;
        RECT 42.720 174.505 43.050 175.305 ;
        RECT 43.220 174.675 43.550 175.475 ;
        RECT 43.850 174.505 44.180 175.305 ;
        RECT 44.825 174.675 45.075 175.475 ;
        RECT 42.720 174.335 45.155 174.505 ;
        RECT 45.345 174.335 45.515 175.475 ;
        RECT 45.685 174.335 46.025 175.305 ;
        RECT 46.310 174.845 46.595 175.305 ;
        RECT 46.765 175.015 47.035 175.475 ;
        RECT 46.310 174.625 47.265 174.845 ;
        RECT 38.835 173.725 39.010 174.335 ;
        RECT 39.705 174.085 39.875 174.335 ;
        RECT 39.180 173.915 39.875 174.085 ;
        RECT 40.050 173.915 40.470 174.115 ;
        RECT 40.640 173.915 40.970 174.115 ;
        RECT 41.140 173.915 41.470 174.115 ;
        RECT 38.835 173.095 39.175 173.725 ;
        RECT 39.345 172.925 39.595 173.725 ;
        RECT 39.785 173.575 41.010 173.745 ;
        RECT 39.785 173.095 40.115 173.575 ;
        RECT 40.285 172.925 40.510 173.385 ;
        RECT 40.680 173.095 41.010 173.575 ;
        RECT 41.640 173.705 41.810 174.335 ;
        RECT 41.995 173.915 42.345 174.165 ;
        RECT 42.515 173.915 42.865 174.165 ;
        RECT 43.050 173.705 43.220 174.335 ;
        RECT 43.390 173.915 43.720 174.115 ;
        RECT 43.890 173.915 44.220 174.115 ;
        RECT 44.390 173.915 44.810 174.115 ;
        RECT 44.985 174.085 45.155 174.335 ;
        RECT 44.985 173.915 45.680 174.085 ;
        RECT 45.850 173.775 46.025 174.335 ;
        RECT 46.195 173.895 46.885 174.455 ;
        RECT 41.640 173.095 42.140 173.705 ;
        RECT 42.720 173.095 43.220 173.705 ;
        RECT 43.850 173.575 45.075 173.745 ;
        RECT 45.795 173.725 46.025 173.775 ;
        RECT 47.055 173.725 47.265 174.625 ;
        RECT 43.850 173.095 44.180 173.575 ;
        RECT 44.350 172.925 44.575 173.385 ;
        RECT 44.745 173.095 45.075 173.575 ;
        RECT 45.265 172.925 45.515 173.725 ;
        RECT 45.685 173.095 46.025 173.725 ;
        RECT 46.310 173.555 47.265 173.725 ;
        RECT 47.435 174.455 47.835 175.305 ;
        RECT 48.025 174.845 48.305 175.305 ;
        RECT 48.825 175.015 49.150 175.475 ;
        RECT 48.025 174.625 49.150 174.845 ;
        RECT 47.435 173.895 48.530 174.455 ;
        RECT 48.700 174.165 49.150 174.625 ;
        RECT 49.320 174.335 49.705 175.305 ;
        RECT 46.310 173.095 46.595 173.555 ;
        RECT 46.765 172.925 47.035 173.385 ;
        RECT 47.435 173.095 47.835 173.895 ;
        RECT 48.700 173.835 49.255 174.165 ;
        RECT 48.700 173.725 49.150 173.835 ;
        RECT 48.025 173.555 49.150 173.725 ;
        RECT 49.425 173.665 49.705 174.335 ;
        RECT 49.875 174.310 50.165 175.475 ;
        RECT 50.335 174.385 52.925 175.475 ;
        RECT 53.095 174.715 53.610 175.125 ;
        RECT 53.845 174.715 54.015 175.475 ;
        RECT 54.185 175.135 56.215 175.305 ;
        RECT 50.335 173.865 51.545 174.385 ;
        RECT 51.715 173.695 52.925 174.215 ;
        RECT 53.095 173.905 53.435 174.715 ;
        RECT 54.185 174.470 54.355 175.135 ;
        RECT 54.750 174.795 55.875 174.965 ;
        RECT 53.605 174.280 54.355 174.470 ;
        RECT 54.525 174.455 55.535 174.625 ;
        RECT 53.095 173.735 54.325 173.905 ;
        RECT 48.025 173.095 48.305 173.555 ;
        RECT 48.825 172.925 49.150 173.385 ;
        RECT 49.320 173.095 49.705 173.665 ;
        RECT 49.875 172.925 50.165 173.650 ;
        RECT 50.335 172.925 52.925 173.695 ;
        RECT 53.370 173.130 53.615 173.735 ;
        RECT 53.835 172.925 54.345 173.460 ;
        RECT 54.525 173.095 54.715 174.455 ;
        RECT 54.885 174.115 55.160 174.255 ;
        RECT 54.885 173.945 55.165 174.115 ;
        RECT 54.885 173.095 55.160 173.945 ;
        RECT 55.365 173.655 55.535 174.455 ;
        RECT 55.705 173.665 55.875 174.795 ;
        RECT 56.045 174.165 56.215 175.135 ;
        RECT 56.385 174.335 56.555 175.475 ;
        RECT 56.725 174.335 57.060 175.305 ;
        RECT 56.045 173.835 56.240 174.165 ;
        RECT 56.465 173.835 56.720 174.165 ;
        RECT 56.465 173.665 56.635 173.835 ;
        RECT 56.890 173.665 57.060 174.335 ;
        RECT 55.705 173.495 56.635 173.665 ;
        RECT 55.705 173.460 55.880 173.495 ;
        RECT 55.350 173.095 55.880 173.460 ;
        RECT 56.305 172.925 56.635 173.325 ;
        RECT 56.805 173.095 57.060 173.665 ;
        RECT 57.240 174.285 57.495 175.165 ;
        RECT 57.665 174.335 57.970 175.475 ;
        RECT 58.310 175.095 58.640 175.475 ;
        RECT 58.820 174.925 58.990 175.215 ;
        RECT 59.160 175.015 59.410 175.475 ;
        RECT 58.190 174.755 58.990 174.925 ;
        RECT 59.580 174.965 60.450 175.305 ;
        RECT 57.240 173.635 57.450 174.285 ;
        RECT 58.190 174.165 58.360 174.755 ;
        RECT 59.580 174.585 59.750 174.965 ;
        RECT 60.685 174.845 60.855 175.305 ;
        RECT 61.025 175.015 61.395 175.475 ;
        RECT 61.690 174.875 61.860 175.215 ;
        RECT 62.030 175.045 62.360 175.475 ;
        RECT 62.595 174.875 62.765 175.215 ;
        RECT 58.530 174.415 59.750 174.585 ;
        RECT 59.920 174.505 60.380 174.795 ;
        RECT 60.685 174.675 61.245 174.845 ;
        RECT 61.690 174.705 62.765 174.875 ;
        RECT 62.935 174.975 63.615 175.305 ;
        RECT 63.830 174.975 64.080 175.305 ;
        RECT 64.250 175.015 64.500 175.475 ;
        RECT 61.075 174.535 61.245 174.675 ;
        RECT 59.920 174.495 60.885 174.505 ;
        RECT 59.580 174.325 59.750 174.415 ;
        RECT 60.210 174.335 60.885 174.495 ;
        RECT 57.620 174.135 58.360 174.165 ;
        RECT 57.620 173.835 58.535 174.135 ;
        RECT 58.210 173.660 58.535 173.835 ;
        RECT 57.240 173.105 57.495 173.635 ;
        RECT 57.665 172.925 57.970 173.385 ;
        RECT 58.215 173.305 58.535 173.660 ;
        RECT 58.705 173.875 59.245 174.245 ;
        RECT 59.580 174.155 59.985 174.325 ;
        RECT 58.705 173.475 58.945 173.875 ;
        RECT 59.425 173.705 59.645 173.985 ;
        RECT 59.115 173.535 59.645 173.705 ;
        RECT 59.115 173.305 59.285 173.535 ;
        RECT 59.815 173.375 59.985 174.155 ;
        RECT 60.155 173.545 60.505 174.165 ;
        RECT 60.675 173.545 60.885 174.335 ;
        RECT 61.075 174.365 62.575 174.535 ;
        RECT 61.075 173.675 61.245 174.365 ;
        RECT 62.935 174.195 63.105 174.975 ;
        RECT 63.910 174.845 64.080 174.975 ;
        RECT 61.415 174.025 63.105 174.195 ;
        RECT 63.275 174.415 63.740 174.805 ;
        RECT 63.910 174.675 64.305 174.845 ;
        RECT 61.415 173.845 61.585 174.025 ;
        RECT 58.215 173.135 59.285 173.305 ;
        RECT 59.455 172.925 59.645 173.365 ;
        RECT 59.815 173.095 60.765 173.375 ;
        RECT 61.075 173.285 61.335 173.675 ;
        RECT 61.755 173.605 62.545 173.855 ;
        RECT 60.985 173.115 61.335 173.285 ;
        RECT 61.545 172.925 61.875 173.385 ;
        RECT 62.750 173.315 62.920 174.025 ;
        RECT 63.275 173.825 63.445 174.415 ;
        RECT 63.090 173.605 63.445 173.825 ;
        RECT 63.615 173.605 63.965 174.225 ;
        RECT 64.135 173.315 64.305 174.675 ;
        RECT 64.670 174.505 64.995 175.290 ;
        RECT 64.475 173.455 64.935 174.505 ;
        RECT 62.750 173.145 63.605 173.315 ;
        RECT 63.810 173.145 64.305 173.315 ;
        RECT 64.475 172.925 64.805 173.285 ;
        RECT 65.165 173.185 65.335 175.305 ;
        RECT 65.505 174.975 65.835 175.475 ;
        RECT 66.005 174.805 66.260 175.305 ;
        RECT 65.510 174.635 66.260 174.805 ;
        RECT 65.510 173.645 65.740 174.635 ;
        RECT 65.910 173.815 66.260 174.465 ;
        RECT 66.435 174.385 68.105 175.475 ;
        RECT 68.285 174.495 68.615 175.305 ;
        RECT 68.785 174.675 69.025 175.475 ;
        RECT 66.435 173.865 67.185 174.385 ;
        RECT 68.285 174.325 69.000 174.495 ;
        RECT 67.355 173.695 68.105 174.215 ;
        RECT 68.280 173.915 68.660 174.155 ;
        RECT 68.830 174.085 69.000 174.325 ;
        RECT 69.205 174.455 69.375 175.305 ;
        RECT 69.545 174.675 69.875 175.475 ;
        RECT 70.045 174.455 70.215 175.305 ;
        RECT 69.205 174.285 70.215 174.455 ;
        RECT 70.385 174.325 70.715 175.475 ;
        RECT 71.040 174.325 71.300 175.475 ;
        RECT 71.475 174.400 71.730 175.305 ;
        RECT 71.900 174.715 72.230 175.475 ;
        RECT 72.445 174.545 72.615 175.305 ;
        RECT 68.830 173.915 69.330 174.085 ;
        RECT 68.830 173.745 69.000 173.915 ;
        RECT 69.720 173.745 70.215 174.285 ;
        RECT 65.510 173.475 66.260 173.645 ;
        RECT 65.505 172.925 65.835 173.305 ;
        RECT 66.005 173.185 66.260 173.475 ;
        RECT 66.435 172.925 68.105 173.695 ;
        RECT 68.365 173.575 69.000 173.745 ;
        RECT 69.205 173.575 70.215 173.745 ;
        RECT 68.365 173.095 68.535 173.575 ;
        RECT 68.715 172.925 68.955 173.405 ;
        RECT 69.205 173.095 69.375 173.575 ;
        RECT 69.545 172.925 69.875 173.405 ;
        RECT 70.045 173.095 70.215 173.575 ;
        RECT 70.385 172.925 70.715 173.725 ;
        RECT 71.040 172.925 71.300 173.765 ;
        RECT 71.475 173.670 71.645 174.400 ;
        RECT 71.900 174.375 72.615 174.545 ;
        RECT 72.875 174.385 75.465 175.475 ;
        RECT 71.900 174.165 72.070 174.375 ;
        RECT 71.815 173.835 72.070 174.165 ;
        RECT 71.475 173.095 71.730 173.670 ;
        RECT 71.900 173.645 72.070 173.835 ;
        RECT 72.350 173.825 72.705 174.195 ;
        RECT 72.875 173.865 74.085 174.385 ;
        RECT 75.635 174.310 75.925 175.475 ;
        RECT 77.015 174.385 80.525 175.475 ;
        RECT 74.255 173.695 75.465 174.215 ;
        RECT 77.015 173.865 78.705 174.385 ;
        RECT 80.695 174.335 81.035 175.305 ;
        RECT 81.205 174.335 81.375 175.475 ;
        RECT 81.645 174.675 81.895 175.475 ;
        RECT 82.540 174.505 82.870 175.305 ;
        RECT 83.170 174.675 83.500 175.475 ;
        RECT 83.670 174.505 84.000 175.305 ;
        RECT 84.840 175.040 90.185 175.475 ;
        RECT 90.360 175.040 95.705 175.475 ;
        RECT 95.880 175.040 101.225 175.475 ;
        RECT 81.565 174.335 84.000 174.505 ;
        RECT 78.875 173.695 80.525 174.215 ;
        RECT 71.900 173.475 72.615 173.645 ;
        RECT 71.900 172.925 72.230 173.305 ;
        RECT 72.445 173.095 72.615 173.475 ;
        RECT 72.875 172.925 75.465 173.695 ;
        RECT 75.635 172.925 75.925 173.650 ;
        RECT 77.015 172.925 80.525 173.695 ;
        RECT 80.695 173.775 80.870 174.335 ;
        RECT 81.565 174.085 81.735 174.335 ;
        RECT 81.040 173.915 81.735 174.085 ;
        RECT 81.910 173.915 82.330 174.115 ;
        RECT 82.500 173.915 82.830 174.115 ;
        RECT 83.000 173.915 83.330 174.115 ;
        RECT 80.695 173.725 80.925 173.775 ;
        RECT 80.695 173.095 81.035 173.725 ;
        RECT 81.205 172.925 81.455 173.725 ;
        RECT 81.645 173.575 82.870 173.745 ;
        RECT 81.645 173.095 81.975 173.575 ;
        RECT 82.145 172.925 82.370 173.385 ;
        RECT 82.540 173.095 82.870 173.575 ;
        RECT 83.500 173.705 83.670 174.335 ;
        RECT 83.855 173.915 84.205 174.165 ;
        RECT 86.430 173.790 86.780 175.040 ;
        RECT 83.500 173.095 84.000 173.705 ;
        RECT 88.260 173.470 88.600 174.300 ;
        RECT 91.950 173.790 92.300 175.040 ;
        RECT 93.780 173.470 94.120 174.300 ;
        RECT 97.470 173.790 97.820 175.040 ;
        RECT 101.395 174.310 101.685 175.475 ;
        RECT 101.855 174.385 103.525 175.475 ;
        RECT 103.900 174.505 104.230 175.305 ;
        RECT 104.400 174.675 104.730 175.475 ;
        RECT 105.030 174.505 105.360 175.305 ;
        RECT 106.005 174.675 106.255 175.475 ;
        RECT 99.300 173.470 99.640 174.300 ;
        RECT 101.855 173.865 102.605 174.385 ;
        RECT 103.900 174.335 106.335 174.505 ;
        RECT 106.525 174.335 106.695 175.475 ;
        RECT 106.865 174.335 107.205 175.305 ;
        RECT 102.775 173.695 103.525 174.215 ;
        RECT 103.695 173.915 104.045 174.165 ;
        RECT 104.230 173.705 104.400 174.335 ;
        RECT 104.570 173.915 104.900 174.115 ;
        RECT 105.070 173.915 105.400 174.115 ;
        RECT 105.570 173.915 105.990 174.115 ;
        RECT 106.165 174.085 106.335 174.335 ;
        RECT 106.165 173.915 106.860 174.085 ;
        RECT 84.840 172.925 90.185 173.470 ;
        RECT 90.360 172.925 95.705 173.470 ;
        RECT 95.880 172.925 101.225 173.470 ;
        RECT 101.395 172.925 101.685 173.650 ;
        RECT 101.855 172.925 103.525 173.695 ;
        RECT 103.900 173.095 104.400 173.705 ;
        RECT 105.030 173.575 106.255 173.745 ;
        RECT 107.030 173.725 107.205 174.335 ;
        RECT 105.030 173.095 105.360 173.575 ;
        RECT 105.530 172.925 105.755 173.385 ;
        RECT 105.925 173.095 106.255 173.575 ;
        RECT 106.445 172.925 106.695 173.725 ;
        RECT 106.865 173.095 107.205 173.725 ;
        RECT 107.375 174.335 107.715 175.305 ;
        RECT 107.885 174.335 108.055 175.475 ;
        RECT 108.325 174.675 108.575 175.475 ;
        RECT 109.220 174.505 109.550 175.305 ;
        RECT 109.850 174.675 110.180 175.475 ;
        RECT 110.350 174.505 110.680 175.305 ;
        RECT 108.245 174.335 110.680 174.505 ;
        RECT 111.055 174.385 112.265 175.475 ;
        RECT 112.440 175.040 117.785 175.475 ;
        RECT 107.375 173.775 107.550 174.335 ;
        RECT 108.245 174.085 108.415 174.335 ;
        RECT 107.720 173.915 108.415 174.085 ;
        RECT 108.590 173.915 109.010 174.115 ;
        RECT 109.180 173.915 109.510 174.115 ;
        RECT 109.680 173.915 110.010 174.115 ;
        RECT 107.375 173.725 107.605 173.775 ;
        RECT 107.375 173.095 107.715 173.725 ;
        RECT 107.885 172.925 108.135 173.725 ;
        RECT 108.325 173.575 109.550 173.745 ;
        RECT 108.325 173.095 108.655 173.575 ;
        RECT 108.825 172.925 109.050 173.385 ;
        RECT 109.220 173.095 109.550 173.575 ;
        RECT 110.180 173.705 110.350 174.335 ;
        RECT 110.535 173.915 110.885 174.165 ;
        RECT 111.055 173.845 111.575 174.385 ;
        RECT 110.180 173.095 110.680 173.705 ;
        RECT 111.745 173.675 112.265 174.215 ;
        RECT 114.030 173.790 114.380 175.040 ;
        RECT 117.995 174.335 118.225 175.475 ;
        RECT 118.395 174.325 118.725 175.305 ;
        RECT 118.895 174.335 119.105 175.475 ;
        RECT 119.335 174.385 120.545 175.475 ;
        RECT 120.720 175.040 126.065 175.475 ;
        RECT 111.055 172.925 112.265 173.675 ;
        RECT 115.860 173.470 116.200 174.300 ;
        RECT 117.975 173.915 118.305 174.165 ;
        RECT 112.440 172.925 117.785 173.470 ;
        RECT 117.995 172.925 118.225 173.745 ;
        RECT 118.475 173.725 118.725 174.325 ;
        RECT 119.335 173.845 119.855 174.385 ;
        RECT 118.395 173.095 118.725 173.725 ;
        RECT 118.895 172.925 119.105 173.745 ;
        RECT 120.025 173.675 120.545 174.215 ;
        RECT 122.310 173.790 122.660 175.040 ;
        RECT 126.235 174.385 127.445 175.475 ;
        RECT 119.335 172.925 120.545 173.675 ;
        RECT 124.140 173.470 124.480 174.300 ;
        RECT 126.235 173.845 126.755 174.385 ;
        RECT 126.925 173.675 127.445 174.215 ;
        RECT 120.720 172.925 126.065 173.470 ;
        RECT 126.235 172.925 127.445 173.675 ;
        RECT 14.370 172.755 127.530 172.925 ;
        RECT 14.455 172.005 15.665 172.755 ;
        RECT 14.455 171.465 14.975 172.005 ;
        RECT 16.755 171.985 20.265 172.755 ;
        RECT 20.440 172.210 25.785 172.755 ;
        RECT 25.960 172.210 31.305 172.755 ;
        RECT 31.480 172.210 36.825 172.755 ;
        RECT 15.145 171.295 15.665 171.835 ;
        RECT 14.455 170.205 15.665 171.295 ;
        RECT 16.755 171.295 18.445 171.815 ;
        RECT 18.615 171.465 20.265 171.985 ;
        RECT 16.755 170.205 20.265 171.295 ;
        RECT 22.030 170.640 22.380 171.890 ;
        RECT 23.860 171.380 24.200 172.210 ;
        RECT 27.550 170.640 27.900 171.890 ;
        RECT 29.380 171.380 29.720 172.210 ;
        RECT 33.070 170.640 33.420 171.890 ;
        RECT 34.900 171.380 35.240 172.210 ;
        RECT 36.995 172.030 37.285 172.755 ;
        RECT 37.455 171.955 37.795 172.585 ;
        RECT 37.965 171.955 38.215 172.755 ;
        RECT 38.405 172.105 38.735 172.585 ;
        RECT 38.905 172.295 39.130 172.755 ;
        RECT 39.300 172.105 39.630 172.585 ;
        RECT 20.440 170.205 25.785 170.640 ;
        RECT 25.960 170.205 31.305 170.640 ;
        RECT 31.480 170.205 36.825 170.640 ;
        RECT 36.995 170.205 37.285 171.370 ;
        RECT 37.455 171.345 37.630 171.955 ;
        RECT 38.405 171.935 39.630 172.105 ;
        RECT 40.260 171.975 40.760 172.585 ;
        RECT 41.595 172.080 41.855 172.585 ;
        RECT 42.035 172.375 42.365 172.755 ;
        RECT 42.545 172.205 42.715 172.585 ;
        RECT 37.800 171.595 38.495 171.765 ;
        RECT 38.325 171.345 38.495 171.595 ;
        RECT 38.670 171.565 39.090 171.765 ;
        RECT 39.260 171.565 39.590 171.765 ;
        RECT 39.760 171.565 40.090 171.765 ;
        RECT 40.260 171.345 40.430 171.975 ;
        RECT 40.615 171.515 40.965 171.765 ;
        RECT 37.455 170.375 37.795 171.345 ;
        RECT 37.965 170.205 38.135 171.345 ;
        RECT 38.325 171.175 40.760 171.345 ;
        RECT 38.405 170.205 38.655 171.005 ;
        RECT 39.300 170.375 39.630 171.175 ;
        RECT 39.930 170.205 40.260 171.005 ;
        RECT 40.430 170.375 40.760 171.175 ;
        RECT 41.595 171.280 41.765 172.080 ;
        RECT 42.050 172.035 42.715 172.205 ;
        RECT 42.050 171.780 42.220 172.035 ;
        RECT 43.895 171.955 44.235 172.585 ;
        RECT 44.405 171.955 44.655 172.755 ;
        RECT 44.845 172.105 45.175 172.585 ;
        RECT 45.345 172.295 45.570 172.755 ;
        RECT 45.740 172.105 46.070 172.585 ;
        RECT 41.935 171.450 42.220 171.780 ;
        RECT 42.455 171.485 42.785 171.855 ;
        RECT 42.050 171.305 42.220 171.450 ;
        RECT 43.895 171.345 44.070 171.955 ;
        RECT 44.845 171.935 46.070 172.105 ;
        RECT 46.700 171.975 47.200 172.585 ;
        RECT 44.240 171.595 44.935 171.765 ;
        RECT 44.765 171.345 44.935 171.595 ;
        RECT 45.110 171.565 45.530 171.765 ;
        RECT 45.700 171.565 46.030 171.765 ;
        RECT 46.200 171.565 46.530 171.765 ;
        RECT 46.700 171.345 46.870 171.975 ;
        RECT 47.575 171.955 47.915 172.585 ;
        RECT 48.085 171.955 48.335 172.755 ;
        RECT 48.525 172.105 48.855 172.585 ;
        RECT 49.025 172.295 49.250 172.755 ;
        RECT 49.420 172.105 49.750 172.585 ;
        RECT 47.055 171.515 47.405 171.765 ;
        RECT 47.575 171.345 47.750 171.955 ;
        RECT 48.525 171.935 49.750 172.105 ;
        RECT 50.380 171.975 50.880 172.585 ;
        RECT 47.920 171.595 48.615 171.765 ;
        RECT 48.445 171.345 48.615 171.595 ;
        RECT 48.790 171.565 49.210 171.765 ;
        RECT 49.380 171.565 49.710 171.765 ;
        RECT 49.880 171.565 50.210 171.765 ;
        RECT 50.380 171.345 50.550 171.975 ;
        RECT 51.255 171.955 51.595 172.585 ;
        RECT 51.765 171.955 52.015 172.755 ;
        RECT 52.205 172.105 52.535 172.585 ;
        RECT 52.705 172.295 52.930 172.755 ;
        RECT 53.100 172.105 53.430 172.585 ;
        RECT 50.735 171.515 51.085 171.765 ;
        RECT 51.255 171.345 51.430 171.955 ;
        RECT 52.205 171.935 53.430 172.105 ;
        RECT 54.060 171.975 54.560 172.585 ;
        RECT 54.935 172.005 56.145 172.755 ;
        RECT 51.600 171.595 52.295 171.765 ;
        RECT 52.125 171.345 52.295 171.595 ;
        RECT 52.470 171.565 52.890 171.765 ;
        RECT 53.060 171.565 53.390 171.765 ;
        RECT 53.560 171.565 53.890 171.765 ;
        RECT 54.060 171.345 54.230 171.975 ;
        RECT 54.415 171.515 54.765 171.765 ;
        RECT 41.595 170.375 41.865 171.280 ;
        RECT 42.050 171.135 42.715 171.305 ;
        RECT 42.035 170.205 42.365 170.965 ;
        RECT 42.545 170.375 42.715 171.135 ;
        RECT 43.895 170.375 44.235 171.345 ;
        RECT 44.405 170.205 44.575 171.345 ;
        RECT 44.765 171.175 47.200 171.345 ;
        RECT 44.845 170.205 45.095 171.005 ;
        RECT 45.740 170.375 46.070 171.175 ;
        RECT 46.370 170.205 46.700 171.005 ;
        RECT 46.870 170.375 47.200 171.175 ;
        RECT 47.575 170.375 47.915 171.345 ;
        RECT 48.085 170.205 48.255 171.345 ;
        RECT 48.445 171.175 50.880 171.345 ;
        RECT 48.525 170.205 48.775 171.005 ;
        RECT 49.420 170.375 49.750 171.175 ;
        RECT 50.050 170.205 50.380 171.005 ;
        RECT 50.550 170.375 50.880 171.175 ;
        RECT 51.255 170.375 51.595 171.345 ;
        RECT 51.765 170.205 51.935 171.345 ;
        RECT 52.125 171.175 54.560 171.345 ;
        RECT 52.205 170.205 52.455 171.005 ;
        RECT 53.100 170.375 53.430 171.175 ;
        RECT 53.730 170.205 54.060 171.005 ;
        RECT 54.230 170.375 54.560 171.175 ;
        RECT 54.935 171.295 55.455 171.835 ;
        RECT 55.625 171.465 56.145 172.005 ;
        RECT 56.315 171.985 59.825 172.755 ;
        RECT 56.315 171.295 58.005 171.815 ;
        RECT 58.175 171.465 59.825 171.985 ;
        RECT 60.055 171.935 60.265 172.755 ;
        RECT 60.435 171.955 60.765 172.585 ;
        RECT 60.435 171.355 60.685 171.955 ;
        RECT 60.935 171.935 61.165 172.755 ;
        RECT 61.465 172.205 61.635 172.585 ;
        RECT 61.815 172.375 62.145 172.755 ;
        RECT 61.465 172.035 62.130 172.205 ;
        RECT 62.325 172.080 62.585 172.585 ;
        RECT 60.855 171.515 61.185 171.765 ;
        RECT 61.395 171.485 61.725 171.855 ;
        RECT 61.960 171.780 62.130 172.035 ;
        RECT 61.960 171.450 62.245 171.780 ;
        RECT 54.935 170.205 56.145 171.295 ;
        RECT 56.315 170.205 59.825 171.295 ;
        RECT 60.055 170.205 60.265 171.345 ;
        RECT 60.435 170.375 60.765 171.355 ;
        RECT 60.935 170.205 61.165 171.345 ;
        RECT 61.960 171.305 62.130 171.450 ;
        RECT 61.465 171.135 62.130 171.305 ;
        RECT 62.415 171.280 62.585 172.080 ;
        RECT 62.755 172.030 63.045 172.755 ;
        RECT 63.675 171.985 65.345 172.755 ;
        RECT 65.520 172.210 70.865 172.755 ;
        RECT 71.040 172.210 76.385 172.755 ;
        RECT 76.560 172.210 81.905 172.755 ;
        RECT 61.465 170.375 61.635 171.135 ;
        RECT 61.815 170.205 62.145 170.965 ;
        RECT 62.315 170.375 62.585 171.280 ;
        RECT 62.755 170.205 63.045 171.370 ;
        RECT 63.675 171.295 64.425 171.815 ;
        RECT 64.595 171.465 65.345 171.985 ;
        RECT 63.675 170.205 65.345 171.295 ;
        RECT 67.110 170.640 67.460 171.890 ;
        RECT 68.940 171.380 69.280 172.210 ;
        RECT 72.630 170.640 72.980 171.890 ;
        RECT 74.460 171.380 74.800 172.210 ;
        RECT 78.150 170.640 78.500 171.890 ;
        RECT 79.980 171.380 80.320 172.210 ;
        RECT 82.165 172.105 82.335 172.585 ;
        RECT 82.515 172.275 82.755 172.755 ;
        RECT 83.005 172.105 83.175 172.585 ;
        RECT 83.345 172.275 83.675 172.755 ;
        RECT 83.845 172.105 84.015 172.585 ;
        RECT 82.165 171.935 82.800 172.105 ;
        RECT 83.005 171.935 84.015 172.105 ;
        RECT 84.185 171.955 84.515 172.755 ;
        RECT 84.950 172.125 85.235 172.585 ;
        RECT 85.405 172.295 85.675 172.755 ;
        RECT 84.950 171.955 85.905 172.125 ;
        RECT 82.630 171.765 82.800 171.935 ;
        RECT 83.515 171.905 84.015 171.935 ;
        RECT 82.080 171.525 82.460 171.765 ;
        RECT 82.630 171.595 83.130 171.765 ;
        RECT 82.630 171.355 82.800 171.595 ;
        RECT 83.520 171.395 84.015 171.905 ;
        RECT 82.085 171.185 82.800 171.355 ;
        RECT 83.005 171.225 84.015 171.395 ;
        RECT 65.520 170.205 70.865 170.640 ;
        RECT 71.040 170.205 76.385 170.640 ;
        RECT 76.560 170.205 81.905 170.640 ;
        RECT 82.085 170.375 82.415 171.185 ;
        RECT 82.585 170.205 82.825 171.005 ;
        RECT 83.005 170.375 83.175 171.225 ;
        RECT 83.345 170.205 83.675 171.005 ;
        RECT 83.845 170.375 84.015 171.225 ;
        RECT 84.185 170.205 84.515 171.355 ;
        RECT 84.835 171.225 85.525 171.785 ;
        RECT 85.695 171.055 85.905 171.955 ;
        RECT 84.950 170.835 85.905 171.055 ;
        RECT 86.075 171.785 86.475 172.585 ;
        RECT 86.665 172.125 86.945 172.585 ;
        RECT 87.465 172.295 87.790 172.755 ;
        RECT 86.665 171.955 87.790 172.125 ;
        RECT 87.960 172.015 88.345 172.585 ;
        RECT 88.515 172.030 88.805 172.755 ;
        RECT 87.340 171.845 87.790 171.955 ;
        RECT 86.075 171.225 87.170 171.785 ;
        RECT 87.340 171.515 87.895 171.845 ;
        RECT 84.950 170.375 85.235 170.835 ;
        RECT 85.405 170.205 85.675 170.665 ;
        RECT 86.075 170.375 86.475 171.225 ;
        RECT 87.340 171.055 87.790 171.515 ;
        RECT 88.065 171.345 88.345 172.015 ;
        RECT 89.475 171.935 89.705 172.755 ;
        RECT 89.875 171.955 90.205 172.585 ;
        RECT 89.455 171.515 89.785 171.765 ;
        RECT 86.665 170.835 87.790 171.055 ;
        RECT 86.665 170.375 86.945 170.835 ;
        RECT 87.465 170.205 87.790 170.665 ;
        RECT 87.960 170.375 88.345 171.345 ;
        RECT 88.515 170.205 88.805 171.370 ;
        RECT 89.955 171.355 90.205 171.955 ;
        RECT 90.375 171.935 90.585 172.755 ;
        RECT 90.820 172.045 91.075 172.575 ;
        RECT 91.245 172.295 91.550 172.755 ;
        RECT 91.795 172.375 92.865 172.545 ;
        RECT 89.475 170.205 89.705 171.345 ;
        RECT 89.875 170.375 90.205 171.355 ;
        RECT 90.820 171.395 91.030 172.045 ;
        RECT 91.795 172.020 92.115 172.375 ;
        RECT 91.790 171.845 92.115 172.020 ;
        RECT 91.200 171.545 92.115 171.845 ;
        RECT 92.285 171.805 92.525 172.205 ;
        RECT 92.695 172.145 92.865 172.375 ;
        RECT 93.035 172.315 93.225 172.755 ;
        RECT 93.395 172.305 94.345 172.585 ;
        RECT 94.565 172.395 94.915 172.565 ;
        RECT 92.695 171.975 93.225 172.145 ;
        RECT 91.200 171.515 91.940 171.545 ;
        RECT 90.375 170.205 90.585 171.345 ;
        RECT 90.820 170.515 91.075 171.395 ;
        RECT 91.245 170.205 91.550 171.345 ;
        RECT 91.770 170.925 91.940 171.515 ;
        RECT 92.285 171.435 92.825 171.805 ;
        RECT 93.005 171.695 93.225 171.975 ;
        RECT 93.395 171.525 93.565 172.305 ;
        RECT 93.160 171.355 93.565 171.525 ;
        RECT 93.735 171.515 94.085 172.135 ;
        RECT 93.160 171.265 93.330 171.355 ;
        RECT 94.255 171.345 94.465 172.135 ;
        RECT 92.110 171.095 93.330 171.265 ;
        RECT 93.790 171.185 94.465 171.345 ;
        RECT 91.770 170.755 92.570 170.925 ;
        RECT 91.890 170.205 92.220 170.585 ;
        RECT 92.400 170.465 92.570 170.755 ;
        RECT 93.160 170.715 93.330 171.095 ;
        RECT 93.500 171.175 94.465 171.185 ;
        RECT 94.655 172.005 94.915 172.395 ;
        RECT 95.125 172.295 95.455 172.755 ;
        RECT 96.330 172.365 97.185 172.535 ;
        RECT 97.390 172.365 97.885 172.535 ;
        RECT 98.055 172.395 98.385 172.755 ;
        RECT 94.655 171.315 94.825 172.005 ;
        RECT 94.995 171.655 95.165 171.835 ;
        RECT 95.335 171.825 96.125 172.075 ;
        RECT 96.330 171.655 96.500 172.365 ;
        RECT 96.670 171.855 97.025 172.075 ;
        RECT 94.995 171.485 96.685 171.655 ;
        RECT 93.500 170.885 93.960 171.175 ;
        RECT 94.655 171.145 96.155 171.315 ;
        RECT 94.655 171.005 94.825 171.145 ;
        RECT 94.265 170.835 94.825 171.005 ;
        RECT 92.740 170.205 92.990 170.665 ;
        RECT 93.160 170.375 94.030 170.715 ;
        RECT 94.265 170.375 94.435 170.835 ;
        RECT 95.270 170.805 96.345 170.975 ;
        RECT 94.605 170.205 94.975 170.665 ;
        RECT 95.270 170.465 95.440 170.805 ;
        RECT 95.610 170.205 95.940 170.635 ;
        RECT 96.175 170.465 96.345 170.805 ;
        RECT 96.515 170.705 96.685 171.485 ;
        RECT 96.855 171.265 97.025 171.855 ;
        RECT 97.195 171.455 97.545 172.075 ;
        RECT 96.855 170.875 97.320 171.265 ;
        RECT 97.715 171.005 97.885 172.365 ;
        RECT 98.055 171.175 98.515 172.225 ;
        RECT 97.490 170.835 97.885 171.005 ;
        RECT 97.490 170.705 97.660 170.835 ;
        RECT 96.515 170.375 97.195 170.705 ;
        RECT 97.410 170.375 97.660 170.705 ;
        RECT 97.830 170.205 98.080 170.665 ;
        RECT 98.250 170.390 98.575 171.175 ;
        RECT 98.745 170.375 98.915 172.495 ;
        RECT 99.085 172.375 99.415 172.755 ;
        RECT 99.585 172.205 99.840 172.495 ;
        RECT 100.940 172.210 106.285 172.755 ;
        RECT 99.090 172.035 99.840 172.205 ;
        RECT 99.090 171.045 99.320 172.035 ;
        RECT 99.490 171.215 99.840 171.865 ;
        RECT 99.090 170.875 99.840 171.045 ;
        RECT 99.085 170.205 99.415 170.705 ;
        RECT 99.585 170.375 99.840 170.875 ;
        RECT 102.530 170.640 102.880 171.890 ;
        RECT 104.360 171.380 104.700 172.210 ;
        RECT 106.515 171.935 106.725 172.755 ;
        RECT 106.895 171.955 107.225 172.585 ;
        RECT 106.895 171.355 107.145 171.955 ;
        RECT 107.395 171.935 107.625 172.755 ;
        RECT 108.040 171.975 108.540 172.585 ;
        RECT 107.315 171.515 107.645 171.765 ;
        RECT 107.835 171.515 108.185 171.765 ;
        RECT 100.940 170.205 106.285 170.640 ;
        RECT 106.515 170.205 106.725 171.345 ;
        RECT 106.895 170.375 107.225 171.355 ;
        RECT 108.370 171.345 108.540 171.975 ;
        RECT 109.170 172.105 109.500 172.585 ;
        RECT 109.670 172.295 109.895 172.755 ;
        RECT 110.065 172.105 110.395 172.585 ;
        RECT 109.170 171.935 110.395 172.105 ;
        RECT 110.585 171.955 110.835 172.755 ;
        RECT 111.005 171.955 111.345 172.585 ;
        RECT 111.515 172.005 112.725 172.755 ;
        RECT 108.710 171.565 109.040 171.765 ;
        RECT 109.210 171.565 109.540 171.765 ;
        RECT 109.710 171.565 110.130 171.765 ;
        RECT 110.305 171.595 111.000 171.765 ;
        RECT 110.305 171.345 110.475 171.595 ;
        RECT 111.170 171.345 111.345 171.955 ;
        RECT 107.395 170.205 107.625 171.345 ;
        RECT 108.040 171.175 110.475 171.345 ;
        RECT 108.040 170.375 108.370 171.175 ;
        RECT 108.540 170.205 108.870 171.005 ;
        RECT 109.170 170.375 109.500 171.175 ;
        RECT 110.145 170.205 110.395 171.005 ;
        RECT 110.665 170.205 110.835 171.345 ;
        RECT 111.005 170.375 111.345 171.345 ;
        RECT 111.515 171.295 112.035 171.835 ;
        RECT 112.205 171.465 112.725 172.005 ;
        RECT 112.935 171.935 113.165 172.755 ;
        RECT 113.335 171.955 113.665 172.585 ;
        RECT 112.915 171.515 113.245 171.765 ;
        RECT 113.415 171.355 113.665 171.955 ;
        RECT 113.835 171.935 114.045 172.755 ;
        RECT 114.275 172.030 114.565 172.755 ;
        RECT 115.660 172.045 115.915 172.575 ;
        RECT 116.085 172.295 116.390 172.755 ;
        RECT 116.635 172.375 117.705 172.545 ;
        RECT 115.660 171.395 115.870 172.045 ;
        RECT 116.635 172.020 116.955 172.375 ;
        RECT 116.630 171.845 116.955 172.020 ;
        RECT 116.040 171.545 116.955 171.845 ;
        RECT 117.125 171.805 117.365 172.205 ;
        RECT 117.535 172.145 117.705 172.375 ;
        RECT 117.875 172.315 118.065 172.755 ;
        RECT 118.235 172.305 119.185 172.585 ;
        RECT 119.405 172.395 119.755 172.565 ;
        RECT 117.535 171.975 118.065 172.145 ;
        RECT 116.040 171.515 116.780 171.545 ;
        RECT 111.515 170.205 112.725 171.295 ;
        RECT 112.935 170.205 113.165 171.345 ;
        RECT 113.335 170.375 113.665 171.355 ;
        RECT 113.835 170.205 114.045 171.345 ;
        RECT 114.275 170.205 114.565 171.370 ;
        RECT 115.660 170.515 115.915 171.395 ;
        RECT 116.085 170.205 116.390 171.345 ;
        RECT 116.610 170.925 116.780 171.515 ;
        RECT 117.125 171.435 117.665 171.805 ;
        RECT 117.845 171.695 118.065 171.975 ;
        RECT 118.235 171.525 118.405 172.305 ;
        RECT 118.000 171.355 118.405 171.525 ;
        RECT 118.575 171.515 118.925 172.135 ;
        RECT 118.000 171.265 118.170 171.355 ;
        RECT 119.095 171.345 119.305 172.135 ;
        RECT 116.950 171.095 118.170 171.265 ;
        RECT 118.630 171.185 119.305 171.345 ;
        RECT 116.610 170.755 117.410 170.925 ;
        RECT 116.730 170.205 117.060 170.585 ;
        RECT 117.240 170.465 117.410 170.755 ;
        RECT 118.000 170.715 118.170 171.095 ;
        RECT 118.340 171.175 119.305 171.185 ;
        RECT 119.495 172.005 119.755 172.395 ;
        RECT 119.965 172.295 120.295 172.755 ;
        RECT 121.170 172.365 122.025 172.535 ;
        RECT 122.230 172.365 122.725 172.535 ;
        RECT 122.895 172.395 123.225 172.755 ;
        RECT 119.495 171.315 119.665 172.005 ;
        RECT 119.835 171.655 120.005 171.835 ;
        RECT 120.175 171.825 120.965 172.075 ;
        RECT 121.170 171.655 121.340 172.365 ;
        RECT 121.510 171.855 121.865 172.075 ;
        RECT 119.835 171.485 121.525 171.655 ;
        RECT 118.340 170.885 118.800 171.175 ;
        RECT 119.495 171.145 120.995 171.315 ;
        RECT 119.495 171.005 119.665 171.145 ;
        RECT 119.105 170.835 119.665 171.005 ;
        RECT 117.580 170.205 117.830 170.665 ;
        RECT 118.000 170.375 118.870 170.715 ;
        RECT 119.105 170.375 119.275 170.835 ;
        RECT 120.110 170.805 121.185 170.975 ;
        RECT 119.445 170.205 119.815 170.665 ;
        RECT 120.110 170.465 120.280 170.805 ;
        RECT 120.450 170.205 120.780 170.635 ;
        RECT 121.015 170.465 121.185 170.805 ;
        RECT 121.355 170.705 121.525 171.485 ;
        RECT 121.695 171.265 121.865 171.855 ;
        RECT 122.035 171.455 122.385 172.075 ;
        RECT 121.695 170.875 122.160 171.265 ;
        RECT 122.555 171.005 122.725 172.365 ;
        RECT 122.895 171.175 123.355 172.225 ;
        RECT 122.330 170.835 122.725 171.005 ;
        RECT 122.330 170.705 122.500 170.835 ;
        RECT 121.355 170.375 122.035 170.705 ;
        RECT 122.250 170.375 122.500 170.705 ;
        RECT 122.670 170.205 122.920 170.665 ;
        RECT 123.090 170.390 123.415 171.175 ;
        RECT 123.585 170.375 123.755 172.495 ;
        RECT 123.925 172.375 124.255 172.755 ;
        RECT 124.425 172.205 124.680 172.495 ;
        RECT 123.930 172.035 124.680 172.205 ;
        RECT 123.930 171.045 124.160 172.035 ;
        RECT 124.855 172.005 126.065 172.755 ;
        RECT 126.235 172.005 127.445 172.755 ;
        RECT 124.330 171.215 124.680 171.865 ;
        RECT 124.855 171.295 125.375 171.835 ;
        RECT 125.545 171.465 126.065 172.005 ;
        RECT 126.235 171.295 126.755 171.835 ;
        RECT 126.925 171.465 127.445 172.005 ;
        RECT 123.930 170.875 124.680 171.045 ;
        RECT 123.925 170.205 124.255 170.705 ;
        RECT 124.425 170.375 124.680 170.875 ;
        RECT 124.855 170.205 126.065 171.295 ;
        RECT 126.235 170.205 127.445 171.295 ;
        RECT 14.370 170.035 127.530 170.205 ;
        RECT 14.455 168.945 15.665 170.035 ;
        RECT 14.455 168.235 14.975 168.775 ;
        RECT 15.145 168.405 15.665 168.945 ;
        RECT 15.835 168.945 18.425 170.035 ;
        RECT 18.600 169.600 23.945 170.035 ;
        RECT 15.835 168.425 17.045 168.945 ;
        RECT 17.215 168.255 18.425 168.775 ;
        RECT 20.190 168.350 20.540 169.600 ;
        RECT 24.115 168.870 24.405 170.035 ;
        RECT 25.035 168.945 26.705 170.035 ;
        RECT 14.455 167.485 15.665 168.235 ;
        RECT 15.835 167.485 18.425 168.255 ;
        RECT 22.020 168.030 22.360 168.860 ;
        RECT 25.035 168.425 25.785 168.945 ;
        RECT 26.915 168.895 27.145 170.035 ;
        RECT 27.315 168.885 27.645 169.865 ;
        RECT 27.815 168.895 28.025 170.035 ;
        RECT 28.715 168.945 32.225 170.035 ;
        RECT 25.955 168.255 26.705 168.775 ;
        RECT 26.895 168.475 27.225 168.725 ;
        RECT 18.600 167.485 23.945 168.030 ;
        RECT 24.115 167.485 24.405 168.210 ;
        RECT 25.035 167.485 26.705 168.255 ;
        RECT 26.915 167.485 27.145 168.305 ;
        RECT 27.395 168.285 27.645 168.885 ;
        RECT 28.715 168.425 30.405 168.945 ;
        RECT 32.455 168.895 32.665 170.035 ;
        RECT 32.835 168.885 33.165 169.865 ;
        RECT 33.335 168.895 33.565 170.035 ;
        RECT 33.775 168.945 34.985 170.035 ;
        RECT 35.245 169.290 35.515 170.035 ;
        RECT 36.145 170.030 42.420 170.035 ;
        RECT 35.685 169.120 35.975 169.860 ;
        RECT 36.145 169.305 36.400 170.030 ;
        RECT 36.585 169.135 36.845 169.860 ;
        RECT 37.015 169.305 37.260 170.030 ;
        RECT 37.445 169.135 37.705 169.860 ;
        RECT 37.875 169.305 38.120 170.030 ;
        RECT 38.305 169.135 38.565 169.860 ;
        RECT 38.735 169.305 38.980 170.030 ;
        RECT 39.150 169.135 39.410 169.860 ;
        RECT 39.580 169.305 39.840 170.030 ;
        RECT 40.010 169.135 40.270 169.860 ;
        RECT 40.440 169.305 40.700 170.030 ;
        RECT 40.870 169.135 41.130 169.860 ;
        RECT 41.300 169.305 41.560 170.030 ;
        RECT 41.730 169.135 41.990 169.860 ;
        RECT 42.160 169.235 42.420 170.030 ;
        RECT 36.585 169.120 41.990 169.135 ;
        RECT 27.315 167.655 27.645 168.285 ;
        RECT 27.815 167.485 28.025 168.305 ;
        RECT 30.575 168.255 32.225 168.775 ;
        RECT 28.715 167.485 32.225 168.255 ;
        RECT 32.455 167.485 32.665 168.305 ;
        RECT 32.835 168.285 33.085 168.885 ;
        RECT 33.255 168.475 33.585 168.725 ;
        RECT 33.775 168.405 34.295 168.945 ;
        RECT 35.245 168.895 41.990 169.120 ;
        RECT 32.835 167.655 33.165 168.285 ;
        RECT 33.335 167.485 33.565 168.305 ;
        RECT 34.465 168.235 34.985 168.775 ;
        RECT 33.775 167.485 34.985 168.235 ;
        RECT 35.245 168.305 36.410 168.895 ;
        RECT 42.590 168.725 42.840 169.860 ;
        RECT 43.020 169.225 43.280 170.035 ;
        RECT 43.455 168.725 43.700 169.865 ;
        RECT 43.880 169.225 44.175 170.035 ;
        RECT 44.360 169.600 49.705 170.035 ;
        RECT 36.580 168.475 43.700 168.725 ;
        RECT 35.245 168.135 41.990 168.305 ;
        RECT 35.245 167.485 35.545 167.965 ;
        RECT 35.715 167.680 35.975 168.135 ;
        RECT 36.145 167.485 36.405 167.965 ;
        RECT 36.585 167.680 36.845 168.135 ;
        RECT 37.015 167.485 37.265 167.965 ;
        RECT 37.445 167.680 37.705 168.135 ;
        RECT 37.875 167.485 38.125 167.965 ;
        RECT 38.305 167.680 38.565 168.135 ;
        RECT 38.735 167.485 38.980 167.965 ;
        RECT 39.150 167.680 39.425 168.135 ;
        RECT 39.595 167.485 39.840 167.965 ;
        RECT 40.010 167.680 40.270 168.135 ;
        RECT 40.440 167.485 40.700 167.965 ;
        RECT 40.870 167.680 41.130 168.135 ;
        RECT 41.300 167.485 41.560 167.965 ;
        RECT 41.730 167.680 41.990 168.135 ;
        RECT 42.160 167.485 42.420 168.045 ;
        RECT 42.590 167.665 42.840 168.475 ;
        RECT 43.020 167.485 43.280 168.010 ;
        RECT 43.450 167.665 43.700 168.475 ;
        RECT 43.870 168.165 44.185 168.725 ;
        RECT 45.950 168.350 46.300 169.600 ;
        RECT 49.875 168.870 50.165 170.035 ;
        RECT 50.335 168.945 51.545 170.035 ;
        RECT 51.720 169.600 57.065 170.035 ;
        RECT 57.240 169.600 62.585 170.035 ;
        RECT 62.760 169.600 68.105 170.035 ;
        RECT 47.780 168.030 48.120 168.860 ;
        RECT 50.335 168.405 50.855 168.945 ;
        RECT 51.025 168.235 51.545 168.775 ;
        RECT 53.310 168.350 53.660 169.600 ;
        RECT 43.880 167.485 44.185 167.995 ;
        RECT 44.360 167.485 49.705 168.030 ;
        RECT 49.875 167.485 50.165 168.210 ;
        RECT 50.335 167.485 51.545 168.235 ;
        RECT 55.140 168.030 55.480 168.860 ;
        RECT 58.830 168.350 59.180 169.600 ;
        RECT 60.660 168.030 61.000 168.860 ;
        RECT 64.350 168.350 64.700 169.600 ;
        RECT 68.280 168.885 68.540 170.035 ;
        RECT 68.715 168.960 68.970 169.865 ;
        RECT 69.140 169.275 69.470 170.035 ;
        RECT 69.685 169.105 69.855 169.865 ;
        RECT 66.180 168.030 66.520 168.860 ;
        RECT 51.720 167.485 57.065 168.030 ;
        RECT 57.240 167.485 62.585 168.030 ;
        RECT 62.760 167.485 68.105 168.030 ;
        RECT 68.280 167.485 68.540 168.325 ;
        RECT 68.715 168.230 68.885 168.960 ;
        RECT 69.140 168.935 69.855 169.105 ;
        RECT 69.140 168.725 69.310 168.935 ;
        RECT 70.120 168.885 70.380 170.035 ;
        RECT 70.555 168.960 70.810 169.865 ;
        RECT 70.980 169.275 71.310 170.035 ;
        RECT 71.525 169.105 71.695 169.865 ;
        RECT 69.055 168.395 69.310 168.725 ;
        RECT 68.715 167.655 68.970 168.230 ;
        RECT 69.140 168.205 69.310 168.395 ;
        RECT 69.590 168.385 69.945 168.755 ;
        RECT 69.140 168.035 69.855 168.205 ;
        RECT 69.140 167.485 69.470 167.865 ;
        RECT 69.685 167.655 69.855 168.035 ;
        RECT 70.120 167.485 70.380 168.325 ;
        RECT 70.555 168.230 70.725 168.960 ;
        RECT 70.980 168.935 71.695 169.105 ;
        RECT 71.955 168.945 75.465 170.035 ;
        RECT 70.980 168.725 71.150 168.935 ;
        RECT 70.895 168.395 71.150 168.725 ;
        RECT 70.555 167.655 70.810 168.230 ;
        RECT 70.980 168.205 71.150 168.395 ;
        RECT 71.430 168.385 71.785 168.755 ;
        RECT 71.955 168.425 73.645 168.945 ;
        RECT 75.635 168.870 75.925 170.035 ;
        RECT 76.095 169.275 76.610 169.685 ;
        RECT 76.845 169.275 77.015 170.035 ;
        RECT 77.185 169.695 79.215 169.865 ;
        RECT 73.815 168.255 75.465 168.775 ;
        RECT 76.095 168.465 76.435 169.275 ;
        RECT 77.185 169.030 77.355 169.695 ;
        RECT 77.750 169.355 78.875 169.525 ;
        RECT 76.605 168.840 77.355 169.030 ;
        RECT 77.525 169.015 78.535 169.185 ;
        RECT 76.095 168.295 77.325 168.465 ;
        RECT 70.980 168.035 71.695 168.205 ;
        RECT 70.980 167.485 71.310 167.865 ;
        RECT 71.525 167.655 71.695 168.035 ;
        RECT 71.955 167.485 75.465 168.255 ;
        RECT 75.635 167.485 75.925 168.210 ;
        RECT 76.370 167.690 76.615 168.295 ;
        RECT 76.835 167.485 77.345 168.020 ;
        RECT 77.525 167.655 77.715 169.015 ;
        RECT 77.885 167.995 78.160 168.815 ;
        RECT 78.365 168.215 78.535 169.015 ;
        RECT 78.705 168.225 78.875 169.355 ;
        RECT 79.045 168.725 79.215 169.695 ;
        RECT 79.385 168.895 79.555 170.035 ;
        RECT 79.725 168.895 80.060 169.865 ;
        RECT 79.045 168.395 79.240 168.725 ;
        RECT 79.465 168.395 79.720 168.725 ;
        RECT 79.465 168.225 79.635 168.395 ;
        RECT 79.890 168.225 80.060 168.895 ;
        RECT 80.610 169.055 80.865 169.725 ;
        RECT 81.045 169.235 81.330 170.035 ;
        RECT 81.510 169.315 81.840 169.825 ;
        RECT 80.610 168.335 80.790 169.055 ;
        RECT 81.510 168.725 81.760 169.315 ;
        RECT 82.110 169.165 82.280 169.775 ;
        RECT 82.450 169.345 82.780 170.035 ;
        RECT 83.010 169.485 83.250 169.775 ;
        RECT 83.450 169.655 83.870 170.035 ;
        RECT 84.050 169.565 84.680 169.815 ;
        RECT 85.150 169.655 85.480 170.035 ;
        RECT 84.050 169.485 84.220 169.565 ;
        RECT 85.650 169.485 85.820 169.775 ;
        RECT 86.000 169.655 86.380 170.035 ;
        RECT 86.620 169.650 87.450 169.820 ;
        RECT 83.010 169.315 84.220 169.485 ;
        RECT 80.960 168.395 81.760 168.725 ;
        RECT 78.705 168.055 79.635 168.225 ;
        RECT 78.705 168.020 78.880 168.055 ;
        RECT 77.885 167.825 78.165 167.995 ;
        RECT 77.885 167.655 78.160 167.825 ;
        RECT 78.350 167.655 78.880 168.020 ;
        RECT 79.305 167.485 79.635 167.885 ;
        RECT 79.805 167.655 80.060 168.225 ;
        RECT 80.525 168.195 80.790 168.335 ;
        RECT 80.525 168.165 80.865 168.195 ;
        RECT 80.610 167.665 80.865 168.165 ;
        RECT 81.045 167.485 81.330 167.945 ;
        RECT 81.510 167.745 81.760 168.395 ;
        RECT 81.960 169.145 82.280 169.165 ;
        RECT 81.960 168.975 83.880 169.145 ;
        RECT 81.960 168.080 82.150 168.975 ;
        RECT 84.050 168.805 84.220 169.315 ;
        RECT 84.390 169.055 84.910 169.365 ;
        RECT 82.320 168.635 84.220 168.805 ;
        RECT 82.320 168.575 82.650 168.635 ;
        RECT 82.800 168.405 83.130 168.465 ;
        RECT 82.470 168.135 83.130 168.405 ;
        RECT 81.960 167.750 82.280 168.080 ;
        RECT 82.460 167.485 83.120 167.965 ;
        RECT 83.320 167.875 83.490 168.635 ;
        RECT 84.390 168.465 84.570 168.875 ;
        RECT 83.660 168.295 83.990 168.415 ;
        RECT 84.740 168.295 84.910 169.055 ;
        RECT 83.660 168.125 84.910 168.295 ;
        RECT 85.080 169.235 86.450 169.485 ;
        RECT 85.080 168.465 85.270 169.235 ;
        RECT 86.200 168.975 86.450 169.235 ;
        RECT 85.440 168.805 85.690 168.965 ;
        RECT 86.620 168.805 86.790 169.650 ;
        RECT 87.685 169.365 87.855 169.865 ;
        RECT 88.025 169.535 88.355 170.035 ;
        RECT 86.960 168.975 87.460 169.355 ;
        RECT 87.685 169.195 88.380 169.365 ;
        RECT 85.440 168.635 86.790 168.805 ;
        RECT 86.370 168.595 86.790 168.635 ;
        RECT 85.080 168.125 85.500 168.465 ;
        RECT 85.790 168.135 86.200 168.465 ;
        RECT 83.320 167.705 84.170 167.875 ;
        RECT 84.730 167.485 85.050 167.945 ;
        RECT 85.250 167.695 85.500 168.125 ;
        RECT 85.790 167.485 86.200 167.925 ;
        RECT 86.370 167.865 86.540 168.595 ;
        RECT 86.710 168.045 87.060 168.415 ;
        RECT 87.240 168.105 87.460 168.975 ;
        RECT 87.630 168.405 88.040 169.025 ;
        RECT 88.210 168.225 88.380 169.195 ;
        RECT 87.685 168.035 88.380 168.225 ;
        RECT 86.370 167.665 87.385 167.865 ;
        RECT 87.685 167.705 87.855 168.035 ;
        RECT 88.025 167.485 88.355 167.865 ;
        RECT 88.570 167.745 88.795 169.865 ;
        RECT 88.965 169.535 89.295 170.035 ;
        RECT 89.465 169.365 89.635 169.865 ;
        RECT 88.970 169.195 89.635 169.365 ;
        RECT 88.970 168.205 89.200 169.195 ;
        RECT 89.370 168.375 89.720 169.025 ;
        RECT 89.895 168.945 91.105 170.035 ;
        RECT 91.275 169.275 91.790 169.685 ;
        RECT 92.025 169.275 92.195 170.035 ;
        RECT 92.365 169.695 94.395 169.865 ;
        RECT 89.895 168.405 90.415 168.945 ;
        RECT 90.585 168.235 91.105 168.775 ;
        RECT 91.275 168.465 91.615 169.275 ;
        RECT 92.365 169.030 92.535 169.695 ;
        RECT 92.930 169.355 94.055 169.525 ;
        RECT 91.785 168.840 92.535 169.030 ;
        RECT 92.705 169.015 93.715 169.185 ;
        RECT 91.275 168.295 92.505 168.465 ;
        RECT 88.970 168.035 89.635 168.205 ;
        RECT 88.965 167.485 89.295 167.865 ;
        RECT 89.465 167.745 89.635 168.035 ;
        RECT 89.895 167.485 91.105 168.235 ;
        RECT 91.550 167.690 91.795 168.295 ;
        RECT 92.015 167.485 92.525 168.020 ;
        RECT 92.705 167.655 92.895 169.015 ;
        RECT 93.065 168.675 93.340 168.815 ;
        RECT 93.065 168.505 93.345 168.675 ;
        RECT 93.065 167.655 93.340 168.505 ;
        RECT 93.545 168.215 93.715 169.015 ;
        RECT 93.885 168.225 94.055 169.355 ;
        RECT 94.225 168.725 94.395 169.695 ;
        RECT 94.565 168.895 94.735 170.035 ;
        RECT 94.905 168.895 95.240 169.865 ;
        RECT 95.965 169.105 96.135 169.865 ;
        RECT 96.315 169.275 96.645 170.035 ;
        RECT 95.965 168.935 96.630 169.105 ;
        RECT 96.815 168.960 97.085 169.865 ;
        RECT 94.225 168.395 94.420 168.725 ;
        RECT 94.645 168.395 94.900 168.725 ;
        RECT 94.645 168.225 94.815 168.395 ;
        RECT 95.070 168.225 95.240 168.895 ;
        RECT 96.460 168.790 96.630 168.935 ;
        RECT 95.895 168.385 96.225 168.755 ;
        RECT 96.460 168.460 96.745 168.790 ;
        RECT 93.885 168.055 94.815 168.225 ;
        RECT 93.885 168.020 94.060 168.055 ;
        RECT 93.530 167.655 94.060 168.020 ;
        RECT 94.485 167.485 94.815 167.885 ;
        RECT 94.985 167.655 95.240 168.225 ;
        RECT 96.460 168.205 96.630 168.460 ;
        RECT 95.965 168.035 96.630 168.205 ;
        RECT 96.915 168.160 97.085 168.960 ;
        RECT 97.715 168.945 101.225 170.035 ;
        RECT 97.715 168.425 99.405 168.945 ;
        RECT 101.395 168.870 101.685 170.035 ;
        RECT 102.780 168.845 103.035 169.725 ;
        RECT 103.205 168.895 103.510 170.035 ;
        RECT 103.850 169.655 104.180 170.035 ;
        RECT 104.360 169.485 104.530 169.775 ;
        RECT 104.700 169.575 104.950 170.035 ;
        RECT 103.730 169.315 104.530 169.485 ;
        RECT 105.120 169.525 105.990 169.865 ;
        RECT 99.575 168.255 101.225 168.775 ;
        RECT 95.965 167.655 96.135 168.035 ;
        RECT 96.315 167.485 96.645 167.865 ;
        RECT 96.825 167.655 97.085 168.160 ;
        RECT 97.715 167.485 101.225 168.255 ;
        RECT 101.395 167.485 101.685 168.210 ;
        RECT 102.780 168.195 102.990 168.845 ;
        RECT 103.730 168.725 103.900 169.315 ;
        RECT 105.120 169.145 105.290 169.525 ;
        RECT 106.225 169.405 106.395 169.865 ;
        RECT 106.565 169.575 106.935 170.035 ;
        RECT 107.230 169.435 107.400 169.775 ;
        RECT 107.570 169.605 107.900 170.035 ;
        RECT 108.135 169.435 108.305 169.775 ;
        RECT 104.070 168.975 105.290 169.145 ;
        RECT 105.460 169.065 105.920 169.355 ;
        RECT 106.225 169.235 106.785 169.405 ;
        RECT 107.230 169.265 108.305 169.435 ;
        RECT 108.475 169.535 109.155 169.865 ;
        RECT 109.370 169.535 109.620 169.865 ;
        RECT 109.790 169.575 110.040 170.035 ;
        RECT 106.615 169.095 106.785 169.235 ;
        RECT 105.460 169.055 106.425 169.065 ;
        RECT 105.120 168.885 105.290 168.975 ;
        RECT 105.750 168.895 106.425 169.055 ;
        RECT 103.160 168.695 103.900 168.725 ;
        RECT 103.160 168.395 104.075 168.695 ;
        RECT 103.750 168.220 104.075 168.395 ;
        RECT 102.780 167.665 103.035 168.195 ;
        RECT 103.205 167.485 103.510 167.945 ;
        RECT 103.755 167.865 104.075 168.220 ;
        RECT 104.245 168.435 104.785 168.805 ;
        RECT 105.120 168.715 105.525 168.885 ;
        RECT 104.245 168.035 104.485 168.435 ;
        RECT 104.965 168.265 105.185 168.545 ;
        RECT 104.655 168.095 105.185 168.265 ;
        RECT 104.655 167.865 104.825 168.095 ;
        RECT 105.355 167.935 105.525 168.715 ;
        RECT 105.695 168.105 106.045 168.725 ;
        RECT 106.215 168.105 106.425 168.895 ;
        RECT 106.615 168.925 108.115 169.095 ;
        RECT 106.615 168.235 106.785 168.925 ;
        RECT 108.475 168.755 108.645 169.535 ;
        RECT 109.450 169.405 109.620 169.535 ;
        RECT 106.955 168.585 108.645 168.755 ;
        RECT 108.815 168.975 109.280 169.365 ;
        RECT 109.450 169.235 109.845 169.405 ;
        RECT 106.955 168.405 107.125 168.585 ;
        RECT 103.755 167.695 104.825 167.865 ;
        RECT 104.995 167.485 105.185 167.925 ;
        RECT 105.355 167.655 106.305 167.935 ;
        RECT 106.615 167.845 106.875 168.235 ;
        RECT 107.295 168.165 108.085 168.415 ;
        RECT 106.525 167.675 106.875 167.845 ;
        RECT 107.085 167.485 107.415 167.945 ;
        RECT 108.290 167.875 108.460 168.585 ;
        RECT 108.815 168.385 108.985 168.975 ;
        RECT 108.630 168.165 108.985 168.385 ;
        RECT 109.155 168.165 109.505 168.785 ;
        RECT 109.675 167.875 109.845 169.235 ;
        RECT 110.210 169.065 110.535 169.850 ;
        RECT 110.015 168.015 110.475 169.065 ;
        RECT 108.290 167.705 109.145 167.875 ;
        RECT 109.350 167.705 109.845 167.875 ;
        RECT 110.015 167.485 110.345 167.845 ;
        RECT 110.705 167.745 110.875 169.865 ;
        RECT 111.045 169.535 111.375 170.035 ;
        RECT 111.545 169.365 111.800 169.865 ;
        RECT 111.050 169.195 111.800 169.365 ;
        RECT 111.050 168.205 111.280 169.195 ;
        RECT 111.450 168.375 111.800 169.025 ;
        RECT 112.440 168.895 112.775 169.865 ;
        RECT 112.945 168.895 113.115 170.035 ;
        RECT 113.285 169.695 115.315 169.865 ;
        RECT 112.440 168.225 112.610 168.895 ;
        RECT 113.285 168.725 113.455 169.695 ;
        RECT 112.780 168.395 113.035 168.725 ;
        RECT 113.260 168.395 113.455 168.725 ;
        RECT 113.625 169.355 114.750 169.525 ;
        RECT 112.865 168.225 113.035 168.395 ;
        RECT 113.625 168.225 113.795 169.355 ;
        RECT 111.050 168.035 111.800 168.205 ;
        RECT 111.045 167.485 111.375 167.865 ;
        RECT 111.545 167.745 111.800 168.035 ;
        RECT 112.440 167.655 112.695 168.225 ;
        RECT 112.865 168.055 113.795 168.225 ;
        RECT 113.965 169.015 114.975 169.185 ;
        RECT 113.965 168.215 114.135 169.015 ;
        RECT 114.340 168.675 114.615 168.815 ;
        RECT 114.335 168.505 114.615 168.675 ;
        RECT 113.620 168.020 113.795 168.055 ;
        RECT 112.865 167.485 113.195 167.885 ;
        RECT 113.620 167.655 114.150 168.020 ;
        RECT 114.340 167.655 114.615 168.505 ;
        RECT 114.785 167.655 114.975 169.015 ;
        RECT 115.145 169.030 115.315 169.695 ;
        RECT 115.485 169.275 115.655 170.035 ;
        RECT 115.890 169.275 116.405 169.685 ;
        RECT 115.145 168.840 115.895 169.030 ;
        RECT 116.065 168.465 116.405 169.275 ;
        RECT 115.175 168.295 116.405 168.465 ;
        RECT 116.575 168.895 116.960 169.865 ;
        RECT 117.130 169.575 117.455 170.035 ;
        RECT 117.975 169.405 118.255 169.865 ;
        RECT 117.130 169.185 118.255 169.405 ;
        RECT 115.155 167.485 115.665 168.020 ;
        RECT 115.885 167.690 116.130 168.295 ;
        RECT 116.575 168.225 116.855 168.895 ;
        RECT 117.130 168.725 117.580 169.185 ;
        RECT 118.445 169.015 118.845 169.865 ;
        RECT 119.245 169.575 119.515 170.035 ;
        RECT 119.685 169.405 119.970 169.865 ;
        RECT 117.025 168.395 117.580 168.725 ;
        RECT 117.750 168.455 118.845 169.015 ;
        RECT 117.130 168.285 117.580 168.395 ;
        RECT 116.575 167.655 116.960 168.225 ;
        RECT 117.130 168.115 118.255 168.285 ;
        RECT 117.130 167.485 117.455 167.945 ;
        RECT 117.975 167.655 118.255 168.115 ;
        RECT 118.445 167.655 118.845 168.455 ;
        RECT 119.015 169.185 119.970 169.405 ;
        RECT 119.015 168.285 119.225 169.185 ;
        RECT 120.345 169.105 120.515 169.865 ;
        RECT 120.695 169.275 121.025 170.035 ;
        RECT 119.395 168.455 120.085 169.015 ;
        RECT 120.345 168.935 121.010 169.105 ;
        RECT 121.195 168.960 121.465 169.865 ;
        RECT 121.640 169.610 121.975 170.035 ;
        RECT 122.145 169.430 122.330 169.835 ;
        RECT 120.840 168.790 121.010 168.935 ;
        RECT 120.275 168.385 120.605 168.755 ;
        RECT 120.840 168.460 121.125 168.790 ;
        RECT 119.015 168.115 119.970 168.285 ;
        RECT 120.840 168.205 121.010 168.460 ;
        RECT 119.245 167.485 119.515 167.945 ;
        RECT 119.685 167.655 119.970 168.115 ;
        RECT 120.345 168.035 121.010 168.205 ;
        RECT 121.295 168.160 121.465 168.960 ;
        RECT 120.345 167.655 120.515 168.035 ;
        RECT 120.695 167.485 121.025 167.865 ;
        RECT 121.205 167.655 121.465 168.160 ;
        RECT 121.665 169.255 122.330 169.430 ;
        RECT 122.535 169.255 122.865 170.035 ;
        RECT 121.665 168.225 122.005 169.255 ;
        RECT 123.035 169.065 123.305 169.835 ;
        RECT 122.175 168.895 123.305 169.065 ;
        RECT 122.175 168.395 122.425 168.895 ;
        RECT 121.665 168.055 122.350 168.225 ;
        RECT 122.605 168.145 122.965 168.725 ;
        RECT 121.640 167.485 121.975 167.885 ;
        RECT 122.145 167.655 122.350 168.055 ;
        RECT 123.135 167.985 123.305 168.895 ;
        RECT 123.475 168.945 126.065 170.035 ;
        RECT 126.235 168.945 127.445 170.035 ;
        RECT 123.475 168.425 124.685 168.945 ;
        RECT 124.855 168.255 126.065 168.775 ;
        RECT 126.235 168.405 126.755 168.945 ;
        RECT 122.560 167.485 122.835 167.965 ;
        RECT 123.045 167.655 123.305 167.985 ;
        RECT 123.475 167.485 126.065 168.255 ;
        RECT 126.925 168.235 127.445 168.775 ;
        RECT 126.235 167.485 127.445 168.235 ;
        RECT 14.370 167.315 127.530 167.485 ;
        RECT 14.455 166.565 15.665 167.315 ;
        RECT 14.455 166.025 14.975 166.565 ;
        RECT 15.835 166.545 17.505 167.315 ;
        RECT 17.680 166.770 23.025 167.315 ;
        RECT 15.145 165.855 15.665 166.395 ;
        RECT 14.455 164.765 15.665 165.855 ;
        RECT 15.835 165.855 16.585 166.375 ;
        RECT 16.755 166.025 17.505 166.545 ;
        RECT 15.835 164.765 17.505 165.855 ;
        RECT 19.270 165.200 19.620 166.450 ;
        RECT 21.100 165.940 21.440 166.770 ;
        RECT 23.200 166.765 23.455 167.055 ;
        RECT 23.625 166.935 23.955 167.315 ;
        RECT 23.200 166.595 23.950 166.765 ;
        RECT 23.200 165.775 23.550 166.425 ;
        RECT 23.720 165.605 23.950 166.595 ;
        RECT 23.200 165.435 23.950 165.605 ;
        RECT 17.680 164.765 23.025 165.200 ;
        RECT 23.200 164.935 23.455 165.435 ;
        RECT 23.625 164.765 23.955 165.265 ;
        RECT 24.125 164.935 24.295 167.055 ;
        RECT 24.655 166.955 24.985 167.315 ;
        RECT 25.155 166.925 25.650 167.095 ;
        RECT 25.855 166.925 26.710 167.095 ;
        RECT 24.525 165.735 24.985 166.785 ;
        RECT 24.465 164.950 24.790 165.735 ;
        RECT 25.155 165.565 25.325 166.925 ;
        RECT 25.495 166.015 25.845 166.635 ;
        RECT 26.015 166.415 26.370 166.635 ;
        RECT 26.015 165.825 26.185 166.415 ;
        RECT 26.540 166.215 26.710 166.925 ;
        RECT 27.585 166.855 27.915 167.315 ;
        RECT 28.125 166.955 28.475 167.125 ;
        RECT 26.915 166.385 27.705 166.635 ;
        RECT 28.125 166.565 28.385 166.955 ;
        RECT 28.695 166.865 29.645 167.145 ;
        RECT 29.815 166.875 30.005 167.315 ;
        RECT 30.175 166.935 31.245 167.105 ;
        RECT 27.875 166.215 28.045 166.395 ;
        RECT 25.155 165.395 25.550 165.565 ;
        RECT 25.720 165.435 26.185 165.825 ;
        RECT 26.355 166.045 28.045 166.215 ;
        RECT 25.380 165.265 25.550 165.395 ;
        RECT 26.355 165.265 26.525 166.045 ;
        RECT 28.215 165.875 28.385 166.565 ;
        RECT 26.885 165.705 28.385 165.875 ;
        RECT 28.575 165.905 28.785 166.695 ;
        RECT 28.955 166.075 29.305 166.695 ;
        RECT 29.475 166.085 29.645 166.865 ;
        RECT 30.175 166.705 30.345 166.935 ;
        RECT 29.815 166.535 30.345 166.705 ;
        RECT 29.815 166.255 30.035 166.535 ;
        RECT 30.515 166.365 30.755 166.765 ;
        RECT 29.475 165.915 29.880 166.085 ;
        RECT 30.215 165.995 30.755 166.365 ;
        RECT 30.925 166.580 31.245 166.935 ;
        RECT 31.490 166.855 31.795 167.315 ;
        RECT 31.965 166.605 32.220 167.135 ;
        RECT 30.925 166.405 31.250 166.580 ;
        RECT 30.925 166.105 31.840 166.405 ;
        RECT 31.100 166.075 31.840 166.105 ;
        RECT 28.575 165.745 29.250 165.905 ;
        RECT 29.710 165.825 29.880 165.915 ;
        RECT 28.575 165.735 29.540 165.745 ;
        RECT 28.215 165.565 28.385 165.705 ;
        RECT 24.960 164.765 25.210 165.225 ;
        RECT 25.380 164.935 25.630 165.265 ;
        RECT 25.845 164.935 26.525 165.265 ;
        RECT 26.695 165.365 27.770 165.535 ;
        RECT 28.215 165.395 28.775 165.565 ;
        RECT 29.080 165.445 29.540 165.735 ;
        RECT 29.710 165.655 30.930 165.825 ;
        RECT 26.695 165.025 26.865 165.365 ;
        RECT 27.100 164.765 27.430 165.195 ;
        RECT 27.600 165.025 27.770 165.365 ;
        RECT 28.065 164.765 28.435 165.225 ;
        RECT 28.605 164.935 28.775 165.395 ;
        RECT 29.710 165.275 29.880 165.655 ;
        RECT 31.100 165.485 31.270 166.075 ;
        RECT 32.010 165.955 32.220 166.605 ;
        RECT 29.010 164.935 29.880 165.275 ;
        RECT 30.470 165.315 31.270 165.485 ;
        RECT 30.050 164.765 30.300 165.225 ;
        RECT 30.470 165.025 30.640 165.315 ;
        RECT 30.820 164.765 31.150 165.145 ;
        RECT 31.490 164.765 31.795 165.905 ;
        RECT 31.965 165.075 32.220 165.955 ;
        RECT 32.395 166.640 32.655 167.145 ;
        RECT 32.835 166.935 33.165 167.315 ;
        RECT 33.345 166.765 33.515 167.145 ;
        RECT 33.875 166.850 34.125 167.315 ;
        RECT 32.395 165.840 32.565 166.640 ;
        RECT 32.850 166.595 33.515 166.765 ;
        RECT 34.295 166.675 34.465 167.145 ;
        RECT 34.715 166.855 34.885 167.315 ;
        RECT 35.135 166.675 35.305 167.145 ;
        RECT 35.555 166.855 35.725 167.315 ;
        RECT 35.975 166.675 36.145 167.145 ;
        RECT 36.515 166.855 36.780 167.315 ;
        RECT 32.850 166.340 33.020 166.595 ;
        RECT 33.775 166.495 36.145 166.675 ;
        RECT 36.995 166.590 37.285 167.315 ;
        RECT 37.495 166.495 37.725 167.315 ;
        RECT 37.895 166.515 38.225 167.145 ;
        RECT 32.735 166.010 33.020 166.340 ;
        RECT 33.255 166.045 33.585 166.415 ;
        RECT 32.850 165.865 33.020 166.010 ;
        RECT 33.775 165.905 34.125 166.495 ;
        RECT 34.295 166.075 36.805 166.325 ;
        RECT 37.475 166.075 37.805 166.325 ;
        RECT 32.395 164.935 32.665 165.840 ;
        RECT 32.850 165.695 33.515 165.865 ;
        RECT 33.775 165.735 36.225 165.905 ;
        RECT 33.775 165.715 34.545 165.735 ;
        RECT 32.835 164.765 33.165 165.525 ;
        RECT 33.345 164.935 33.515 165.695 ;
        RECT 33.875 164.765 34.045 165.225 ;
        RECT 34.215 164.935 34.545 165.715 ;
        RECT 34.715 164.765 34.885 165.565 ;
        RECT 35.055 164.935 35.385 165.735 ;
        RECT 35.555 164.765 35.725 165.565 ;
        RECT 35.895 164.935 36.225 165.735 ;
        RECT 36.485 164.765 36.780 165.905 ;
        RECT 36.995 164.765 37.285 165.930 ;
        RECT 37.975 165.915 38.225 166.515 ;
        RECT 38.395 166.495 38.605 167.315 ;
        RECT 38.950 166.685 39.235 167.145 ;
        RECT 39.405 166.855 39.675 167.315 ;
        RECT 38.950 166.515 39.905 166.685 ;
        RECT 37.495 164.765 37.725 165.905 ;
        RECT 37.895 164.935 38.225 165.915 ;
        RECT 38.395 164.765 38.605 165.905 ;
        RECT 38.835 165.785 39.525 166.345 ;
        RECT 39.695 165.615 39.905 166.515 ;
        RECT 38.950 165.395 39.905 165.615 ;
        RECT 40.075 166.345 40.475 167.145 ;
        RECT 40.665 166.685 40.945 167.145 ;
        RECT 41.465 166.855 41.790 167.315 ;
        RECT 40.665 166.515 41.790 166.685 ;
        RECT 41.960 166.575 42.345 167.145 ;
        RECT 41.340 166.405 41.790 166.515 ;
        RECT 40.075 165.785 41.170 166.345 ;
        RECT 41.340 166.075 41.895 166.405 ;
        RECT 38.950 164.935 39.235 165.395 ;
        RECT 39.405 164.765 39.675 165.225 ;
        RECT 40.075 164.935 40.475 165.785 ;
        RECT 41.340 165.615 41.790 166.075 ;
        RECT 42.065 165.905 42.345 166.575 ;
        RECT 40.665 165.395 41.790 165.615 ;
        RECT 40.665 164.935 40.945 165.395 ;
        RECT 41.465 164.765 41.790 165.225 ;
        RECT 41.960 164.935 42.345 165.905 ;
        RECT 42.515 166.575 42.900 167.145 ;
        RECT 43.070 166.855 43.395 167.315 ;
        RECT 43.915 166.685 44.195 167.145 ;
        RECT 42.515 165.905 42.795 166.575 ;
        RECT 43.070 166.515 44.195 166.685 ;
        RECT 43.070 166.405 43.520 166.515 ;
        RECT 42.965 166.075 43.520 166.405 ;
        RECT 44.385 166.345 44.785 167.145 ;
        RECT 45.185 166.855 45.455 167.315 ;
        RECT 45.625 166.685 45.910 167.145 ;
        RECT 42.515 164.935 42.900 165.905 ;
        RECT 43.070 165.615 43.520 166.075 ;
        RECT 43.690 165.785 44.785 166.345 ;
        RECT 43.070 165.395 44.195 165.615 ;
        RECT 43.070 164.765 43.395 165.225 ;
        RECT 43.915 164.935 44.195 165.395 ;
        RECT 44.385 164.935 44.785 165.785 ;
        RECT 44.955 166.515 45.910 166.685 ;
        RECT 47.120 166.605 47.375 167.135 ;
        RECT 47.545 166.855 47.850 167.315 ;
        RECT 48.095 166.935 49.165 167.105 ;
        RECT 44.955 165.615 45.165 166.515 ;
        RECT 45.335 165.785 46.025 166.345 ;
        RECT 47.120 165.955 47.330 166.605 ;
        RECT 48.095 166.580 48.415 166.935 ;
        RECT 48.090 166.405 48.415 166.580 ;
        RECT 47.500 166.105 48.415 166.405 ;
        RECT 48.585 166.365 48.825 166.765 ;
        RECT 48.995 166.705 49.165 166.935 ;
        RECT 49.335 166.875 49.525 167.315 ;
        RECT 49.695 166.865 50.645 167.145 ;
        RECT 50.865 166.955 51.215 167.125 ;
        RECT 48.995 166.535 49.525 166.705 ;
        RECT 47.500 166.075 48.240 166.105 ;
        RECT 44.955 165.395 45.910 165.615 ;
        RECT 45.185 164.765 45.455 165.225 ;
        RECT 45.625 164.935 45.910 165.395 ;
        RECT 47.120 165.075 47.375 165.955 ;
        RECT 47.545 164.765 47.850 165.905 ;
        RECT 48.070 165.485 48.240 166.075 ;
        RECT 48.585 165.995 49.125 166.365 ;
        RECT 49.305 166.255 49.525 166.535 ;
        RECT 49.695 166.085 49.865 166.865 ;
        RECT 49.460 165.915 49.865 166.085 ;
        RECT 50.035 166.075 50.385 166.695 ;
        RECT 49.460 165.825 49.630 165.915 ;
        RECT 50.555 165.905 50.765 166.695 ;
        RECT 48.410 165.655 49.630 165.825 ;
        RECT 50.090 165.745 50.765 165.905 ;
        RECT 48.070 165.315 48.870 165.485 ;
        RECT 48.190 164.765 48.520 165.145 ;
        RECT 48.700 165.025 48.870 165.315 ;
        RECT 49.460 165.275 49.630 165.655 ;
        RECT 49.800 165.735 50.765 165.745 ;
        RECT 50.955 166.565 51.215 166.955 ;
        RECT 51.425 166.855 51.755 167.315 ;
        RECT 52.630 166.925 53.485 167.095 ;
        RECT 53.690 166.925 54.185 167.095 ;
        RECT 54.355 166.955 54.685 167.315 ;
        RECT 50.955 165.875 51.125 166.565 ;
        RECT 51.295 166.215 51.465 166.395 ;
        RECT 51.635 166.385 52.425 166.635 ;
        RECT 52.630 166.215 52.800 166.925 ;
        RECT 52.970 166.415 53.325 166.635 ;
        RECT 51.295 166.045 52.985 166.215 ;
        RECT 49.800 165.445 50.260 165.735 ;
        RECT 50.955 165.705 52.455 165.875 ;
        RECT 50.955 165.565 51.125 165.705 ;
        RECT 50.565 165.395 51.125 165.565 ;
        RECT 49.040 164.765 49.290 165.225 ;
        RECT 49.460 164.935 50.330 165.275 ;
        RECT 50.565 164.935 50.735 165.395 ;
        RECT 51.570 165.365 52.645 165.535 ;
        RECT 50.905 164.765 51.275 165.225 ;
        RECT 51.570 165.025 51.740 165.365 ;
        RECT 51.910 164.765 52.240 165.195 ;
        RECT 52.475 165.025 52.645 165.365 ;
        RECT 52.815 165.265 52.985 166.045 ;
        RECT 53.155 165.825 53.325 166.415 ;
        RECT 53.495 166.015 53.845 166.635 ;
        RECT 53.155 165.435 53.620 165.825 ;
        RECT 54.015 165.565 54.185 166.925 ;
        RECT 54.355 165.735 54.815 166.785 ;
        RECT 53.790 165.395 54.185 165.565 ;
        RECT 53.790 165.265 53.960 165.395 ;
        RECT 52.815 164.935 53.495 165.265 ;
        RECT 53.710 164.935 53.960 165.265 ;
        RECT 54.130 164.765 54.380 165.225 ;
        RECT 54.550 164.950 54.875 165.735 ;
        RECT 55.045 164.935 55.215 167.055 ;
        RECT 55.385 166.935 55.715 167.315 ;
        RECT 55.885 166.765 56.140 167.055 ;
        RECT 55.390 166.595 56.140 166.765 ;
        RECT 55.390 165.605 55.620 166.595 ;
        RECT 56.315 166.545 57.985 167.315 ;
        RECT 55.790 165.775 56.140 166.425 ;
        RECT 56.315 165.855 57.065 166.375 ;
        RECT 57.235 166.025 57.985 166.545 ;
        RECT 58.215 166.495 58.425 167.315 ;
        RECT 58.595 166.515 58.925 167.145 ;
        RECT 58.595 165.915 58.845 166.515 ;
        RECT 59.095 166.495 59.325 167.315 ;
        RECT 60.145 166.515 60.475 167.315 ;
        RECT 60.645 166.665 60.815 167.145 ;
        RECT 60.985 166.835 61.315 167.315 ;
        RECT 61.485 166.665 61.655 167.145 ;
        RECT 61.905 166.835 62.145 167.315 ;
        RECT 62.325 166.665 62.495 167.145 ;
        RECT 60.645 166.495 61.655 166.665 ;
        RECT 61.860 166.495 62.495 166.665 ;
        RECT 62.755 166.590 63.045 167.315 ;
        RECT 63.215 166.545 64.885 167.315 ;
        RECT 65.115 166.835 65.395 167.315 ;
        RECT 65.565 166.665 65.825 167.055 ;
        RECT 66.000 166.835 66.255 167.315 ;
        RECT 66.425 166.665 66.720 167.055 ;
        RECT 66.900 166.835 67.175 167.315 ;
        RECT 67.345 166.815 67.645 167.145 ;
        RECT 59.015 166.075 59.345 166.325 ;
        RECT 60.645 166.295 61.140 166.495 ;
        RECT 61.860 166.325 62.030 166.495 ;
        RECT 60.645 166.125 61.145 166.295 ;
        RECT 61.530 166.155 62.030 166.325 ;
        RECT 60.645 165.955 61.140 166.125 ;
        RECT 55.390 165.435 56.140 165.605 ;
        RECT 55.385 164.765 55.715 165.265 ;
        RECT 55.885 164.935 56.140 165.435 ;
        RECT 56.315 164.765 57.985 165.855 ;
        RECT 58.215 164.765 58.425 165.905 ;
        RECT 58.595 164.935 58.925 165.915 ;
        RECT 59.095 164.765 59.325 165.905 ;
        RECT 60.145 164.765 60.475 165.915 ;
        RECT 60.645 165.785 61.655 165.955 ;
        RECT 60.645 164.935 60.815 165.785 ;
        RECT 60.985 164.765 61.315 165.565 ;
        RECT 61.485 164.935 61.655 165.785 ;
        RECT 61.860 165.915 62.030 166.155 ;
        RECT 62.200 166.085 62.580 166.325 ;
        RECT 61.860 165.745 62.575 165.915 ;
        RECT 61.835 164.765 62.075 165.565 ;
        RECT 62.245 164.935 62.575 165.745 ;
        RECT 62.755 164.765 63.045 165.930 ;
        RECT 63.215 165.855 63.965 166.375 ;
        RECT 64.135 166.025 64.885 166.545 ;
        RECT 65.070 166.495 66.720 166.665 ;
        RECT 65.070 165.985 65.475 166.495 ;
        RECT 65.645 166.155 66.785 166.325 ;
        RECT 63.215 164.765 64.885 165.855 ;
        RECT 65.070 165.815 65.825 165.985 ;
        RECT 65.110 164.765 65.395 165.635 ;
        RECT 65.565 165.565 65.825 165.815 ;
        RECT 66.615 165.905 66.785 166.155 ;
        RECT 66.955 166.075 67.305 166.645 ;
        RECT 67.475 165.905 67.645 166.815 ;
        RECT 66.615 165.735 67.645 165.905 ;
        RECT 65.565 165.395 66.685 165.565 ;
        RECT 65.565 164.935 65.825 165.395 ;
        RECT 66.000 164.765 66.255 165.225 ;
        RECT 66.425 164.935 66.685 165.395 ;
        RECT 66.855 164.765 67.165 165.565 ;
        RECT 67.335 164.935 67.645 165.735 ;
        RECT 67.815 166.815 68.115 167.145 ;
        RECT 68.285 166.835 68.560 167.315 ;
        RECT 67.815 165.905 67.985 166.815 ;
        RECT 68.740 166.665 69.035 167.055 ;
        RECT 69.205 166.835 69.460 167.315 ;
        RECT 69.635 166.665 69.895 167.055 ;
        RECT 70.065 166.835 70.345 167.315 ;
        RECT 70.585 166.785 70.915 167.145 ;
        RECT 71.085 166.955 71.415 167.315 ;
        RECT 71.615 166.785 71.945 167.145 ;
        RECT 68.155 166.075 68.505 166.645 ;
        RECT 68.740 166.495 70.390 166.665 ;
        RECT 70.585 166.575 71.945 166.785 ;
        RECT 72.455 166.555 73.165 167.145 ;
        RECT 68.675 166.155 69.815 166.325 ;
        RECT 68.675 165.905 68.845 166.155 ;
        RECT 69.985 165.985 70.390 166.495 ;
        RECT 72.935 166.465 73.165 166.555 ;
        RECT 73.335 166.545 75.005 167.315 ;
        RECT 70.575 166.075 70.885 166.405 ;
        RECT 71.095 166.075 71.470 166.405 ;
        RECT 71.790 166.075 72.285 166.405 ;
        RECT 67.815 165.735 68.845 165.905 ;
        RECT 69.635 165.815 70.390 165.985 ;
        RECT 67.815 164.935 68.125 165.735 ;
        RECT 69.635 165.565 69.895 165.815 ;
        RECT 68.295 164.765 68.605 165.565 ;
        RECT 68.775 165.395 69.895 165.565 ;
        RECT 68.775 164.935 69.035 165.395 ;
        RECT 69.205 164.765 69.460 165.225 ;
        RECT 69.635 164.935 69.895 165.395 ;
        RECT 70.065 164.765 70.350 165.635 ;
        RECT 70.585 164.765 70.915 165.825 ;
        RECT 71.095 165.150 71.265 166.075 ;
        RECT 71.435 165.585 71.765 165.805 ;
        RECT 71.960 165.785 72.285 166.075 ;
        RECT 72.460 165.785 72.790 166.325 ;
        RECT 72.960 165.585 73.165 166.465 ;
        RECT 71.435 165.355 73.165 165.585 ;
        RECT 71.435 164.955 71.765 165.355 ;
        RECT 71.935 164.765 72.265 165.125 ;
        RECT 72.465 164.935 73.165 165.355 ;
        RECT 73.335 165.855 74.085 166.375 ;
        RECT 74.255 166.025 75.005 166.545 ;
        RECT 75.550 166.605 75.805 167.135 ;
        RECT 75.985 166.855 76.270 167.315 ;
        RECT 73.335 164.765 75.005 165.855 ;
        RECT 75.550 165.745 75.730 166.605 ;
        RECT 76.450 166.405 76.700 167.055 ;
        RECT 75.900 166.075 76.700 166.405 ;
        RECT 75.550 165.275 75.805 165.745 ;
        RECT 75.465 165.105 75.805 165.275 ;
        RECT 75.550 165.075 75.805 165.105 ;
        RECT 75.985 164.765 76.270 165.565 ;
        RECT 76.450 165.485 76.700 166.075 ;
        RECT 76.900 166.720 77.220 167.050 ;
        RECT 77.400 166.835 78.060 167.315 ;
        RECT 78.260 166.925 79.110 167.095 ;
        RECT 76.900 165.825 77.090 166.720 ;
        RECT 77.410 166.395 78.070 166.665 ;
        RECT 77.740 166.335 78.070 166.395 ;
        RECT 77.260 166.165 77.590 166.225 ;
        RECT 78.260 166.165 78.430 166.925 ;
        RECT 79.670 166.855 79.990 167.315 ;
        RECT 80.190 166.675 80.440 167.105 ;
        RECT 80.730 166.875 81.140 167.315 ;
        RECT 81.310 166.935 82.325 167.135 ;
        RECT 78.600 166.505 79.850 166.675 ;
        RECT 78.600 166.385 78.930 166.505 ;
        RECT 77.260 165.995 79.160 166.165 ;
        RECT 76.900 165.655 78.820 165.825 ;
        RECT 76.900 165.635 77.220 165.655 ;
        RECT 76.450 164.975 76.780 165.485 ;
        RECT 77.050 165.025 77.220 165.635 ;
        RECT 78.990 165.485 79.160 165.995 ;
        RECT 79.330 165.925 79.510 166.335 ;
        RECT 79.680 165.745 79.850 166.505 ;
        RECT 77.390 164.765 77.720 165.455 ;
        RECT 77.950 165.315 79.160 165.485 ;
        RECT 79.330 165.435 79.850 165.745 ;
        RECT 80.020 166.335 80.440 166.675 ;
        RECT 80.730 166.335 81.140 166.665 ;
        RECT 80.020 165.565 80.210 166.335 ;
        RECT 81.310 166.205 81.480 166.935 ;
        RECT 82.625 166.765 82.795 167.095 ;
        RECT 82.965 166.935 83.295 167.315 ;
        RECT 81.650 166.385 82.000 166.755 ;
        RECT 81.310 166.165 81.730 166.205 ;
        RECT 80.380 165.995 81.730 166.165 ;
        RECT 80.380 165.835 80.630 165.995 ;
        RECT 81.140 165.565 81.390 165.825 ;
        RECT 80.020 165.315 81.390 165.565 ;
        RECT 77.950 165.025 78.190 165.315 ;
        RECT 78.990 165.235 79.160 165.315 ;
        RECT 78.390 164.765 78.810 165.145 ;
        RECT 78.990 164.985 79.620 165.235 ;
        RECT 80.090 164.765 80.420 165.145 ;
        RECT 80.590 165.025 80.760 165.315 ;
        RECT 81.560 165.150 81.730 165.995 ;
        RECT 82.180 165.825 82.400 166.695 ;
        RECT 82.625 166.575 83.320 166.765 ;
        RECT 81.900 165.445 82.400 165.825 ;
        RECT 82.570 165.775 82.980 166.395 ;
        RECT 83.150 165.605 83.320 166.575 ;
        RECT 82.625 165.435 83.320 165.605 ;
        RECT 80.940 164.765 81.320 165.145 ;
        RECT 81.560 164.980 82.390 165.150 ;
        RECT 82.625 164.935 82.795 165.435 ;
        RECT 82.965 164.765 83.295 165.265 ;
        RECT 83.510 164.935 83.735 167.055 ;
        RECT 83.905 166.935 84.235 167.315 ;
        RECT 84.405 166.765 84.575 167.055 ;
        RECT 83.910 166.595 84.575 166.765 ;
        RECT 83.910 165.605 84.140 166.595 ;
        RECT 84.895 166.495 85.105 167.315 ;
        RECT 85.275 166.515 85.605 167.145 ;
        RECT 84.310 165.775 84.660 166.425 ;
        RECT 85.275 165.915 85.525 166.515 ;
        RECT 85.775 166.495 86.005 167.315 ;
        RECT 86.275 166.495 86.485 167.315 ;
        RECT 86.655 166.515 86.985 167.145 ;
        RECT 85.695 166.075 86.025 166.325 ;
        RECT 86.655 165.915 86.905 166.515 ;
        RECT 87.155 166.495 87.385 167.315 ;
        RECT 88.515 166.590 88.805 167.315 ;
        RECT 89.435 166.545 92.945 167.315 ;
        RECT 87.075 166.075 87.405 166.325 ;
        RECT 83.910 165.435 84.575 165.605 ;
        RECT 83.905 164.765 84.235 165.265 ;
        RECT 84.405 164.935 84.575 165.435 ;
        RECT 84.895 164.765 85.105 165.905 ;
        RECT 85.275 164.935 85.605 165.915 ;
        RECT 85.775 164.765 86.005 165.905 ;
        RECT 86.275 164.765 86.485 165.905 ;
        RECT 86.655 164.935 86.985 165.915 ;
        RECT 87.155 164.765 87.385 165.905 ;
        RECT 88.515 164.765 88.805 165.930 ;
        RECT 89.435 165.855 91.125 166.375 ;
        RECT 91.295 166.025 92.945 166.545 ;
        RECT 93.390 166.505 93.635 167.110 ;
        RECT 93.855 166.780 94.365 167.315 ;
        RECT 93.115 166.335 94.345 166.505 ;
        RECT 89.435 164.765 92.945 165.855 ;
        RECT 93.115 165.525 93.455 166.335 ;
        RECT 93.625 165.770 94.375 165.960 ;
        RECT 93.115 165.115 93.630 165.525 ;
        RECT 93.865 164.765 94.035 165.525 ;
        RECT 94.205 165.105 94.375 165.770 ;
        RECT 94.545 165.785 94.735 167.145 ;
        RECT 94.905 166.295 95.180 167.145 ;
        RECT 95.370 166.780 95.900 167.145 ;
        RECT 96.325 166.915 96.655 167.315 ;
        RECT 95.725 166.745 95.900 166.780 ;
        RECT 94.905 166.125 95.185 166.295 ;
        RECT 94.905 165.985 95.180 166.125 ;
        RECT 95.385 165.785 95.555 166.585 ;
        RECT 94.545 165.615 95.555 165.785 ;
        RECT 95.725 166.575 96.655 166.745 ;
        RECT 96.825 166.575 97.080 167.145 ;
        RECT 95.725 165.445 95.895 166.575 ;
        RECT 96.485 166.405 96.655 166.575 ;
        RECT 94.770 165.275 95.895 165.445 ;
        RECT 96.065 166.075 96.260 166.405 ;
        RECT 96.485 166.075 96.740 166.405 ;
        RECT 96.065 165.105 96.235 166.075 ;
        RECT 96.910 165.905 97.080 166.575 ;
        RECT 97.630 166.605 97.885 167.135 ;
        RECT 98.065 166.855 98.350 167.315 ;
        RECT 97.630 165.955 97.810 166.605 ;
        RECT 98.530 166.405 98.780 167.055 ;
        RECT 97.980 166.075 98.780 166.405 ;
        RECT 94.205 164.935 96.235 165.105 ;
        RECT 96.405 164.765 96.575 165.905 ;
        RECT 96.745 164.935 97.080 165.905 ;
        RECT 97.545 165.785 97.810 165.955 ;
        RECT 97.630 165.745 97.810 165.785 ;
        RECT 97.630 165.075 97.885 165.745 ;
        RECT 98.065 164.765 98.350 165.565 ;
        RECT 98.530 165.485 98.780 166.075 ;
        RECT 98.980 166.720 99.300 167.050 ;
        RECT 99.480 166.835 100.140 167.315 ;
        RECT 100.340 166.925 101.190 167.095 ;
        RECT 98.980 165.825 99.170 166.720 ;
        RECT 99.490 166.395 100.150 166.665 ;
        RECT 99.820 166.335 100.150 166.395 ;
        RECT 99.340 166.165 99.670 166.225 ;
        RECT 100.340 166.165 100.510 166.925 ;
        RECT 101.750 166.855 102.070 167.315 ;
        RECT 102.270 166.675 102.520 167.105 ;
        RECT 102.810 166.875 103.220 167.315 ;
        RECT 103.390 166.935 104.405 167.135 ;
        RECT 100.680 166.505 101.930 166.675 ;
        RECT 100.680 166.385 101.010 166.505 ;
        RECT 99.340 165.995 101.240 166.165 ;
        RECT 98.980 165.655 100.900 165.825 ;
        RECT 98.980 165.635 99.300 165.655 ;
        RECT 98.530 164.975 98.860 165.485 ;
        RECT 99.130 165.025 99.300 165.635 ;
        RECT 101.070 165.485 101.240 165.995 ;
        RECT 101.410 165.925 101.590 166.335 ;
        RECT 101.760 165.745 101.930 166.505 ;
        RECT 99.470 164.765 99.800 165.455 ;
        RECT 100.030 165.315 101.240 165.485 ;
        RECT 101.410 165.435 101.930 165.745 ;
        RECT 102.100 166.335 102.520 166.675 ;
        RECT 102.810 166.335 103.220 166.665 ;
        RECT 102.100 165.565 102.290 166.335 ;
        RECT 103.390 166.205 103.560 166.935 ;
        RECT 104.705 166.765 104.875 167.095 ;
        RECT 105.045 166.935 105.375 167.315 ;
        RECT 103.730 166.385 104.080 166.755 ;
        RECT 103.390 166.165 103.810 166.205 ;
        RECT 102.460 165.995 103.810 166.165 ;
        RECT 102.460 165.835 102.710 165.995 ;
        RECT 103.220 165.565 103.470 165.825 ;
        RECT 102.100 165.315 103.470 165.565 ;
        RECT 100.030 165.025 100.270 165.315 ;
        RECT 101.070 165.235 101.240 165.315 ;
        RECT 100.470 164.765 100.890 165.145 ;
        RECT 101.070 164.985 101.700 165.235 ;
        RECT 102.170 164.765 102.500 165.145 ;
        RECT 102.670 165.025 102.840 165.315 ;
        RECT 103.640 165.150 103.810 165.995 ;
        RECT 104.260 165.825 104.480 166.695 ;
        RECT 104.705 166.575 105.400 166.765 ;
        RECT 103.980 165.445 104.480 165.825 ;
        RECT 104.650 165.775 105.060 166.395 ;
        RECT 105.230 165.605 105.400 166.575 ;
        RECT 104.705 165.435 105.400 165.605 ;
        RECT 103.020 164.765 103.400 165.145 ;
        RECT 103.640 164.980 104.470 165.150 ;
        RECT 104.705 164.935 104.875 165.435 ;
        RECT 105.045 164.765 105.375 165.265 ;
        RECT 105.590 164.935 105.815 167.055 ;
        RECT 105.985 166.935 106.315 167.315 ;
        RECT 106.485 166.765 106.655 167.055 ;
        RECT 105.990 166.595 106.655 166.765 ;
        RECT 107.030 166.685 107.315 167.145 ;
        RECT 107.485 166.855 107.755 167.315 ;
        RECT 105.990 165.605 106.220 166.595 ;
        RECT 107.030 166.515 107.985 166.685 ;
        RECT 106.390 165.775 106.740 166.425 ;
        RECT 106.915 165.785 107.605 166.345 ;
        RECT 107.775 165.615 107.985 166.515 ;
        RECT 105.990 165.435 106.655 165.605 ;
        RECT 105.985 164.765 106.315 165.265 ;
        RECT 106.485 164.935 106.655 165.435 ;
        RECT 107.030 165.395 107.985 165.615 ;
        RECT 108.155 166.345 108.555 167.145 ;
        RECT 108.745 166.685 109.025 167.145 ;
        RECT 109.545 166.855 109.870 167.315 ;
        RECT 108.745 166.515 109.870 166.685 ;
        RECT 110.040 166.575 110.425 167.145 ;
        RECT 109.420 166.405 109.870 166.515 ;
        RECT 108.155 165.785 109.250 166.345 ;
        RECT 109.420 166.075 109.975 166.405 ;
        RECT 107.030 164.935 107.315 165.395 ;
        RECT 107.485 164.765 107.755 165.225 ;
        RECT 108.155 164.935 108.555 165.785 ;
        RECT 109.420 165.615 109.870 166.075 ;
        RECT 110.145 165.905 110.425 166.575 ;
        RECT 110.710 166.685 110.995 167.145 ;
        RECT 111.165 166.855 111.435 167.315 ;
        RECT 110.710 166.515 111.665 166.685 ;
        RECT 108.745 165.395 109.870 165.615 ;
        RECT 108.745 164.935 109.025 165.395 ;
        RECT 109.545 164.765 109.870 165.225 ;
        RECT 110.040 164.935 110.425 165.905 ;
        RECT 110.595 165.785 111.285 166.345 ;
        RECT 111.455 165.615 111.665 166.515 ;
        RECT 110.710 165.395 111.665 165.615 ;
        RECT 111.835 166.345 112.235 167.145 ;
        RECT 112.425 166.685 112.705 167.145 ;
        RECT 113.225 166.855 113.550 167.315 ;
        RECT 112.425 166.515 113.550 166.685 ;
        RECT 113.720 166.575 114.105 167.145 ;
        RECT 114.275 166.590 114.565 167.315 ;
        RECT 115.660 166.605 115.915 167.135 ;
        RECT 116.085 166.855 116.390 167.315 ;
        RECT 116.635 166.935 117.705 167.105 ;
        RECT 113.100 166.405 113.550 166.515 ;
        RECT 111.835 165.785 112.930 166.345 ;
        RECT 113.100 166.075 113.655 166.405 ;
        RECT 110.710 164.935 110.995 165.395 ;
        RECT 111.165 164.765 111.435 165.225 ;
        RECT 111.835 164.935 112.235 165.785 ;
        RECT 113.100 165.615 113.550 166.075 ;
        RECT 113.825 165.905 114.105 166.575 ;
        RECT 115.660 165.955 115.870 166.605 ;
        RECT 116.635 166.580 116.955 166.935 ;
        RECT 116.630 166.405 116.955 166.580 ;
        RECT 116.040 166.105 116.955 166.405 ;
        RECT 117.125 166.365 117.365 166.765 ;
        RECT 117.535 166.705 117.705 166.935 ;
        RECT 117.875 166.875 118.065 167.315 ;
        RECT 118.235 166.865 119.185 167.145 ;
        RECT 119.405 166.955 119.755 167.125 ;
        RECT 117.535 166.535 118.065 166.705 ;
        RECT 116.040 166.075 116.780 166.105 ;
        RECT 112.425 165.395 113.550 165.615 ;
        RECT 112.425 164.935 112.705 165.395 ;
        RECT 113.225 164.765 113.550 165.225 ;
        RECT 113.720 164.935 114.105 165.905 ;
        RECT 114.275 164.765 114.565 165.930 ;
        RECT 115.660 165.075 115.915 165.955 ;
        RECT 116.085 164.765 116.390 165.905 ;
        RECT 116.610 165.485 116.780 166.075 ;
        RECT 117.125 165.995 117.665 166.365 ;
        RECT 117.845 166.255 118.065 166.535 ;
        RECT 118.235 166.085 118.405 166.865 ;
        RECT 118.000 165.915 118.405 166.085 ;
        RECT 118.575 166.075 118.925 166.695 ;
        RECT 118.000 165.825 118.170 165.915 ;
        RECT 119.095 165.905 119.305 166.695 ;
        RECT 116.950 165.655 118.170 165.825 ;
        RECT 118.630 165.745 119.305 165.905 ;
        RECT 116.610 165.315 117.410 165.485 ;
        RECT 116.730 164.765 117.060 165.145 ;
        RECT 117.240 165.025 117.410 165.315 ;
        RECT 118.000 165.275 118.170 165.655 ;
        RECT 118.340 165.735 119.305 165.745 ;
        RECT 119.495 166.565 119.755 166.955 ;
        RECT 119.965 166.855 120.295 167.315 ;
        RECT 121.170 166.925 122.025 167.095 ;
        RECT 122.230 166.925 122.725 167.095 ;
        RECT 122.895 166.955 123.225 167.315 ;
        RECT 119.495 165.875 119.665 166.565 ;
        RECT 119.835 166.215 120.005 166.395 ;
        RECT 120.175 166.385 120.965 166.635 ;
        RECT 121.170 166.215 121.340 166.925 ;
        RECT 121.510 166.415 121.865 166.635 ;
        RECT 119.835 166.045 121.525 166.215 ;
        RECT 118.340 165.445 118.800 165.735 ;
        RECT 119.495 165.705 120.995 165.875 ;
        RECT 119.495 165.565 119.665 165.705 ;
        RECT 119.105 165.395 119.665 165.565 ;
        RECT 117.580 164.765 117.830 165.225 ;
        RECT 118.000 164.935 118.870 165.275 ;
        RECT 119.105 164.935 119.275 165.395 ;
        RECT 120.110 165.365 121.185 165.535 ;
        RECT 119.445 164.765 119.815 165.225 ;
        RECT 120.110 165.025 120.280 165.365 ;
        RECT 120.450 164.765 120.780 165.195 ;
        RECT 121.015 165.025 121.185 165.365 ;
        RECT 121.355 165.265 121.525 166.045 ;
        RECT 121.695 165.825 121.865 166.415 ;
        RECT 122.035 166.015 122.385 166.635 ;
        RECT 121.695 165.435 122.160 165.825 ;
        RECT 122.555 165.565 122.725 166.925 ;
        RECT 122.895 165.735 123.355 166.785 ;
        RECT 122.330 165.395 122.725 165.565 ;
        RECT 122.330 165.265 122.500 165.395 ;
        RECT 121.355 164.935 122.035 165.265 ;
        RECT 122.250 164.935 122.500 165.265 ;
        RECT 122.670 164.765 122.920 165.225 ;
        RECT 123.090 164.950 123.415 165.735 ;
        RECT 123.585 164.935 123.755 167.055 ;
        RECT 123.925 166.935 124.255 167.315 ;
        RECT 124.425 166.765 124.680 167.055 ;
        RECT 123.930 166.595 124.680 166.765 ;
        RECT 123.930 165.605 124.160 166.595 ;
        RECT 124.855 166.565 126.065 167.315 ;
        RECT 126.235 166.565 127.445 167.315 ;
        RECT 124.330 165.775 124.680 166.425 ;
        RECT 124.855 165.855 125.375 166.395 ;
        RECT 125.545 166.025 126.065 166.565 ;
        RECT 126.235 165.855 126.755 166.395 ;
        RECT 126.925 166.025 127.445 166.565 ;
        RECT 123.930 165.435 124.680 165.605 ;
        RECT 123.925 164.765 124.255 165.265 ;
        RECT 124.425 164.935 124.680 165.435 ;
        RECT 124.855 164.765 126.065 165.855 ;
        RECT 126.235 164.765 127.445 165.855 ;
        RECT 14.370 164.595 127.530 164.765 ;
        RECT 14.455 163.505 15.665 164.595 ;
        RECT 14.455 162.795 14.975 163.335 ;
        RECT 15.145 162.965 15.665 163.505 ;
        RECT 15.835 163.505 18.425 164.595 ;
        RECT 18.600 164.160 23.945 164.595 ;
        RECT 15.835 162.985 17.045 163.505 ;
        RECT 17.215 162.815 18.425 163.335 ;
        RECT 20.190 162.910 20.540 164.160 ;
        RECT 24.115 163.430 24.405 164.595 ;
        RECT 25.495 163.520 25.765 164.425 ;
        RECT 25.935 163.835 26.265 164.595 ;
        RECT 26.445 163.665 26.615 164.425 ;
        RECT 26.880 163.925 27.135 164.425 ;
        RECT 27.305 164.095 27.635 164.595 ;
        RECT 26.880 163.755 27.630 163.925 ;
        RECT 14.455 162.045 15.665 162.795 ;
        RECT 15.835 162.045 18.425 162.815 ;
        RECT 22.020 162.590 22.360 163.420 ;
        RECT 18.600 162.045 23.945 162.590 ;
        RECT 24.115 162.045 24.405 162.770 ;
        RECT 25.495 162.720 25.665 163.520 ;
        RECT 25.950 163.495 26.615 163.665 ;
        RECT 25.950 163.350 26.120 163.495 ;
        RECT 25.835 163.020 26.120 163.350 ;
        RECT 25.950 162.765 26.120 163.020 ;
        RECT 26.355 162.945 26.685 163.315 ;
        RECT 26.880 162.935 27.230 163.585 ;
        RECT 27.400 162.765 27.630 163.755 ;
        RECT 25.495 162.215 25.755 162.720 ;
        RECT 25.950 162.595 26.615 162.765 ;
        RECT 25.935 162.045 26.265 162.425 ;
        RECT 26.445 162.215 26.615 162.595 ;
        RECT 26.880 162.595 27.630 162.765 ;
        RECT 26.880 162.305 27.135 162.595 ;
        RECT 27.305 162.045 27.635 162.425 ;
        RECT 27.805 162.305 27.975 164.425 ;
        RECT 28.145 163.625 28.470 164.410 ;
        RECT 28.640 164.135 28.890 164.595 ;
        RECT 29.060 164.095 29.310 164.425 ;
        RECT 29.525 164.095 30.205 164.425 ;
        RECT 29.060 163.965 29.230 164.095 ;
        RECT 28.835 163.795 29.230 163.965 ;
        RECT 28.205 162.575 28.665 163.625 ;
        RECT 28.835 162.435 29.005 163.795 ;
        RECT 29.400 163.535 29.865 163.925 ;
        RECT 29.175 162.725 29.525 163.345 ;
        RECT 29.695 162.945 29.865 163.535 ;
        RECT 30.035 163.315 30.205 164.095 ;
        RECT 30.375 163.995 30.545 164.335 ;
        RECT 30.780 164.165 31.110 164.595 ;
        RECT 31.280 163.995 31.450 164.335 ;
        RECT 31.745 164.135 32.115 164.595 ;
        RECT 30.375 163.825 31.450 163.995 ;
        RECT 32.285 163.965 32.455 164.425 ;
        RECT 32.690 164.085 33.560 164.425 ;
        RECT 33.730 164.135 33.980 164.595 ;
        RECT 31.895 163.795 32.455 163.965 ;
        RECT 31.895 163.655 32.065 163.795 ;
        RECT 30.565 163.485 32.065 163.655 ;
        RECT 32.760 163.625 33.220 163.915 ;
        RECT 30.035 163.145 31.725 163.315 ;
        RECT 29.695 162.725 30.050 162.945 ;
        RECT 30.220 162.435 30.390 163.145 ;
        RECT 30.595 162.725 31.385 162.975 ;
        RECT 31.555 162.965 31.725 163.145 ;
        RECT 31.895 162.795 32.065 163.485 ;
        RECT 28.335 162.045 28.665 162.405 ;
        RECT 28.835 162.265 29.330 162.435 ;
        RECT 29.535 162.265 30.390 162.435 ;
        RECT 31.265 162.045 31.595 162.505 ;
        RECT 31.805 162.405 32.065 162.795 ;
        RECT 32.255 163.615 33.220 163.625 ;
        RECT 33.390 163.705 33.560 164.085 ;
        RECT 34.150 164.045 34.320 164.335 ;
        RECT 34.500 164.215 34.830 164.595 ;
        RECT 34.150 163.875 34.950 164.045 ;
        RECT 32.255 163.455 32.930 163.615 ;
        RECT 33.390 163.535 34.610 163.705 ;
        RECT 32.255 162.665 32.465 163.455 ;
        RECT 33.390 163.445 33.560 163.535 ;
        RECT 32.635 162.665 32.985 163.285 ;
        RECT 33.155 163.275 33.560 163.445 ;
        RECT 33.155 162.495 33.325 163.275 ;
        RECT 33.495 162.825 33.715 163.105 ;
        RECT 33.895 162.995 34.435 163.365 ;
        RECT 34.780 163.285 34.950 163.875 ;
        RECT 35.170 163.455 35.475 164.595 ;
        RECT 35.645 163.405 35.900 164.285 ;
        RECT 34.780 163.255 35.520 163.285 ;
        RECT 33.495 162.655 34.025 162.825 ;
        RECT 31.805 162.235 32.155 162.405 ;
        RECT 32.375 162.215 33.325 162.495 ;
        RECT 33.495 162.045 33.685 162.485 ;
        RECT 33.855 162.425 34.025 162.655 ;
        RECT 34.195 162.595 34.435 162.995 ;
        RECT 34.605 162.955 35.520 163.255 ;
        RECT 34.605 162.780 34.930 162.955 ;
        RECT 34.605 162.425 34.925 162.780 ;
        RECT 35.690 162.755 35.900 163.405 ;
        RECT 33.855 162.255 34.925 162.425 ;
        RECT 35.170 162.045 35.475 162.505 ;
        RECT 35.645 162.225 35.900 162.755 ;
        RECT 36.080 163.405 36.335 164.285 ;
        RECT 36.505 163.455 36.810 164.595 ;
        RECT 37.150 164.215 37.480 164.595 ;
        RECT 37.660 164.045 37.830 164.335 ;
        RECT 38.000 164.135 38.250 164.595 ;
        RECT 37.030 163.875 37.830 164.045 ;
        RECT 38.420 164.085 39.290 164.425 ;
        RECT 36.080 162.755 36.290 163.405 ;
        RECT 37.030 163.285 37.200 163.875 ;
        RECT 38.420 163.705 38.590 164.085 ;
        RECT 39.525 163.965 39.695 164.425 ;
        RECT 39.865 164.135 40.235 164.595 ;
        RECT 40.530 163.995 40.700 164.335 ;
        RECT 40.870 164.165 41.200 164.595 ;
        RECT 41.435 163.995 41.605 164.335 ;
        RECT 37.370 163.535 38.590 163.705 ;
        RECT 38.760 163.625 39.220 163.915 ;
        RECT 39.525 163.795 40.085 163.965 ;
        RECT 40.530 163.825 41.605 163.995 ;
        RECT 41.775 164.095 42.455 164.425 ;
        RECT 42.670 164.095 42.920 164.425 ;
        RECT 43.090 164.135 43.340 164.595 ;
        RECT 39.915 163.655 40.085 163.795 ;
        RECT 38.760 163.615 39.725 163.625 ;
        RECT 38.420 163.445 38.590 163.535 ;
        RECT 39.050 163.455 39.725 163.615 ;
        RECT 36.460 163.255 37.200 163.285 ;
        RECT 36.460 162.955 37.375 163.255 ;
        RECT 37.050 162.780 37.375 162.955 ;
        RECT 36.080 162.225 36.335 162.755 ;
        RECT 36.505 162.045 36.810 162.505 ;
        RECT 37.055 162.425 37.375 162.780 ;
        RECT 37.545 162.995 38.085 163.365 ;
        RECT 38.420 163.275 38.825 163.445 ;
        RECT 37.545 162.595 37.785 162.995 ;
        RECT 38.265 162.825 38.485 163.105 ;
        RECT 37.955 162.655 38.485 162.825 ;
        RECT 37.955 162.425 38.125 162.655 ;
        RECT 38.655 162.495 38.825 163.275 ;
        RECT 38.995 162.665 39.345 163.285 ;
        RECT 39.515 162.665 39.725 163.455 ;
        RECT 39.915 163.485 41.415 163.655 ;
        RECT 39.915 162.795 40.085 163.485 ;
        RECT 41.775 163.315 41.945 164.095 ;
        RECT 42.750 163.965 42.920 164.095 ;
        RECT 40.255 163.145 41.945 163.315 ;
        RECT 42.115 163.535 42.580 163.925 ;
        RECT 42.750 163.795 43.145 163.965 ;
        RECT 40.255 162.965 40.425 163.145 ;
        RECT 37.055 162.255 38.125 162.425 ;
        RECT 38.295 162.045 38.485 162.485 ;
        RECT 38.655 162.215 39.605 162.495 ;
        RECT 39.915 162.405 40.175 162.795 ;
        RECT 40.595 162.725 41.385 162.975 ;
        RECT 39.825 162.235 40.175 162.405 ;
        RECT 40.385 162.045 40.715 162.505 ;
        RECT 41.590 162.435 41.760 163.145 ;
        RECT 42.115 162.945 42.285 163.535 ;
        RECT 41.930 162.725 42.285 162.945 ;
        RECT 42.455 162.725 42.805 163.345 ;
        RECT 42.975 162.435 43.145 163.795 ;
        RECT 43.510 163.625 43.835 164.410 ;
        RECT 43.315 162.575 43.775 163.625 ;
        RECT 41.590 162.265 42.445 162.435 ;
        RECT 42.650 162.265 43.145 162.435 ;
        RECT 43.315 162.045 43.645 162.405 ;
        RECT 44.005 162.305 44.175 164.425 ;
        RECT 44.345 164.095 44.675 164.595 ;
        RECT 44.845 163.925 45.100 164.425 ;
        RECT 44.350 163.755 45.100 163.925 ;
        RECT 46.310 163.965 46.595 164.425 ;
        RECT 46.765 164.135 47.035 164.595 ;
        RECT 44.350 162.765 44.580 163.755 ;
        RECT 46.310 163.745 47.265 163.965 ;
        RECT 44.750 162.935 45.100 163.585 ;
        RECT 46.195 163.015 46.885 163.575 ;
        RECT 47.055 162.845 47.265 163.745 ;
        RECT 44.350 162.595 45.100 162.765 ;
        RECT 44.345 162.045 44.675 162.425 ;
        RECT 44.845 162.305 45.100 162.595 ;
        RECT 46.310 162.675 47.265 162.845 ;
        RECT 47.435 163.575 47.835 164.425 ;
        RECT 48.025 163.965 48.305 164.425 ;
        RECT 48.825 164.135 49.150 164.595 ;
        RECT 48.025 163.745 49.150 163.965 ;
        RECT 47.435 163.015 48.530 163.575 ;
        RECT 48.700 163.285 49.150 163.745 ;
        RECT 49.320 163.455 49.705 164.425 ;
        RECT 46.310 162.215 46.595 162.675 ;
        RECT 46.765 162.045 47.035 162.505 ;
        RECT 47.435 162.215 47.835 163.015 ;
        RECT 48.700 162.955 49.255 163.285 ;
        RECT 48.700 162.845 49.150 162.955 ;
        RECT 48.025 162.675 49.150 162.845 ;
        RECT 49.425 162.785 49.705 163.455 ;
        RECT 49.875 163.430 50.165 164.595 ;
        RECT 50.395 163.455 50.605 164.595 ;
        RECT 50.775 163.445 51.105 164.425 ;
        RECT 51.275 163.455 51.505 164.595 ;
        RECT 51.715 163.505 53.385 164.595 ;
        RECT 53.645 163.665 53.815 164.425 ;
        RECT 53.995 163.835 54.325 164.595 ;
        RECT 48.025 162.215 48.305 162.675 ;
        RECT 48.825 162.045 49.150 162.505 ;
        RECT 49.320 162.215 49.705 162.785 ;
        RECT 49.875 162.045 50.165 162.770 ;
        RECT 50.395 162.045 50.605 162.865 ;
        RECT 50.775 162.845 51.025 163.445 ;
        RECT 51.195 163.035 51.525 163.285 ;
        RECT 51.715 162.985 52.465 163.505 ;
        RECT 53.645 163.495 54.310 163.665 ;
        RECT 54.495 163.520 54.765 164.425 ;
        RECT 54.140 163.350 54.310 163.495 ;
        RECT 50.775 162.215 51.105 162.845 ;
        RECT 51.275 162.045 51.505 162.865 ;
        RECT 52.635 162.815 53.385 163.335 ;
        RECT 53.575 162.945 53.905 163.315 ;
        RECT 54.140 163.020 54.425 163.350 ;
        RECT 51.715 162.045 53.385 162.815 ;
        RECT 54.140 162.765 54.310 163.020 ;
        RECT 53.645 162.595 54.310 162.765 ;
        RECT 54.595 162.720 54.765 163.520 ;
        RECT 53.645 162.215 53.815 162.595 ;
        RECT 53.995 162.045 54.325 162.425 ;
        RECT 54.505 162.215 54.765 162.720 ;
        RECT 54.940 163.405 55.195 164.285 ;
        RECT 55.365 163.455 55.670 164.595 ;
        RECT 56.010 164.215 56.340 164.595 ;
        RECT 56.520 164.045 56.690 164.335 ;
        RECT 56.860 164.135 57.110 164.595 ;
        RECT 55.890 163.875 56.690 164.045 ;
        RECT 57.280 164.085 58.150 164.425 ;
        RECT 54.940 162.755 55.150 163.405 ;
        RECT 55.890 163.285 56.060 163.875 ;
        RECT 57.280 163.705 57.450 164.085 ;
        RECT 58.385 163.965 58.555 164.425 ;
        RECT 58.725 164.135 59.095 164.595 ;
        RECT 59.390 163.995 59.560 164.335 ;
        RECT 59.730 164.165 60.060 164.595 ;
        RECT 60.295 163.995 60.465 164.335 ;
        RECT 56.230 163.535 57.450 163.705 ;
        RECT 57.620 163.625 58.080 163.915 ;
        RECT 58.385 163.795 58.945 163.965 ;
        RECT 59.390 163.825 60.465 163.995 ;
        RECT 60.635 164.095 61.315 164.425 ;
        RECT 61.530 164.095 61.780 164.425 ;
        RECT 61.950 164.135 62.200 164.595 ;
        RECT 58.775 163.655 58.945 163.795 ;
        RECT 57.620 163.615 58.585 163.625 ;
        RECT 57.280 163.445 57.450 163.535 ;
        RECT 57.910 163.455 58.585 163.615 ;
        RECT 55.320 163.255 56.060 163.285 ;
        RECT 55.320 162.955 56.235 163.255 ;
        RECT 55.910 162.780 56.235 162.955 ;
        RECT 54.940 162.225 55.195 162.755 ;
        RECT 55.365 162.045 55.670 162.505 ;
        RECT 55.915 162.425 56.235 162.780 ;
        RECT 56.405 162.995 56.945 163.365 ;
        RECT 57.280 163.275 57.685 163.445 ;
        RECT 56.405 162.595 56.645 162.995 ;
        RECT 57.125 162.825 57.345 163.105 ;
        RECT 56.815 162.655 57.345 162.825 ;
        RECT 56.815 162.425 56.985 162.655 ;
        RECT 57.515 162.495 57.685 163.275 ;
        RECT 57.855 162.665 58.205 163.285 ;
        RECT 58.375 162.665 58.585 163.455 ;
        RECT 58.775 163.485 60.275 163.655 ;
        RECT 58.775 162.795 58.945 163.485 ;
        RECT 60.635 163.315 60.805 164.095 ;
        RECT 61.610 163.965 61.780 164.095 ;
        RECT 59.115 163.145 60.805 163.315 ;
        RECT 60.975 163.535 61.440 163.925 ;
        RECT 61.610 163.795 62.005 163.965 ;
        RECT 59.115 162.965 59.285 163.145 ;
        RECT 55.915 162.255 56.985 162.425 ;
        RECT 57.155 162.045 57.345 162.485 ;
        RECT 57.515 162.215 58.465 162.495 ;
        RECT 58.775 162.405 59.035 162.795 ;
        RECT 59.455 162.725 60.245 162.975 ;
        RECT 58.685 162.235 59.035 162.405 ;
        RECT 59.245 162.045 59.575 162.505 ;
        RECT 60.450 162.435 60.620 163.145 ;
        RECT 60.975 162.945 61.145 163.535 ;
        RECT 60.790 162.725 61.145 162.945 ;
        RECT 61.315 162.725 61.665 163.345 ;
        RECT 61.835 162.435 62.005 163.795 ;
        RECT 62.370 163.625 62.695 164.410 ;
        RECT 62.175 162.575 62.635 163.625 ;
        RECT 60.450 162.265 61.305 162.435 ;
        RECT 61.510 162.265 62.005 162.435 ;
        RECT 62.175 162.045 62.505 162.405 ;
        RECT 62.865 162.305 63.035 164.425 ;
        RECT 63.205 164.095 63.535 164.595 ;
        RECT 63.705 163.925 63.960 164.425 ;
        RECT 63.210 163.755 63.960 163.925 ;
        RECT 63.210 162.765 63.440 163.755 ;
        RECT 63.610 162.935 63.960 163.585 ;
        RECT 64.285 163.445 64.615 164.595 ;
        RECT 64.785 163.575 64.955 164.425 ;
        RECT 65.125 163.795 65.455 164.595 ;
        RECT 65.625 163.575 65.795 164.425 ;
        RECT 65.975 163.795 66.215 164.595 ;
        RECT 66.385 163.615 66.715 164.425 ;
        RECT 66.950 163.725 67.235 164.595 ;
        RECT 67.405 163.965 67.665 164.425 ;
        RECT 67.840 164.135 68.095 164.595 ;
        RECT 68.265 163.965 68.525 164.425 ;
        RECT 67.405 163.795 68.525 163.965 ;
        RECT 68.695 163.795 69.005 164.595 ;
        RECT 64.785 163.405 65.795 163.575 ;
        RECT 66.000 163.445 66.715 163.615 ;
        RECT 67.405 163.545 67.665 163.795 ;
        RECT 69.175 163.625 69.485 164.425 ;
        RECT 70.120 164.160 75.465 164.595 ;
        RECT 64.785 162.895 65.280 163.405 ;
        RECT 66.000 163.205 66.170 163.445 ;
        RECT 66.910 163.375 67.665 163.545 ;
        RECT 68.455 163.455 69.485 163.625 ;
        RECT 65.670 163.035 66.170 163.205 ;
        RECT 66.340 163.035 66.720 163.275 ;
        RECT 64.785 162.865 65.285 162.895 ;
        RECT 66.000 162.865 66.170 163.035 ;
        RECT 66.910 162.865 67.315 163.375 ;
        RECT 68.455 163.205 68.625 163.455 ;
        RECT 67.485 163.035 68.625 163.205 ;
        RECT 63.210 162.595 63.960 162.765 ;
        RECT 63.205 162.045 63.535 162.425 ;
        RECT 63.705 162.305 63.960 162.595 ;
        RECT 64.285 162.045 64.615 162.845 ;
        RECT 64.785 162.695 65.795 162.865 ;
        RECT 66.000 162.695 66.635 162.865 ;
        RECT 66.910 162.695 68.560 162.865 ;
        RECT 68.795 162.715 69.145 163.285 ;
        RECT 64.785 162.215 64.955 162.695 ;
        RECT 65.125 162.045 65.455 162.525 ;
        RECT 65.625 162.215 65.795 162.695 ;
        RECT 66.045 162.045 66.285 162.525 ;
        RECT 66.465 162.215 66.635 162.695 ;
        RECT 66.955 162.045 67.235 162.525 ;
        RECT 67.405 162.305 67.665 162.695 ;
        RECT 67.840 162.045 68.095 162.525 ;
        RECT 68.265 162.305 68.560 162.695 ;
        RECT 69.315 162.545 69.485 163.455 ;
        RECT 71.710 162.910 72.060 164.160 ;
        RECT 75.635 163.430 75.925 164.595 ;
        RECT 76.095 163.505 77.765 164.595 ;
        RECT 77.935 163.835 78.450 164.245 ;
        RECT 78.685 163.835 78.855 164.595 ;
        RECT 79.025 164.255 81.055 164.425 ;
        RECT 73.540 162.590 73.880 163.420 ;
        RECT 76.095 162.985 76.845 163.505 ;
        RECT 77.015 162.815 77.765 163.335 ;
        RECT 77.935 163.025 78.275 163.835 ;
        RECT 79.025 163.590 79.195 164.255 ;
        RECT 79.590 163.915 80.715 164.085 ;
        RECT 78.445 163.400 79.195 163.590 ;
        RECT 79.365 163.575 80.375 163.745 ;
        RECT 77.935 162.855 79.165 163.025 ;
        RECT 68.740 162.045 69.015 162.525 ;
        RECT 69.185 162.215 69.485 162.545 ;
        RECT 70.120 162.045 75.465 162.590 ;
        RECT 75.635 162.045 75.925 162.770 ;
        RECT 76.095 162.045 77.765 162.815 ;
        RECT 78.210 162.250 78.455 162.855 ;
        RECT 78.675 162.045 79.185 162.580 ;
        RECT 79.365 162.215 79.555 163.575 ;
        RECT 79.725 162.555 80.000 163.375 ;
        RECT 80.205 162.775 80.375 163.575 ;
        RECT 80.545 162.785 80.715 163.915 ;
        RECT 80.885 163.285 81.055 164.255 ;
        RECT 81.225 163.455 81.395 164.595 ;
        RECT 81.565 163.455 81.900 164.425 ;
        RECT 82.165 163.665 82.335 164.425 ;
        RECT 82.515 163.835 82.845 164.595 ;
        RECT 82.165 163.495 82.830 163.665 ;
        RECT 83.015 163.520 83.285 164.425 ;
        RECT 80.885 162.955 81.080 163.285 ;
        RECT 81.305 162.955 81.560 163.285 ;
        RECT 81.305 162.785 81.475 162.955 ;
        RECT 81.730 162.785 81.900 163.455 ;
        RECT 82.660 163.350 82.830 163.495 ;
        RECT 82.095 162.945 82.425 163.315 ;
        RECT 82.660 163.020 82.945 163.350 ;
        RECT 80.545 162.615 81.475 162.785 ;
        RECT 80.545 162.580 80.720 162.615 ;
        RECT 79.725 162.385 80.005 162.555 ;
        RECT 79.725 162.215 80.000 162.385 ;
        RECT 80.190 162.215 80.720 162.580 ;
        RECT 81.145 162.045 81.475 162.445 ;
        RECT 81.645 162.215 81.900 162.785 ;
        RECT 82.660 162.765 82.830 163.020 ;
        RECT 82.165 162.595 82.830 162.765 ;
        RECT 83.115 162.720 83.285 163.520 ;
        RECT 83.455 163.505 85.125 164.595 ;
        RECT 85.385 163.665 85.555 164.425 ;
        RECT 85.735 163.835 86.065 164.595 ;
        RECT 83.455 162.985 84.205 163.505 ;
        RECT 85.385 163.495 86.050 163.665 ;
        RECT 86.235 163.520 86.505 164.425 ;
        RECT 86.680 164.160 92.025 164.595 ;
        RECT 85.880 163.350 86.050 163.495 ;
        RECT 84.375 162.815 85.125 163.335 ;
        RECT 85.315 162.945 85.645 163.315 ;
        RECT 85.880 163.020 86.165 163.350 ;
        RECT 82.165 162.215 82.335 162.595 ;
        RECT 82.515 162.045 82.845 162.425 ;
        RECT 83.025 162.215 83.285 162.720 ;
        RECT 83.455 162.045 85.125 162.815 ;
        RECT 85.880 162.765 86.050 163.020 ;
        RECT 85.385 162.595 86.050 162.765 ;
        RECT 86.335 162.720 86.505 163.520 ;
        RECT 88.270 162.910 88.620 164.160 ;
        RECT 92.285 163.850 92.555 164.595 ;
        RECT 93.185 164.590 99.460 164.595 ;
        RECT 92.725 163.680 93.015 164.420 ;
        RECT 93.185 163.865 93.440 164.590 ;
        RECT 93.625 163.695 93.885 164.420 ;
        RECT 94.055 163.865 94.300 164.590 ;
        RECT 94.485 163.695 94.745 164.420 ;
        RECT 94.915 163.865 95.160 164.590 ;
        RECT 95.345 163.695 95.605 164.420 ;
        RECT 95.775 163.865 96.020 164.590 ;
        RECT 96.190 163.695 96.450 164.420 ;
        RECT 96.620 163.865 96.880 164.590 ;
        RECT 97.050 163.695 97.310 164.420 ;
        RECT 97.480 163.865 97.740 164.590 ;
        RECT 97.910 163.695 98.170 164.420 ;
        RECT 98.340 163.865 98.600 164.590 ;
        RECT 98.770 163.695 99.030 164.420 ;
        RECT 99.200 163.795 99.460 164.590 ;
        RECT 93.625 163.680 99.030 163.695 ;
        RECT 92.285 163.455 99.030 163.680 ;
        RECT 85.385 162.215 85.555 162.595 ;
        RECT 85.735 162.045 86.065 162.425 ;
        RECT 86.245 162.215 86.505 162.720 ;
        RECT 90.100 162.590 90.440 163.420 ;
        RECT 92.285 162.865 93.450 163.455 ;
        RECT 99.630 163.285 99.880 164.420 ;
        RECT 100.060 163.785 100.320 164.595 ;
        RECT 100.495 163.285 100.740 164.425 ;
        RECT 100.920 163.785 101.215 164.595 ;
        RECT 101.395 163.430 101.685 164.595 ;
        RECT 101.855 163.835 102.370 164.245 ;
        RECT 102.605 163.835 102.775 164.595 ;
        RECT 102.945 164.255 104.975 164.425 ;
        RECT 93.620 163.035 100.740 163.285 ;
        RECT 92.285 162.695 99.030 162.865 ;
        RECT 86.680 162.045 92.025 162.590 ;
        RECT 92.285 162.045 92.585 162.525 ;
        RECT 92.755 162.240 93.015 162.695 ;
        RECT 93.185 162.045 93.445 162.525 ;
        RECT 93.625 162.240 93.885 162.695 ;
        RECT 94.055 162.045 94.305 162.525 ;
        RECT 94.485 162.240 94.745 162.695 ;
        RECT 94.915 162.045 95.165 162.525 ;
        RECT 95.345 162.240 95.605 162.695 ;
        RECT 95.775 162.045 96.020 162.525 ;
        RECT 96.190 162.240 96.465 162.695 ;
        RECT 96.635 162.045 96.880 162.525 ;
        RECT 97.050 162.240 97.310 162.695 ;
        RECT 97.480 162.045 97.740 162.525 ;
        RECT 97.910 162.240 98.170 162.695 ;
        RECT 98.340 162.045 98.600 162.525 ;
        RECT 98.770 162.240 99.030 162.695 ;
        RECT 99.200 162.045 99.460 162.605 ;
        RECT 99.630 162.225 99.880 163.035 ;
        RECT 100.060 162.045 100.320 162.570 ;
        RECT 100.490 162.225 100.740 163.035 ;
        RECT 100.910 162.725 101.225 163.285 ;
        RECT 101.855 163.025 102.195 163.835 ;
        RECT 102.945 163.590 103.115 164.255 ;
        RECT 103.510 163.915 104.635 164.085 ;
        RECT 102.365 163.400 103.115 163.590 ;
        RECT 103.285 163.575 104.295 163.745 ;
        RECT 101.855 162.855 103.085 163.025 ;
        RECT 100.920 162.045 101.225 162.555 ;
        RECT 101.395 162.045 101.685 162.770 ;
        RECT 102.130 162.250 102.375 162.855 ;
        RECT 102.595 162.045 103.105 162.580 ;
        RECT 103.285 162.215 103.475 163.575 ;
        RECT 103.645 162.895 103.920 163.375 ;
        RECT 103.645 162.725 103.925 162.895 ;
        RECT 104.125 162.775 104.295 163.575 ;
        RECT 104.465 162.785 104.635 163.915 ;
        RECT 104.805 163.285 104.975 164.255 ;
        RECT 105.145 163.455 105.315 164.595 ;
        RECT 105.485 163.455 105.820 164.425 ;
        RECT 104.805 162.955 105.000 163.285 ;
        RECT 105.225 162.955 105.480 163.285 ;
        RECT 105.225 162.785 105.395 162.955 ;
        RECT 105.650 162.785 105.820 163.455 ;
        RECT 103.645 162.215 103.920 162.725 ;
        RECT 104.465 162.615 105.395 162.785 ;
        RECT 104.465 162.580 104.640 162.615 ;
        RECT 104.110 162.215 104.640 162.580 ;
        RECT 105.065 162.045 105.395 162.445 ;
        RECT 105.565 162.215 105.820 162.785 ;
        RECT 106.460 163.455 106.795 164.425 ;
        RECT 106.965 163.455 107.135 164.595 ;
        RECT 107.305 164.255 109.335 164.425 ;
        RECT 106.460 162.785 106.630 163.455 ;
        RECT 107.305 163.285 107.475 164.255 ;
        RECT 106.800 162.955 107.055 163.285 ;
        RECT 107.280 162.955 107.475 163.285 ;
        RECT 107.645 163.915 108.770 164.085 ;
        RECT 106.885 162.785 107.055 162.955 ;
        RECT 107.645 162.785 107.815 163.915 ;
        RECT 106.460 162.215 106.715 162.785 ;
        RECT 106.885 162.615 107.815 162.785 ;
        RECT 107.985 163.575 108.995 163.745 ;
        RECT 107.985 162.775 108.155 163.575 ;
        RECT 107.640 162.580 107.815 162.615 ;
        RECT 106.885 162.045 107.215 162.445 ;
        RECT 107.640 162.215 108.170 162.580 ;
        RECT 108.360 162.555 108.635 163.375 ;
        RECT 108.355 162.385 108.635 162.555 ;
        RECT 108.360 162.215 108.635 162.385 ;
        RECT 108.805 162.215 108.995 163.575 ;
        RECT 109.165 163.590 109.335 164.255 ;
        RECT 109.505 163.835 109.675 164.595 ;
        RECT 109.910 163.835 110.425 164.245 ;
        RECT 109.165 163.400 109.915 163.590 ;
        RECT 110.085 163.025 110.425 163.835 ;
        RECT 110.745 163.445 111.075 164.595 ;
        RECT 111.245 163.575 111.415 164.425 ;
        RECT 111.585 163.795 111.915 164.595 ;
        RECT 112.085 163.575 112.255 164.425 ;
        RECT 112.435 163.795 112.675 164.595 ;
        RECT 112.845 163.615 113.175 164.425 ;
        RECT 109.195 162.855 110.425 163.025 ;
        RECT 111.245 163.405 112.255 163.575 ;
        RECT 112.460 163.445 113.175 163.615 ;
        RECT 111.245 162.895 111.740 163.405 ;
        RECT 112.460 163.205 112.630 163.445 ;
        RECT 113.360 163.405 113.615 164.285 ;
        RECT 113.785 163.455 114.090 164.595 ;
        RECT 114.430 164.215 114.760 164.595 ;
        RECT 114.940 164.045 115.110 164.335 ;
        RECT 115.280 164.135 115.530 164.595 ;
        RECT 114.310 163.875 115.110 164.045 ;
        RECT 115.700 164.085 116.570 164.425 ;
        RECT 112.130 163.035 112.630 163.205 ;
        RECT 112.800 163.035 113.180 163.275 ;
        RECT 111.245 162.865 111.745 162.895 ;
        RECT 112.460 162.865 112.630 163.035 ;
        RECT 109.175 162.045 109.685 162.580 ;
        RECT 109.905 162.250 110.150 162.855 ;
        RECT 110.745 162.045 111.075 162.845 ;
        RECT 111.245 162.695 112.255 162.865 ;
        RECT 112.460 162.695 113.095 162.865 ;
        RECT 111.245 162.215 111.415 162.695 ;
        RECT 111.585 162.045 111.915 162.525 ;
        RECT 112.085 162.215 112.255 162.695 ;
        RECT 112.505 162.045 112.745 162.525 ;
        RECT 112.925 162.215 113.095 162.695 ;
        RECT 113.360 162.755 113.570 163.405 ;
        RECT 114.310 163.285 114.480 163.875 ;
        RECT 115.700 163.705 115.870 164.085 ;
        RECT 116.805 163.965 116.975 164.425 ;
        RECT 117.145 164.135 117.515 164.595 ;
        RECT 117.810 163.995 117.980 164.335 ;
        RECT 118.150 164.165 118.480 164.595 ;
        RECT 118.715 163.995 118.885 164.335 ;
        RECT 114.650 163.535 115.870 163.705 ;
        RECT 116.040 163.625 116.500 163.915 ;
        RECT 116.805 163.795 117.365 163.965 ;
        RECT 117.810 163.825 118.885 163.995 ;
        RECT 119.055 164.095 119.735 164.425 ;
        RECT 119.950 164.095 120.200 164.425 ;
        RECT 120.370 164.135 120.620 164.595 ;
        RECT 117.195 163.655 117.365 163.795 ;
        RECT 116.040 163.615 117.005 163.625 ;
        RECT 115.700 163.445 115.870 163.535 ;
        RECT 116.330 163.455 117.005 163.615 ;
        RECT 113.740 163.255 114.480 163.285 ;
        RECT 113.740 162.955 114.655 163.255 ;
        RECT 114.330 162.780 114.655 162.955 ;
        RECT 113.360 162.225 113.615 162.755 ;
        RECT 113.785 162.045 114.090 162.505 ;
        RECT 114.335 162.425 114.655 162.780 ;
        RECT 114.825 162.995 115.365 163.365 ;
        RECT 115.700 163.275 116.105 163.445 ;
        RECT 114.825 162.595 115.065 162.995 ;
        RECT 115.545 162.825 115.765 163.105 ;
        RECT 115.235 162.655 115.765 162.825 ;
        RECT 115.235 162.425 115.405 162.655 ;
        RECT 115.935 162.495 116.105 163.275 ;
        RECT 116.275 162.665 116.625 163.285 ;
        RECT 116.795 162.665 117.005 163.455 ;
        RECT 117.195 163.485 118.695 163.655 ;
        RECT 117.195 162.795 117.365 163.485 ;
        RECT 119.055 163.315 119.225 164.095 ;
        RECT 120.030 163.965 120.200 164.095 ;
        RECT 117.535 163.145 119.225 163.315 ;
        RECT 119.395 163.535 119.860 163.925 ;
        RECT 120.030 163.795 120.425 163.965 ;
        RECT 117.535 162.965 117.705 163.145 ;
        RECT 114.335 162.255 115.405 162.425 ;
        RECT 115.575 162.045 115.765 162.485 ;
        RECT 115.935 162.215 116.885 162.495 ;
        RECT 117.195 162.405 117.455 162.795 ;
        RECT 117.875 162.725 118.665 162.975 ;
        RECT 117.105 162.235 117.455 162.405 ;
        RECT 117.665 162.045 117.995 162.505 ;
        RECT 118.870 162.435 119.040 163.145 ;
        RECT 119.395 162.945 119.565 163.535 ;
        RECT 119.210 162.725 119.565 162.945 ;
        RECT 119.735 162.725 120.085 163.345 ;
        RECT 120.255 162.435 120.425 163.795 ;
        RECT 120.790 163.625 121.115 164.410 ;
        RECT 120.595 162.575 121.055 163.625 ;
        RECT 118.870 162.265 119.725 162.435 ;
        RECT 119.930 162.265 120.425 162.435 ;
        RECT 120.595 162.045 120.925 162.405 ;
        RECT 121.285 162.305 121.455 164.425 ;
        RECT 121.625 164.095 121.955 164.595 ;
        RECT 122.125 163.925 122.380 164.425 ;
        RECT 121.630 163.755 122.380 163.925 ;
        RECT 121.630 162.765 121.860 163.755 ;
        RECT 122.030 162.935 122.380 163.585 ;
        RECT 122.555 163.520 122.825 164.425 ;
        RECT 122.995 163.835 123.325 164.595 ;
        RECT 123.505 163.665 123.675 164.425 ;
        RECT 121.630 162.595 122.380 162.765 ;
        RECT 121.625 162.045 121.955 162.425 ;
        RECT 122.125 162.305 122.380 162.595 ;
        RECT 122.555 162.720 122.725 163.520 ;
        RECT 123.010 163.495 123.675 163.665 ;
        RECT 124.395 163.505 126.065 164.595 ;
        RECT 126.235 163.505 127.445 164.595 ;
        RECT 123.010 163.350 123.180 163.495 ;
        RECT 122.895 163.020 123.180 163.350 ;
        RECT 123.010 162.765 123.180 163.020 ;
        RECT 123.415 162.945 123.745 163.315 ;
        RECT 124.395 162.985 125.145 163.505 ;
        RECT 125.315 162.815 126.065 163.335 ;
        RECT 126.235 162.965 126.755 163.505 ;
        RECT 122.555 162.215 122.815 162.720 ;
        RECT 123.010 162.595 123.675 162.765 ;
        RECT 122.995 162.045 123.325 162.425 ;
        RECT 123.505 162.215 123.675 162.595 ;
        RECT 124.395 162.045 126.065 162.815 ;
        RECT 126.925 162.795 127.445 163.335 ;
        RECT 126.235 162.045 127.445 162.795 ;
        RECT 14.370 161.875 127.530 162.045 ;
        RECT 14.455 161.125 15.665 161.875 ;
        RECT 14.455 160.585 14.975 161.125 ;
        RECT 15.835 161.105 17.505 161.875 ;
        RECT 15.145 160.415 15.665 160.955 ;
        RECT 14.455 159.325 15.665 160.415 ;
        RECT 15.835 160.415 16.585 160.935 ;
        RECT 16.755 160.585 17.505 161.105 ;
        RECT 18.050 161.165 18.305 161.695 ;
        RECT 18.485 161.415 18.770 161.875 ;
        RECT 15.835 159.325 17.505 160.415 ;
        RECT 18.050 160.305 18.230 161.165 ;
        RECT 18.950 160.965 19.200 161.615 ;
        RECT 18.400 160.635 19.200 160.965 ;
        RECT 18.050 159.835 18.305 160.305 ;
        RECT 17.965 159.665 18.305 159.835 ;
        RECT 18.050 159.635 18.305 159.665 ;
        RECT 18.485 159.325 18.770 160.125 ;
        RECT 18.950 160.045 19.200 160.635 ;
        RECT 19.400 161.280 19.720 161.610 ;
        RECT 19.900 161.395 20.560 161.875 ;
        RECT 20.760 161.485 21.610 161.655 ;
        RECT 19.400 160.385 19.590 161.280 ;
        RECT 19.910 160.955 20.570 161.225 ;
        RECT 20.240 160.895 20.570 160.955 ;
        RECT 19.760 160.725 20.090 160.785 ;
        RECT 20.760 160.725 20.930 161.485 ;
        RECT 22.170 161.415 22.490 161.875 ;
        RECT 22.690 161.235 22.940 161.665 ;
        RECT 23.230 161.435 23.640 161.875 ;
        RECT 23.810 161.495 24.825 161.695 ;
        RECT 21.100 161.065 22.350 161.235 ;
        RECT 21.100 160.945 21.430 161.065 ;
        RECT 19.760 160.555 21.660 160.725 ;
        RECT 19.400 160.215 21.320 160.385 ;
        RECT 19.400 160.195 19.720 160.215 ;
        RECT 18.950 159.535 19.280 160.045 ;
        RECT 19.550 159.585 19.720 160.195 ;
        RECT 21.490 160.045 21.660 160.555 ;
        RECT 21.830 160.485 22.010 160.895 ;
        RECT 22.180 160.305 22.350 161.065 ;
        RECT 19.890 159.325 20.220 160.015 ;
        RECT 20.450 159.875 21.660 160.045 ;
        RECT 21.830 159.995 22.350 160.305 ;
        RECT 22.520 160.895 22.940 161.235 ;
        RECT 23.230 160.895 23.640 161.225 ;
        RECT 22.520 160.125 22.710 160.895 ;
        RECT 23.810 160.765 23.980 161.495 ;
        RECT 25.125 161.325 25.295 161.655 ;
        RECT 25.465 161.495 25.795 161.875 ;
        RECT 24.150 160.945 24.500 161.315 ;
        RECT 23.810 160.725 24.230 160.765 ;
        RECT 22.880 160.555 24.230 160.725 ;
        RECT 22.880 160.395 23.130 160.555 ;
        RECT 23.640 160.125 23.890 160.385 ;
        RECT 22.520 159.875 23.890 160.125 ;
        RECT 20.450 159.585 20.690 159.875 ;
        RECT 21.490 159.795 21.660 159.875 ;
        RECT 20.890 159.325 21.310 159.705 ;
        RECT 21.490 159.545 22.120 159.795 ;
        RECT 22.590 159.325 22.920 159.705 ;
        RECT 23.090 159.585 23.260 159.875 ;
        RECT 24.060 159.710 24.230 160.555 ;
        RECT 24.680 160.385 24.900 161.255 ;
        RECT 25.125 161.135 25.820 161.325 ;
        RECT 24.400 160.005 24.900 160.385 ;
        RECT 25.070 160.335 25.480 160.955 ;
        RECT 25.650 160.165 25.820 161.135 ;
        RECT 25.125 159.995 25.820 160.165 ;
        RECT 23.440 159.325 23.820 159.705 ;
        RECT 24.060 159.540 24.890 159.710 ;
        RECT 25.125 159.495 25.295 159.995 ;
        RECT 25.465 159.325 25.795 159.825 ;
        RECT 26.010 159.495 26.235 161.615 ;
        RECT 26.405 161.495 26.735 161.875 ;
        RECT 26.905 161.325 27.075 161.615 ;
        RECT 26.410 161.155 27.075 161.325 ;
        RECT 26.410 160.165 26.640 161.155 ;
        RECT 27.340 161.135 27.595 161.705 ;
        RECT 27.765 161.475 28.095 161.875 ;
        RECT 28.520 161.340 29.050 161.705 ;
        RECT 28.520 161.305 28.695 161.340 ;
        RECT 27.765 161.135 28.695 161.305 ;
        RECT 29.240 161.195 29.515 161.705 ;
        RECT 26.810 160.335 27.160 160.985 ;
        RECT 27.340 160.465 27.510 161.135 ;
        RECT 27.765 160.965 27.935 161.135 ;
        RECT 27.680 160.635 27.935 160.965 ;
        RECT 28.160 160.635 28.355 160.965 ;
        RECT 26.410 159.995 27.075 160.165 ;
        RECT 26.405 159.325 26.735 159.825 ;
        RECT 26.905 159.495 27.075 159.995 ;
        RECT 27.340 159.495 27.675 160.465 ;
        RECT 27.845 159.325 28.015 160.465 ;
        RECT 28.185 159.665 28.355 160.635 ;
        RECT 28.525 160.005 28.695 161.135 ;
        RECT 28.865 160.345 29.035 161.145 ;
        RECT 29.235 161.025 29.515 161.195 ;
        RECT 29.240 160.545 29.515 161.025 ;
        RECT 29.685 160.345 29.875 161.705 ;
        RECT 30.055 161.340 30.565 161.875 ;
        RECT 30.785 161.065 31.030 161.670 ;
        RECT 31.475 161.125 32.685 161.875 ;
        RECT 30.075 160.895 31.305 161.065 ;
        RECT 28.865 160.175 29.875 160.345 ;
        RECT 30.045 160.330 30.795 160.520 ;
        RECT 28.525 159.835 29.650 160.005 ;
        RECT 30.045 159.665 30.215 160.330 ;
        RECT 30.965 160.085 31.305 160.895 ;
        RECT 28.185 159.495 30.215 159.665 ;
        RECT 30.385 159.325 30.555 160.085 ;
        RECT 30.790 159.675 31.305 160.085 ;
        RECT 31.475 160.415 31.995 160.955 ;
        RECT 32.165 160.585 32.685 161.125 ;
        RECT 32.860 161.135 33.115 161.705 ;
        RECT 33.285 161.475 33.615 161.875 ;
        RECT 34.040 161.340 34.570 161.705 ;
        RECT 34.040 161.305 34.215 161.340 ;
        RECT 33.285 161.135 34.215 161.305 ;
        RECT 34.760 161.195 35.035 161.705 ;
        RECT 32.860 160.465 33.030 161.135 ;
        RECT 33.285 160.965 33.455 161.135 ;
        RECT 33.200 160.635 33.455 160.965 ;
        RECT 33.680 160.635 33.875 160.965 ;
        RECT 31.475 159.325 32.685 160.415 ;
        RECT 32.860 159.495 33.195 160.465 ;
        RECT 33.365 159.325 33.535 160.465 ;
        RECT 33.705 159.665 33.875 160.635 ;
        RECT 34.045 160.005 34.215 161.135 ;
        RECT 34.385 160.345 34.555 161.145 ;
        RECT 34.755 161.025 35.035 161.195 ;
        RECT 34.760 160.545 35.035 161.025 ;
        RECT 35.205 160.345 35.395 161.705 ;
        RECT 35.575 161.340 36.085 161.875 ;
        RECT 36.305 161.065 36.550 161.670 ;
        RECT 36.995 161.150 37.285 161.875 ;
        RECT 37.915 161.105 39.585 161.875 ;
        RECT 35.595 160.895 36.825 161.065 ;
        RECT 34.385 160.175 35.395 160.345 ;
        RECT 35.565 160.330 36.315 160.520 ;
        RECT 34.045 159.835 35.170 160.005 ;
        RECT 35.565 159.665 35.735 160.330 ;
        RECT 36.485 160.085 36.825 160.895 ;
        RECT 33.705 159.495 35.735 159.665 ;
        RECT 35.905 159.325 36.075 160.085 ;
        RECT 36.310 159.675 36.825 160.085 ;
        RECT 36.995 159.325 37.285 160.490 ;
        RECT 37.915 160.415 38.665 160.935 ;
        RECT 38.835 160.585 39.585 161.105 ;
        RECT 39.870 161.245 40.155 161.705 ;
        RECT 40.325 161.415 40.595 161.875 ;
        RECT 39.870 161.075 40.825 161.245 ;
        RECT 37.915 159.325 39.585 160.415 ;
        RECT 39.755 160.345 40.445 160.905 ;
        RECT 40.615 160.175 40.825 161.075 ;
        RECT 39.870 159.955 40.825 160.175 ;
        RECT 40.995 160.905 41.395 161.705 ;
        RECT 41.585 161.245 41.865 161.705 ;
        RECT 42.385 161.415 42.710 161.875 ;
        RECT 41.585 161.075 42.710 161.245 ;
        RECT 42.880 161.135 43.265 161.705 ;
        RECT 42.260 160.965 42.710 161.075 ;
        RECT 40.995 160.345 42.090 160.905 ;
        RECT 42.260 160.635 42.815 160.965 ;
        RECT 39.870 159.495 40.155 159.955 ;
        RECT 40.325 159.325 40.595 159.785 ;
        RECT 40.995 159.495 41.395 160.345 ;
        RECT 42.260 160.175 42.710 160.635 ;
        RECT 42.985 160.465 43.265 161.135 ;
        RECT 41.585 159.955 42.710 160.175 ;
        RECT 41.585 159.495 41.865 159.955 ;
        RECT 42.385 159.325 42.710 159.785 ;
        RECT 42.880 159.495 43.265 160.465 ;
        RECT 43.440 161.135 43.695 161.705 ;
        RECT 43.865 161.475 44.195 161.875 ;
        RECT 44.620 161.340 45.150 161.705 ;
        RECT 45.340 161.535 45.615 161.705 ;
        RECT 45.335 161.365 45.615 161.535 ;
        RECT 44.620 161.305 44.795 161.340 ;
        RECT 43.865 161.135 44.795 161.305 ;
        RECT 43.440 160.465 43.610 161.135 ;
        RECT 43.865 160.965 44.035 161.135 ;
        RECT 43.780 160.635 44.035 160.965 ;
        RECT 44.260 160.635 44.455 160.965 ;
        RECT 43.440 159.495 43.775 160.465 ;
        RECT 43.945 159.325 44.115 160.465 ;
        RECT 44.285 159.665 44.455 160.635 ;
        RECT 44.625 160.005 44.795 161.135 ;
        RECT 44.965 160.345 45.135 161.145 ;
        RECT 45.340 160.545 45.615 161.365 ;
        RECT 45.785 160.345 45.975 161.705 ;
        RECT 46.155 161.340 46.665 161.875 ;
        RECT 46.885 161.065 47.130 161.670 ;
        RECT 47.575 161.200 47.835 161.705 ;
        RECT 48.015 161.495 48.345 161.875 ;
        RECT 48.525 161.325 48.695 161.705 ;
        RECT 46.175 160.895 47.405 161.065 ;
        RECT 44.965 160.175 45.975 160.345 ;
        RECT 46.145 160.330 46.895 160.520 ;
        RECT 44.625 159.835 45.750 160.005 ;
        RECT 46.145 159.665 46.315 160.330 ;
        RECT 47.065 160.085 47.405 160.895 ;
        RECT 44.285 159.495 46.315 159.665 ;
        RECT 46.485 159.325 46.655 160.085 ;
        RECT 46.890 159.675 47.405 160.085 ;
        RECT 47.575 160.400 47.745 161.200 ;
        RECT 48.030 161.155 48.695 161.325 ;
        RECT 48.030 160.900 48.200 161.155 ;
        RECT 48.960 161.135 49.215 161.705 ;
        RECT 49.385 161.475 49.715 161.875 ;
        RECT 50.140 161.340 50.670 161.705 ;
        RECT 50.140 161.305 50.315 161.340 ;
        RECT 49.385 161.135 50.315 161.305 ;
        RECT 47.915 160.570 48.200 160.900 ;
        RECT 48.435 160.605 48.765 160.975 ;
        RECT 48.030 160.425 48.200 160.570 ;
        RECT 48.960 160.465 49.130 161.135 ;
        RECT 49.385 160.965 49.555 161.135 ;
        RECT 49.300 160.635 49.555 160.965 ;
        RECT 49.780 160.635 49.975 160.965 ;
        RECT 47.575 159.495 47.845 160.400 ;
        RECT 48.030 160.255 48.695 160.425 ;
        RECT 48.015 159.325 48.345 160.085 ;
        RECT 48.525 159.495 48.695 160.255 ;
        RECT 48.960 159.495 49.295 160.465 ;
        RECT 49.465 159.325 49.635 160.465 ;
        RECT 49.805 159.665 49.975 160.635 ;
        RECT 50.145 160.005 50.315 161.135 ;
        RECT 50.485 160.345 50.655 161.145 ;
        RECT 50.860 160.855 51.135 161.705 ;
        RECT 50.855 160.685 51.135 160.855 ;
        RECT 50.860 160.545 51.135 160.685 ;
        RECT 51.305 160.345 51.495 161.705 ;
        RECT 51.675 161.340 52.185 161.875 ;
        RECT 52.405 161.065 52.650 161.670 ;
        RECT 53.370 161.065 53.615 161.670 ;
        RECT 53.835 161.340 54.345 161.875 ;
        RECT 51.695 160.895 52.925 161.065 ;
        RECT 50.485 160.175 51.495 160.345 ;
        RECT 51.665 160.330 52.415 160.520 ;
        RECT 50.145 159.835 51.270 160.005 ;
        RECT 51.665 159.665 51.835 160.330 ;
        RECT 52.585 160.085 52.925 160.895 ;
        RECT 49.805 159.495 51.835 159.665 ;
        RECT 52.005 159.325 52.175 160.085 ;
        RECT 52.410 159.675 52.925 160.085 ;
        RECT 53.095 160.895 54.325 161.065 ;
        RECT 53.095 160.085 53.435 160.895 ;
        RECT 53.605 160.330 54.355 160.520 ;
        RECT 53.095 159.675 53.610 160.085 ;
        RECT 53.845 159.325 54.015 160.085 ;
        RECT 54.185 159.665 54.355 160.330 ;
        RECT 54.525 160.345 54.715 161.705 ;
        RECT 54.885 161.535 55.160 161.705 ;
        RECT 54.885 161.365 55.165 161.535 ;
        RECT 54.885 160.545 55.160 161.365 ;
        RECT 55.350 161.340 55.880 161.705 ;
        RECT 56.305 161.475 56.635 161.875 ;
        RECT 55.705 161.305 55.880 161.340 ;
        RECT 55.365 160.345 55.535 161.145 ;
        RECT 54.525 160.175 55.535 160.345 ;
        RECT 55.705 161.135 56.635 161.305 ;
        RECT 56.805 161.135 57.060 161.705 ;
        RECT 55.705 160.005 55.875 161.135 ;
        RECT 56.465 160.965 56.635 161.135 ;
        RECT 54.750 159.835 55.875 160.005 ;
        RECT 56.045 160.635 56.240 160.965 ;
        RECT 56.465 160.635 56.720 160.965 ;
        RECT 56.045 159.665 56.215 160.635 ;
        RECT 56.890 160.465 57.060 161.135 ;
        RECT 57.695 161.105 59.365 161.875 ;
        RECT 59.625 161.325 59.795 161.705 ;
        RECT 59.975 161.495 60.305 161.875 ;
        RECT 59.625 161.155 60.290 161.325 ;
        RECT 60.485 161.200 60.745 161.705 ;
        RECT 54.185 159.495 56.215 159.665 ;
        RECT 56.385 159.325 56.555 160.465 ;
        RECT 56.725 159.495 57.060 160.465 ;
        RECT 57.695 160.415 58.445 160.935 ;
        RECT 58.615 160.585 59.365 161.105 ;
        RECT 59.555 160.605 59.885 160.975 ;
        RECT 60.120 160.900 60.290 161.155 ;
        RECT 60.120 160.570 60.405 160.900 ;
        RECT 60.120 160.425 60.290 160.570 ;
        RECT 57.695 159.325 59.365 160.415 ;
        RECT 59.625 160.255 60.290 160.425 ;
        RECT 60.575 160.400 60.745 161.200 ;
        RECT 60.915 161.105 62.585 161.875 ;
        RECT 62.755 161.150 63.045 161.875 ;
        RECT 63.215 161.125 64.425 161.875 ;
        RECT 59.625 159.495 59.795 160.255 ;
        RECT 59.975 159.325 60.305 160.085 ;
        RECT 60.475 159.495 60.745 160.400 ;
        RECT 60.915 160.415 61.665 160.935 ;
        RECT 61.835 160.585 62.585 161.105 ;
        RECT 60.915 159.325 62.585 160.415 ;
        RECT 62.755 159.325 63.045 160.490 ;
        RECT 63.215 160.415 63.735 160.955 ;
        RECT 63.905 160.585 64.425 161.125 ;
        RECT 64.600 161.035 64.860 161.875 ;
        RECT 65.035 161.130 65.290 161.705 ;
        RECT 65.460 161.495 65.790 161.875 ;
        RECT 66.005 161.325 66.175 161.705 ;
        RECT 65.460 161.155 66.175 161.325 ;
        RECT 63.215 159.325 64.425 160.415 ;
        RECT 64.600 159.325 64.860 160.475 ;
        RECT 65.035 160.400 65.205 161.130 ;
        RECT 65.460 160.965 65.630 161.155 ;
        RECT 66.440 161.035 66.700 161.875 ;
        RECT 66.875 161.130 67.130 161.705 ;
        RECT 67.300 161.495 67.630 161.875 ;
        RECT 67.845 161.325 68.015 161.705 ;
        RECT 67.300 161.155 68.015 161.325 ;
        RECT 68.365 161.325 68.535 161.705 ;
        RECT 68.750 161.495 69.080 161.875 ;
        RECT 68.365 161.155 69.080 161.325 ;
        RECT 65.375 160.635 65.630 160.965 ;
        RECT 65.460 160.425 65.630 160.635 ;
        RECT 65.910 160.605 66.265 160.975 ;
        RECT 65.035 159.495 65.290 160.400 ;
        RECT 65.460 160.255 66.175 160.425 ;
        RECT 65.460 159.325 65.790 160.085 ;
        RECT 66.005 159.495 66.175 160.255 ;
        RECT 66.440 159.325 66.700 160.475 ;
        RECT 66.875 160.400 67.045 161.130 ;
        RECT 67.300 160.965 67.470 161.155 ;
        RECT 67.215 160.635 67.470 160.965 ;
        RECT 67.300 160.425 67.470 160.635 ;
        RECT 67.750 160.605 68.105 160.975 ;
        RECT 68.275 160.605 68.630 160.975 ;
        RECT 68.910 160.965 69.080 161.155 ;
        RECT 69.250 161.130 69.505 161.705 ;
        RECT 68.910 160.635 69.165 160.965 ;
        RECT 68.910 160.425 69.080 160.635 ;
        RECT 66.875 159.495 67.130 160.400 ;
        RECT 67.300 160.255 68.015 160.425 ;
        RECT 67.300 159.325 67.630 160.085 ;
        RECT 67.845 159.495 68.015 160.255 ;
        RECT 68.365 160.255 69.080 160.425 ;
        RECT 69.335 160.400 69.505 161.130 ;
        RECT 69.680 161.035 69.940 161.875 ;
        RECT 70.205 161.325 70.375 161.705 ;
        RECT 70.590 161.495 70.920 161.875 ;
        RECT 70.205 161.155 70.920 161.325 ;
        RECT 70.115 160.605 70.470 160.975 ;
        RECT 70.750 160.965 70.920 161.155 ;
        RECT 71.090 161.130 71.345 161.705 ;
        RECT 70.750 160.635 71.005 160.965 ;
        RECT 68.365 159.495 68.535 160.255 ;
        RECT 68.750 159.325 69.080 160.085 ;
        RECT 69.250 159.495 69.505 160.400 ;
        RECT 69.680 159.325 69.940 160.475 ;
        RECT 70.750 160.425 70.920 160.635 ;
        RECT 70.205 160.255 70.920 160.425 ;
        RECT 71.175 160.400 71.345 161.130 ;
        RECT 71.520 161.035 71.780 161.875 ;
        RECT 72.415 161.105 75.005 161.875 ;
        RECT 75.180 161.330 80.525 161.875 ;
        RECT 70.205 159.495 70.375 160.255 ;
        RECT 70.590 159.325 70.920 160.085 ;
        RECT 71.090 159.495 71.345 160.400 ;
        RECT 71.520 159.325 71.780 160.475 ;
        RECT 72.415 160.415 73.625 160.935 ;
        RECT 73.795 160.585 75.005 161.105 ;
        RECT 72.415 159.325 75.005 160.415 ;
        RECT 76.770 159.760 77.120 161.010 ;
        RECT 78.600 160.500 78.940 161.330 ;
        RECT 80.755 161.055 80.965 161.875 ;
        RECT 81.135 161.075 81.465 161.705 ;
        RECT 81.135 160.475 81.385 161.075 ;
        RECT 81.635 161.055 81.865 161.875 ;
        RECT 82.350 161.065 82.595 161.670 ;
        RECT 82.815 161.340 83.325 161.875 ;
        RECT 82.075 160.895 83.305 161.065 ;
        RECT 81.555 160.635 81.885 160.885 ;
        RECT 75.180 159.325 80.525 159.760 ;
        RECT 80.755 159.325 80.965 160.465 ;
        RECT 81.135 159.495 81.465 160.475 ;
        RECT 81.635 159.325 81.865 160.465 ;
        RECT 82.075 160.085 82.415 160.895 ;
        RECT 82.585 160.330 83.335 160.520 ;
        RECT 82.075 159.675 82.590 160.085 ;
        RECT 82.825 159.325 82.995 160.085 ;
        RECT 83.165 159.665 83.335 160.330 ;
        RECT 83.505 160.345 83.695 161.705 ;
        RECT 83.865 161.195 84.140 161.705 ;
        RECT 84.330 161.340 84.860 161.705 ;
        RECT 85.285 161.475 85.615 161.875 ;
        RECT 84.685 161.305 84.860 161.340 ;
        RECT 83.865 161.025 84.145 161.195 ;
        RECT 83.865 160.545 84.140 161.025 ;
        RECT 84.345 160.345 84.515 161.145 ;
        RECT 83.505 160.175 84.515 160.345 ;
        RECT 84.685 161.135 85.615 161.305 ;
        RECT 85.785 161.135 86.040 161.705 ;
        RECT 86.305 161.325 86.475 161.705 ;
        RECT 86.655 161.495 86.985 161.875 ;
        RECT 86.305 161.155 86.970 161.325 ;
        RECT 87.165 161.200 87.425 161.705 ;
        RECT 84.685 160.005 84.855 161.135 ;
        RECT 85.445 160.965 85.615 161.135 ;
        RECT 83.730 159.835 84.855 160.005 ;
        RECT 85.025 160.635 85.220 160.965 ;
        RECT 85.445 160.635 85.700 160.965 ;
        RECT 85.025 159.665 85.195 160.635 ;
        RECT 85.870 160.465 86.040 161.135 ;
        RECT 86.235 160.605 86.565 160.975 ;
        RECT 86.800 160.900 86.970 161.155 ;
        RECT 83.165 159.495 85.195 159.665 ;
        RECT 85.365 159.325 85.535 160.465 ;
        RECT 85.705 159.495 86.040 160.465 ;
        RECT 86.800 160.570 87.085 160.900 ;
        RECT 86.800 160.425 86.970 160.570 ;
        RECT 86.305 160.255 86.970 160.425 ;
        RECT 87.255 160.400 87.425 161.200 ;
        RECT 88.515 161.150 88.805 161.875 ;
        RECT 89.810 161.535 90.065 161.695 ;
        RECT 89.725 161.365 90.065 161.535 ;
        RECT 90.245 161.415 90.530 161.875 ;
        RECT 89.810 161.165 90.065 161.365 ;
        RECT 86.305 159.495 86.475 160.255 ;
        RECT 86.655 159.325 86.985 160.085 ;
        RECT 87.155 159.495 87.425 160.400 ;
        RECT 88.515 159.325 88.805 160.490 ;
        RECT 89.810 160.305 89.990 161.165 ;
        RECT 90.710 160.965 90.960 161.615 ;
        RECT 90.160 160.635 90.960 160.965 ;
        RECT 89.810 159.635 90.065 160.305 ;
        RECT 90.245 159.325 90.530 160.125 ;
        RECT 90.710 160.045 90.960 160.635 ;
        RECT 91.160 161.280 91.480 161.610 ;
        RECT 91.660 161.395 92.320 161.875 ;
        RECT 92.520 161.485 93.370 161.655 ;
        RECT 91.160 160.385 91.350 161.280 ;
        RECT 91.670 160.955 92.330 161.225 ;
        RECT 92.000 160.895 92.330 160.955 ;
        RECT 91.520 160.725 91.850 160.785 ;
        RECT 92.520 160.725 92.690 161.485 ;
        RECT 93.930 161.415 94.250 161.875 ;
        RECT 94.450 161.235 94.700 161.665 ;
        RECT 94.990 161.435 95.400 161.875 ;
        RECT 95.570 161.495 96.585 161.695 ;
        RECT 92.860 161.065 94.110 161.235 ;
        RECT 92.860 160.945 93.190 161.065 ;
        RECT 91.520 160.555 93.420 160.725 ;
        RECT 91.160 160.215 93.080 160.385 ;
        RECT 91.160 160.195 91.480 160.215 ;
        RECT 90.710 159.535 91.040 160.045 ;
        RECT 91.310 159.585 91.480 160.195 ;
        RECT 93.250 160.045 93.420 160.555 ;
        RECT 93.590 160.485 93.770 160.895 ;
        RECT 93.940 160.305 94.110 161.065 ;
        RECT 91.650 159.325 91.980 160.015 ;
        RECT 92.210 159.875 93.420 160.045 ;
        RECT 93.590 159.995 94.110 160.305 ;
        RECT 94.280 160.895 94.700 161.235 ;
        RECT 94.990 160.895 95.400 161.225 ;
        RECT 94.280 160.125 94.470 160.895 ;
        RECT 95.570 160.765 95.740 161.495 ;
        RECT 96.885 161.325 97.055 161.655 ;
        RECT 97.225 161.495 97.555 161.875 ;
        RECT 95.910 160.945 96.260 161.315 ;
        RECT 95.570 160.725 95.990 160.765 ;
        RECT 94.640 160.555 95.990 160.725 ;
        RECT 94.640 160.395 94.890 160.555 ;
        RECT 95.400 160.125 95.650 160.385 ;
        RECT 94.280 159.875 95.650 160.125 ;
        RECT 92.210 159.585 92.450 159.875 ;
        RECT 93.250 159.795 93.420 159.875 ;
        RECT 92.650 159.325 93.070 159.705 ;
        RECT 93.250 159.545 93.880 159.795 ;
        RECT 94.350 159.325 94.680 159.705 ;
        RECT 94.850 159.585 95.020 159.875 ;
        RECT 95.820 159.710 95.990 160.555 ;
        RECT 96.440 160.385 96.660 161.255 ;
        RECT 96.885 161.135 97.580 161.325 ;
        RECT 96.160 160.005 96.660 160.385 ;
        RECT 96.830 160.335 97.240 160.955 ;
        RECT 97.410 160.165 97.580 161.135 ;
        RECT 96.885 159.995 97.580 160.165 ;
        RECT 95.200 159.325 95.580 159.705 ;
        RECT 95.820 159.540 96.650 159.710 ;
        RECT 96.885 159.495 97.055 159.995 ;
        RECT 97.225 159.325 97.555 159.825 ;
        RECT 97.770 159.495 97.995 161.615 ;
        RECT 98.165 161.495 98.495 161.875 ;
        RECT 98.665 161.325 98.835 161.615 ;
        RECT 99.195 161.410 99.445 161.875 ;
        RECT 98.170 161.155 98.835 161.325 ;
        RECT 99.615 161.235 99.785 161.705 ;
        RECT 100.035 161.415 100.205 161.875 ;
        RECT 100.455 161.235 100.625 161.705 ;
        RECT 100.875 161.415 101.045 161.875 ;
        RECT 101.295 161.235 101.465 161.705 ;
        RECT 101.835 161.415 102.100 161.875 ;
        RECT 98.170 160.165 98.400 161.155 ;
        RECT 99.095 161.055 101.465 161.235 ;
        RECT 102.430 161.245 102.715 161.705 ;
        RECT 102.885 161.415 103.155 161.875 ;
        RECT 102.430 161.075 103.385 161.245 ;
        RECT 98.570 160.335 98.920 160.985 ;
        RECT 99.095 160.465 99.445 161.055 ;
        RECT 99.615 160.635 102.125 160.885 ;
        RECT 99.095 160.295 101.545 160.465 ;
        RECT 99.095 160.275 99.865 160.295 ;
        RECT 98.170 159.995 98.835 160.165 ;
        RECT 98.165 159.325 98.495 159.825 ;
        RECT 98.665 159.495 98.835 159.995 ;
        RECT 99.195 159.325 99.365 159.785 ;
        RECT 99.535 159.495 99.865 160.275 ;
        RECT 100.035 159.325 100.205 160.125 ;
        RECT 100.375 159.495 100.705 160.295 ;
        RECT 100.875 159.325 101.045 160.125 ;
        RECT 101.215 159.495 101.545 160.295 ;
        RECT 101.805 159.325 102.100 160.465 ;
        RECT 102.315 160.345 103.005 160.905 ;
        RECT 103.175 160.175 103.385 161.075 ;
        RECT 102.430 159.955 103.385 160.175 ;
        RECT 103.555 160.905 103.955 161.705 ;
        RECT 104.145 161.245 104.425 161.705 ;
        RECT 104.945 161.415 105.270 161.875 ;
        RECT 104.145 161.075 105.270 161.245 ;
        RECT 105.440 161.135 105.825 161.705 ;
        RECT 104.820 160.965 105.270 161.075 ;
        RECT 103.555 160.345 104.650 160.905 ;
        RECT 104.820 160.635 105.375 160.965 ;
        RECT 102.430 159.495 102.715 159.955 ;
        RECT 102.885 159.325 103.155 159.785 ;
        RECT 103.555 159.495 103.955 160.345 ;
        RECT 104.820 160.175 105.270 160.635 ;
        RECT 105.545 160.465 105.825 161.135 ;
        RECT 106.570 161.245 106.855 161.705 ;
        RECT 107.025 161.415 107.295 161.875 ;
        RECT 106.570 161.075 107.525 161.245 ;
        RECT 104.145 159.955 105.270 160.175 ;
        RECT 104.145 159.495 104.425 159.955 ;
        RECT 104.945 159.325 105.270 159.785 ;
        RECT 105.440 159.495 105.825 160.465 ;
        RECT 106.455 160.345 107.145 160.905 ;
        RECT 107.315 160.175 107.525 161.075 ;
        RECT 106.570 159.955 107.525 160.175 ;
        RECT 107.695 160.905 108.095 161.705 ;
        RECT 108.285 161.245 108.565 161.705 ;
        RECT 109.085 161.415 109.410 161.875 ;
        RECT 108.285 161.075 109.410 161.245 ;
        RECT 109.580 161.135 109.965 161.705 ;
        RECT 108.960 160.965 109.410 161.075 ;
        RECT 107.695 160.345 108.790 160.905 ;
        RECT 108.960 160.635 109.515 160.965 ;
        RECT 106.570 159.495 106.855 159.955 ;
        RECT 107.025 159.325 107.295 159.785 ;
        RECT 107.695 159.495 108.095 160.345 ;
        RECT 108.960 160.175 109.410 160.635 ;
        RECT 109.685 160.465 109.965 161.135 ;
        RECT 110.410 161.065 110.655 161.670 ;
        RECT 110.875 161.340 111.385 161.875 ;
        RECT 108.285 159.955 109.410 160.175 ;
        RECT 108.285 159.495 108.565 159.955 ;
        RECT 109.085 159.325 109.410 159.785 ;
        RECT 109.580 159.495 109.965 160.465 ;
        RECT 110.135 160.895 111.365 161.065 ;
        RECT 110.135 160.085 110.475 160.895 ;
        RECT 110.645 160.330 111.395 160.520 ;
        RECT 110.135 159.675 110.650 160.085 ;
        RECT 110.885 159.325 111.055 160.085 ;
        RECT 111.225 159.665 111.395 160.330 ;
        RECT 111.565 160.345 111.755 161.705 ;
        RECT 111.925 160.855 112.200 161.705 ;
        RECT 112.390 161.340 112.920 161.705 ;
        RECT 113.345 161.475 113.675 161.875 ;
        RECT 112.745 161.305 112.920 161.340 ;
        RECT 111.925 160.685 112.205 160.855 ;
        RECT 111.925 160.545 112.200 160.685 ;
        RECT 112.405 160.345 112.575 161.145 ;
        RECT 111.565 160.175 112.575 160.345 ;
        RECT 112.745 161.135 113.675 161.305 ;
        RECT 113.845 161.135 114.100 161.705 ;
        RECT 114.275 161.150 114.565 161.875 ;
        RECT 112.745 160.005 112.915 161.135 ;
        RECT 113.505 160.965 113.675 161.135 ;
        RECT 111.790 159.835 112.915 160.005 ;
        RECT 113.085 160.635 113.280 160.965 ;
        RECT 113.505 160.635 113.760 160.965 ;
        RECT 113.085 159.665 113.255 160.635 ;
        RECT 113.930 160.465 114.100 161.135 ;
        RECT 115.010 161.065 115.255 161.670 ;
        RECT 115.475 161.340 115.985 161.875 ;
        RECT 114.735 160.895 115.965 161.065 ;
        RECT 111.225 159.495 113.255 159.665 ;
        RECT 113.425 159.325 113.595 160.465 ;
        RECT 113.765 159.495 114.100 160.465 ;
        RECT 114.275 159.325 114.565 160.490 ;
        RECT 114.735 160.085 115.075 160.895 ;
        RECT 115.245 160.330 115.995 160.520 ;
        RECT 114.735 159.675 115.250 160.085 ;
        RECT 115.485 159.325 115.655 160.085 ;
        RECT 115.825 159.665 115.995 160.330 ;
        RECT 116.165 160.345 116.355 161.705 ;
        RECT 116.525 161.535 116.800 161.705 ;
        RECT 116.525 161.365 116.805 161.535 ;
        RECT 116.525 160.545 116.800 161.365 ;
        RECT 116.990 161.340 117.520 161.705 ;
        RECT 117.945 161.475 118.275 161.875 ;
        RECT 117.345 161.305 117.520 161.340 ;
        RECT 117.005 160.345 117.175 161.145 ;
        RECT 116.165 160.175 117.175 160.345 ;
        RECT 117.345 161.135 118.275 161.305 ;
        RECT 118.445 161.135 118.700 161.705 ;
        RECT 117.345 160.005 117.515 161.135 ;
        RECT 118.105 160.965 118.275 161.135 ;
        RECT 116.390 159.835 117.515 160.005 ;
        RECT 117.685 160.635 117.880 160.965 ;
        RECT 118.105 160.635 118.360 160.965 ;
        RECT 117.685 159.665 117.855 160.635 ;
        RECT 118.530 160.465 118.700 161.135 ;
        RECT 118.915 161.055 119.145 161.875 ;
        RECT 119.315 161.075 119.645 161.705 ;
        RECT 118.895 160.635 119.225 160.885 ;
        RECT 119.395 160.475 119.645 161.075 ;
        RECT 119.815 161.055 120.025 161.875 ;
        RECT 120.805 161.325 120.975 161.705 ;
        RECT 121.155 161.495 121.485 161.875 ;
        RECT 120.805 161.155 121.470 161.325 ;
        RECT 121.665 161.200 121.925 161.705 ;
        RECT 120.735 160.605 121.065 160.975 ;
        RECT 121.300 160.900 121.470 161.155 ;
        RECT 115.825 159.495 117.855 159.665 ;
        RECT 118.025 159.325 118.195 160.465 ;
        RECT 118.365 159.495 118.700 160.465 ;
        RECT 118.915 159.325 119.145 160.465 ;
        RECT 119.315 159.495 119.645 160.475 ;
        RECT 121.300 160.570 121.585 160.900 ;
        RECT 119.815 159.325 120.025 160.465 ;
        RECT 121.300 160.425 121.470 160.570 ;
        RECT 120.805 160.255 121.470 160.425 ;
        RECT 121.755 160.400 121.925 161.200 ;
        RECT 122.555 161.105 126.065 161.875 ;
        RECT 126.235 161.125 127.445 161.875 ;
        RECT 120.805 159.495 120.975 160.255 ;
        RECT 121.155 159.325 121.485 160.085 ;
        RECT 121.655 159.495 121.925 160.400 ;
        RECT 122.555 160.415 124.245 160.935 ;
        RECT 124.415 160.585 126.065 161.105 ;
        RECT 126.235 160.415 126.755 160.955 ;
        RECT 126.925 160.585 127.445 161.125 ;
        RECT 122.555 159.325 126.065 160.415 ;
        RECT 126.235 159.325 127.445 160.415 ;
        RECT 14.370 159.155 127.530 159.325 ;
        RECT 14.455 158.065 15.665 159.155 ;
        RECT 14.455 157.355 14.975 157.895 ;
        RECT 15.145 157.525 15.665 158.065 ;
        RECT 15.835 158.065 17.045 159.155 ;
        RECT 15.835 157.525 16.355 158.065 ;
        RECT 17.275 158.015 17.485 159.155 ;
        RECT 17.655 158.005 17.985 158.985 ;
        RECT 18.155 158.015 18.385 159.155 ;
        RECT 18.635 158.015 18.865 159.155 ;
        RECT 19.035 158.005 19.365 158.985 ;
        RECT 19.535 158.015 19.745 159.155 ;
        RECT 19.975 158.395 20.490 158.805 ;
        RECT 20.725 158.395 20.895 159.155 ;
        RECT 21.065 158.815 23.095 158.985 ;
        RECT 16.525 157.355 17.045 157.895 ;
        RECT 14.455 156.605 15.665 157.355 ;
        RECT 15.835 156.605 17.045 157.355 ;
        RECT 17.275 156.605 17.485 157.425 ;
        RECT 17.655 157.405 17.905 158.005 ;
        RECT 18.075 157.595 18.405 157.845 ;
        RECT 18.615 157.595 18.945 157.845 ;
        RECT 17.655 156.775 17.985 157.405 ;
        RECT 18.155 156.605 18.385 157.425 ;
        RECT 18.635 156.605 18.865 157.425 ;
        RECT 19.115 157.405 19.365 158.005 ;
        RECT 19.975 157.585 20.315 158.395 ;
        RECT 21.065 158.150 21.235 158.815 ;
        RECT 21.630 158.475 22.755 158.645 ;
        RECT 20.485 157.960 21.235 158.150 ;
        RECT 21.405 158.135 22.415 158.305 ;
        RECT 19.035 156.775 19.365 157.405 ;
        RECT 19.535 156.605 19.745 157.425 ;
        RECT 19.975 157.415 21.205 157.585 ;
        RECT 20.250 156.810 20.495 157.415 ;
        RECT 20.715 156.605 21.225 157.140 ;
        RECT 21.405 156.775 21.595 158.135 ;
        RECT 21.765 157.115 22.040 157.935 ;
        RECT 22.245 157.335 22.415 158.135 ;
        RECT 22.585 157.345 22.755 158.475 ;
        RECT 22.925 157.845 23.095 158.815 ;
        RECT 23.265 158.015 23.435 159.155 ;
        RECT 23.605 158.015 23.940 158.985 ;
        RECT 22.925 157.515 23.120 157.845 ;
        RECT 23.345 157.515 23.600 157.845 ;
        RECT 23.345 157.345 23.515 157.515 ;
        RECT 23.770 157.345 23.940 158.015 ;
        RECT 24.115 157.990 24.405 159.155 ;
        RECT 24.665 158.225 24.835 158.985 ;
        RECT 25.015 158.395 25.345 159.155 ;
        RECT 24.665 158.055 25.330 158.225 ;
        RECT 25.515 158.080 25.785 158.985 ;
        RECT 25.160 157.910 25.330 158.055 ;
        RECT 24.595 157.505 24.925 157.875 ;
        RECT 25.160 157.580 25.445 157.910 ;
        RECT 22.585 157.175 23.515 157.345 ;
        RECT 22.585 157.140 22.760 157.175 ;
        RECT 21.765 156.945 22.045 157.115 ;
        RECT 21.765 156.775 22.040 156.945 ;
        RECT 22.230 156.775 22.760 157.140 ;
        RECT 23.185 156.605 23.515 157.005 ;
        RECT 23.685 156.775 23.940 157.345 ;
        RECT 24.115 156.605 24.405 157.330 ;
        RECT 25.160 157.325 25.330 157.580 ;
        RECT 24.665 157.155 25.330 157.325 ;
        RECT 25.615 157.280 25.785 158.080 ;
        RECT 25.955 158.065 27.625 159.155 ;
        RECT 27.910 158.525 28.195 158.985 ;
        RECT 28.365 158.695 28.635 159.155 ;
        RECT 27.910 158.305 28.865 158.525 ;
        RECT 25.955 157.545 26.705 158.065 ;
        RECT 26.875 157.375 27.625 157.895 ;
        RECT 27.795 157.575 28.485 158.135 ;
        RECT 28.655 157.405 28.865 158.305 ;
        RECT 24.665 156.775 24.835 157.155 ;
        RECT 25.015 156.605 25.345 156.985 ;
        RECT 25.525 156.775 25.785 157.280 ;
        RECT 25.955 156.605 27.625 157.375 ;
        RECT 27.910 157.235 28.865 157.405 ;
        RECT 29.035 158.135 29.435 158.985 ;
        RECT 29.625 158.525 29.905 158.985 ;
        RECT 30.425 158.695 30.750 159.155 ;
        RECT 29.625 158.305 30.750 158.525 ;
        RECT 29.035 157.575 30.130 158.135 ;
        RECT 30.300 157.845 30.750 158.305 ;
        RECT 30.920 158.015 31.305 158.985 ;
        RECT 31.590 158.525 31.875 158.985 ;
        RECT 32.045 158.695 32.315 159.155 ;
        RECT 31.590 158.305 32.545 158.525 ;
        RECT 27.910 156.775 28.195 157.235 ;
        RECT 28.365 156.605 28.635 157.065 ;
        RECT 29.035 156.775 29.435 157.575 ;
        RECT 30.300 157.515 30.855 157.845 ;
        RECT 30.300 157.405 30.750 157.515 ;
        RECT 29.625 157.235 30.750 157.405 ;
        RECT 31.025 157.345 31.305 158.015 ;
        RECT 31.475 157.575 32.165 158.135 ;
        RECT 32.335 157.405 32.545 158.305 ;
        RECT 29.625 156.775 29.905 157.235 ;
        RECT 30.425 156.605 30.750 157.065 ;
        RECT 30.920 156.775 31.305 157.345 ;
        RECT 31.590 157.235 32.545 157.405 ;
        RECT 32.715 158.135 33.115 158.985 ;
        RECT 33.305 158.525 33.585 158.985 ;
        RECT 34.105 158.695 34.430 159.155 ;
        RECT 33.305 158.305 34.430 158.525 ;
        RECT 32.715 157.575 33.810 158.135 ;
        RECT 33.980 157.845 34.430 158.305 ;
        RECT 34.600 158.015 34.985 158.985 ;
        RECT 31.590 156.775 31.875 157.235 ;
        RECT 32.045 156.605 32.315 157.065 ;
        RECT 32.715 156.775 33.115 157.575 ;
        RECT 33.980 157.515 34.535 157.845 ;
        RECT 33.980 157.405 34.430 157.515 ;
        RECT 33.305 157.235 34.430 157.405 ;
        RECT 34.705 157.345 34.985 158.015 ;
        RECT 35.155 158.065 38.665 159.155 ;
        RECT 39.040 158.185 39.370 158.985 ;
        RECT 39.540 158.355 39.870 159.155 ;
        RECT 40.170 158.185 40.500 158.985 ;
        RECT 41.145 158.355 41.395 159.155 ;
        RECT 35.155 157.545 36.845 158.065 ;
        RECT 39.040 158.015 41.475 158.185 ;
        RECT 41.665 158.015 41.835 159.155 ;
        RECT 42.005 158.015 42.345 158.985 ;
        RECT 42.720 158.185 43.050 158.985 ;
        RECT 43.220 158.355 43.550 159.155 ;
        RECT 43.850 158.185 44.180 158.985 ;
        RECT 44.825 158.355 45.075 159.155 ;
        RECT 42.720 158.015 45.155 158.185 ;
        RECT 45.345 158.015 45.515 159.155 ;
        RECT 45.685 158.015 46.025 158.985 ;
        RECT 46.310 158.525 46.595 158.985 ;
        RECT 46.765 158.695 47.035 159.155 ;
        RECT 46.310 158.305 47.265 158.525 ;
        RECT 37.015 157.375 38.665 157.895 ;
        RECT 38.835 157.595 39.185 157.845 ;
        RECT 39.370 157.385 39.540 158.015 ;
        RECT 39.710 157.595 40.040 157.795 ;
        RECT 40.210 157.595 40.540 157.795 ;
        RECT 40.710 157.595 41.130 157.795 ;
        RECT 41.305 157.765 41.475 158.015 ;
        RECT 41.305 157.595 42.000 157.765 ;
        RECT 33.305 156.775 33.585 157.235 ;
        RECT 34.105 156.605 34.430 157.065 ;
        RECT 34.600 156.775 34.985 157.345 ;
        RECT 35.155 156.605 38.665 157.375 ;
        RECT 39.040 156.775 39.540 157.385 ;
        RECT 40.170 157.255 41.395 157.425 ;
        RECT 42.170 157.405 42.345 158.015 ;
        RECT 42.515 157.595 42.865 157.845 ;
        RECT 40.170 156.775 40.500 157.255 ;
        RECT 40.670 156.605 40.895 157.065 ;
        RECT 41.065 156.775 41.395 157.255 ;
        RECT 41.585 156.605 41.835 157.405 ;
        RECT 42.005 156.775 42.345 157.405 ;
        RECT 43.050 157.385 43.220 158.015 ;
        RECT 43.390 157.595 43.720 157.795 ;
        RECT 43.890 157.595 44.220 157.795 ;
        RECT 44.390 157.595 44.810 157.795 ;
        RECT 44.985 157.765 45.155 158.015 ;
        RECT 44.985 157.595 45.680 157.765 ;
        RECT 42.720 156.775 43.220 157.385 ;
        RECT 43.850 157.255 45.075 157.425 ;
        RECT 45.850 157.405 46.025 158.015 ;
        RECT 46.195 157.575 46.885 158.135 ;
        RECT 47.055 157.405 47.265 158.305 ;
        RECT 43.850 156.775 44.180 157.255 ;
        RECT 44.350 156.605 44.575 157.065 ;
        RECT 44.745 156.775 45.075 157.255 ;
        RECT 45.265 156.605 45.515 157.405 ;
        RECT 45.685 156.775 46.025 157.405 ;
        RECT 46.310 157.235 47.265 157.405 ;
        RECT 47.435 158.135 47.835 158.985 ;
        RECT 48.025 158.525 48.305 158.985 ;
        RECT 48.825 158.695 49.150 159.155 ;
        RECT 48.025 158.305 49.150 158.525 ;
        RECT 47.435 157.575 48.530 158.135 ;
        RECT 48.700 157.845 49.150 158.305 ;
        RECT 49.320 158.015 49.705 158.985 ;
        RECT 46.310 156.775 46.595 157.235 ;
        RECT 46.765 156.605 47.035 157.065 ;
        RECT 47.435 156.775 47.835 157.575 ;
        RECT 48.700 157.515 49.255 157.845 ;
        RECT 48.700 157.405 49.150 157.515 ;
        RECT 48.025 157.235 49.150 157.405 ;
        RECT 49.425 157.345 49.705 158.015 ;
        RECT 49.875 157.990 50.165 159.155 ;
        RECT 50.335 158.015 50.675 158.985 ;
        RECT 50.845 158.015 51.015 159.155 ;
        RECT 51.285 158.355 51.535 159.155 ;
        RECT 52.180 158.185 52.510 158.985 ;
        RECT 52.810 158.355 53.140 159.155 ;
        RECT 53.310 158.185 53.640 158.985 ;
        RECT 54.480 158.720 59.825 159.155 ;
        RECT 51.205 158.015 53.640 158.185 ;
        RECT 48.025 156.775 48.305 157.235 ;
        RECT 48.825 156.605 49.150 157.065 ;
        RECT 49.320 156.775 49.705 157.345 ;
        RECT 50.335 157.405 50.510 158.015 ;
        RECT 51.205 157.765 51.375 158.015 ;
        RECT 50.680 157.595 51.375 157.765 ;
        RECT 51.550 157.595 51.970 157.795 ;
        RECT 52.140 157.595 52.470 157.795 ;
        RECT 52.640 157.595 52.970 157.795 ;
        RECT 49.875 156.605 50.165 157.330 ;
        RECT 50.335 156.775 50.675 157.405 ;
        RECT 50.845 156.605 51.095 157.405 ;
        RECT 51.285 157.255 52.510 157.425 ;
        RECT 51.285 156.775 51.615 157.255 ;
        RECT 51.785 156.605 52.010 157.065 ;
        RECT 52.180 156.775 52.510 157.255 ;
        RECT 53.140 157.385 53.310 158.015 ;
        RECT 53.495 157.595 53.845 157.845 ;
        RECT 56.070 157.470 56.420 158.720 ;
        RECT 60.055 158.015 60.265 159.155 ;
        RECT 60.435 158.005 60.765 158.985 ;
        RECT 60.935 158.015 61.165 159.155 ;
        RECT 61.525 158.005 61.855 159.155 ;
        RECT 62.025 158.135 62.195 158.985 ;
        RECT 62.365 158.355 62.695 159.155 ;
        RECT 62.865 158.135 63.035 158.985 ;
        RECT 63.215 158.355 63.455 159.155 ;
        RECT 63.625 158.175 63.955 158.985 ;
        RECT 53.140 156.775 53.640 157.385 ;
        RECT 57.900 157.150 58.240 157.980 ;
        RECT 54.480 156.605 59.825 157.150 ;
        RECT 60.055 156.605 60.265 157.425 ;
        RECT 60.435 157.405 60.685 158.005 ;
        RECT 62.025 157.965 63.035 158.135 ;
        RECT 63.240 158.005 63.955 158.175 ;
        RECT 64.595 158.065 68.105 159.155 ;
        RECT 68.365 158.225 68.535 158.985 ;
        RECT 68.750 158.395 69.080 159.155 ;
        RECT 60.855 157.595 61.185 157.845 ;
        RECT 62.025 157.795 62.520 157.965 ;
        RECT 62.025 157.625 62.525 157.795 ;
        RECT 63.240 157.765 63.410 158.005 ;
        RECT 62.025 157.425 62.520 157.625 ;
        RECT 62.910 157.595 63.410 157.765 ;
        RECT 63.580 157.595 63.960 157.835 ;
        RECT 63.240 157.425 63.410 157.595 ;
        RECT 64.595 157.545 66.285 158.065 ;
        RECT 68.365 158.055 69.080 158.225 ;
        RECT 69.250 158.080 69.505 158.985 ;
        RECT 60.435 156.775 60.765 157.405 ;
        RECT 60.935 156.605 61.165 157.425 ;
        RECT 61.525 156.605 61.855 157.405 ;
        RECT 62.025 157.255 63.035 157.425 ;
        RECT 63.240 157.255 63.875 157.425 ;
        RECT 66.455 157.375 68.105 157.895 ;
        RECT 68.275 157.505 68.630 157.875 ;
        RECT 68.910 157.845 69.080 158.055 ;
        RECT 68.910 157.515 69.165 157.845 ;
        RECT 62.025 156.775 62.195 157.255 ;
        RECT 62.365 156.605 62.695 157.085 ;
        RECT 62.865 156.775 63.035 157.255 ;
        RECT 63.285 156.605 63.525 157.085 ;
        RECT 63.705 156.775 63.875 157.255 ;
        RECT 64.595 156.605 68.105 157.375 ;
        RECT 68.910 157.325 69.080 157.515 ;
        RECT 69.335 157.350 69.505 158.080 ;
        RECT 69.680 158.005 69.940 159.155 ;
        RECT 70.205 158.225 70.375 158.985 ;
        RECT 70.590 158.395 70.920 159.155 ;
        RECT 70.205 158.055 70.920 158.225 ;
        RECT 71.090 158.080 71.345 158.985 ;
        RECT 70.115 157.505 70.470 157.875 ;
        RECT 70.750 157.845 70.920 158.055 ;
        RECT 70.750 157.515 71.005 157.845 ;
        RECT 68.365 157.155 69.080 157.325 ;
        RECT 68.365 156.775 68.535 157.155 ;
        RECT 68.750 156.605 69.080 156.985 ;
        RECT 69.250 156.775 69.505 157.350 ;
        RECT 69.680 156.605 69.940 157.445 ;
        RECT 70.750 157.325 70.920 157.515 ;
        RECT 71.175 157.350 71.345 158.080 ;
        RECT 71.520 158.005 71.780 159.155 ;
        RECT 72.160 158.185 72.490 158.985 ;
        RECT 72.660 158.355 72.990 159.155 ;
        RECT 73.290 158.185 73.620 158.985 ;
        RECT 74.265 158.355 74.515 159.155 ;
        RECT 72.160 158.015 74.595 158.185 ;
        RECT 74.785 158.015 74.955 159.155 ;
        RECT 75.125 158.015 75.465 158.985 ;
        RECT 71.955 157.595 72.305 157.845 ;
        RECT 70.205 157.155 70.920 157.325 ;
        RECT 70.205 156.775 70.375 157.155 ;
        RECT 70.590 156.605 70.920 156.985 ;
        RECT 71.090 156.775 71.345 157.350 ;
        RECT 71.520 156.605 71.780 157.445 ;
        RECT 72.490 157.385 72.660 158.015 ;
        RECT 72.830 157.595 73.160 157.795 ;
        RECT 73.330 157.595 73.660 157.795 ;
        RECT 73.830 157.595 74.250 157.795 ;
        RECT 74.425 157.765 74.595 158.015 ;
        RECT 74.425 157.595 75.120 157.765 ;
        RECT 72.160 156.775 72.660 157.385 ;
        RECT 73.290 157.255 74.515 157.425 ;
        RECT 75.290 157.405 75.465 158.015 ;
        RECT 75.635 157.990 75.925 159.155 ;
        RECT 76.760 158.185 77.090 158.985 ;
        RECT 77.260 158.355 77.590 159.155 ;
        RECT 77.890 158.185 78.220 158.985 ;
        RECT 78.865 158.355 79.115 159.155 ;
        RECT 76.760 158.015 79.195 158.185 ;
        RECT 79.385 158.015 79.555 159.155 ;
        RECT 79.725 158.015 80.065 158.985 ;
        RECT 81.070 158.815 81.325 158.845 ;
        RECT 80.985 158.645 81.325 158.815 ;
        RECT 76.555 157.595 76.905 157.845 ;
        RECT 73.290 156.775 73.620 157.255 ;
        RECT 73.790 156.605 74.015 157.065 ;
        RECT 74.185 156.775 74.515 157.255 ;
        RECT 74.705 156.605 74.955 157.405 ;
        RECT 75.125 156.775 75.465 157.405 ;
        RECT 77.090 157.385 77.260 158.015 ;
        RECT 77.430 157.595 77.760 157.795 ;
        RECT 77.930 157.595 78.260 157.795 ;
        RECT 78.430 157.595 78.850 157.795 ;
        RECT 79.025 157.765 79.195 158.015 ;
        RECT 79.025 157.595 79.720 157.765 ;
        RECT 75.635 156.605 75.925 157.330 ;
        RECT 76.760 156.775 77.260 157.385 ;
        RECT 77.890 157.255 79.115 157.425 ;
        RECT 79.890 157.405 80.065 158.015 ;
        RECT 77.890 156.775 78.220 157.255 ;
        RECT 78.390 156.605 78.615 157.065 ;
        RECT 78.785 156.775 79.115 157.255 ;
        RECT 79.305 156.605 79.555 157.405 ;
        RECT 79.725 156.775 80.065 157.405 ;
        RECT 81.070 158.175 81.325 158.645 ;
        RECT 81.505 158.355 81.790 159.155 ;
        RECT 81.970 158.435 82.300 158.945 ;
        RECT 81.070 157.315 81.250 158.175 ;
        RECT 81.970 157.845 82.220 158.435 ;
        RECT 82.570 158.285 82.740 158.895 ;
        RECT 82.910 158.465 83.240 159.155 ;
        RECT 83.470 158.605 83.710 158.895 ;
        RECT 83.910 158.775 84.330 159.155 ;
        RECT 84.510 158.685 85.140 158.935 ;
        RECT 85.610 158.775 85.940 159.155 ;
        RECT 84.510 158.605 84.680 158.685 ;
        RECT 86.110 158.605 86.280 158.895 ;
        RECT 86.460 158.775 86.840 159.155 ;
        RECT 87.080 158.770 87.910 158.940 ;
        RECT 83.470 158.435 84.680 158.605 ;
        RECT 81.420 157.515 82.220 157.845 ;
        RECT 81.070 156.785 81.325 157.315 ;
        RECT 81.505 156.605 81.790 157.065 ;
        RECT 81.970 156.865 82.220 157.515 ;
        RECT 82.420 158.265 82.740 158.285 ;
        RECT 82.420 158.095 84.340 158.265 ;
        RECT 82.420 157.200 82.610 158.095 ;
        RECT 84.510 157.925 84.680 158.435 ;
        RECT 84.850 158.175 85.370 158.485 ;
        RECT 82.780 157.755 84.680 157.925 ;
        RECT 82.780 157.695 83.110 157.755 ;
        RECT 83.260 157.525 83.590 157.585 ;
        RECT 82.930 157.255 83.590 157.525 ;
        RECT 82.420 156.870 82.740 157.200 ;
        RECT 82.920 156.605 83.580 157.085 ;
        RECT 83.780 156.995 83.950 157.755 ;
        RECT 84.850 157.585 85.030 157.995 ;
        RECT 84.120 157.415 84.450 157.535 ;
        RECT 85.200 157.415 85.370 158.175 ;
        RECT 84.120 157.245 85.370 157.415 ;
        RECT 85.540 158.355 86.910 158.605 ;
        RECT 85.540 157.585 85.730 158.355 ;
        RECT 86.660 158.095 86.910 158.355 ;
        RECT 85.900 157.925 86.150 158.085 ;
        RECT 87.080 157.925 87.250 158.770 ;
        RECT 88.145 158.485 88.315 158.985 ;
        RECT 88.485 158.655 88.815 159.155 ;
        RECT 87.420 158.095 87.920 158.475 ;
        RECT 88.145 158.315 88.840 158.485 ;
        RECT 85.900 157.755 87.250 157.925 ;
        RECT 86.830 157.715 87.250 157.755 ;
        RECT 85.540 157.245 85.960 157.585 ;
        RECT 86.250 157.255 86.660 157.585 ;
        RECT 83.780 156.825 84.630 156.995 ;
        RECT 85.190 156.605 85.510 157.065 ;
        RECT 85.710 156.815 85.960 157.245 ;
        RECT 86.250 156.605 86.660 157.045 ;
        RECT 86.830 156.985 87.000 157.715 ;
        RECT 87.170 157.165 87.520 157.535 ;
        RECT 87.700 157.225 87.920 158.095 ;
        RECT 88.090 157.525 88.500 158.145 ;
        RECT 88.670 157.345 88.840 158.315 ;
        RECT 88.145 157.155 88.840 157.345 ;
        RECT 86.830 156.785 87.845 156.985 ;
        RECT 88.145 156.825 88.315 157.155 ;
        RECT 88.485 156.605 88.815 156.985 ;
        RECT 89.030 156.865 89.255 158.985 ;
        RECT 89.425 158.655 89.755 159.155 ;
        RECT 89.925 158.485 90.095 158.985 ;
        RECT 89.430 158.315 90.095 158.485 ;
        RECT 89.430 157.325 89.660 158.315 ;
        RECT 89.830 157.495 90.180 158.145 ;
        RECT 90.815 158.065 92.485 159.155 ;
        RECT 90.815 157.545 91.565 158.065 ;
        RECT 92.695 158.015 92.925 159.155 ;
        RECT 93.095 158.005 93.425 158.985 ;
        RECT 93.595 158.015 93.805 159.155 ;
        RECT 94.495 158.065 96.165 159.155 ;
        RECT 96.425 158.225 96.595 158.985 ;
        RECT 96.775 158.395 97.105 159.155 ;
        RECT 91.735 157.375 92.485 157.895 ;
        RECT 92.675 157.595 93.005 157.845 ;
        RECT 89.430 157.155 90.095 157.325 ;
        RECT 89.425 156.605 89.755 156.985 ;
        RECT 89.925 156.865 90.095 157.155 ;
        RECT 90.815 156.605 92.485 157.375 ;
        RECT 92.695 156.605 92.925 157.425 ;
        RECT 93.175 157.405 93.425 158.005 ;
        RECT 94.495 157.545 95.245 158.065 ;
        RECT 96.425 158.055 97.090 158.225 ;
        RECT 97.275 158.080 97.545 158.985 ;
        RECT 96.920 157.910 97.090 158.055 ;
        RECT 93.095 156.775 93.425 157.405 ;
        RECT 93.595 156.605 93.805 157.425 ;
        RECT 95.415 157.375 96.165 157.895 ;
        RECT 96.355 157.505 96.685 157.875 ;
        RECT 96.920 157.580 97.205 157.910 ;
        RECT 94.495 156.605 96.165 157.375 ;
        RECT 96.920 157.325 97.090 157.580 ;
        RECT 96.425 157.155 97.090 157.325 ;
        RECT 97.375 157.280 97.545 158.080 ;
        RECT 97.715 158.065 99.385 159.155 ;
        RECT 97.715 157.545 98.465 158.065 ;
        RECT 99.595 158.015 99.825 159.155 ;
        RECT 99.995 158.005 100.325 158.985 ;
        RECT 100.495 158.015 100.705 159.155 ;
        RECT 98.635 157.375 99.385 157.895 ;
        RECT 99.575 157.595 99.905 157.845 ;
        RECT 96.425 156.775 96.595 157.155 ;
        RECT 96.775 156.605 97.105 156.985 ;
        RECT 97.285 156.775 97.545 157.280 ;
        RECT 97.715 156.605 99.385 157.375 ;
        RECT 99.595 156.605 99.825 157.425 ;
        RECT 100.075 157.405 100.325 158.005 ;
        RECT 101.395 157.990 101.685 159.155 ;
        RECT 102.315 158.065 103.985 159.155 ;
        RECT 104.155 158.080 104.425 158.985 ;
        RECT 104.595 158.395 104.925 159.155 ;
        RECT 105.105 158.225 105.275 158.985 ;
        RECT 102.315 157.545 103.065 158.065 ;
        RECT 99.995 156.775 100.325 157.405 ;
        RECT 100.495 156.605 100.705 157.425 ;
        RECT 103.235 157.375 103.985 157.895 ;
        RECT 101.395 156.605 101.685 157.330 ;
        RECT 102.315 156.605 103.985 157.375 ;
        RECT 104.155 157.280 104.325 158.080 ;
        RECT 104.610 158.055 105.275 158.225 ;
        RECT 105.625 158.225 105.795 158.985 ;
        RECT 105.975 158.395 106.305 159.155 ;
        RECT 105.625 158.055 106.290 158.225 ;
        RECT 106.475 158.080 106.745 158.985 ;
        RECT 104.610 157.910 104.780 158.055 ;
        RECT 104.495 157.580 104.780 157.910 ;
        RECT 106.120 157.910 106.290 158.055 ;
        RECT 104.610 157.325 104.780 157.580 ;
        RECT 105.015 157.505 105.345 157.875 ;
        RECT 105.555 157.505 105.885 157.875 ;
        RECT 106.120 157.580 106.405 157.910 ;
        RECT 106.120 157.325 106.290 157.580 ;
        RECT 104.155 156.775 104.415 157.280 ;
        RECT 104.610 157.155 105.275 157.325 ;
        RECT 104.595 156.605 104.925 156.985 ;
        RECT 105.105 156.775 105.275 157.155 ;
        RECT 105.625 157.155 106.290 157.325 ;
        RECT 106.575 157.280 106.745 158.080 ;
        RECT 105.625 156.775 105.795 157.155 ;
        RECT 105.975 156.605 106.305 156.985 ;
        RECT 106.485 156.775 106.745 157.280 ;
        RECT 107.835 158.015 108.175 158.985 ;
        RECT 108.345 158.015 108.515 159.155 ;
        RECT 108.785 158.355 109.035 159.155 ;
        RECT 109.680 158.185 110.010 158.985 ;
        RECT 110.310 158.355 110.640 159.155 ;
        RECT 110.810 158.185 111.140 158.985 ;
        RECT 108.705 158.015 111.140 158.185 ;
        RECT 112.435 158.065 115.945 159.155 ;
        RECT 116.230 158.525 116.515 158.985 ;
        RECT 116.685 158.695 116.955 159.155 ;
        RECT 116.230 158.305 117.185 158.525 ;
        RECT 107.835 157.405 108.010 158.015 ;
        RECT 108.705 157.765 108.875 158.015 ;
        RECT 108.180 157.595 108.875 157.765 ;
        RECT 109.050 157.595 109.470 157.795 ;
        RECT 109.640 157.595 109.970 157.795 ;
        RECT 110.140 157.595 110.470 157.795 ;
        RECT 107.835 156.775 108.175 157.405 ;
        RECT 108.345 156.605 108.595 157.405 ;
        RECT 108.785 157.255 110.010 157.425 ;
        RECT 108.785 156.775 109.115 157.255 ;
        RECT 109.285 156.605 109.510 157.065 ;
        RECT 109.680 156.775 110.010 157.255 ;
        RECT 110.640 157.385 110.810 158.015 ;
        RECT 110.995 157.595 111.345 157.845 ;
        RECT 112.435 157.545 114.125 158.065 ;
        RECT 110.640 156.775 111.140 157.385 ;
        RECT 114.295 157.375 115.945 157.895 ;
        RECT 116.115 157.575 116.805 158.135 ;
        RECT 116.975 157.405 117.185 158.305 ;
        RECT 112.435 156.605 115.945 157.375 ;
        RECT 116.230 157.235 117.185 157.405 ;
        RECT 117.355 158.135 117.755 158.985 ;
        RECT 117.945 158.525 118.225 158.985 ;
        RECT 118.745 158.695 119.070 159.155 ;
        RECT 117.945 158.305 119.070 158.525 ;
        RECT 117.355 157.575 118.450 158.135 ;
        RECT 118.620 157.845 119.070 158.305 ;
        RECT 119.240 158.015 119.625 158.985 ;
        RECT 120.720 158.720 126.065 159.155 ;
        RECT 116.230 156.775 116.515 157.235 ;
        RECT 116.685 156.605 116.955 157.065 ;
        RECT 117.355 156.775 117.755 157.575 ;
        RECT 118.620 157.515 119.175 157.845 ;
        RECT 118.620 157.405 119.070 157.515 ;
        RECT 117.945 157.235 119.070 157.405 ;
        RECT 119.345 157.345 119.625 158.015 ;
        RECT 122.310 157.470 122.660 158.720 ;
        RECT 126.235 158.065 127.445 159.155 ;
        RECT 117.945 156.775 118.225 157.235 ;
        RECT 118.745 156.605 119.070 157.065 ;
        RECT 119.240 156.775 119.625 157.345 ;
        RECT 124.140 157.150 124.480 157.980 ;
        RECT 126.235 157.525 126.755 158.065 ;
        RECT 126.925 157.355 127.445 157.895 ;
        RECT 120.720 156.605 126.065 157.150 ;
        RECT 126.235 156.605 127.445 157.355 ;
        RECT 14.370 156.435 127.530 156.605 ;
        RECT 14.455 155.685 15.665 156.435 ;
        RECT 17.130 156.095 17.385 156.255 ;
        RECT 17.045 155.925 17.385 156.095 ;
        RECT 17.565 155.975 17.850 156.435 ;
        RECT 17.130 155.725 17.385 155.925 ;
        RECT 14.455 155.145 14.975 155.685 ;
        RECT 15.145 154.975 15.665 155.515 ;
        RECT 14.455 153.885 15.665 154.975 ;
        RECT 17.130 154.865 17.310 155.725 ;
        RECT 18.030 155.525 18.280 156.175 ;
        RECT 17.480 155.195 18.280 155.525 ;
        RECT 17.130 154.195 17.385 154.865 ;
        RECT 17.565 153.885 17.850 154.685 ;
        RECT 18.030 154.605 18.280 155.195 ;
        RECT 18.480 155.840 18.800 156.170 ;
        RECT 18.980 155.955 19.640 156.435 ;
        RECT 19.840 156.045 20.690 156.215 ;
        RECT 18.480 154.945 18.670 155.840 ;
        RECT 18.990 155.515 19.650 155.785 ;
        RECT 19.320 155.455 19.650 155.515 ;
        RECT 18.840 155.285 19.170 155.345 ;
        RECT 19.840 155.285 20.010 156.045 ;
        RECT 21.250 155.975 21.570 156.435 ;
        RECT 21.770 155.795 22.020 156.225 ;
        RECT 22.310 155.995 22.720 156.435 ;
        RECT 22.890 156.055 23.905 156.255 ;
        RECT 20.180 155.625 21.430 155.795 ;
        RECT 20.180 155.505 20.510 155.625 ;
        RECT 18.840 155.115 20.740 155.285 ;
        RECT 18.480 154.775 20.400 154.945 ;
        RECT 18.480 154.755 18.800 154.775 ;
        RECT 18.030 154.095 18.360 154.605 ;
        RECT 18.630 154.145 18.800 154.755 ;
        RECT 20.570 154.605 20.740 155.115 ;
        RECT 20.910 155.045 21.090 155.455 ;
        RECT 21.260 154.865 21.430 155.625 ;
        RECT 18.970 153.885 19.300 154.575 ;
        RECT 19.530 154.435 20.740 154.605 ;
        RECT 20.910 154.555 21.430 154.865 ;
        RECT 21.600 155.455 22.020 155.795 ;
        RECT 22.310 155.455 22.720 155.785 ;
        RECT 21.600 154.685 21.790 155.455 ;
        RECT 22.890 155.325 23.060 156.055 ;
        RECT 24.205 155.885 24.375 156.215 ;
        RECT 24.545 156.055 24.875 156.435 ;
        RECT 23.230 155.505 23.580 155.875 ;
        RECT 22.890 155.285 23.310 155.325 ;
        RECT 21.960 155.115 23.310 155.285 ;
        RECT 21.960 154.955 22.210 155.115 ;
        RECT 22.720 154.685 22.970 154.945 ;
        RECT 21.600 154.435 22.970 154.685 ;
        RECT 19.530 154.145 19.770 154.435 ;
        RECT 20.570 154.355 20.740 154.435 ;
        RECT 19.970 153.885 20.390 154.265 ;
        RECT 20.570 154.105 21.200 154.355 ;
        RECT 21.670 153.885 22.000 154.265 ;
        RECT 22.170 154.145 22.340 154.435 ;
        RECT 23.140 154.270 23.310 155.115 ;
        RECT 23.760 154.945 23.980 155.815 ;
        RECT 24.205 155.695 24.900 155.885 ;
        RECT 23.480 154.565 23.980 154.945 ;
        RECT 24.150 154.895 24.560 155.515 ;
        RECT 24.730 154.725 24.900 155.695 ;
        RECT 24.205 154.555 24.900 154.725 ;
        RECT 22.520 153.885 22.900 154.265 ;
        RECT 23.140 154.100 23.970 154.270 ;
        RECT 24.205 154.055 24.375 154.555 ;
        RECT 24.545 153.885 24.875 154.385 ;
        RECT 25.090 154.055 25.315 156.175 ;
        RECT 25.485 156.055 25.815 156.435 ;
        RECT 25.985 155.885 26.155 156.175 ;
        RECT 25.490 155.715 26.155 155.885 ;
        RECT 26.415 155.760 26.675 156.265 ;
        RECT 26.855 156.055 27.185 156.435 ;
        RECT 27.365 155.885 27.535 156.265 ;
        RECT 25.490 154.725 25.720 155.715 ;
        RECT 25.890 154.895 26.240 155.545 ;
        RECT 26.415 154.960 26.585 155.760 ;
        RECT 26.870 155.715 27.535 155.885 ;
        RECT 26.870 155.460 27.040 155.715 ;
        RECT 27.795 155.685 29.005 156.435 ;
        RECT 26.755 155.130 27.040 155.460 ;
        RECT 27.275 155.165 27.605 155.535 ;
        RECT 26.870 154.985 27.040 155.130 ;
        RECT 25.490 154.555 26.155 154.725 ;
        RECT 25.485 153.885 25.815 154.385 ;
        RECT 25.985 154.055 26.155 154.555 ;
        RECT 26.415 154.055 26.685 154.960 ;
        RECT 26.870 154.815 27.535 154.985 ;
        RECT 26.855 153.885 27.185 154.645 ;
        RECT 27.365 154.055 27.535 154.815 ;
        RECT 27.795 154.975 28.315 155.515 ;
        RECT 28.485 155.145 29.005 155.685 ;
        RECT 29.175 155.665 32.685 156.435 ;
        RECT 29.175 154.975 30.865 155.495 ;
        RECT 31.035 155.145 32.685 155.665 ;
        RECT 33.130 155.625 33.375 156.230 ;
        RECT 33.595 155.900 34.105 156.435 ;
        RECT 32.855 155.455 34.085 155.625 ;
        RECT 27.795 153.885 29.005 154.975 ;
        RECT 29.175 153.885 32.685 154.975 ;
        RECT 32.855 154.645 33.195 155.455 ;
        RECT 33.365 154.890 34.115 155.080 ;
        RECT 32.855 154.235 33.370 154.645 ;
        RECT 33.605 153.885 33.775 154.645 ;
        RECT 33.945 154.225 34.115 154.890 ;
        RECT 34.285 154.905 34.475 156.265 ;
        RECT 34.645 156.095 34.920 156.265 ;
        RECT 34.645 155.925 34.925 156.095 ;
        RECT 34.645 155.105 34.920 155.925 ;
        RECT 35.110 155.900 35.640 156.265 ;
        RECT 36.065 156.035 36.395 156.435 ;
        RECT 35.465 155.865 35.640 155.900 ;
        RECT 35.125 154.905 35.295 155.705 ;
        RECT 34.285 154.735 35.295 154.905 ;
        RECT 35.465 155.695 36.395 155.865 ;
        RECT 36.565 155.695 36.820 156.265 ;
        RECT 36.995 155.710 37.285 156.435 ;
        RECT 35.465 154.565 35.635 155.695 ;
        RECT 36.225 155.525 36.395 155.695 ;
        RECT 34.510 154.395 35.635 154.565 ;
        RECT 35.805 155.195 36.000 155.525 ;
        RECT 36.225 155.195 36.480 155.525 ;
        RECT 35.805 154.225 35.975 155.195 ;
        RECT 36.650 155.025 36.820 155.695 ;
        RECT 37.915 155.665 39.585 156.435 ;
        RECT 33.945 154.055 35.975 154.225 ;
        RECT 36.145 153.885 36.315 155.025 ;
        RECT 36.485 154.055 36.820 155.025 ;
        RECT 36.995 153.885 37.285 155.050 ;
        RECT 37.915 154.975 38.665 155.495 ;
        RECT 38.835 155.145 39.585 155.665 ;
        RECT 39.755 155.635 40.095 156.265 ;
        RECT 40.265 155.635 40.515 156.435 ;
        RECT 40.705 155.785 41.035 156.265 ;
        RECT 41.205 155.975 41.430 156.435 ;
        RECT 41.600 155.785 41.930 156.265 ;
        RECT 39.755 155.025 39.930 155.635 ;
        RECT 40.705 155.615 41.930 155.785 ;
        RECT 42.560 155.655 43.060 156.265 ;
        RECT 40.100 155.275 40.795 155.445 ;
        RECT 40.625 155.025 40.795 155.275 ;
        RECT 40.970 155.245 41.390 155.445 ;
        RECT 41.560 155.245 41.890 155.445 ;
        RECT 42.060 155.245 42.390 155.445 ;
        RECT 42.560 155.025 42.730 155.655 ;
        RECT 43.435 155.635 43.775 156.265 ;
        RECT 43.945 155.635 44.195 156.435 ;
        RECT 44.385 155.785 44.715 156.265 ;
        RECT 44.885 155.975 45.110 156.435 ;
        RECT 45.280 155.785 45.610 156.265 ;
        RECT 42.915 155.195 43.265 155.445 ;
        RECT 43.435 155.025 43.610 155.635 ;
        RECT 44.385 155.615 45.610 155.785 ;
        RECT 46.240 155.655 46.740 156.265 ;
        RECT 43.780 155.275 44.475 155.445 ;
        RECT 44.305 155.025 44.475 155.275 ;
        RECT 44.650 155.245 45.070 155.445 ;
        RECT 45.240 155.245 45.570 155.445 ;
        RECT 45.740 155.245 46.070 155.445 ;
        RECT 46.240 155.025 46.410 155.655 ;
        RECT 47.115 155.635 47.455 156.265 ;
        RECT 47.625 155.635 47.875 156.435 ;
        RECT 48.065 155.785 48.395 156.265 ;
        RECT 48.565 155.975 48.790 156.435 ;
        RECT 48.960 155.785 49.290 156.265 ;
        RECT 46.595 155.195 46.945 155.445 ;
        RECT 47.115 155.025 47.290 155.635 ;
        RECT 48.065 155.615 49.290 155.785 ;
        RECT 49.920 155.655 50.420 156.265 ;
        RECT 51.255 155.665 52.925 156.435 ;
        RECT 47.460 155.275 48.155 155.445 ;
        RECT 47.985 155.025 48.155 155.275 ;
        RECT 48.330 155.245 48.750 155.445 ;
        RECT 48.920 155.245 49.250 155.445 ;
        RECT 49.420 155.245 49.750 155.445 ;
        RECT 49.920 155.025 50.090 155.655 ;
        RECT 50.275 155.195 50.625 155.445 ;
        RECT 37.915 153.885 39.585 154.975 ;
        RECT 39.755 154.055 40.095 155.025 ;
        RECT 40.265 153.885 40.435 155.025 ;
        RECT 40.625 154.855 43.060 155.025 ;
        RECT 40.705 153.885 40.955 154.685 ;
        RECT 41.600 154.055 41.930 154.855 ;
        RECT 42.230 153.885 42.560 154.685 ;
        RECT 42.730 154.055 43.060 154.855 ;
        RECT 43.435 154.055 43.775 155.025 ;
        RECT 43.945 153.885 44.115 155.025 ;
        RECT 44.305 154.855 46.740 155.025 ;
        RECT 44.385 153.885 44.635 154.685 ;
        RECT 45.280 154.055 45.610 154.855 ;
        RECT 45.910 153.885 46.240 154.685 ;
        RECT 46.410 154.055 46.740 154.855 ;
        RECT 47.115 154.055 47.455 155.025 ;
        RECT 47.625 153.885 47.795 155.025 ;
        RECT 47.985 154.855 50.420 155.025 ;
        RECT 48.065 153.885 48.315 154.685 ;
        RECT 48.960 154.055 49.290 154.855 ;
        RECT 49.590 153.885 49.920 154.685 ;
        RECT 50.090 154.055 50.420 154.855 ;
        RECT 51.255 154.975 52.005 155.495 ;
        RECT 52.175 155.145 52.925 155.665 ;
        RECT 53.470 155.725 53.725 156.255 ;
        RECT 53.905 155.975 54.190 156.435 ;
        RECT 51.255 153.885 52.925 154.975 ;
        RECT 53.470 154.865 53.650 155.725 ;
        RECT 54.370 155.525 54.620 156.175 ;
        RECT 53.820 155.195 54.620 155.525 ;
        RECT 53.470 154.395 53.725 154.865 ;
        RECT 53.385 154.225 53.725 154.395 ;
        RECT 53.470 154.195 53.725 154.225 ;
        RECT 53.905 153.885 54.190 154.685 ;
        RECT 54.370 154.605 54.620 155.195 ;
        RECT 54.820 155.840 55.140 156.170 ;
        RECT 55.320 155.955 55.980 156.435 ;
        RECT 56.180 156.045 57.030 156.215 ;
        RECT 54.820 154.945 55.010 155.840 ;
        RECT 55.330 155.515 55.990 155.785 ;
        RECT 55.660 155.455 55.990 155.515 ;
        RECT 55.180 155.285 55.510 155.345 ;
        RECT 56.180 155.285 56.350 156.045 ;
        RECT 57.590 155.975 57.910 156.435 ;
        RECT 58.110 155.795 58.360 156.225 ;
        RECT 58.650 155.995 59.060 156.435 ;
        RECT 59.230 156.055 60.245 156.255 ;
        RECT 56.520 155.625 57.770 155.795 ;
        RECT 56.520 155.505 56.850 155.625 ;
        RECT 55.180 155.115 57.080 155.285 ;
        RECT 54.820 154.775 56.740 154.945 ;
        RECT 54.820 154.755 55.140 154.775 ;
        RECT 54.370 154.095 54.700 154.605 ;
        RECT 54.970 154.145 55.140 154.755 ;
        RECT 56.910 154.605 57.080 155.115 ;
        RECT 57.250 155.045 57.430 155.455 ;
        RECT 57.600 154.865 57.770 155.625 ;
        RECT 55.310 153.885 55.640 154.575 ;
        RECT 55.870 154.435 57.080 154.605 ;
        RECT 57.250 154.555 57.770 154.865 ;
        RECT 57.940 155.455 58.360 155.795 ;
        RECT 58.650 155.455 59.060 155.785 ;
        RECT 57.940 154.685 58.130 155.455 ;
        RECT 59.230 155.325 59.400 156.055 ;
        RECT 60.545 155.885 60.715 156.215 ;
        RECT 60.885 156.055 61.215 156.435 ;
        RECT 59.570 155.505 59.920 155.875 ;
        RECT 59.230 155.285 59.650 155.325 ;
        RECT 58.300 155.115 59.650 155.285 ;
        RECT 58.300 154.955 58.550 155.115 ;
        RECT 59.060 154.685 59.310 154.945 ;
        RECT 57.940 154.435 59.310 154.685 ;
        RECT 55.870 154.145 56.110 154.435 ;
        RECT 56.910 154.355 57.080 154.435 ;
        RECT 56.310 153.885 56.730 154.265 ;
        RECT 56.910 154.105 57.540 154.355 ;
        RECT 58.010 153.885 58.340 154.265 ;
        RECT 58.510 154.145 58.680 154.435 ;
        RECT 59.480 154.270 59.650 155.115 ;
        RECT 60.100 154.945 60.320 155.815 ;
        RECT 60.545 155.695 61.240 155.885 ;
        RECT 59.820 154.565 60.320 154.945 ;
        RECT 60.490 154.895 60.900 155.515 ;
        RECT 61.070 154.725 61.240 155.695 ;
        RECT 60.545 154.555 61.240 154.725 ;
        RECT 58.860 153.885 59.240 154.265 ;
        RECT 59.480 154.100 60.310 154.270 ;
        RECT 60.545 154.055 60.715 154.555 ;
        RECT 60.885 153.885 61.215 154.385 ;
        RECT 61.430 154.055 61.655 156.175 ;
        RECT 61.825 156.055 62.155 156.435 ;
        RECT 62.325 155.885 62.495 156.175 ;
        RECT 61.830 155.715 62.495 155.885 ;
        RECT 61.830 154.725 62.060 155.715 ;
        RECT 62.755 155.710 63.045 156.435 ;
        RECT 63.675 155.665 65.345 156.435 ;
        RECT 65.605 155.955 65.905 156.435 ;
        RECT 66.075 155.785 66.335 156.240 ;
        RECT 66.505 155.955 66.765 156.435 ;
        RECT 66.945 155.785 67.205 156.240 ;
        RECT 67.375 155.955 67.625 156.435 ;
        RECT 67.805 155.785 68.065 156.240 ;
        RECT 68.235 155.955 68.485 156.435 ;
        RECT 68.665 155.785 68.925 156.240 ;
        RECT 69.095 155.955 69.340 156.435 ;
        RECT 69.510 155.785 69.785 156.240 ;
        RECT 69.955 155.955 70.200 156.435 ;
        RECT 70.370 155.785 70.630 156.240 ;
        RECT 70.800 155.955 71.060 156.435 ;
        RECT 71.230 155.785 71.490 156.240 ;
        RECT 71.660 155.955 71.920 156.435 ;
        RECT 72.090 155.785 72.350 156.240 ;
        RECT 72.520 155.875 72.780 156.435 ;
        RECT 62.230 154.895 62.580 155.545 ;
        RECT 61.830 154.555 62.495 154.725 ;
        RECT 61.825 153.885 62.155 154.385 ;
        RECT 62.325 154.055 62.495 154.555 ;
        RECT 62.755 153.885 63.045 155.050 ;
        RECT 63.675 154.975 64.425 155.495 ;
        RECT 64.595 155.145 65.345 155.665 ;
        RECT 65.605 155.615 72.350 155.785 ;
        RECT 65.605 155.075 66.770 155.615 ;
        RECT 72.950 155.445 73.200 156.255 ;
        RECT 73.380 155.910 73.640 156.435 ;
        RECT 73.810 155.445 74.060 156.255 ;
        RECT 74.240 155.925 74.545 156.435 ;
        RECT 66.940 155.195 74.060 155.445 ;
        RECT 74.230 155.195 74.545 155.755 ;
        RECT 74.715 155.665 76.385 156.435 ;
        RECT 65.575 155.025 66.770 155.075 ;
        RECT 63.675 153.885 65.345 154.975 ;
        RECT 65.575 154.905 72.350 155.025 ;
        RECT 65.605 154.800 72.350 154.905 ;
        RECT 65.605 153.885 65.875 154.630 ;
        RECT 66.045 154.060 66.335 154.800 ;
        RECT 66.945 154.785 72.350 154.800 ;
        RECT 66.505 153.890 66.760 154.615 ;
        RECT 66.945 154.060 67.205 154.785 ;
        RECT 67.375 153.890 67.620 154.615 ;
        RECT 67.805 154.060 68.065 154.785 ;
        RECT 68.235 153.890 68.480 154.615 ;
        RECT 68.665 154.060 68.925 154.785 ;
        RECT 69.095 153.890 69.340 154.615 ;
        RECT 69.510 154.060 69.770 154.785 ;
        RECT 69.940 153.890 70.200 154.615 ;
        RECT 70.370 154.060 70.630 154.785 ;
        RECT 70.800 153.890 71.060 154.615 ;
        RECT 71.230 154.060 71.490 154.785 ;
        RECT 71.660 153.890 71.920 154.615 ;
        RECT 72.090 154.060 72.350 154.785 ;
        RECT 72.520 153.890 72.780 154.685 ;
        RECT 72.950 154.060 73.200 155.195 ;
        RECT 66.505 153.885 72.780 153.890 ;
        RECT 73.380 153.885 73.640 154.695 ;
        RECT 73.815 154.055 74.060 155.195 ;
        RECT 74.715 154.975 75.465 155.495 ;
        RECT 75.635 155.145 76.385 155.665 ;
        RECT 76.555 155.635 76.895 156.265 ;
        RECT 77.065 155.635 77.315 156.435 ;
        RECT 77.505 155.785 77.835 156.265 ;
        RECT 78.005 155.975 78.230 156.435 ;
        RECT 78.400 155.785 78.730 156.265 ;
        RECT 76.555 155.025 76.730 155.635 ;
        RECT 77.505 155.615 78.730 155.785 ;
        RECT 79.360 155.655 79.860 156.265 ;
        RECT 76.900 155.275 77.595 155.445 ;
        RECT 77.425 155.025 77.595 155.275 ;
        RECT 77.770 155.245 78.190 155.445 ;
        RECT 78.360 155.245 78.690 155.445 ;
        RECT 78.860 155.245 79.190 155.445 ;
        RECT 79.360 155.025 79.530 155.655 ;
        RECT 80.235 155.635 80.575 156.265 ;
        RECT 80.745 155.635 80.995 156.435 ;
        RECT 81.185 155.785 81.515 156.265 ;
        RECT 81.685 155.975 81.910 156.435 ;
        RECT 82.080 155.785 82.410 156.265 ;
        RECT 79.715 155.195 80.065 155.445 ;
        RECT 80.235 155.025 80.410 155.635 ;
        RECT 81.185 155.615 82.410 155.785 ;
        RECT 83.040 155.655 83.540 156.265 ;
        RECT 84.835 155.665 88.345 156.435 ;
        RECT 88.515 155.710 88.805 156.435 ;
        RECT 88.975 155.665 91.565 156.435 ;
        RECT 91.740 155.890 97.085 156.435 ;
        RECT 80.580 155.275 81.275 155.445 ;
        RECT 81.105 155.025 81.275 155.275 ;
        RECT 81.450 155.245 81.870 155.445 ;
        RECT 82.040 155.245 82.370 155.445 ;
        RECT 82.540 155.245 82.870 155.445 ;
        RECT 83.040 155.025 83.210 155.655 ;
        RECT 83.395 155.195 83.745 155.445 ;
        RECT 74.240 153.885 74.535 154.695 ;
        RECT 74.715 153.885 76.385 154.975 ;
        RECT 76.555 154.055 76.895 155.025 ;
        RECT 77.065 153.885 77.235 155.025 ;
        RECT 77.425 154.855 79.860 155.025 ;
        RECT 77.505 153.885 77.755 154.685 ;
        RECT 78.400 154.055 78.730 154.855 ;
        RECT 79.030 153.885 79.360 154.685 ;
        RECT 79.530 154.055 79.860 154.855 ;
        RECT 80.235 154.055 80.575 155.025 ;
        RECT 80.745 153.885 80.915 155.025 ;
        RECT 81.105 154.855 83.540 155.025 ;
        RECT 81.185 153.885 81.435 154.685 ;
        RECT 82.080 154.055 82.410 154.855 ;
        RECT 82.710 153.885 83.040 154.685 ;
        RECT 83.210 154.055 83.540 154.855 ;
        RECT 84.835 154.975 86.525 155.495 ;
        RECT 86.695 155.145 88.345 155.665 ;
        RECT 84.835 153.885 88.345 154.975 ;
        RECT 88.515 153.885 88.805 155.050 ;
        RECT 88.975 154.975 90.185 155.495 ;
        RECT 90.355 155.145 91.565 155.665 ;
        RECT 88.975 153.885 91.565 154.975 ;
        RECT 93.330 154.320 93.680 155.570 ;
        RECT 95.160 155.060 95.500 155.890 ;
        RECT 97.460 155.655 97.960 156.265 ;
        RECT 97.255 155.195 97.605 155.445 ;
        RECT 97.790 155.025 97.960 155.655 ;
        RECT 98.590 155.785 98.920 156.265 ;
        RECT 99.090 155.975 99.315 156.435 ;
        RECT 99.485 155.785 99.815 156.265 ;
        RECT 98.590 155.615 99.815 155.785 ;
        RECT 100.005 155.635 100.255 156.435 ;
        RECT 100.425 155.635 100.765 156.265 ;
        RECT 101.395 155.665 103.065 156.435 ;
        RECT 98.130 155.245 98.460 155.445 ;
        RECT 98.630 155.245 98.960 155.445 ;
        RECT 99.130 155.245 99.550 155.445 ;
        RECT 99.725 155.275 100.420 155.445 ;
        RECT 99.725 155.025 99.895 155.275 ;
        RECT 100.590 155.025 100.765 155.635 ;
        RECT 97.460 154.855 99.895 155.025 ;
        RECT 91.740 153.885 97.085 154.320 ;
        RECT 97.460 154.055 97.790 154.855 ;
        RECT 97.960 153.885 98.290 154.685 ;
        RECT 98.590 154.055 98.920 154.855 ;
        RECT 99.565 153.885 99.815 154.685 ;
        RECT 100.085 153.885 100.255 155.025 ;
        RECT 100.425 154.055 100.765 155.025 ;
        RECT 101.395 154.975 102.145 155.495 ;
        RECT 102.315 155.145 103.065 155.665 ;
        RECT 103.235 155.635 103.575 156.265 ;
        RECT 103.745 155.635 103.995 156.435 ;
        RECT 104.185 155.785 104.515 156.265 ;
        RECT 104.685 155.975 104.910 156.435 ;
        RECT 105.080 155.785 105.410 156.265 ;
        RECT 103.235 155.025 103.410 155.635 ;
        RECT 104.185 155.615 105.410 155.785 ;
        RECT 106.040 155.655 106.540 156.265 ;
        RECT 107.120 155.655 107.620 156.265 ;
        RECT 103.580 155.275 104.275 155.445 ;
        RECT 104.105 155.025 104.275 155.275 ;
        RECT 104.450 155.245 104.870 155.445 ;
        RECT 105.040 155.245 105.370 155.445 ;
        RECT 105.540 155.245 105.870 155.445 ;
        RECT 106.040 155.025 106.210 155.655 ;
        RECT 106.395 155.195 106.745 155.445 ;
        RECT 106.915 155.195 107.265 155.445 ;
        RECT 107.450 155.025 107.620 155.655 ;
        RECT 108.250 155.785 108.580 156.265 ;
        RECT 108.750 155.975 108.975 156.435 ;
        RECT 109.145 155.785 109.475 156.265 ;
        RECT 108.250 155.615 109.475 155.785 ;
        RECT 109.665 155.635 109.915 156.435 ;
        RECT 110.085 155.635 110.425 156.265 ;
        RECT 110.595 155.665 114.105 156.435 ;
        RECT 114.275 155.710 114.565 156.435 ;
        RECT 114.735 155.685 115.945 156.435 ;
        RECT 107.790 155.245 108.120 155.445 ;
        RECT 108.290 155.245 108.620 155.445 ;
        RECT 108.790 155.245 109.210 155.445 ;
        RECT 109.385 155.275 110.080 155.445 ;
        RECT 109.385 155.025 109.555 155.275 ;
        RECT 110.250 155.025 110.425 155.635 ;
        RECT 101.395 153.885 103.065 154.975 ;
        RECT 103.235 154.055 103.575 155.025 ;
        RECT 103.745 153.885 103.915 155.025 ;
        RECT 104.105 154.855 106.540 155.025 ;
        RECT 104.185 153.885 104.435 154.685 ;
        RECT 105.080 154.055 105.410 154.855 ;
        RECT 105.710 153.885 106.040 154.685 ;
        RECT 106.210 154.055 106.540 154.855 ;
        RECT 107.120 154.855 109.555 155.025 ;
        RECT 107.120 154.055 107.450 154.855 ;
        RECT 107.620 153.885 107.950 154.685 ;
        RECT 108.250 154.055 108.580 154.855 ;
        RECT 109.225 153.885 109.475 154.685 ;
        RECT 109.745 153.885 109.915 155.025 ;
        RECT 110.085 154.055 110.425 155.025 ;
        RECT 110.595 154.975 112.285 155.495 ;
        RECT 112.455 155.145 114.105 155.665 ;
        RECT 110.595 153.885 114.105 154.975 ;
        RECT 114.275 153.885 114.565 155.050 ;
        RECT 114.735 154.975 115.255 155.515 ;
        RECT 115.425 155.145 115.945 155.685 ;
        RECT 116.205 155.785 116.375 156.265 ;
        RECT 116.555 155.955 116.795 156.435 ;
        RECT 117.045 155.785 117.215 156.265 ;
        RECT 117.385 155.955 117.715 156.435 ;
        RECT 117.885 155.785 118.055 156.265 ;
        RECT 116.205 155.615 116.840 155.785 ;
        RECT 117.045 155.615 118.055 155.785 ;
        RECT 118.225 155.635 118.555 156.435 ;
        RECT 118.875 155.665 120.545 156.435 ;
        RECT 120.720 155.890 126.065 156.435 ;
        RECT 116.670 155.445 116.840 155.615 ;
        RECT 116.120 155.205 116.500 155.445 ;
        RECT 116.670 155.275 117.170 155.445 ;
        RECT 116.670 155.035 116.840 155.275 ;
        RECT 117.560 155.075 118.055 155.615 ;
        RECT 114.735 153.885 115.945 154.975 ;
        RECT 116.125 154.865 116.840 155.035 ;
        RECT 117.045 154.905 118.055 155.075 ;
        RECT 116.125 154.055 116.455 154.865 ;
        RECT 116.625 153.885 116.865 154.685 ;
        RECT 117.045 154.055 117.215 154.905 ;
        RECT 117.385 153.885 117.715 154.685 ;
        RECT 117.885 154.055 118.055 154.905 ;
        RECT 118.225 153.885 118.555 155.035 ;
        RECT 118.875 154.975 119.625 155.495 ;
        RECT 119.795 155.145 120.545 155.665 ;
        RECT 118.875 153.885 120.545 154.975 ;
        RECT 122.310 154.320 122.660 155.570 ;
        RECT 124.140 155.060 124.480 155.890 ;
        RECT 126.235 155.685 127.445 156.435 ;
        RECT 126.235 154.975 126.755 155.515 ;
        RECT 126.925 155.145 127.445 155.685 ;
        RECT 120.720 153.885 126.065 154.320 ;
        RECT 126.235 153.885 127.445 154.975 ;
        RECT 14.370 153.715 127.530 153.885 ;
        RECT 14.455 152.625 15.665 153.715 ;
        RECT 14.455 151.915 14.975 152.455 ;
        RECT 15.145 152.085 15.665 152.625 ;
        RECT 16.295 152.625 19.805 153.715 ;
        RECT 19.975 152.955 20.490 153.365 ;
        RECT 20.725 152.955 20.895 153.715 ;
        RECT 21.065 153.375 23.095 153.545 ;
        RECT 16.295 152.105 17.985 152.625 ;
        RECT 18.155 151.935 19.805 152.455 ;
        RECT 19.975 152.145 20.315 152.955 ;
        RECT 21.065 152.710 21.235 153.375 ;
        RECT 21.630 153.035 22.755 153.205 ;
        RECT 20.485 152.520 21.235 152.710 ;
        RECT 21.405 152.695 22.415 152.865 ;
        RECT 19.975 151.975 21.205 152.145 ;
        RECT 14.455 151.165 15.665 151.915 ;
        RECT 16.295 151.165 19.805 151.935 ;
        RECT 20.250 151.370 20.495 151.975 ;
        RECT 20.715 151.165 21.225 151.700 ;
        RECT 21.405 151.335 21.595 152.695 ;
        RECT 21.765 151.675 22.040 152.495 ;
        RECT 22.245 151.895 22.415 152.695 ;
        RECT 22.585 151.905 22.755 153.035 ;
        RECT 22.925 152.405 23.095 153.375 ;
        RECT 23.265 152.575 23.435 153.715 ;
        RECT 23.605 152.575 23.940 153.545 ;
        RECT 22.925 152.075 23.120 152.405 ;
        RECT 23.345 152.075 23.600 152.405 ;
        RECT 23.345 151.905 23.515 152.075 ;
        RECT 23.770 151.905 23.940 152.575 ;
        RECT 24.115 152.550 24.405 153.715 ;
        RECT 24.575 152.625 25.785 153.715 ;
        RECT 25.955 152.625 29.465 153.715 ;
        RECT 30.010 152.735 30.265 153.405 ;
        RECT 30.445 152.915 30.730 153.715 ;
        RECT 30.910 152.995 31.240 153.505 ;
        RECT 24.575 152.085 25.095 152.625 ;
        RECT 25.265 151.915 25.785 152.455 ;
        RECT 25.955 152.105 27.645 152.625 ;
        RECT 27.815 151.935 29.465 152.455 ;
        RECT 22.585 151.735 23.515 151.905 ;
        RECT 22.585 151.700 22.760 151.735 ;
        RECT 21.765 151.505 22.045 151.675 ;
        RECT 21.765 151.335 22.040 151.505 ;
        RECT 22.230 151.335 22.760 151.700 ;
        RECT 23.185 151.165 23.515 151.565 ;
        RECT 23.685 151.335 23.940 151.905 ;
        RECT 24.115 151.165 24.405 151.890 ;
        RECT 24.575 151.165 25.785 151.915 ;
        RECT 25.955 151.165 29.465 151.935 ;
        RECT 30.010 151.875 30.190 152.735 ;
        RECT 30.910 152.405 31.160 152.995 ;
        RECT 31.510 152.845 31.680 153.455 ;
        RECT 31.850 153.025 32.180 153.715 ;
        RECT 32.410 153.165 32.650 153.455 ;
        RECT 32.850 153.335 33.270 153.715 ;
        RECT 33.450 153.245 34.080 153.495 ;
        RECT 34.550 153.335 34.880 153.715 ;
        RECT 33.450 153.165 33.620 153.245 ;
        RECT 35.050 153.165 35.220 153.455 ;
        RECT 35.400 153.335 35.780 153.715 ;
        RECT 36.020 153.330 36.850 153.500 ;
        RECT 32.410 152.995 33.620 153.165 ;
        RECT 30.360 152.075 31.160 152.405 ;
        RECT 30.010 151.675 30.265 151.875 ;
        RECT 29.925 151.505 30.265 151.675 ;
        RECT 30.010 151.345 30.265 151.505 ;
        RECT 30.445 151.165 30.730 151.625 ;
        RECT 30.910 151.425 31.160 152.075 ;
        RECT 31.360 152.825 31.680 152.845 ;
        RECT 31.360 152.655 33.280 152.825 ;
        RECT 31.360 151.760 31.550 152.655 ;
        RECT 33.450 152.485 33.620 152.995 ;
        RECT 33.790 152.735 34.310 153.045 ;
        RECT 31.720 152.315 33.620 152.485 ;
        RECT 31.720 152.255 32.050 152.315 ;
        RECT 32.200 152.085 32.530 152.145 ;
        RECT 31.870 151.815 32.530 152.085 ;
        RECT 31.360 151.430 31.680 151.760 ;
        RECT 31.860 151.165 32.520 151.645 ;
        RECT 32.720 151.555 32.890 152.315 ;
        RECT 33.790 152.145 33.970 152.555 ;
        RECT 33.060 151.975 33.390 152.095 ;
        RECT 34.140 151.975 34.310 152.735 ;
        RECT 33.060 151.805 34.310 151.975 ;
        RECT 34.480 152.915 35.850 153.165 ;
        RECT 34.480 152.145 34.670 152.915 ;
        RECT 35.600 152.655 35.850 152.915 ;
        RECT 34.840 152.485 35.090 152.645 ;
        RECT 36.020 152.485 36.190 153.330 ;
        RECT 37.085 153.045 37.255 153.545 ;
        RECT 37.425 153.215 37.755 153.715 ;
        RECT 36.360 152.655 36.860 153.035 ;
        RECT 37.085 152.875 37.780 153.045 ;
        RECT 34.840 152.315 36.190 152.485 ;
        RECT 35.770 152.275 36.190 152.315 ;
        RECT 34.480 151.805 34.900 152.145 ;
        RECT 35.190 151.815 35.600 152.145 ;
        RECT 32.720 151.385 33.570 151.555 ;
        RECT 34.130 151.165 34.450 151.625 ;
        RECT 34.650 151.375 34.900 151.805 ;
        RECT 35.190 151.165 35.600 151.605 ;
        RECT 35.770 151.545 35.940 152.275 ;
        RECT 36.110 151.725 36.460 152.095 ;
        RECT 36.640 151.785 36.860 152.655 ;
        RECT 37.030 152.085 37.440 152.705 ;
        RECT 37.610 151.905 37.780 152.875 ;
        RECT 37.085 151.715 37.780 151.905 ;
        RECT 35.770 151.345 36.785 151.545 ;
        RECT 37.085 151.385 37.255 151.715 ;
        RECT 37.425 151.165 37.755 151.545 ;
        RECT 37.970 151.425 38.195 153.545 ;
        RECT 38.365 153.215 38.695 153.715 ;
        RECT 38.865 153.045 39.035 153.545 ;
        RECT 38.370 152.875 39.035 153.045 ;
        RECT 38.370 151.885 38.600 152.875 ;
        RECT 38.770 152.055 39.120 152.705 ;
        RECT 39.295 152.575 39.635 153.545 ;
        RECT 39.805 152.575 39.975 153.715 ;
        RECT 40.245 152.915 40.495 153.715 ;
        RECT 41.140 152.745 41.470 153.545 ;
        RECT 41.770 152.915 42.100 153.715 ;
        RECT 42.270 152.745 42.600 153.545 ;
        RECT 40.165 152.575 42.600 152.745 ;
        RECT 42.975 152.625 44.185 153.715 ;
        RECT 44.360 153.280 49.705 153.715 ;
        RECT 39.295 151.965 39.470 152.575 ;
        RECT 40.165 152.325 40.335 152.575 ;
        RECT 39.640 152.155 40.335 152.325 ;
        RECT 40.510 152.155 40.930 152.355 ;
        RECT 41.100 152.155 41.430 152.355 ;
        RECT 41.600 152.155 41.930 152.355 ;
        RECT 38.370 151.715 39.035 151.885 ;
        RECT 38.365 151.165 38.695 151.545 ;
        RECT 38.865 151.425 39.035 151.715 ;
        RECT 39.295 151.335 39.635 151.965 ;
        RECT 39.805 151.165 40.055 151.965 ;
        RECT 40.245 151.815 41.470 151.985 ;
        RECT 40.245 151.335 40.575 151.815 ;
        RECT 40.745 151.165 40.970 151.625 ;
        RECT 41.140 151.335 41.470 151.815 ;
        RECT 42.100 151.945 42.270 152.575 ;
        RECT 42.455 152.155 42.805 152.405 ;
        RECT 42.975 152.085 43.495 152.625 ;
        RECT 42.100 151.335 42.600 151.945 ;
        RECT 43.665 151.915 44.185 152.455 ;
        RECT 45.950 152.030 46.300 153.280 ;
        RECT 49.875 152.550 50.165 153.715 ;
        RECT 51.260 153.280 56.605 153.715 ;
        RECT 42.975 151.165 44.185 151.915 ;
        RECT 47.780 151.710 48.120 152.540 ;
        RECT 52.850 152.030 53.200 153.280 ;
        RECT 56.815 152.575 57.045 153.715 ;
        RECT 57.215 152.565 57.545 153.545 ;
        RECT 57.715 152.575 57.925 153.715 ;
        RECT 58.530 152.735 58.785 153.405 ;
        RECT 58.965 152.915 59.250 153.715 ;
        RECT 59.430 152.995 59.760 153.505 ;
        RECT 44.360 151.165 49.705 151.710 ;
        RECT 49.875 151.165 50.165 151.890 ;
        RECT 54.680 151.710 55.020 152.540 ;
        RECT 56.795 152.155 57.125 152.405 ;
        RECT 51.260 151.165 56.605 151.710 ;
        RECT 56.815 151.165 57.045 151.985 ;
        RECT 57.295 151.965 57.545 152.565 ;
        RECT 57.215 151.335 57.545 151.965 ;
        RECT 57.715 151.165 57.925 151.985 ;
        RECT 58.530 151.875 58.710 152.735 ;
        RECT 59.430 152.405 59.680 152.995 ;
        RECT 60.030 152.845 60.200 153.455 ;
        RECT 60.370 153.025 60.700 153.715 ;
        RECT 60.930 153.165 61.170 153.455 ;
        RECT 61.370 153.335 61.790 153.715 ;
        RECT 61.970 153.245 62.600 153.495 ;
        RECT 63.070 153.335 63.400 153.715 ;
        RECT 61.970 153.165 62.140 153.245 ;
        RECT 63.570 153.165 63.740 153.455 ;
        RECT 63.920 153.335 64.300 153.715 ;
        RECT 64.540 153.330 65.370 153.500 ;
        RECT 60.930 152.995 62.140 153.165 ;
        RECT 58.880 152.075 59.680 152.405 ;
        RECT 58.530 151.675 58.785 151.875 ;
        RECT 58.445 151.505 58.785 151.675 ;
        RECT 58.530 151.345 58.785 151.505 ;
        RECT 58.965 151.165 59.250 151.625 ;
        RECT 59.430 151.425 59.680 152.075 ;
        RECT 59.880 152.825 60.200 152.845 ;
        RECT 59.880 152.655 61.800 152.825 ;
        RECT 59.880 151.760 60.070 152.655 ;
        RECT 61.970 152.485 62.140 152.995 ;
        RECT 62.310 152.735 62.830 153.045 ;
        RECT 60.240 152.315 62.140 152.485 ;
        RECT 60.240 152.255 60.570 152.315 ;
        RECT 60.720 152.085 61.050 152.145 ;
        RECT 60.390 151.815 61.050 152.085 ;
        RECT 59.880 151.430 60.200 151.760 ;
        RECT 60.380 151.165 61.040 151.645 ;
        RECT 61.240 151.555 61.410 152.315 ;
        RECT 62.310 152.145 62.490 152.555 ;
        RECT 61.580 151.975 61.910 152.095 ;
        RECT 62.660 151.975 62.830 152.735 ;
        RECT 61.580 151.805 62.830 151.975 ;
        RECT 63.000 152.915 64.370 153.165 ;
        RECT 63.000 152.145 63.190 152.915 ;
        RECT 64.120 152.655 64.370 152.915 ;
        RECT 63.360 152.485 63.610 152.645 ;
        RECT 64.540 152.485 64.710 153.330 ;
        RECT 65.605 153.045 65.775 153.545 ;
        RECT 65.945 153.215 66.275 153.715 ;
        RECT 64.880 152.655 65.380 153.035 ;
        RECT 65.605 152.875 66.300 153.045 ;
        RECT 63.360 152.315 64.710 152.485 ;
        RECT 64.290 152.275 64.710 152.315 ;
        RECT 63.000 151.805 63.420 152.145 ;
        RECT 63.710 151.815 64.120 152.145 ;
        RECT 61.240 151.385 62.090 151.555 ;
        RECT 62.650 151.165 62.970 151.625 ;
        RECT 63.170 151.375 63.420 151.805 ;
        RECT 63.710 151.165 64.120 151.605 ;
        RECT 64.290 151.545 64.460 152.275 ;
        RECT 64.630 151.725 64.980 152.095 ;
        RECT 65.160 151.785 65.380 152.655 ;
        RECT 65.550 152.085 65.960 152.705 ;
        RECT 66.130 151.905 66.300 152.875 ;
        RECT 65.605 151.715 66.300 151.905 ;
        RECT 64.290 151.345 65.305 151.545 ;
        RECT 65.605 151.385 65.775 151.715 ;
        RECT 65.945 151.165 66.275 151.545 ;
        RECT 66.490 151.425 66.715 153.545 ;
        RECT 66.885 153.215 67.215 153.715 ;
        RECT 67.385 153.045 67.555 153.545 ;
        RECT 66.890 152.875 67.555 153.045 ;
        RECT 66.890 151.885 67.120 152.875 ;
        RECT 67.290 152.055 67.640 152.705 ;
        RECT 68.275 152.625 70.865 153.715 ;
        RECT 71.125 152.785 71.295 153.545 ;
        RECT 71.510 152.955 71.840 153.715 ;
        RECT 68.275 152.105 69.485 152.625 ;
        RECT 71.125 152.615 71.840 152.785 ;
        RECT 72.010 152.640 72.265 153.545 ;
        RECT 69.655 151.935 70.865 152.455 ;
        RECT 71.035 152.065 71.390 152.435 ;
        RECT 71.670 152.405 71.840 152.615 ;
        RECT 71.670 152.075 71.925 152.405 ;
        RECT 66.890 151.715 67.555 151.885 ;
        RECT 66.885 151.165 67.215 151.545 ;
        RECT 67.385 151.425 67.555 151.715 ;
        RECT 68.275 151.165 70.865 151.935 ;
        RECT 71.670 151.885 71.840 152.075 ;
        RECT 72.095 151.910 72.265 152.640 ;
        RECT 72.440 152.565 72.700 153.715 ;
        RECT 72.885 152.655 73.215 153.715 ;
        RECT 73.395 152.405 73.565 153.375 ;
        RECT 73.735 153.125 74.065 153.525 ;
        RECT 74.235 153.355 74.565 153.715 ;
        RECT 74.765 153.125 75.465 153.545 ;
        RECT 73.735 152.895 75.465 153.125 ;
        RECT 73.735 152.675 74.065 152.895 ;
        RECT 74.260 152.405 74.585 152.695 ;
        RECT 72.875 152.075 73.185 152.405 ;
        RECT 73.395 152.075 73.770 152.405 ;
        RECT 74.090 152.075 74.585 152.405 ;
        RECT 74.760 152.155 75.090 152.695 ;
        RECT 71.125 151.715 71.840 151.885 ;
        RECT 71.125 151.335 71.295 151.715 ;
        RECT 71.510 151.165 71.840 151.545 ;
        RECT 72.010 151.335 72.265 151.910 ;
        RECT 72.440 151.165 72.700 152.005 ;
        RECT 75.260 151.925 75.465 152.895 ;
        RECT 75.635 152.550 75.925 153.715 ;
        RECT 77.015 152.625 80.525 153.715 ;
        RECT 80.700 153.280 86.045 153.715 ;
        RECT 77.015 152.105 78.705 152.625 ;
        RECT 78.875 151.935 80.525 152.455 ;
        RECT 82.290 152.030 82.640 153.280 ;
        RECT 86.590 152.735 86.845 153.405 ;
        RECT 87.025 152.915 87.310 153.715 ;
        RECT 87.490 152.995 87.820 153.505 ;
        RECT 72.885 151.695 74.245 151.905 ;
        RECT 72.885 151.335 73.215 151.695 ;
        RECT 73.385 151.165 73.715 151.525 ;
        RECT 73.915 151.335 74.245 151.695 ;
        RECT 74.755 151.335 75.465 151.925 ;
        RECT 75.635 151.165 75.925 151.890 ;
        RECT 77.015 151.165 80.525 151.935 ;
        RECT 84.120 151.710 84.460 152.540 ;
        RECT 86.590 151.875 86.770 152.735 ;
        RECT 87.490 152.405 87.740 152.995 ;
        RECT 88.090 152.845 88.260 153.455 ;
        RECT 88.430 153.025 88.760 153.715 ;
        RECT 88.990 153.165 89.230 153.455 ;
        RECT 89.430 153.335 89.850 153.715 ;
        RECT 90.030 153.245 90.660 153.495 ;
        RECT 91.130 153.335 91.460 153.715 ;
        RECT 90.030 153.165 90.200 153.245 ;
        RECT 91.630 153.165 91.800 153.455 ;
        RECT 91.980 153.335 92.360 153.715 ;
        RECT 92.600 153.330 93.430 153.500 ;
        RECT 88.990 152.995 90.200 153.165 ;
        RECT 86.940 152.075 87.740 152.405 ;
        RECT 80.700 151.165 86.045 151.710 ;
        RECT 86.590 151.675 86.845 151.875 ;
        RECT 86.505 151.505 86.845 151.675 ;
        RECT 86.590 151.345 86.845 151.505 ;
        RECT 87.025 151.165 87.310 151.625 ;
        RECT 87.490 151.425 87.740 152.075 ;
        RECT 87.940 152.825 88.260 152.845 ;
        RECT 87.940 152.655 89.860 152.825 ;
        RECT 87.940 151.760 88.130 152.655 ;
        RECT 90.030 152.485 90.200 152.995 ;
        RECT 90.370 152.735 90.890 153.045 ;
        RECT 88.300 152.315 90.200 152.485 ;
        RECT 88.300 152.255 88.630 152.315 ;
        RECT 88.780 152.085 89.110 152.145 ;
        RECT 88.450 151.815 89.110 152.085 ;
        RECT 87.940 151.430 88.260 151.760 ;
        RECT 88.440 151.165 89.100 151.645 ;
        RECT 89.300 151.555 89.470 152.315 ;
        RECT 90.370 152.145 90.550 152.555 ;
        RECT 89.640 151.975 89.970 152.095 ;
        RECT 90.720 151.975 90.890 152.735 ;
        RECT 89.640 151.805 90.890 151.975 ;
        RECT 91.060 152.915 92.430 153.165 ;
        RECT 91.060 152.145 91.250 152.915 ;
        RECT 92.180 152.655 92.430 152.915 ;
        RECT 91.420 152.485 91.670 152.645 ;
        RECT 92.600 152.485 92.770 153.330 ;
        RECT 93.665 153.045 93.835 153.545 ;
        RECT 94.005 153.215 94.335 153.715 ;
        RECT 92.940 152.655 93.440 153.035 ;
        RECT 93.665 152.875 94.360 153.045 ;
        RECT 91.420 152.315 92.770 152.485 ;
        RECT 92.350 152.275 92.770 152.315 ;
        RECT 91.060 151.805 91.480 152.145 ;
        RECT 91.770 151.815 92.180 152.145 ;
        RECT 89.300 151.385 90.150 151.555 ;
        RECT 90.710 151.165 91.030 151.625 ;
        RECT 91.230 151.375 91.480 151.805 ;
        RECT 91.770 151.165 92.180 151.605 ;
        RECT 92.350 151.545 92.520 152.275 ;
        RECT 92.690 151.725 93.040 152.095 ;
        RECT 93.220 151.785 93.440 152.655 ;
        RECT 93.610 152.085 94.020 152.705 ;
        RECT 94.190 151.905 94.360 152.875 ;
        RECT 93.665 151.715 94.360 151.905 ;
        RECT 92.350 151.345 93.365 151.545 ;
        RECT 93.665 151.385 93.835 151.715 ;
        RECT 94.005 151.165 94.335 151.545 ;
        RECT 94.550 151.425 94.775 153.545 ;
        RECT 94.945 153.215 95.275 153.715 ;
        RECT 95.445 153.045 95.615 153.545 ;
        RECT 95.880 153.280 101.225 153.715 ;
        RECT 94.950 152.875 95.615 153.045 ;
        RECT 94.950 151.885 95.180 152.875 ;
        RECT 95.350 152.055 95.700 152.705 ;
        RECT 97.470 152.030 97.820 153.280 ;
        RECT 101.395 152.550 101.685 153.715 ;
        RECT 102.315 152.575 102.585 153.545 ;
        RECT 102.795 152.915 103.075 153.715 ;
        RECT 103.245 153.205 104.900 153.495 ;
        RECT 103.310 152.865 104.900 153.035 ;
        RECT 103.310 152.745 103.480 152.865 ;
        RECT 102.755 152.575 103.480 152.745 ;
        RECT 94.950 151.715 95.615 151.885 ;
        RECT 94.945 151.165 95.275 151.545 ;
        RECT 95.445 151.425 95.615 151.715 ;
        RECT 99.300 151.710 99.640 152.540 ;
        RECT 95.880 151.165 101.225 151.710 ;
        RECT 101.395 151.165 101.685 151.890 ;
        RECT 102.315 151.840 102.485 152.575 ;
        RECT 102.755 152.405 102.925 152.575 ;
        RECT 103.670 152.525 104.385 152.695 ;
        RECT 104.580 152.575 104.900 152.865 ;
        RECT 105.075 152.575 105.415 153.545 ;
        RECT 105.585 152.575 105.755 153.715 ;
        RECT 106.025 152.915 106.275 153.715 ;
        RECT 106.920 152.745 107.250 153.545 ;
        RECT 107.550 152.915 107.880 153.715 ;
        RECT 108.050 152.745 108.380 153.545 ;
        RECT 105.945 152.575 108.380 152.745 ;
        RECT 108.755 152.575 109.095 153.545 ;
        RECT 109.265 152.575 109.435 153.715 ;
        RECT 109.705 152.915 109.955 153.715 ;
        RECT 110.600 152.745 110.930 153.545 ;
        RECT 111.230 152.915 111.560 153.715 ;
        RECT 111.730 152.745 112.060 153.545 ;
        RECT 112.900 153.280 118.245 153.715 ;
        RECT 109.625 152.575 112.060 152.745 ;
        RECT 102.655 152.075 102.925 152.405 ;
        RECT 103.095 152.075 103.500 152.405 ;
        RECT 103.670 152.075 104.380 152.525 ;
        RECT 102.755 151.905 102.925 152.075 ;
        RECT 102.315 151.495 102.585 151.840 ;
        RECT 102.755 151.735 104.365 151.905 ;
        RECT 104.550 151.835 104.900 152.405 ;
        RECT 105.075 151.965 105.250 152.575 ;
        RECT 105.945 152.325 106.115 152.575 ;
        RECT 105.420 152.155 106.115 152.325 ;
        RECT 106.290 152.155 106.710 152.355 ;
        RECT 106.880 152.155 107.210 152.355 ;
        RECT 107.380 152.155 107.710 152.355 ;
        RECT 102.775 151.165 103.155 151.565 ;
        RECT 103.325 151.385 103.495 151.735 ;
        RECT 103.665 151.165 103.995 151.565 ;
        RECT 104.195 151.385 104.365 151.735 ;
        RECT 104.565 151.165 104.895 151.665 ;
        RECT 105.075 151.335 105.415 151.965 ;
        RECT 105.585 151.165 105.835 151.965 ;
        RECT 106.025 151.815 107.250 151.985 ;
        RECT 106.025 151.335 106.355 151.815 ;
        RECT 106.525 151.165 106.750 151.625 ;
        RECT 106.920 151.335 107.250 151.815 ;
        RECT 107.880 151.945 108.050 152.575 ;
        RECT 108.235 152.155 108.585 152.405 ;
        RECT 108.755 152.015 108.930 152.575 ;
        RECT 109.625 152.325 109.795 152.575 ;
        RECT 109.100 152.155 109.795 152.325 ;
        RECT 109.970 152.155 110.390 152.355 ;
        RECT 110.560 152.155 110.890 152.355 ;
        RECT 111.060 152.155 111.390 152.355 ;
        RECT 108.755 151.965 108.985 152.015 ;
        RECT 107.880 151.335 108.380 151.945 ;
        RECT 108.755 151.335 109.095 151.965 ;
        RECT 109.265 151.165 109.515 151.965 ;
        RECT 109.705 151.815 110.930 151.985 ;
        RECT 109.705 151.335 110.035 151.815 ;
        RECT 110.205 151.165 110.430 151.625 ;
        RECT 110.600 151.335 110.930 151.815 ;
        RECT 111.560 151.945 111.730 152.575 ;
        RECT 111.915 152.155 112.265 152.405 ;
        RECT 114.490 152.030 114.840 153.280 ;
        RECT 118.475 152.575 118.685 153.715 ;
        RECT 118.855 152.565 119.185 153.545 ;
        RECT 119.355 152.575 119.585 153.715 ;
        RECT 120.345 152.785 120.515 153.545 ;
        RECT 120.695 152.955 121.025 153.715 ;
        RECT 120.345 152.615 121.010 152.785 ;
        RECT 121.195 152.640 121.465 153.545 ;
        RECT 111.560 151.335 112.060 151.945 ;
        RECT 116.320 151.710 116.660 152.540 ;
        RECT 112.900 151.165 118.245 151.710 ;
        RECT 118.475 151.165 118.685 151.985 ;
        RECT 118.855 151.965 119.105 152.565 ;
        RECT 120.840 152.470 121.010 152.615 ;
        RECT 119.275 152.155 119.605 152.405 ;
        RECT 120.275 152.065 120.605 152.435 ;
        RECT 120.840 152.140 121.125 152.470 ;
        RECT 118.855 151.335 119.185 151.965 ;
        RECT 119.355 151.165 119.585 151.985 ;
        RECT 120.840 151.885 121.010 152.140 ;
        RECT 120.345 151.715 121.010 151.885 ;
        RECT 121.295 151.840 121.465 152.640 ;
        RECT 122.555 152.625 126.065 153.715 ;
        RECT 126.235 152.625 127.445 153.715 ;
        RECT 122.555 152.105 124.245 152.625 ;
        RECT 124.415 151.935 126.065 152.455 ;
        RECT 126.235 152.085 126.755 152.625 ;
        RECT 120.345 151.335 120.515 151.715 ;
        RECT 120.695 151.165 121.025 151.545 ;
        RECT 121.205 151.335 121.465 151.840 ;
        RECT 122.555 151.165 126.065 151.935 ;
        RECT 126.925 151.915 127.445 152.455 ;
        RECT 126.235 151.165 127.445 151.915 ;
        RECT 14.370 150.995 127.530 151.165 ;
        RECT 14.455 150.245 15.665 150.995 ;
        RECT 16.670 150.285 16.925 150.815 ;
        RECT 17.105 150.535 17.390 150.995 ;
        RECT 14.455 149.705 14.975 150.245 ;
        RECT 15.145 149.535 15.665 150.075 ;
        RECT 16.670 149.635 16.850 150.285 ;
        RECT 17.570 150.085 17.820 150.735 ;
        RECT 17.020 149.755 17.820 150.085 ;
        RECT 14.455 148.445 15.665 149.535 ;
        RECT 16.585 149.465 16.850 149.635 ;
        RECT 16.670 149.425 16.850 149.465 ;
        RECT 16.670 148.755 16.925 149.425 ;
        RECT 17.105 148.445 17.390 149.245 ;
        RECT 17.570 149.165 17.820 149.755 ;
        RECT 18.020 150.400 18.340 150.730 ;
        RECT 18.520 150.515 19.180 150.995 ;
        RECT 19.380 150.605 20.230 150.775 ;
        RECT 18.020 149.505 18.210 150.400 ;
        RECT 18.530 150.075 19.190 150.345 ;
        RECT 18.860 150.015 19.190 150.075 ;
        RECT 18.380 149.845 18.710 149.905 ;
        RECT 19.380 149.845 19.550 150.605 ;
        RECT 20.790 150.535 21.110 150.995 ;
        RECT 21.310 150.355 21.560 150.785 ;
        RECT 21.850 150.555 22.260 150.995 ;
        RECT 22.430 150.615 23.445 150.815 ;
        RECT 19.720 150.185 20.970 150.355 ;
        RECT 19.720 150.065 20.050 150.185 ;
        RECT 18.380 149.675 20.280 149.845 ;
        RECT 18.020 149.335 19.940 149.505 ;
        RECT 18.020 149.315 18.340 149.335 ;
        RECT 17.570 148.655 17.900 149.165 ;
        RECT 18.170 148.705 18.340 149.315 ;
        RECT 20.110 149.165 20.280 149.675 ;
        RECT 20.450 149.605 20.630 150.015 ;
        RECT 20.800 149.425 20.970 150.185 ;
        RECT 18.510 148.445 18.840 149.135 ;
        RECT 19.070 148.995 20.280 149.165 ;
        RECT 20.450 149.115 20.970 149.425 ;
        RECT 21.140 150.015 21.560 150.355 ;
        RECT 21.850 150.015 22.260 150.345 ;
        RECT 21.140 149.245 21.330 150.015 ;
        RECT 22.430 149.885 22.600 150.615 ;
        RECT 23.745 150.445 23.915 150.775 ;
        RECT 24.085 150.615 24.415 150.995 ;
        RECT 22.770 150.065 23.120 150.435 ;
        RECT 22.430 149.845 22.850 149.885 ;
        RECT 21.500 149.675 22.850 149.845 ;
        RECT 21.500 149.515 21.750 149.675 ;
        RECT 22.260 149.245 22.510 149.505 ;
        RECT 21.140 148.995 22.510 149.245 ;
        RECT 19.070 148.705 19.310 148.995 ;
        RECT 20.110 148.915 20.280 148.995 ;
        RECT 19.510 148.445 19.930 148.825 ;
        RECT 20.110 148.665 20.740 148.915 ;
        RECT 21.210 148.445 21.540 148.825 ;
        RECT 21.710 148.705 21.880 148.995 ;
        RECT 22.680 148.830 22.850 149.675 ;
        RECT 23.300 149.505 23.520 150.375 ;
        RECT 23.745 150.255 24.440 150.445 ;
        RECT 23.020 149.125 23.520 149.505 ;
        RECT 23.690 149.455 24.100 150.075 ;
        RECT 24.270 149.285 24.440 150.255 ;
        RECT 23.745 149.115 24.440 149.285 ;
        RECT 22.060 148.445 22.440 148.825 ;
        RECT 22.680 148.660 23.510 148.830 ;
        RECT 23.745 148.615 23.915 149.115 ;
        RECT 24.085 148.445 24.415 148.945 ;
        RECT 24.630 148.615 24.855 150.735 ;
        RECT 25.025 150.615 25.355 150.995 ;
        RECT 25.525 150.445 25.695 150.735 ;
        RECT 25.030 150.275 25.695 150.445 ;
        RECT 25.030 149.285 25.260 150.275 ;
        RECT 25.955 150.245 27.165 150.995 ;
        RECT 27.340 150.450 32.685 150.995 ;
        RECT 25.430 149.455 25.780 150.105 ;
        RECT 25.955 149.535 26.475 150.075 ;
        RECT 26.645 149.705 27.165 150.245 ;
        RECT 25.030 149.115 25.695 149.285 ;
        RECT 25.025 148.445 25.355 148.945 ;
        RECT 25.525 148.615 25.695 149.115 ;
        RECT 25.955 148.445 27.165 149.535 ;
        RECT 28.930 148.880 29.280 150.130 ;
        RECT 30.760 149.620 31.100 150.450 ;
        RECT 32.895 150.175 33.125 150.995 ;
        RECT 33.295 150.195 33.625 150.825 ;
        RECT 32.875 149.755 33.205 150.005 ;
        RECT 33.375 149.595 33.625 150.195 ;
        RECT 33.795 150.175 34.005 150.995 ;
        RECT 34.235 150.245 35.445 150.995 ;
        RECT 35.705 150.445 35.875 150.825 ;
        RECT 36.055 150.615 36.385 150.995 ;
        RECT 35.705 150.275 36.370 150.445 ;
        RECT 36.565 150.320 36.825 150.825 ;
        RECT 27.340 148.445 32.685 148.880 ;
        RECT 32.895 148.445 33.125 149.585 ;
        RECT 33.295 148.615 33.625 149.595 ;
        RECT 33.795 148.445 34.005 149.585 ;
        RECT 34.235 149.535 34.755 150.075 ;
        RECT 34.925 149.705 35.445 150.245 ;
        RECT 35.635 149.725 35.965 150.095 ;
        RECT 36.200 150.020 36.370 150.275 ;
        RECT 36.200 149.690 36.485 150.020 ;
        RECT 36.200 149.545 36.370 149.690 ;
        RECT 34.235 148.445 35.445 149.535 ;
        RECT 35.705 149.375 36.370 149.545 ;
        RECT 36.655 149.520 36.825 150.320 ;
        RECT 36.995 150.270 37.285 150.995 ;
        RECT 37.455 150.225 40.965 150.995 ;
        RECT 35.705 148.615 35.875 149.375 ;
        RECT 36.055 148.445 36.385 149.205 ;
        RECT 36.555 148.615 36.825 149.520 ;
        RECT 36.995 148.445 37.285 149.610 ;
        RECT 37.455 149.535 39.145 150.055 ;
        RECT 39.315 149.705 40.965 150.225 ;
        RECT 41.135 150.195 41.475 150.825 ;
        RECT 41.645 150.195 41.895 150.995 ;
        RECT 42.085 150.345 42.415 150.825 ;
        RECT 42.585 150.535 42.810 150.995 ;
        RECT 42.980 150.345 43.310 150.825 ;
        RECT 41.135 149.585 41.310 150.195 ;
        RECT 42.085 150.175 43.310 150.345 ;
        RECT 43.940 150.215 44.440 150.825 ;
        RECT 44.815 150.225 48.325 150.995 ;
        RECT 48.505 150.495 48.835 150.995 ;
        RECT 49.035 150.425 49.205 150.775 ;
        RECT 49.405 150.595 49.735 150.995 ;
        RECT 49.905 150.425 50.075 150.775 ;
        RECT 50.245 150.595 50.625 150.995 ;
        RECT 41.480 149.835 42.175 150.005 ;
        RECT 42.005 149.585 42.175 149.835 ;
        RECT 42.350 149.805 42.770 150.005 ;
        RECT 42.940 149.805 43.270 150.005 ;
        RECT 43.440 149.805 43.770 150.005 ;
        RECT 43.940 149.585 44.110 150.215 ;
        RECT 44.295 149.755 44.645 150.005 ;
        RECT 37.455 148.445 40.965 149.535 ;
        RECT 41.135 148.615 41.475 149.585 ;
        RECT 41.645 148.445 41.815 149.585 ;
        RECT 42.005 149.415 44.440 149.585 ;
        RECT 42.085 148.445 42.335 149.245 ;
        RECT 42.980 148.615 43.310 149.415 ;
        RECT 43.610 148.445 43.940 149.245 ;
        RECT 44.110 148.615 44.440 149.415 ;
        RECT 44.815 149.535 46.505 150.055 ;
        RECT 46.675 149.705 48.325 150.225 ;
        RECT 48.500 149.755 48.850 150.325 ;
        RECT 49.035 150.255 50.645 150.425 ;
        RECT 50.815 150.320 51.085 150.665 ;
        RECT 50.475 150.085 50.645 150.255 ;
        RECT 44.815 148.445 48.325 149.535 ;
        RECT 48.500 149.295 48.820 149.585 ;
        RECT 49.020 149.465 49.730 150.085 ;
        RECT 49.900 149.755 50.305 150.085 ;
        RECT 50.475 149.755 50.745 150.085 ;
        RECT 50.475 149.585 50.645 149.755 ;
        RECT 50.915 149.585 51.085 150.320 ;
        RECT 49.920 149.415 50.645 149.585 ;
        RECT 49.920 149.295 50.090 149.415 ;
        RECT 48.500 149.125 50.090 149.295 ;
        RECT 48.500 148.665 50.155 148.955 ;
        RECT 50.325 148.445 50.605 149.245 ;
        RECT 50.815 148.615 51.085 149.585 ;
        RECT 51.255 150.195 51.595 150.825 ;
        RECT 51.765 150.195 52.015 150.995 ;
        RECT 52.205 150.345 52.535 150.825 ;
        RECT 52.705 150.535 52.930 150.995 ;
        RECT 53.100 150.345 53.430 150.825 ;
        RECT 51.255 149.585 51.430 150.195 ;
        RECT 52.205 150.175 53.430 150.345 ;
        RECT 54.060 150.215 54.560 150.825 ;
        RECT 54.935 150.225 56.605 150.995 ;
        RECT 51.600 149.835 52.295 150.005 ;
        RECT 52.125 149.585 52.295 149.835 ;
        RECT 52.470 149.805 52.890 150.005 ;
        RECT 53.060 149.805 53.390 150.005 ;
        RECT 53.560 149.805 53.890 150.005 ;
        RECT 54.060 149.585 54.230 150.215 ;
        RECT 54.415 149.755 54.765 150.005 ;
        RECT 51.255 148.615 51.595 149.585 ;
        RECT 51.765 148.445 51.935 149.585 ;
        RECT 52.125 149.415 54.560 149.585 ;
        RECT 52.205 148.445 52.455 149.245 ;
        RECT 53.100 148.615 53.430 149.415 ;
        RECT 53.730 148.445 54.060 149.245 ;
        RECT 54.230 148.615 54.560 149.415 ;
        RECT 54.935 149.535 55.685 150.055 ;
        RECT 55.855 149.705 56.605 150.225 ;
        RECT 57.050 150.185 57.295 150.790 ;
        RECT 57.515 150.460 58.025 150.995 ;
        RECT 56.775 150.015 58.005 150.185 ;
        RECT 54.935 148.445 56.605 149.535 ;
        RECT 56.775 149.205 57.115 150.015 ;
        RECT 57.285 149.450 58.035 149.640 ;
        RECT 56.775 148.795 57.290 149.205 ;
        RECT 57.525 148.445 57.695 149.205 ;
        RECT 57.865 148.785 58.035 149.450 ;
        RECT 58.205 149.465 58.395 150.825 ;
        RECT 58.565 149.975 58.840 150.825 ;
        RECT 59.030 150.460 59.560 150.825 ;
        RECT 59.985 150.595 60.315 150.995 ;
        RECT 59.385 150.425 59.560 150.460 ;
        RECT 58.565 149.805 58.845 149.975 ;
        RECT 58.565 149.665 58.840 149.805 ;
        RECT 59.045 149.465 59.215 150.265 ;
        RECT 58.205 149.295 59.215 149.465 ;
        RECT 59.385 150.255 60.315 150.425 ;
        RECT 60.485 150.255 60.740 150.825 ;
        RECT 59.385 149.125 59.555 150.255 ;
        RECT 60.145 150.085 60.315 150.255 ;
        RECT 58.430 148.955 59.555 149.125 ;
        RECT 59.725 149.755 59.920 150.085 ;
        RECT 60.145 149.755 60.400 150.085 ;
        RECT 59.725 148.785 59.895 149.755 ;
        RECT 60.570 149.585 60.740 150.255 ;
        RECT 57.865 148.615 59.895 148.785 ;
        RECT 60.065 148.445 60.235 149.585 ;
        RECT 60.405 148.615 60.740 149.585 ;
        RECT 61.375 150.320 61.635 150.825 ;
        RECT 61.815 150.615 62.145 150.995 ;
        RECT 62.325 150.445 62.495 150.825 ;
        RECT 61.375 149.520 61.545 150.320 ;
        RECT 61.830 150.275 62.495 150.445 ;
        RECT 61.830 150.020 62.000 150.275 ;
        RECT 62.755 150.270 63.045 150.995 ;
        RECT 63.765 150.445 63.935 150.825 ;
        RECT 64.115 150.615 64.445 150.995 ;
        RECT 63.765 150.275 64.430 150.445 ;
        RECT 64.625 150.320 64.885 150.825 ;
        RECT 61.715 149.690 62.000 150.020 ;
        RECT 62.235 149.725 62.565 150.095 ;
        RECT 63.695 149.725 64.025 150.095 ;
        RECT 64.260 150.020 64.430 150.275 ;
        RECT 61.830 149.545 62.000 149.690 ;
        RECT 64.260 149.690 64.545 150.020 ;
        RECT 61.375 148.615 61.645 149.520 ;
        RECT 61.830 149.375 62.495 149.545 ;
        RECT 61.815 148.445 62.145 149.205 ;
        RECT 62.325 148.615 62.495 149.375 ;
        RECT 62.755 148.445 63.045 149.610 ;
        RECT 64.260 149.545 64.430 149.690 ;
        RECT 63.765 149.375 64.430 149.545 ;
        RECT 64.715 149.520 64.885 150.320 ;
        RECT 65.515 150.225 67.185 150.995 ;
        RECT 67.445 150.445 67.615 150.825 ;
        RECT 67.830 150.615 68.160 150.995 ;
        RECT 67.445 150.275 68.160 150.445 ;
        RECT 63.765 148.615 63.935 149.375 ;
        RECT 64.115 148.445 64.445 149.205 ;
        RECT 64.615 148.615 64.885 149.520 ;
        RECT 65.515 149.535 66.265 150.055 ;
        RECT 66.435 149.705 67.185 150.225 ;
        RECT 67.355 149.725 67.710 150.095 ;
        RECT 67.990 150.085 68.160 150.275 ;
        RECT 68.330 150.250 68.585 150.825 ;
        RECT 67.990 149.755 68.245 150.085 ;
        RECT 67.990 149.545 68.160 149.755 ;
        RECT 65.515 148.445 67.185 149.535 ;
        RECT 67.445 149.375 68.160 149.545 ;
        RECT 68.415 149.520 68.585 150.250 ;
        RECT 68.760 150.155 69.020 150.995 ;
        RECT 69.200 150.155 69.460 150.995 ;
        RECT 69.635 150.250 69.890 150.825 ;
        RECT 70.060 150.615 70.390 150.995 ;
        RECT 70.605 150.445 70.775 150.825 ;
        RECT 71.095 150.515 71.375 150.995 ;
        RECT 70.060 150.275 70.775 150.445 ;
        RECT 71.545 150.345 71.805 150.735 ;
        RECT 71.980 150.515 72.235 150.995 ;
        RECT 72.405 150.345 72.700 150.735 ;
        RECT 72.880 150.515 73.155 150.995 ;
        RECT 73.325 150.495 73.625 150.825 ;
        RECT 67.445 148.615 67.615 149.375 ;
        RECT 67.830 148.445 68.160 149.205 ;
        RECT 68.330 148.615 68.585 149.520 ;
        RECT 68.760 148.445 69.020 149.595 ;
        RECT 69.200 148.445 69.460 149.595 ;
        RECT 69.635 149.520 69.805 150.250 ;
        RECT 70.060 150.085 70.230 150.275 ;
        RECT 71.050 150.175 72.700 150.345 ;
        RECT 69.975 149.755 70.230 150.085 ;
        RECT 70.060 149.545 70.230 149.755 ;
        RECT 70.510 149.725 70.865 150.095 ;
        RECT 71.050 149.665 71.455 150.175 ;
        RECT 71.625 149.835 72.765 150.005 ;
        RECT 69.635 148.615 69.890 149.520 ;
        RECT 70.060 149.375 70.775 149.545 ;
        RECT 71.050 149.495 71.805 149.665 ;
        RECT 70.060 148.445 70.390 149.205 ;
        RECT 70.605 148.615 70.775 149.375 ;
        RECT 71.090 148.445 71.375 149.315 ;
        RECT 71.545 149.245 71.805 149.495 ;
        RECT 72.595 149.585 72.765 149.835 ;
        RECT 72.935 149.755 73.285 150.325 ;
        RECT 73.455 149.585 73.625 150.495 ;
        RECT 72.595 149.415 73.625 149.585 ;
        RECT 71.545 149.075 72.665 149.245 ;
        RECT 71.545 148.615 71.805 149.075 ;
        RECT 71.980 148.445 72.235 148.905 ;
        RECT 72.405 148.615 72.665 149.075 ;
        RECT 72.835 148.445 73.145 149.245 ;
        RECT 73.315 148.615 73.625 149.415 ;
        RECT 74.715 150.495 75.015 150.825 ;
        RECT 75.185 150.515 75.460 150.995 ;
        RECT 74.715 149.585 74.885 150.495 ;
        RECT 75.640 150.345 75.935 150.735 ;
        RECT 76.105 150.515 76.360 150.995 ;
        RECT 76.535 150.345 76.795 150.735 ;
        RECT 76.965 150.515 77.245 150.995 ;
        RECT 75.055 149.755 75.405 150.325 ;
        RECT 75.640 150.175 77.290 150.345 ;
        RECT 75.575 149.835 76.715 150.005 ;
        RECT 75.575 149.585 75.745 149.835 ;
        RECT 76.885 149.665 77.290 150.175 ;
        RECT 74.715 149.415 75.745 149.585 ;
        RECT 76.535 149.495 77.290 149.665 ;
        RECT 77.475 150.320 77.745 150.665 ;
        RECT 77.935 150.595 78.315 150.995 ;
        RECT 78.485 150.425 78.655 150.775 ;
        RECT 78.825 150.595 79.155 150.995 ;
        RECT 79.355 150.425 79.525 150.775 ;
        RECT 79.725 150.495 80.055 150.995 ;
        RECT 77.475 149.585 77.645 150.320 ;
        RECT 77.915 150.255 79.525 150.425 ;
        RECT 77.915 150.085 78.085 150.255 ;
        RECT 77.815 149.755 78.085 150.085 ;
        RECT 78.255 149.755 78.660 150.085 ;
        RECT 77.915 149.585 78.085 149.755 ;
        RECT 78.830 149.635 79.540 150.085 ;
        RECT 79.710 149.755 80.060 150.325 ;
        RECT 80.695 150.225 84.205 150.995 ;
        RECT 74.715 148.615 75.025 149.415 ;
        RECT 76.535 149.245 76.795 149.495 ;
        RECT 75.195 148.445 75.505 149.245 ;
        RECT 75.675 149.075 76.795 149.245 ;
        RECT 75.675 148.615 75.935 149.075 ;
        RECT 76.105 148.445 76.360 148.905 ;
        RECT 76.535 148.615 76.795 149.075 ;
        RECT 76.965 148.445 77.250 149.315 ;
        RECT 77.475 148.615 77.745 149.585 ;
        RECT 77.915 149.415 78.640 149.585 ;
        RECT 78.830 149.465 79.545 149.635 ;
        RECT 78.470 149.295 78.640 149.415 ;
        RECT 79.740 149.295 80.060 149.585 ;
        RECT 77.955 148.445 78.235 149.245 ;
        RECT 78.470 149.125 80.060 149.295 ;
        RECT 80.695 149.535 82.385 150.055 ;
        RECT 82.555 149.705 84.205 150.225 ;
        RECT 84.650 150.185 84.895 150.790 ;
        RECT 85.115 150.460 85.625 150.995 ;
        RECT 84.375 150.015 85.605 150.185 ;
        RECT 78.405 148.665 80.060 148.955 ;
        RECT 80.695 148.445 84.205 149.535 ;
        RECT 84.375 149.205 84.715 150.015 ;
        RECT 84.885 149.450 85.635 149.640 ;
        RECT 84.375 148.795 84.890 149.205 ;
        RECT 85.125 148.445 85.295 149.205 ;
        RECT 85.465 148.785 85.635 149.450 ;
        RECT 85.805 149.465 85.995 150.825 ;
        RECT 86.165 149.975 86.440 150.825 ;
        RECT 86.630 150.460 87.160 150.825 ;
        RECT 87.585 150.595 87.915 150.995 ;
        RECT 86.985 150.425 87.160 150.460 ;
        RECT 86.165 149.805 86.445 149.975 ;
        RECT 86.165 149.665 86.440 149.805 ;
        RECT 86.645 149.465 86.815 150.265 ;
        RECT 85.805 149.295 86.815 149.465 ;
        RECT 86.985 150.255 87.915 150.425 ;
        RECT 88.085 150.255 88.340 150.825 ;
        RECT 88.515 150.270 88.805 150.995 ;
        RECT 86.985 149.125 87.155 150.255 ;
        RECT 87.745 150.085 87.915 150.255 ;
        RECT 86.030 148.955 87.155 149.125 ;
        RECT 87.325 149.755 87.520 150.085 ;
        RECT 87.745 149.755 88.000 150.085 ;
        RECT 87.325 148.785 87.495 149.755 ;
        RECT 88.170 149.585 88.340 150.255 ;
        RECT 89.495 150.175 89.705 150.995 ;
        RECT 89.875 150.195 90.205 150.825 ;
        RECT 85.465 148.615 87.495 148.785 ;
        RECT 87.665 148.445 87.835 149.585 ;
        RECT 88.005 148.615 88.340 149.585 ;
        RECT 88.515 148.445 88.805 149.610 ;
        RECT 89.875 149.595 90.125 150.195 ;
        RECT 90.375 150.175 90.605 150.995 ;
        RECT 91.825 150.445 91.995 150.825 ;
        RECT 92.175 150.615 92.505 150.995 ;
        RECT 91.825 150.275 92.490 150.445 ;
        RECT 92.685 150.320 92.945 150.825 ;
        RECT 90.295 149.755 90.625 150.005 ;
        RECT 91.755 149.725 92.085 150.095 ;
        RECT 92.320 150.020 92.490 150.275 ;
        RECT 92.320 149.690 92.605 150.020 ;
        RECT 89.495 148.445 89.705 149.585 ;
        RECT 89.875 148.615 90.205 149.595 ;
        RECT 90.375 148.445 90.605 149.585 ;
        RECT 92.320 149.545 92.490 149.690 ;
        RECT 91.825 149.375 92.490 149.545 ;
        RECT 92.775 149.520 92.945 150.320 ;
        RECT 93.175 150.175 93.385 150.995 ;
        RECT 93.555 150.195 93.885 150.825 ;
        RECT 93.555 149.595 93.805 150.195 ;
        RECT 94.055 150.175 94.285 150.995 ;
        RECT 94.495 150.225 96.165 150.995 ;
        RECT 93.975 149.755 94.305 150.005 ;
        RECT 91.825 148.615 91.995 149.375 ;
        RECT 92.175 148.445 92.505 149.205 ;
        RECT 92.675 148.615 92.945 149.520 ;
        RECT 93.175 148.445 93.385 149.585 ;
        RECT 93.555 148.615 93.885 149.595 ;
        RECT 94.055 148.445 94.285 149.585 ;
        RECT 94.495 149.535 95.245 150.055 ;
        RECT 95.415 149.705 96.165 150.225 ;
        RECT 96.340 150.285 96.595 150.815 ;
        RECT 96.765 150.535 97.070 150.995 ;
        RECT 97.315 150.615 98.385 150.785 ;
        RECT 96.340 149.635 96.550 150.285 ;
        RECT 97.315 150.260 97.635 150.615 ;
        RECT 97.310 150.085 97.635 150.260 ;
        RECT 96.720 149.785 97.635 150.085 ;
        RECT 97.805 150.045 98.045 150.445 ;
        RECT 98.215 150.385 98.385 150.615 ;
        RECT 98.555 150.555 98.745 150.995 ;
        RECT 98.915 150.545 99.865 150.825 ;
        RECT 100.085 150.635 100.435 150.805 ;
        RECT 98.215 150.215 98.745 150.385 ;
        RECT 96.720 149.755 97.460 149.785 ;
        RECT 94.495 148.445 96.165 149.535 ;
        RECT 96.340 148.755 96.595 149.635 ;
        RECT 96.765 148.445 97.070 149.585 ;
        RECT 97.290 149.165 97.460 149.755 ;
        RECT 97.805 149.675 98.345 150.045 ;
        RECT 98.525 149.935 98.745 150.215 ;
        RECT 98.915 149.765 99.085 150.545 ;
        RECT 98.680 149.595 99.085 149.765 ;
        RECT 99.255 149.755 99.605 150.375 ;
        RECT 98.680 149.505 98.850 149.595 ;
        RECT 99.775 149.585 99.985 150.375 ;
        RECT 97.630 149.335 98.850 149.505 ;
        RECT 99.310 149.425 99.985 149.585 ;
        RECT 97.290 148.995 98.090 149.165 ;
        RECT 97.410 148.445 97.740 148.825 ;
        RECT 97.920 148.705 98.090 148.995 ;
        RECT 98.680 148.955 98.850 149.335 ;
        RECT 99.020 149.415 99.985 149.425 ;
        RECT 100.175 150.245 100.435 150.635 ;
        RECT 100.645 150.535 100.975 150.995 ;
        RECT 101.850 150.605 102.705 150.775 ;
        RECT 102.910 150.605 103.405 150.775 ;
        RECT 103.575 150.635 103.905 150.995 ;
        RECT 100.175 149.555 100.345 150.245 ;
        RECT 100.515 149.895 100.685 150.075 ;
        RECT 100.855 150.065 101.645 150.315 ;
        RECT 101.850 149.895 102.020 150.605 ;
        RECT 102.190 150.095 102.545 150.315 ;
        RECT 100.515 149.725 102.205 149.895 ;
        RECT 99.020 149.125 99.480 149.415 ;
        RECT 100.175 149.385 101.675 149.555 ;
        RECT 100.175 149.245 100.345 149.385 ;
        RECT 99.785 149.075 100.345 149.245 ;
        RECT 98.260 148.445 98.510 148.905 ;
        RECT 98.680 148.615 99.550 148.955 ;
        RECT 99.785 148.615 99.955 149.075 ;
        RECT 100.790 149.045 101.865 149.215 ;
        RECT 100.125 148.445 100.495 148.905 ;
        RECT 100.790 148.705 100.960 149.045 ;
        RECT 101.130 148.445 101.460 148.875 ;
        RECT 101.695 148.705 101.865 149.045 ;
        RECT 102.035 148.945 102.205 149.725 ;
        RECT 102.375 149.505 102.545 150.095 ;
        RECT 102.715 149.695 103.065 150.315 ;
        RECT 102.375 149.115 102.840 149.505 ;
        RECT 103.235 149.245 103.405 150.605 ;
        RECT 103.575 149.415 104.035 150.465 ;
        RECT 103.010 149.075 103.405 149.245 ;
        RECT 103.010 148.945 103.180 149.075 ;
        RECT 102.035 148.615 102.715 148.945 ;
        RECT 102.930 148.615 103.180 148.945 ;
        RECT 103.350 148.445 103.600 148.905 ;
        RECT 103.770 148.630 104.095 149.415 ;
        RECT 104.265 148.615 104.435 150.735 ;
        RECT 104.605 150.615 104.935 150.995 ;
        RECT 105.105 150.445 105.360 150.735 ;
        RECT 104.610 150.275 105.360 150.445 ;
        RECT 104.610 149.285 104.840 150.275 ;
        RECT 105.535 150.245 106.745 150.995 ;
        RECT 105.010 149.455 105.360 150.105 ;
        RECT 105.535 149.535 106.055 150.075 ;
        RECT 106.225 149.705 106.745 150.245 ;
        RECT 106.915 150.195 107.255 150.825 ;
        RECT 107.425 150.195 107.675 150.995 ;
        RECT 107.865 150.345 108.195 150.825 ;
        RECT 108.365 150.535 108.590 150.995 ;
        RECT 108.760 150.345 109.090 150.825 ;
        RECT 106.915 149.585 107.090 150.195 ;
        RECT 107.865 150.175 109.090 150.345 ;
        RECT 109.720 150.215 110.220 150.825 ;
        RECT 110.710 150.365 110.995 150.825 ;
        RECT 111.165 150.535 111.435 150.995 ;
        RECT 107.260 149.835 107.955 150.005 ;
        RECT 107.785 149.585 107.955 149.835 ;
        RECT 108.130 149.805 108.550 150.005 ;
        RECT 108.720 149.805 109.050 150.005 ;
        RECT 109.220 149.805 109.550 150.005 ;
        RECT 109.720 149.585 109.890 150.215 ;
        RECT 110.710 150.195 111.665 150.365 ;
        RECT 110.075 149.755 110.425 150.005 ;
        RECT 104.610 149.115 105.360 149.285 ;
        RECT 104.605 148.445 104.935 148.945 ;
        RECT 105.105 148.615 105.360 149.115 ;
        RECT 105.535 148.445 106.745 149.535 ;
        RECT 106.915 148.615 107.255 149.585 ;
        RECT 107.425 148.445 107.595 149.585 ;
        RECT 107.785 149.415 110.220 149.585 ;
        RECT 110.595 149.465 111.285 150.025 ;
        RECT 107.865 148.445 108.115 149.245 ;
        RECT 108.760 148.615 109.090 149.415 ;
        RECT 109.390 148.445 109.720 149.245 ;
        RECT 109.890 148.615 110.220 149.415 ;
        RECT 111.455 149.295 111.665 150.195 ;
        RECT 110.710 149.075 111.665 149.295 ;
        RECT 111.835 150.025 112.235 150.825 ;
        RECT 112.425 150.365 112.705 150.825 ;
        RECT 113.225 150.535 113.550 150.995 ;
        RECT 112.425 150.195 113.550 150.365 ;
        RECT 113.720 150.255 114.105 150.825 ;
        RECT 114.275 150.270 114.565 150.995 ;
        RECT 115.660 150.285 115.915 150.815 ;
        RECT 116.085 150.535 116.390 150.995 ;
        RECT 116.635 150.615 117.705 150.785 ;
        RECT 113.100 150.085 113.550 150.195 ;
        RECT 111.835 149.465 112.930 150.025 ;
        RECT 113.100 149.755 113.655 150.085 ;
        RECT 110.710 148.615 110.995 149.075 ;
        RECT 111.165 148.445 111.435 148.905 ;
        RECT 111.835 148.615 112.235 149.465 ;
        RECT 113.100 149.295 113.550 149.755 ;
        RECT 113.825 149.585 114.105 150.255 ;
        RECT 115.660 149.635 115.870 150.285 ;
        RECT 116.635 150.260 116.955 150.615 ;
        RECT 116.630 150.085 116.955 150.260 ;
        RECT 116.040 149.785 116.955 150.085 ;
        RECT 117.125 150.045 117.365 150.445 ;
        RECT 117.535 150.385 117.705 150.615 ;
        RECT 117.875 150.555 118.065 150.995 ;
        RECT 118.235 150.545 119.185 150.825 ;
        RECT 119.405 150.635 119.755 150.805 ;
        RECT 117.535 150.215 118.065 150.385 ;
        RECT 116.040 149.755 116.780 149.785 ;
        RECT 112.425 149.075 113.550 149.295 ;
        RECT 112.425 148.615 112.705 149.075 ;
        RECT 113.225 148.445 113.550 148.905 ;
        RECT 113.720 148.615 114.105 149.585 ;
        RECT 114.275 148.445 114.565 149.610 ;
        RECT 115.660 148.755 115.915 149.635 ;
        RECT 116.085 148.445 116.390 149.585 ;
        RECT 116.610 149.165 116.780 149.755 ;
        RECT 117.125 149.675 117.665 150.045 ;
        RECT 117.845 149.935 118.065 150.215 ;
        RECT 118.235 149.765 118.405 150.545 ;
        RECT 118.000 149.595 118.405 149.765 ;
        RECT 118.575 149.755 118.925 150.375 ;
        RECT 118.000 149.505 118.170 149.595 ;
        RECT 119.095 149.585 119.305 150.375 ;
        RECT 116.950 149.335 118.170 149.505 ;
        RECT 118.630 149.425 119.305 149.585 ;
        RECT 116.610 148.995 117.410 149.165 ;
        RECT 116.730 148.445 117.060 148.825 ;
        RECT 117.240 148.705 117.410 148.995 ;
        RECT 118.000 148.955 118.170 149.335 ;
        RECT 118.340 149.415 119.305 149.425 ;
        RECT 119.495 150.245 119.755 150.635 ;
        RECT 119.965 150.535 120.295 150.995 ;
        RECT 121.170 150.605 122.025 150.775 ;
        RECT 122.230 150.605 122.725 150.775 ;
        RECT 122.895 150.635 123.225 150.995 ;
        RECT 119.495 149.555 119.665 150.245 ;
        RECT 119.835 149.895 120.005 150.075 ;
        RECT 120.175 150.065 120.965 150.315 ;
        RECT 121.170 149.895 121.340 150.605 ;
        RECT 121.510 150.095 121.865 150.315 ;
        RECT 119.835 149.725 121.525 149.895 ;
        RECT 118.340 149.125 118.800 149.415 ;
        RECT 119.495 149.385 120.995 149.555 ;
        RECT 119.495 149.245 119.665 149.385 ;
        RECT 119.105 149.075 119.665 149.245 ;
        RECT 117.580 148.445 117.830 148.905 ;
        RECT 118.000 148.615 118.870 148.955 ;
        RECT 119.105 148.615 119.275 149.075 ;
        RECT 120.110 149.045 121.185 149.215 ;
        RECT 119.445 148.445 119.815 148.905 ;
        RECT 120.110 148.705 120.280 149.045 ;
        RECT 120.450 148.445 120.780 148.875 ;
        RECT 121.015 148.705 121.185 149.045 ;
        RECT 121.355 148.945 121.525 149.725 ;
        RECT 121.695 149.505 121.865 150.095 ;
        RECT 122.035 149.695 122.385 150.315 ;
        RECT 121.695 149.115 122.160 149.505 ;
        RECT 122.555 149.245 122.725 150.605 ;
        RECT 122.895 149.415 123.355 150.465 ;
        RECT 122.330 149.075 122.725 149.245 ;
        RECT 122.330 148.945 122.500 149.075 ;
        RECT 121.355 148.615 122.035 148.945 ;
        RECT 122.250 148.615 122.500 148.945 ;
        RECT 122.670 148.445 122.920 148.905 ;
        RECT 123.090 148.630 123.415 149.415 ;
        RECT 123.585 148.615 123.755 150.735 ;
        RECT 123.925 150.615 124.255 150.995 ;
        RECT 124.425 150.445 124.680 150.735 ;
        RECT 123.930 150.275 124.680 150.445 ;
        RECT 123.930 149.285 124.160 150.275 ;
        RECT 124.855 150.245 126.065 150.995 ;
        RECT 126.235 150.245 127.445 150.995 ;
        RECT 124.330 149.455 124.680 150.105 ;
        RECT 124.855 149.535 125.375 150.075 ;
        RECT 125.545 149.705 126.065 150.245 ;
        RECT 126.235 149.535 126.755 150.075 ;
        RECT 126.925 149.705 127.445 150.245 ;
        RECT 123.930 149.115 124.680 149.285 ;
        RECT 123.925 148.445 124.255 148.945 ;
        RECT 124.425 148.615 124.680 149.115 ;
        RECT 124.855 148.445 126.065 149.535 ;
        RECT 126.235 148.445 127.445 149.535 ;
        RECT 14.370 148.275 127.530 148.445 ;
        RECT 14.455 147.185 15.665 148.275 ;
        RECT 14.455 146.475 14.975 147.015 ;
        RECT 15.145 146.645 15.665 147.185 ;
        RECT 16.295 147.185 19.805 148.275 ;
        RECT 19.975 147.515 20.490 147.925 ;
        RECT 20.725 147.515 20.895 148.275 ;
        RECT 21.065 147.935 23.095 148.105 ;
        RECT 16.295 146.665 17.985 147.185 ;
        RECT 18.155 146.495 19.805 147.015 ;
        RECT 19.975 146.705 20.315 147.515 ;
        RECT 21.065 147.270 21.235 147.935 ;
        RECT 21.630 147.595 22.755 147.765 ;
        RECT 20.485 147.080 21.235 147.270 ;
        RECT 21.405 147.255 22.415 147.425 ;
        RECT 19.975 146.535 21.205 146.705 ;
        RECT 14.455 145.725 15.665 146.475 ;
        RECT 16.295 145.725 19.805 146.495 ;
        RECT 20.250 145.930 20.495 146.535 ;
        RECT 20.715 145.725 21.225 146.260 ;
        RECT 21.405 145.895 21.595 147.255 ;
        RECT 21.765 146.575 22.040 147.055 ;
        RECT 21.765 146.405 22.045 146.575 ;
        RECT 22.245 146.455 22.415 147.255 ;
        RECT 22.585 146.465 22.755 147.595 ;
        RECT 22.925 146.965 23.095 147.935 ;
        RECT 23.265 147.135 23.435 148.275 ;
        RECT 23.605 147.135 23.940 148.105 ;
        RECT 22.925 146.635 23.120 146.965 ;
        RECT 23.345 146.635 23.600 146.965 ;
        RECT 23.345 146.465 23.515 146.635 ;
        RECT 23.770 146.465 23.940 147.135 ;
        RECT 24.115 147.110 24.405 148.275 ;
        RECT 24.575 147.200 24.845 148.105 ;
        RECT 25.015 147.515 25.345 148.275 ;
        RECT 25.525 147.345 25.695 148.105 ;
        RECT 21.765 145.895 22.040 146.405 ;
        RECT 22.585 146.295 23.515 146.465 ;
        RECT 22.585 146.260 22.760 146.295 ;
        RECT 22.230 145.895 22.760 146.260 ;
        RECT 23.185 145.725 23.515 146.125 ;
        RECT 23.685 145.895 23.940 146.465 ;
        RECT 24.115 145.725 24.405 146.450 ;
        RECT 24.575 146.400 24.745 147.200 ;
        RECT 25.030 147.175 25.695 147.345 ;
        RECT 25.955 147.185 27.625 148.275 ;
        RECT 27.885 147.345 28.055 148.105 ;
        RECT 28.235 147.515 28.565 148.275 ;
        RECT 25.030 147.030 25.200 147.175 ;
        RECT 24.915 146.700 25.200 147.030 ;
        RECT 25.030 146.445 25.200 146.700 ;
        RECT 25.435 146.625 25.765 146.995 ;
        RECT 25.955 146.665 26.705 147.185 ;
        RECT 27.885 147.175 28.550 147.345 ;
        RECT 28.735 147.200 29.005 148.105 ;
        RECT 28.380 147.030 28.550 147.175 ;
        RECT 26.875 146.495 27.625 147.015 ;
        RECT 27.815 146.625 28.145 146.995 ;
        RECT 28.380 146.700 28.665 147.030 ;
        RECT 24.575 145.895 24.835 146.400 ;
        RECT 25.030 146.275 25.695 146.445 ;
        RECT 25.015 145.725 25.345 146.105 ;
        RECT 25.525 145.895 25.695 146.275 ;
        RECT 25.955 145.725 27.625 146.495 ;
        RECT 28.380 146.445 28.550 146.700 ;
        RECT 27.885 146.275 28.550 146.445 ;
        RECT 28.835 146.400 29.005 147.200 ;
        RECT 27.885 145.895 28.055 146.275 ;
        RECT 28.235 145.725 28.565 146.105 ;
        RECT 28.745 145.895 29.005 146.400 ;
        RECT 29.180 147.135 29.515 148.105 ;
        RECT 29.685 147.135 29.855 148.275 ;
        RECT 30.025 147.935 32.055 148.105 ;
        RECT 29.180 146.465 29.350 147.135 ;
        RECT 30.025 146.965 30.195 147.935 ;
        RECT 29.520 146.635 29.775 146.965 ;
        RECT 30.000 146.635 30.195 146.965 ;
        RECT 30.365 147.595 31.490 147.765 ;
        RECT 29.605 146.465 29.775 146.635 ;
        RECT 30.365 146.465 30.535 147.595 ;
        RECT 29.180 145.895 29.435 146.465 ;
        RECT 29.605 146.295 30.535 146.465 ;
        RECT 30.705 147.255 31.715 147.425 ;
        RECT 30.705 146.455 30.875 147.255 ;
        RECT 31.080 146.915 31.355 147.055 ;
        RECT 31.075 146.745 31.355 146.915 ;
        RECT 30.360 146.260 30.535 146.295 ;
        RECT 29.605 145.725 29.935 146.125 ;
        RECT 30.360 145.895 30.890 146.260 ;
        RECT 31.080 145.895 31.355 146.745 ;
        RECT 31.525 145.895 31.715 147.255 ;
        RECT 31.885 147.270 32.055 147.935 ;
        RECT 32.225 147.515 32.395 148.275 ;
        RECT 32.630 147.515 33.145 147.925 ;
        RECT 31.885 147.080 32.635 147.270 ;
        RECT 32.805 146.705 33.145 147.515 ;
        RECT 31.915 146.535 33.145 146.705 ;
        RECT 33.775 147.185 35.445 148.275 ;
        RECT 35.820 147.305 36.150 148.105 ;
        RECT 36.320 147.475 36.650 148.275 ;
        RECT 36.950 147.305 37.280 148.105 ;
        RECT 37.925 147.475 38.175 148.275 ;
        RECT 33.775 146.665 34.525 147.185 ;
        RECT 35.820 147.135 38.255 147.305 ;
        RECT 38.445 147.135 38.615 148.275 ;
        RECT 38.785 147.135 39.125 148.105 ;
        RECT 31.895 145.725 32.405 146.260 ;
        RECT 32.625 145.930 32.870 146.535 ;
        RECT 34.695 146.495 35.445 147.015 ;
        RECT 35.615 146.715 35.965 146.965 ;
        RECT 36.150 146.505 36.320 147.135 ;
        RECT 36.490 146.715 36.820 146.915 ;
        RECT 36.990 146.715 37.320 146.915 ;
        RECT 37.490 146.715 37.910 146.915 ;
        RECT 38.085 146.885 38.255 147.135 ;
        RECT 38.085 146.715 38.780 146.885 ;
        RECT 33.775 145.725 35.445 146.495 ;
        RECT 35.820 145.895 36.320 146.505 ;
        RECT 36.950 146.375 38.175 146.545 ;
        RECT 38.950 146.525 39.125 147.135 ;
        RECT 36.950 145.895 37.280 146.375 ;
        RECT 37.450 145.725 37.675 146.185 ;
        RECT 37.845 145.895 38.175 146.375 ;
        RECT 38.365 145.725 38.615 146.525 ;
        RECT 38.785 145.895 39.125 146.525 ;
        RECT 39.295 147.135 39.635 148.105 ;
        RECT 39.805 147.135 39.975 148.275 ;
        RECT 40.245 147.475 40.495 148.275 ;
        RECT 41.140 147.305 41.470 148.105 ;
        RECT 41.770 147.475 42.100 148.275 ;
        RECT 42.270 147.305 42.600 148.105 ;
        RECT 40.165 147.135 42.600 147.305 ;
        RECT 43.435 147.185 46.945 148.275 ;
        RECT 47.120 147.765 48.775 148.055 ;
        RECT 47.120 147.425 48.710 147.595 ;
        RECT 48.945 147.475 49.225 148.275 ;
        RECT 39.295 146.575 39.470 147.135 ;
        RECT 40.165 146.885 40.335 147.135 ;
        RECT 39.640 146.715 40.335 146.885 ;
        RECT 40.510 146.715 40.930 146.915 ;
        RECT 41.100 146.715 41.430 146.915 ;
        RECT 41.600 146.715 41.930 146.915 ;
        RECT 39.295 146.525 39.525 146.575 ;
        RECT 39.295 145.895 39.635 146.525 ;
        RECT 39.805 145.725 40.055 146.525 ;
        RECT 40.245 146.375 41.470 146.545 ;
        RECT 40.245 145.895 40.575 146.375 ;
        RECT 40.745 145.725 40.970 146.185 ;
        RECT 41.140 145.895 41.470 146.375 ;
        RECT 42.100 146.505 42.270 147.135 ;
        RECT 42.455 146.715 42.805 146.965 ;
        RECT 43.435 146.665 45.125 147.185 ;
        RECT 47.120 147.135 47.440 147.425 ;
        RECT 48.540 147.305 48.710 147.425 ;
        RECT 42.100 145.895 42.600 146.505 ;
        RECT 45.295 146.495 46.945 147.015 ;
        RECT 43.435 145.725 46.945 146.495 ;
        RECT 47.120 146.395 47.470 146.965 ;
        RECT 47.640 146.635 48.350 147.255 ;
        RECT 48.540 147.135 49.265 147.305 ;
        RECT 49.435 147.135 49.705 148.105 ;
        RECT 49.095 146.965 49.265 147.135 ;
        RECT 48.520 146.635 48.925 146.965 ;
        RECT 49.095 146.635 49.365 146.965 ;
        RECT 49.095 146.465 49.265 146.635 ;
        RECT 47.655 146.295 49.265 146.465 ;
        RECT 49.535 146.400 49.705 147.135 ;
        RECT 49.875 147.110 50.165 148.275 ;
        RECT 50.795 147.200 51.065 148.105 ;
        RECT 51.235 147.515 51.565 148.275 ;
        RECT 51.745 147.345 51.915 148.105 ;
        RECT 47.125 145.725 47.455 146.225 ;
        RECT 47.655 145.945 47.825 146.295 ;
        RECT 48.025 145.725 48.355 146.125 ;
        RECT 48.525 145.945 48.695 146.295 ;
        RECT 48.865 145.725 49.245 146.125 ;
        RECT 49.435 146.055 49.705 146.400 ;
        RECT 49.875 145.725 50.165 146.450 ;
        RECT 50.795 146.400 50.965 147.200 ;
        RECT 51.250 147.175 51.915 147.345 ;
        RECT 51.250 147.030 51.420 147.175 ;
        RECT 51.135 146.700 51.420 147.030 ;
        RECT 53.095 147.135 53.435 148.105 ;
        RECT 53.605 147.135 53.775 148.275 ;
        RECT 54.045 147.475 54.295 148.275 ;
        RECT 54.940 147.305 55.270 148.105 ;
        RECT 55.570 147.475 55.900 148.275 ;
        RECT 56.070 147.305 56.400 148.105 ;
        RECT 53.965 147.135 56.400 147.305 ;
        RECT 56.775 147.185 59.365 148.275 ;
        RECT 59.535 147.515 60.050 147.925 ;
        RECT 60.285 147.515 60.455 148.275 ;
        RECT 60.625 147.935 62.655 148.105 ;
        RECT 51.250 146.445 51.420 146.700 ;
        RECT 51.655 146.625 51.985 146.995 ;
        RECT 53.095 146.525 53.270 147.135 ;
        RECT 53.965 146.885 54.135 147.135 ;
        RECT 53.440 146.715 54.135 146.885 ;
        RECT 54.310 146.715 54.730 146.915 ;
        RECT 54.900 146.715 55.230 146.915 ;
        RECT 55.400 146.715 55.730 146.915 ;
        RECT 50.795 145.895 51.055 146.400 ;
        RECT 51.250 146.275 51.915 146.445 ;
        RECT 51.235 145.725 51.565 146.105 ;
        RECT 51.745 145.895 51.915 146.275 ;
        RECT 53.095 145.895 53.435 146.525 ;
        RECT 53.605 145.725 53.855 146.525 ;
        RECT 54.045 146.375 55.270 146.545 ;
        RECT 54.045 145.895 54.375 146.375 ;
        RECT 54.545 145.725 54.770 146.185 ;
        RECT 54.940 145.895 55.270 146.375 ;
        RECT 55.900 146.505 56.070 147.135 ;
        RECT 56.255 146.715 56.605 146.965 ;
        RECT 56.775 146.665 57.985 147.185 ;
        RECT 55.900 145.895 56.400 146.505 ;
        RECT 58.155 146.495 59.365 147.015 ;
        RECT 59.535 146.705 59.875 147.515 ;
        RECT 60.625 147.270 60.795 147.935 ;
        RECT 61.190 147.595 62.315 147.765 ;
        RECT 60.045 147.080 60.795 147.270 ;
        RECT 60.965 147.255 61.975 147.425 ;
        RECT 59.535 146.535 60.765 146.705 ;
        RECT 56.775 145.725 59.365 146.495 ;
        RECT 59.810 145.930 60.055 146.535 ;
        RECT 60.275 145.725 60.785 146.260 ;
        RECT 60.965 145.895 61.155 147.255 ;
        RECT 61.325 146.235 61.600 147.055 ;
        RECT 61.805 146.455 61.975 147.255 ;
        RECT 62.145 146.465 62.315 147.595 ;
        RECT 62.485 146.965 62.655 147.935 ;
        RECT 62.825 147.135 62.995 148.275 ;
        RECT 63.165 147.135 63.500 148.105 ;
        RECT 62.485 146.635 62.680 146.965 ;
        RECT 62.905 146.635 63.160 146.965 ;
        RECT 62.905 146.465 63.075 146.635 ;
        RECT 63.330 146.465 63.500 147.135 ;
        RECT 63.675 147.185 64.885 148.275 ;
        RECT 65.060 147.840 70.405 148.275 ;
        RECT 63.675 146.645 64.195 147.185 ;
        RECT 64.365 146.475 64.885 147.015 ;
        RECT 66.650 146.590 67.000 147.840 ;
        RECT 70.580 147.125 70.840 148.275 ;
        RECT 71.015 147.200 71.270 148.105 ;
        RECT 71.440 147.515 71.770 148.275 ;
        RECT 71.985 147.345 72.155 148.105 ;
        RECT 62.145 146.295 63.075 146.465 ;
        RECT 62.145 146.260 62.320 146.295 ;
        RECT 61.325 146.065 61.605 146.235 ;
        RECT 61.325 145.895 61.600 146.065 ;
        RECT 61.790 145.895 62.320 146.260 ;
        RECT 62.745 145.725 63.075 146.125 ;
        RECT 63.245 145.895 63.500 146.465 ;
        RECT 63.675 145.725 64.885 146.475 ;
        RECT 68.480 146.270 68.820 147.100 ;
        RECT 65.060 145.725 70.405 146.270 ;
        RECT 70.580 145.725 70.840 146.565 ;
        RECT 71.015 146.470 71.185 147.200 ;
        RECT 71.440 147.175 72.155 147.345 ;
        RECT 72.505 147.345 72.675 148.105 ;
        RECT 72.890 147.515 73.220 148.275 ;
        RECT 72.505 147.175 73.220 147.345 ;
        RECT 73.390 147.200 73.645 148.105 ;
        RECT 71.440 146.965 71.610 147.175 ;
        RECT 71.355 146.635 71.610 146.965 ;
        RECT 71.015 145.895 71.270 146.470 ;
        RECT 71.440 146.445 71.610 146.635 ;
        RECT 71.890 146.625 72.245 146.995 ;
        RECT 72.415 146.625 72.770 146.995 ;
        RECT 73.050 146.965 73.220 147.175 ;
        RECT 73.050 146.635 73.305 146.965 ;
        RECT 73.050 146.445 73.220 146.635 ;
        RECT 73.475 146.470 73.645 147.200 ;
        RECT 73.820 147.125 74.080 148.275 ;
        RECT 74.255 147.185 75.465 148.275 ;
        RECT 74.255 146.645 74.775 147.185 ;
        RECT 75.635 147.110 75.925 148.275 ;
        RECT 76.300 147.305 76.630 148.105 ;
        RECT 76.800 147.475 77.130 148.275 ;
        RECT 77.430 147.305 77.760 148.105 ;
        RECT 78.405 147.475 78.655 148.275 ;
        RECT 76.300 147.135 78.735 147.305 ;
        RECT 78.925 147.135 79.095 148.275 ;
        RECT 79.265 147.135 79.605 148.105 ;
        RECT 71.440 146.275 72.155 146.445 ;
        RECT 71.440 145.725 71.770 146.105 ;
        RECT 71.985 145.895 72.155 146.275 ;
        RECT 72.505 146.275 73.220 146.445 ;
        RECT 72.505 145.895 72.675 146.275 ;
        RECT 72.890 145.725 73.220 146.105 ;
        RECT 73.390 145.895 73.645 146.470 ;
        RECT 73.820 145.725 74.080 146.565 ;
        RECT 74.945 146.475 75.465 147.015 ;
        RECT 76.095 146.715 76.445 146.965 ;
        RECT 76.630 146.505 76.800 147.135 ;
        RECT 76.970 146.715 77.300 146.915 ;
        RECT 77.470 146.715 77.800 146.915 ;
        RECT 77.970 146.715 78.390 146.915 ;
        RECT 78.565 146.885 78.735 147.135 ;
        RECT 78.565 146.715 79.260 146.885 ;
        RECT 74.255 145.725 75.465 146.475 ;
        RECT 75.635 145.725 75.925 146.450 ;
        RECT 76.300 145.895 76.800 146.505 ;
        RECT 77.430 146.375 78.655 146.545 ;
        RECT 79.430 146.525 79.605 147.135 ;
        RECT 77.430 145.895 77.760 146.375 ;
        RECT 77.930 145.725 78.155 146.185 ;
        RECT 78.325 145.895 78.655 146.375 ;
        RECT 78.845 145.725 79.095 146.525 ;
        RECT 79.265 145.895 79.605 146.525 ;
        RECT 79.775 147.135 80.115 148.105 ;
        RECT 80.285 147.135 80.455 148.275 ;
        RECT 80.725 147.475 80.975 148.275 ;
        RECT 81.620 147.305 81.950 148.105 ;
        RECT 82.250 147.475 82.580 148.275 ;
        RECT 82.750 147.305 83.080 148.105 ;
        RECT 80.645 147.135 83.080 147.305 ;
        RECT 83.455 147.185 84.665 148.275 ;
        RECT 85.210 147.295 85.465 147.965 ;
        RECT 85.645 147.475 85.930 148.275 ;
        RECT 86.110 147.555 86.440 148.065 ;
        RECT 79.775 146.525 79.950 147.135 ;
        RECT 80.645 146.885 80.815 147.135 ;
        RECT 80.120 146.715 80.815 146.885 ;
        RECT 80.990 146.715 81.410 146.915 ;
        RECT 81.580 146.715 81.910 146.915 ;
        RECT 82.080 146.715 82.410 146.915 ;
        RECT 79.775 145.895 80.115 146.525 ;
        RECT 80.285 145.725 80.535 146.525 ;
        RECT 80.725 146.375 81.950 146.545 ;
        RECT 80.725 145.895 81.055 146.375 ;
        RECT 81.225 145.725 81.450 146.185 ;
        RECT 81.620 145.895 81.950 146.375 ;
        RECT 82.580 146.505 82.750 147.135 ;
        RECT 82.935 146.715 83.285 146.965 ;
        RECT 83.455 146.645 83.975 147.185 ;
        RECT 82.580 145.895 83.080 146.505 ;
        RECT 84.145 146.475 84.665 147.015 ;
        RECT 83.455 145.725 84.665 146.475 ;
        RECT 85.210 146.435 85.390 147.295 ;
        RECT 86.110 146.965 86.360 147.555 ;
        RECT 86.710 147.405 86.880 148.015 ;
        RECT 87.050 147.585 87.380 148.275 ;
        RECT 87.610 147.725 87.850 148.015 ;
        RECT 88.050 147.895 88.470 148.275 ;
        RECT 88.650 147.805 89.280 148.055 ;
        RECT 89.750 147.895 90.080 148.275 ;
        RECT 88.650 147.725 88.820 147.805 ;
        RECT 90.250 147.725 90.420 148.015 ;
        RECT 90.600 147.895 90.980 148.275 ;
        RECT 91.220 147.890 92.050 148.060 ;
        RECT 87.610 147.555 88.820 147.725 ;
        RECT 85.560 146.635 86.360 146.965 ;
        RECT 85.210 146.235 85.465 146.435 ;
        RECT 85.125 146.065 85.465 146.235 ;
        RECT 85.210 145.905 85.465 146.065 ;
        RECT 85.645 145.725 85.930 146.185 ;
        RECT 86.110 145.985 86.360 146.635 ;
        RECT 86.560 147.385 86.880 147.405 ;
        RECT 86.560 147.215 88.480 147.385 ;
        RECT 86.560 146.320 86.750 147.215 ;
        RECT 88.650 147.045 88.820 147.555 ;
        RECT 88.990 147.295 89.510 147.605 ;
        RECT 86.920 146.875 88.820 147.045 ;
        RECT 86.920 146.815 87.250 146.875 ;
        RECT 87.400 146.645 87.730 146.705 ;
        RECT 87.070 146.375 87.730 146.645 ;
        RECT 86.560 145.990 86.880 146.320 ;
        RECT 87.060 145.725 87.720 146.205 ;
        RECT 87.920 146.115 88.090 146.875 ;
        RECT 88.990 146.705 89.170 147.115 ;
        RECT 88.260 146.535 88.590 146.655 ;
        RECT 89.340 146.535 89.510 147.295 ;
        RECT 88.260 146.365 89.510 146.535 ;
        RECT 89.680 147.475 91.050 147.725 ;
        RECT 89.680 146.705 89.870 147.475 ;
        RECT 90.800 147.215 91.050 147.475 ;
        RECT 90.040 147.045 90.290 147.205 ;
        RECT 91.220 147.045 91.390 147.890 ;
        RECT 92.285 147.605 92.455 148.105 ;
        RECT 92.625 147.775 92.955 148.275 ;
        RECT 91.560 147.215 92.060 147.595 ;
        RECT 92.285 147.435 92.980 147.605 ;
        RECT 90.040 146.875 91.390 147.045 ;
        RECT 90.970 146.835 91.390 146.875 ;
        RECT 89.680 146.365 90.100 146.705 ;
        RECT 90.390 146.375 90.800 146.705 ;
        RECT 87.920 145.945 88.770 146.115 ;
        RECT 89.330 145.725 89.650 146.185 ;
        RECT 89.850 145.935 90.100 146.365 ;
        RECT 90.390 145.725 90.800 146.165 ;
        RECT 90.970 146.105 91.140 146.835 ;
        RECT 91.310 146.285 91.660 146.655 ;
        RECT 91.840 146.345 92.060 147.215 ;
        RECT 92.230 146.645 92.640 147.265 ;
        RECT 92.810 146.465 92.980 147.435 ;
        RECT 92.285 146.275 92.980 146.465 ;
        RECT 90.970 145.905 91.985 146.105 ;
        RECT 92.285 145.945 92.455 146.275 ;
        RECT 92.625 145.725 92.955 146.105 ;
        RECT 93.170 145.985 93.395 148.105 ;
        RECT 93.565 147.775 93.895 148.275 ;
        RECT 94.065 147.605 94.235 148.105 ;
        RECT 93.570 147.435 94.235 147.605 ;
        RECT 93.570 146.445 93.800 147.435 ;
        RECT 93.970 146.615 94.320 147.265 ;
        RECT 94.995 147.135 95.225 148.275 ;
        RECT 95.395 147.125 95.725 148.105 ;
        RECT 95.895 147.135 96.105 148.275 ;
        RECT 96.335 147.515 96.850 147.925 ;
        RECT 97.085 147.515 97.255 148.275 ;
        RECT 97.425 147.935 99.455 148.105 ;
        RECT 94.975 146.715 95.305 146.965 ;
        RECT 93.570 146.275 94.235 146.445 ;
        RECT 93.565 145.725 93.895 146.105 ;
        RECT 94.065 145.985 94.235 146.275 ;
        RECT 94.995 145.725 95.225 146.545 ;
        RECT 95.475 146.525 95.725 147.125 ;
        RECT 96.335 146.705 96.675 147.515 ;
        RECT 97.425 147.270 97.595 147.935 ;
        RECT 97.990 147.595 99.115 147.765 ;
        RECT 96.845 147.080 97.595 147.270 ;
        RECT 97.765 147.255 98.775 147.425 ;
        RECT 95.395 145.895 95.725 146.525 ;
        RECT 95.895 145.725 96.105 146.545 ;
        RECT 96.335 146.535 97.565 146.705 ;
        RECT 96.610 145.930 96.855 146.535 ;
        RECT 97.075 145.725 97.585 146.260 ;
        RECT 97.765 145.895 97.955 147.255 ;
        RECT 98.125 146.915 98.400 147.055 ;
        RECT 98.125 146.745 98.405 146.915 ;
        RECT 98.125 145.895 98.400 146.745 ;
        RECT 98.605 146.455 98.775 147.255 ;
        RECT 98.945 146.465 99.115 147.595 ;
        RECT 99.285 146.965 99.455 147.935 ;
        RECT 99.625 147.135 99.795 148.275 ;
        RECT 99.965 147.135 100.300 148.105 ;
        RECT 99.285 146.635 99.480 146.965 ;
        RECT 99.705 146.635 99.960 146.965 ;
        RECT 99.705 146.465 99.875 146.635 ;
        RECT 100.130 146.465 100.300 147.135 ;
        RECT 101.395 147.110 101.685 148.275 ;
        RECT 101.945 147.345 102.115 148.105 ;
        RECT 102.295 147.515 102.625 148.275 ;
        RECT 101.945 147.175 102.610 147.345 ;
        RECT 102.795 147.200 103.065 148.105 ;
        RECT 102.440 147.030 102.610 147.175 ;
        RECT 101.875 146.625 102.205 146.995 ;
        RECT 102.440 146.700 102.725 147.030 ;
        RECT 98.945 146.295 99.875 146.465 ;
        RECT 98.945 146.260 99.120 146.295 ;
        RECT 98.590 145.895 99.120 146.260 ;
        RECT 99.545 145.725 99.875 146.125 ;
        RECT 100.045 145.895 100.300 146.465 ;
        RECT 101.395 145.725 101.685 146.450 ;
        RECT 102.440 146.445 102.610 146.700 ;
        RECT 101.945 146.275 102.610 146.445 ;
        RECT 102.895 146.400 103.065 147.200 ;
        RECT 101.945 145.895 102.115 146.275 ;
        RECT 102.295 145.725 102.625 146.105 ;
        RECT 102.805 145.895 103.065 146.400 ;
        RECT 103.695 147.135 103.965 148.105 ;
        RECT 104.175 147.475 104.455 148.275 ;
        RECT 104.625 147.765 106.280 148.055 ;
        RECT 104.690 147.425 106.280 147.595 ;
        RECT 104.690 147.305 104.860 147.425 ;
        RECT 104.135 147.135 104.860 147.305 ;
        RECT 103.695 146.400 103.865 147.135 ;
        RECT 104.135 146.965 104.305 147.135 ;
        RECT 105.050 147.085 105.765 147.255 ;
        RECT 105.960 147.135 106.280 147.425 ;
        RECT 106.455 147.135 106.795 148.105 ;
        RECT 106.965 147.135 107.135 148.275 ;
        RECT 107.405 147.475 107.655 148.275 ;
        RECT 108.300 147.305 108.630 148.105 ;
        RECT 108.930 147.475 109.260 148.275 ;
        RECT 109.430 147.305 109.760 148.105 ;
        RECT 107.325 147.135 109.760 147.305 ;
        RECT 110.135 147.185 111.805 148.275 ;
        RECT 111.975 147.515 112.490 147.925 ;
        RECT 112.725 147.515 112.895 148.275 ;
        RECT 113.065 147.935 115.095 148.105 ;
        RECT 104.035 146.635 104.305 146.965 ;
        RECT 104.475 146.635 104.880 146.965 ;
        RECT 105.050 146.635 105.760 147.085 ;
        RECT 104.135 146.465 104.305 146.635 ;
        RECT 103.695 146.055 103.965 146.400 ;
        RECT 104.135 146.295 105.745 146.465 ;
        RECT 105.930 146.395 106.280 146.965 ;
        RECT 106.455 146.575 106.630 147.135 ;
        RECT 107.325 146.885 107.495 147.135 ;
        RECT 106.800 146.715 107.495 146.885 ;
        RECT 107.670 146.715 108.090 146.915 ;
        RECT 108.260 146.715 108.590 146.915 ;
        RECT 108.760 146.715 109.090 146.915 ;
        RECT 106.455 146.525 106.685 146.575 ;
        RECT 104.155 145.725 104.535 146.125 ;
        RECT 104.705 145.945 104.875 146.295 ;
        RECT 105.045 145.725 105.375 146.125 ;
        RECT 105.575 145.945 105.745 146.295 ;
        RECT 105.945 145.725 106.275 146.225 ;
        RECT 106.455 145.895 106.795 146.525 ;
        RECT 106.965 145.725 107.215 146.525 ;
        RECT 107.405 146.375 108.630 146.545 ;
        RECT 107.405 145.895 107.735 146.375 ;
        RECT 107.905 145.725 108.130 146.185 ;
        RECT 108.300 145.895 108.630 146.375 ;
        RECT 109.260 146.505 109.430 147.135 ;
        RECT 109.615 146.715 109.965 146.965 ;
        RECT 110.135 146.665 110.885 147.185 ;
        RECT 109.260 145.895 109.760 146.505 ;
        RECT 111.055 146.495 111.805 147.015 ;
        RECT 111.975 146.705 112.315 147.515 ;
        RECT 113.065 147.270 113.235 147.935 ;
        RECT 113.630 147.595 114.755 147.765 ;
        RECT 112.485 147.080 113.235 147.270 ;
        RECT 113.405 147.255 114.415 147.425 ;
        RECT 111.975 146.535 113.205 146.705 ;
        RECT 110.135 145.725 111.805 146.495 ;
        RECT 112.250 145.930 112.495 146.535 ;
        RECT 112.715 145.725 113.225 146.260 ;
        RECT 113.405 145.895 113.595 147.255 ;
        RECT 113.765 146.915 114.040 147.055 ;
        RECT 113.765 146.745 114.045 146.915 ;
        RECT 113.765 145.895 114.040 146.745 ;
        RECT 114.245 146.455 114.415 147.255 ;
        RECT 114.585 146.465 114.755 147.595 ;
        RECT 114.925 146.965 115.095 147.935 ;
        RECT 115.265 147.135 115.435 148.275 ;
        RECT 115.605 147.135 115.940 148.105 ;
        RECT 114.925 146.635 115.120 146.965 ;
        RECT 115.345 146.635 115.600 146.965 ;
        RECT 115.345 146.465 115.515 146.635 ;
        RECT 115.770 146.465 115.940 147.135 ;
        RECT 116.490 147.295 116.745 147.965 ;
        RECT 116.925 147.475 117.210 148.275 ;
        RECT 117.390 147.555 117.720 148.065 ;
        RECT 116.490 146.575 116.670 147.295 ;
        RECT 117.390 146.965 117.640 147.555 ;
        RECT 117.990 147.405 118.160 148.015 ;
        RECT 118.330 147.585 118.660 148.275 ;
        RECT 118.890 147.725 119.130 148.015 ;
        RECT 119.330 147.895 119.750 148.275 ;
        RECT 119.930 147.805 120.560 148.055 ;
        RECT 121.030 147.895 121.360 148.275 ;
        RECT 119.930 147.725 120.100 147.805 ;
        RECT 121.530 147.725 121.700 148.015 ;
        RECT 121.880 147.895 122.260 148.275 ;
        RECT 122.500 147.890 123.330 148.060 ;
        RECT 118.890 147.555 120.100 147.725 ;
        RECT 116.840 146.635 117.640 146.965 ;
        RECT 114.585 146.295 115.515 146.465 ;
        RECT 114.585 146.260 114.760 146.295 ;
        RECT 114.230 145.895 114.760 146.260 ;
        RECT 115.185 145.725 115.515 146.125 ;
        RECT 115.685 145.895 115.940 146.465 ;
        RECT 116.405 146.435 116.670 146.575 ;
        RECT 116.405 146.405 116.745 146.435 ;
        RECT 116.490 145.905 116.745 146.405 ;
        RECT 116.925 145.725 117.210 146.185 ;
        RECT 117.390 145.985 117.640 146.635 ;
        RECT 117.840 147.385 118.160 147.405 ;
        RECT 117.840 147.215 119.760 147.385 ;
        RECT 117.840 146.320 118.030 147.215 ;
        RECT 119.930 147.045 120.100 147.555 ;
        RECT 120.270 147.295 120.790 147.605 ;
        RECT 118.200 146.875 120.100 147.045 ;
        RECT 118.200 146.815 118.530 146.875 ;
        RECT 118.680 146.645 119.010 146.705 ;
        RECT 118.350 146.375 119.010 146.645 ;
        RECT 117.840 145.990 118.160 146.320 ;
        RECT 118.340 145.725 119.000 146.205 ;
        RECT 119.200 146.115 119.370 146.875 ;
        RECT 120.270 146.705 120.450 147.115 ;
        RECT 119.540 146.535 119.870 146.655 ;
        RECT 120.620 146.535 120.790 147.295 ;
        RECT 119.540 146.365 120.790 146.535 ;
        RECT 120.960 147.475 122.330 147.725 ;
        RECT 120.960 146.705 121.150 147.475 ;
        RECT 122.080 147.215 122.330 147.475 ;
        RECT 121.320 147.045 121.570 147.205 ;
        RECT 122.500 147.045 122.670 147.890 ;
        RECT 123.565 147.605 123.735 148.105 ;
        RECT 123.905 147.775 124.235 148.275 ;
        RECT 122.840 147.215 123.340 147.595 ;
        RECT 123.565 147.435 124.260 147.605 ;
        RECT 121.320 146.875 122.670 147.045 ;
        RECT 122.250 146.835 122.670 146.875 ;
        RECT 120.960 146.365 121.380 146.705 ;
        RECT 121.670 146.375 122.080 146.705 ;
        RECT 119.200 145.945 120.050 146.115 ;
        RECT 120.610 145.725 120.930 146.185 ;
        RECT 121.130 145.935 121.380 146.365 ;
        RECT 121.670 145.725 122.080 146.165 ;
        RECT 122.250 146.105 122.420 146.835 ;
        RECT 122.590 146.285 122.940 146.655 ;
        RECT 123.120 146.345 123.340 147.215 ;
        RECT 123.510 146.645 123.920 147.265 ;
        RECT 124.090 146.465 124.260 147.435 ;
        RECT 123.565 146.275 124.260 146.465 ;
        RECT 122.250 145.905 123.265 146.105 ;
        RECT 123.565 145.945 123.735 146.275 ;
        RECT 123.905 145.725 124.235 146.105 ;
        RECT 124.450 145.985 124.675 148.105 ;
        RECT 124.845 147.775 125.175 148.275 ;
        RECT 125.345 147.605 125.515 148.105 ;
        RECT 124.850 147.435 125.515 147.605 ;
        RECT 124.850 146.445 125.080 147.435 ;
        RECT 125.250 146.615 125.600 147.265 ;
        RECT 126.235 147.185 127.445 148.275 ;
        RECT 126.235 146.645 126.755 147.185 ;
        RECT 126.925 146.475 127.445 147.015 ;
        RECT 124.850 146.275 125.515 146.445 ;
        RECT 124.845 145.725 125.175 146.105 ;
        RECT 125.345 145.985 125.515 146.275 ;
        RECT 126.235 145.725 127.445 146.475 ;
        RECT 14.370 145.555 127.530 145.725 ;
        RECT 14.455 144.805 15.665 145.555 ;
        RECT 14.455 144.265 14.975 144.805 ;
        RECT 15.835 144.785 19.345 145.555 ;
        RECT 15.145 144.095 15.665 144.635 ;
        RECT 14.455 143.005 15.665 144.095 ;
        RECT 15.835 144.095 17.525 144.615 ;
        RECT 17.695 144.265 19.345 144.785 ;
        RECT 19.555 144.735 19.785 145.555 ;
        RECT 19.955 144.755 20.285 145.385 ;
        RECT 19.535 144.315 19.865 144.565 ;
        RECT 20.035 144.155 20.285 144.755 ;
        RECT 20.455 144.735 20.665 145.555 ;
        RECT 20.935 144.735 21.165 145.555 ;
        RECT 21.335 144.755 21.665 145.385 ;
        RECT 20.915 144.315 21.245 144.565 ;
        RECT 21.415 144.155 21.665 144.755 ;
        RECT 21.835 144.735 22.045 145.555 ;
        RECT 22.650 145.215 22.905 145.375 ;
        RECT 22.565 145.045 22.905 145.215 ;
        RECT 23.085 145.095 23.370 145.555 ;
        RECT 22.650 144.845 22.905 145.045 ;
        RECT 15.835 143.005 19.345 144.095 ;
        RECT 19.555 143.005 19.785 144.145 ;
        RECT 19.955 143.175 20.285 144.155 ;
        RECT 20.455 143.005 20.665 144.145 ;
        RECT 20.935 143.005 21.165 144.145 ;
        RECT 21.335 143.175 21.665 144.155 ;
        RECT 21.835 143.005 22.045 144.145 ;
        RECT 22.650 143.985 22.830 144.845 ;
        RECT 23.550 144.645 23.800 145.295 ;
        RECT 23.000 144.315 23.800 144.645 ;
        RECT 22.650 143.315 22.905 143.985 ;
        RECT 23.085 143.005 23.370 143.805 ;
        RECT 23.550 143.725 23.800 144.315 ;
        RECT 24.000 144.960 24.320 145.290 ;
        RECT 24.500 145.075 25.160 145.555 ;
        RECT 25.360 145.165 26.210 145.335 ;
        RECT 24.000 144.065 24.190 144.960 ;
        RECT 24.510 144.635 25.170 144.905 ;
        RECT 24.840 144.575 25.170 144.635 ;
        RECT 24.360 144.405 24.690 144.465 ;
        RECT 25.360 144.405 25.530 145.165 ;
        RECT 26.770 145.095 27.090 145.555 ;
        RECT 27.290 144.915 27.540 145.345 ;
        RECT 27.830 145.115 28.240 145.555 ;
        RECT 28.410 145.175 29.425 145.375 ;
        RECT 25.700 144.745 26.950 144.915 ;
        RECT 25.700 144.625 26.030 144.745 ;
        RECT 24.360 144.235 26.260 144.405 ;
        RECT 24.000 143.895 25.920 144.065 ;
        RECT 24.000 143.875 24.320 143.895 ;
        RECT 23.550 143.215 23.880 143.725 ;
        RECT 24.150 143.265 24.320 143.875 ;
        RECT 26.090 143.725 26.260 144.235 ;
        RECT 26.430 144.165 26.610 144.575 ;
        RECT 26.780 143.985 26.950 144.745 ;
        RECT 24.490 143.005 24.820 143.695 ;
        RECT 25.050 143.555 26.260 143.725 ;
        RECT 26.430 143.675 26.950 143.985 ;
        RECT 27.120 144.575 27.540 144.915 ;
        RECT 27.830 144.575 28.240 144.905 ;
        RECT 27.120 143.805 27.310 144.575 ;
        RECT 28.410 144.445 28.580 145.175 ;
        RECT 29.725 145.005 29.895 145.335 ;
        RECT 30.065 145.175 30.395 145.555 ;
        RECT 28.750 144.625 29.100 144.995 ;
        RECT 28.410 144.405 28.830 144.445 ;
        RECT 27.480 144.235 28.830 144.405 ;
        RECT 27.480 144.075 27.730 144.235 ;
        RECT 28.240 143.805 28.490 144.065 ;
        RECT 27.120 143.555 28.490 143.805 ;
        RECT 25.050 143.265 25.290 143.555 ;
        RECT 26.090 143.475 26.260 143.555 ;
        RECT 25.490 143.005 25.910 143.385 ;
        RECT 26.090 143.225 26.720 143.475 ;
        RECT 27.190 143.005 27.520 143.385 ;
        RECT 27.690 143.265 27.860 143.555 ;
        RECT 28.660 143.390 28.830 144.235 ;
        RECT 29.280 144.065 29.500 144.935 ;
        RECT 29.725 144.815 30.420 145.005 ;
        RECT 29.000 143.685 29.500 144.065 ;
        RECT 29.670 144.015 30.080 144.635 ;
        RECT 30.250 143.845 30.420 144.815 ;
        RECT 29.725 143.675 30.420 143.845 ;
        RECT 28.040 143.005 28.420 143.385 ;
        RECT 28.660 143.220 29.490 143.390 ;
        RECT 29.725 143.175 29.895 143.675 ;
        RECT 30.065 143.005 30.395 143.505 ;
        RECT 30.610 143.175 30.835 145.295 ;
        RECT 31.005 145.175 31.335 145.555 ;
        RECT 31.505 145.005 31.675 145.295 ;
        RECT 31.010 144.835 31.675 145.005 ;
        RECT 31.010 143.845 31.240 144.835 ;
        RECT 31.935 144.805 33.145 145.555 ;
        RECT 31.410 144.015 31.760 144.665 ;
        RECT 31.935 144.095 32.455 144.635 ;
        RECT 32.625 144.265 33.145 144.805 ;
        RECT 33.315 144.785 36.825 145.555 ;
        RECT 36.995 144.830 37.285 145.555 ;
        RECT 37.915 144.785 40.505 145.555 ;
        RECT 33.315 144.095 35.005 144.615 ;
        RECT 35.175 144.265 36.825 144.785 ;
        RECT 31.010 143.675 31.675 143.845 ;
        RECT 31.005 143.005 31.335 143.505 ;
        RECT 31.505 143.175 31.675 143.675 ;
        RECT 31.935 143.005 33.145 144.095 ;
        RECT 33.315 143.005 36.825 144.095 ;
        RECT 36.995 143.005 37.285 144.170 ;
        RECT 37.915 144.095 39.125 144.615 ;
        RECT 39.295 144.265 40.505 144.785 ;
        RECT 40.715 144.735 40.945 145.555 ;
        RECT 41.115 144.755 41.445 145.385 ;
        RECT 40.695 144.315 41.025 144.565 ;
        RECT 41.195 144.155 41.445 144.755 ;
        RECT 41.615 144.735 41.825 145.555 ;
        RECT 42.430 144.845 42.685 145.375 ;
        RECT 42.865 145.095 43.150 145.555 ;
        RECT 42.430 144.195 42.610 144.845 ;
        RECT 43.330 144.645 43.580 145.295 ;
        RECT 42.780 144.315 43.580 144.645 ;
        RECT 37.915 143.005 40.505 144.095 ;
        RECT 40.715 143.005 40.945 144.145 ;
        RECT 41.115 143.175 41.445 144.155 ;
        RECT 41.615 143.005 41.825 144.145 ;
        RECT 42.345 144.025 42.610 144.195 ;
        RECT 42.430 143.985 42.610 144.025 ;
        RECT 42.430 143.315 42.685 143.985 ;
        RECT 42.865 143.005 43.150 143.805 ;
        RECT 43.330 143.725 43.580 144.315 ;
        RECT 43.780 144.960 44.100 145.290 ;
        RECT 44.280 145.075 44.940 145.555 ;
        RECT 45.140 145.165 45.990 145.335 ;
        RECT 43.780 144.065 43.970 144.960 ;
        RECT 44.290 144.635 44.950 144.905 ;
        RECT 44.620 144.575 44.950 144.635 ;
        RECT 44.140 144.405 44.470 144.465 ;
        RECT 45.140 144.405 45.310 145.165 ;
        RECT 46.550 145.095 46.870 145.555 ;
        RECT 47.070 144.915 47.320 145.345 ;
        RECT 47.610 145.115 48.020 145.555 ;
        RECT 48.190 145.175 49.205 145.375 ;
        RECT 45.480 144.745 46.730 144.915 ;
        RECT 45.480 144.625 45.810 144.745 ;
        RECT 44.140 144.235 46.040 144.405 ;
        RECT 43.780 143.895 45.700 144.065 ;
        RECT 43.780 143.875 44.100 143.895 ;
        RECT 43.330 143.215 43.660 143.725 ;
        RECT 43.930 143.265 44.100 143.875 ;
        RECT 45.870 143.725 46.040 144.235 ;
        RECT 46.210 144.165 46.390 144.575 ;
        RECT 46.560 143.985 46.730 144.745 ;
        RECT 44.270 143.005 44.600 143.695 ;
        RECT 44.830 143.555 46.040 143.725 ;
        RECT 46.210 143.675 46.730 143.985 ;
        RECT 46.900 144.575 47.320 144.915 ;
        RECT 47.610 144.575 48.020 144.905 ;
        RECT 46.900 143.805 47.090 144.575 ;
        RECT 48.190 144.445 48.360 145.175 ;
        RECT 49.505 145.005 49.675 145.335 ;
        RECT 49.845 145.175 50.175 145.555 ;
        RECT 48.530 144.625 48.880 144.995 ;
        RECT 48.190 144.405 48.610 144.445 ;
        RECT 47.260 144.235 48.610 144.405 ;
        RECT 47.260 144.075 47.510 144.235 ;
        RECT 48.020 143.805 48.270 144.065 ;
        RECT 46.900 143.555 48.270 143.805 ;
        RECT 44.830 143.265 45.070 143.555 ;
        RECT 45.870 143.475 46.040 143.555 ;
        RECT 45.270 143.005 45.690 143.385 ;
        RECT 45.870 143.225 46.500 143.475 ;
        RECT 46.970 143.005 47.300 143.385 ;
        RECT 47.470 143.265 47.640 143.555 ;
        RECT 48.440 143.390 48.610 144.235 ;
        RECT 49.060 144.065 49.280 144.935 ;
        RECT 49.505 144.815 50.200 145.005 ;
        RECT 48.780 143.685 49.280 144.065 ;
        RECT 49.450 144.015 49.860 144.635 ;
        RECT 50.030 143.845 50.200 144.815 ;
        RECT 49.505 143.675 50.200 143.845 ;
        RECT 47.820 143.005 48.200 143.385 ;
        RECT 48.440 143.220 49.270 143.390 ;
        RECT 49.505 143.175 49.675 143.675 ;
        RECT 49.845 143.005 50.175 143.505 ;
        RECT 50.390 143.175 50.615 145.295 ;
        RECT 50.785 145.175 51.115 145.555 ;
        RECT 51.285 145.005 51.455 145.295 ;
        RECT 50.790 144.835 51.455 145.005 ;
        RECT 50.790 143.845 51.020 144.835 ;
        RECT 51.720 144.815 51.975 145.385 ;
        RECT 52.145 145.155 52.475 145.555 ;
        RECT 52.900 145.020 53.430 145.385 ;
        RECT 53.620 145.215 53.895 145.385 ;
        RECT 53.615 145.045 53.895 145.215 ;
        RECT 52.900 144.985 53.075 145.020 ;
        RECT 52.145 144.815 53.075 144.985 ;
        RECT 51.190 144.015 51.540 144.665 ;
        RECT 51.720 144.145 51.890 144.815 ;
        RECT 52.145 144.645 52.315 144.815 ;
        RECT 52.060 144.315 52.315 144.645 ;
        RECT 52.540 144.315 52.735 144.645 ;
        RECT 50.790 143.675 51.455 143.845 ;
        RECT 50.785 143.005 51.115 143.505 ;
        RECT 51.285 143.175 51.455 143.675 ;
        RECT 51.720 143.175 52.055 144.145 ;
        RECT 52.225 143.005 52.395 144.145 ;
        RECT 52.565 143.345 52.735 144.315 ;
        RECT 52.905 143.685 53.075 144.815 ;
        RECT 53.245 144.025 53.415 144.825 ;
        RECT 53.620 144.225 53.895 145.045 ;
        RECT 54.065 144.025 54.255 145.385 ;
        RECT 54.435 145.020 54.945 145.555 ;
        RECT 55.165 144.745 55.410 145.350 ;
        RECT 56.315 144.785 57.985 145.555 ;
        RECT 54.455 144.575 55.685 144.745 ;
        RECT 53.245 143.855 54.255 144.025 ;
        RECT 54.425 144.010 55.175 144.200 ;
        RECT 52.905 143.515 54.030 143.685 ;
        RECT 54.425 143.345 54.595 144.010 ;
        RECT 55.345 143.765 55.685 144.575 ;
        RECT 52.565 143.175 54.595 143.345 ;
        RECT 54.765 143.005 54.935 143.765 ;
        RECT 55.170 143.355 55.685 143.765 ;
        RECT 56.315 144.095 57.065 144.615 ;
        RECT 57.235 144.265 57.985 144.785 ;
        RECT 58.195 144.735 58.425 145.555 ;
        RECT 58.595 144.755 58.925 145.385 ;
        RECT 58.175 144.315 58.505 144.565 ;
        RECT 58.675 144.155 58.925 144.755 ;
        RECT 59.095 144.735 59.305 145.555 ;
        RECT 59.995 144.785 62.585 145.555 ;
        RECT 62.755 144.830 63.045 145.555 ;
        RECT 56.315 143.005 57.985 144.095 ;
        RECT 58.195 143.005 58.425 144.145 ;
        RECT 58.595 143.175 58.925 144.155 ;
        RECT 59.095 143.005 59.305 144.145 ;
        RECT 59.995 144.095 61.205 144.615 ;
        RECT 61.375 144.265 62.585 144.785 ;
        RECT 63.950 144.745 64.195 145.350 ;
        RECT 64.415 145.020 64.925 145.555 ;
        RECT 63.675 144.575 64.905 144.745 ;
        RECT 59.995 143.005 62.585 144.095 ;
        RECT 62.755 143.005 63.045 144.170 ;
        RECT 63.675 143.765 64.015 144.575 ;
        RECT 64.185 144.010 64.935 144.200 ;
        RECT 63.675 143.355 64.190 143.765 ;
        RECT 64.425 143.005 64.595 143.765 ;
        RECT 64.765 143.345 64.935 144.010 ;
        RECT 65.105 144.025 65.295 145.385 ;
        RECT 65.465 144.535 65.740 145.385 ;
        RECT 65.930 145.020 66.460 145.385 ;
        RECT 66.885 145.155 67.215 145.555 ;
        RECT 66.285 144.985 66.460 145.020 ;
        RECT 65.465 144.365 65.745 144.535 ;
        RECT 65.465 144.225 65.740 144.365 ;
        RECT 65.945 144.025 66.115 144.825 ;
        RECT 65.105 143.855 66.115 144.025 ;
        RECT 66.285 144.815 67.215 144.985 ;
        RECT 67.385 144.815 67.640 145.385 ;
        RECT 68.280 145.010 73.625 145.555 ;
        RECT 73.800 145.010 79.145 145.555 ;
        RECT 79.325 145.055 79.655 145.555 ;
        RECT 66.285 143.685 66.455 144.815 ;
        RECT 67.045 144.645 67.215 144.815 ;
        RECT 65.330 143.515 66.455 143.685 ;
        RECT 66.625 144.315 66.820 144.645 ;
        RECT 67.045 144.315 67.300 144.645 ;
        RECT 66.625 143.345 66.795 144.315 ;
        RECT 67.470 144.145 67.640 144.815 ;
        RECT 64.765 143.175 66.795 143.345 ;
        RECT 66.965 143.005 67.135 144.145 ;
        RECT 67.305 143.175 67.640 144.145 ;
        RECT 69.870 143.440 70.220 144.690 ;
        RECT 71.700 144.180 72.040 145.010 ;
        RECT 75.390 143.440 75.740 144.690 ;
        RECT 77.220 144.180 77.560 145.010 ;
        RECT 79.855 144.985 80.025 145.335 ;
        RECT 80.225 145.155 80.555 145.555 ;
        RECT 80.725 144.985 80.895 145.335 ;
        RECT 81.065 145.155 81.445 145.555 ;
        RECT 79.320 144.315 79.670 144.885 ;
        RECT 79.855 144.815 81.465 144.985 ;
        RECT 81.635 144.880 81.905 145.225 ;
        RECT 81.295 144.645 81.465 144.815 ;
        RECT 79.320 143.855 79.640 144.145 ;
        RECT 79.840 144.025 80.550 144.645 ;
        RECT 80.720 144.315 81.125 144.645 ;
        RECT 81.295 144.315 81.565 144.645 ;
        RECT 81.295 144.145 81.465 144.315 ;
        RECT 81.735 144.145 81.905 144.880 ;
        RECT 82.535 144.785 84.205 145.555 ;
        RECT 80.740 143.975 81.465 144.145 ;
        RECT 80.740 143.855 80.910 143.975 ;
        RECT 79.320 143.685 80.910 143.855 ;
        RECT 68.280 143.005 73.625 143.440 ;
        RECT 73.800 143.005 79.145 143.440 ;
        RECT 79.320 143.225 80.975 143.515 ;
        RECT 81.145 143.005 81.425 143.805 ;
        RECT 81.635 143.175 81.905 144.145 ;
        RECT 82.535 144.095 83.285 144.615 ;
        RECT 83.455 144.265 84.205 144.785 ;
        RECT 84.650 144.745 84.895 145.350 ;
        RECT 85.115 145.020 85.625 145.555 ;
        RECT 84.375 144.575 85.605 144.745 ;
        RECT 82.535 143.005 84.205 144.095 ;
        RECT 84.375 143.765 84.715 144.575 ;
        RECT 84.885 144.010 85.635 144.200 ;
        RECT 84.375 143.355 84.890 143.765 ;
        RECT 85.125 143.005 85.295 143.765 ;
        RECT 85.465 143.345 85.635 144.010 ;
        RECT 85.805 144.025 85.995 145.385 ;
        RECT 86.165 144.535 86.440 145.385 ;
        RECT 86.630 145.020 87.160 145.385 ;
        RECT 87.585 145.155 87.915 145.555 ;
        RECT 86.985 144.985 87.160 145.020 ;
        RECT 86.165 144.365 86.445 144.535 ;
        RECT 86.165 144.225 86.440 144.365 ;
        RECT 86.645 144.025 86.815 144.825 ;
        RECT 85.805 143.855 86.815 144.025 ;
        RECT 86.985 144.815 87.915 144.985 ;
        RECT 88.085 144.815 88.340 145.385 ;
        RECT 88.515 144.830 88.805 145.555 ;
        RECT 89.985 145.005 90.155 145.385 ;
        RECT 90.335 145.175 90.665 145.555 ;
        RECT 89.985 144.835 90.650 145.005 ;
        RECT 90.845 144.880 91.105 145.385 ;
        RECT 86.985 143.685 87.155 144.815 ;
        RECT 87.745 144.645 87.915 144.815 ;
        RECT 86.030 143.515 87.155 143.685 ;
        RECT 87.325 144.315 87.520 144.645 ;
        RECT 87.745 144.315 88.000 144.645 ;
        RECT 87.325 143.345 87.495 144.315 ;
        RECT 88.170 144.145 88.340 144.815 ;
        RECT 89.915 144.285 90.245 144.655 ;
        RECT 90.480 144.580 90.650 144.835 ;
        RECT 90.480 144.250 90.765 144.580 ;
        RECT 85.465 143.175 87.495 143.345 ;
        RECT 87.665 143.005 87.835 144.145 ;
        RECT 88.005 143.175 88.340 144.145 ;
        RECT 88.515 143.005 88.805 144.170 ;
        RECT 90.480 144.105 90.650 144.250 ;
        RECT 89.985 143.935 90.650 144.105 ;
        RECT 90.935 144.080 91.105 144.880 ;
        RECT 91.735 144.785 93.405 145.555 ;
        RECT 89.985 143.175 90.155 143.935 ;
        RECT 90.335 143.005 90.665 143.765 ;
        RECT 90.835 143.175 91.105 144.080 ;
        RECT 91.735 144.095 92.485 144.615 ;
        RECT 92.655 144.265 93.405 144.785 ;
        RECT 93.690 144.925 93.975 145.385 ;
        RECT 94.145 145.095 94.415 145.555 ;
        RECT 93.690 144.755 94.645 144.925 ;
        RECT 91.735 143.005 93.405 144.095 ;
        RECT 93.575 144.025 94.265 144.585 ;
        RECT 94.435 143.855 94.645 144.755 ;
        RECT 93.690 143.635 94.645 143.855 ;
        RECT 94.815 144.585 95.215 145.385 ;
        RECT 95.405 144.925 95.685 145.385 ;
        RECT 96.205 145.095 96.530 145.555 ;
        RECT 95.405 144.755 96.530 144.925 ;
        RECT 96.700 144.815 97.085 145.385 ;
        RECT 96.080 144.645 96.530 144.755 ;
        RECT 94.815 144.025 95.910 144.585 ;
        RECT 96.080 144.315 96.635 144.645 ;
        RECT 93.690 143.175 93.975 143.635 ;
        RECT 94.145 143.005 94.415 143.465 ;
        RECT 94.815 143.175 95.215 144.025 ;
        RECT 96.080 143.855 96.530 144.315 ;
        RECT 96.805 144.145 97.085 144.815 ;
        RECT 97.715 144.785 101.225 145.555 ;
        RECT 101.400 145.010 106.745 145.555 ;
        RECT 106.925 145.055 107.255 145.555 ;
        RECT 95.405 143.635 96.530 143.855 ;
        RECT 95.405 143.175 95.685 143.635 ;
        RECT 96.205 143.005 96.530 143.465 ;
        RECT 96.700 143.175 97.085 144.145 ;
        RECT 97.715 144.095 99.405 144.615 ;
        RECT 99.575 144.265 101.225 144.785 ;
        RECT 97.715 143.005 101.225 144.095 ;
        RECT 102.990 143.440 103.340 144.690 ;
        RECT 104.820 144.180 105.160 145.010 ;
        RECT 107.455 144.985 107.625 145.335 ;
        RECT 107.825 145.155 108.155 145.555 ;
        RECT 108.325 144.985 108.495 145.335 ;
        RECT 108.665 145.155 109.045 145.555 ;
        RECT 106.920 144.315 107.270 144.885 ;
        RECT 107.455 144.815 109.065 144.985 ;
        RECT 109.235 144.880 109.505 145.225 ;
        RECT 108.895 144.645 109.065 144.815 ;
        RECT 106.920 143.855 107.240 144.145 ;
        RECT 107.440 144.025 108.150 144.645 ;
        RECT 108.320 144.315 108.725 144.645 ;
        RECT 108.895 144.315 109.165 144.645 ;
        RECT 108.895 144.145 109.065 144.315 ;
        RECT 109.335 144.145 109.505 144.880 ;
        RECT 108.340 143.975 109.065 144.145 ;
        RECT 108.340 143.855 108.510 143.975 ;
        RECT 106.920 143.685 108.510 143.855 ;
        RECT 101.400 143.005 106.745 143.440 ;
        RECT 106.920 143.225 108.575 143.515 ;
        RECT 108.745 143.005 109.025 143.805 ;
        RECT 109.235 143.175 109.505 144.145 ;
        RECT 109.675 144.755 110.015 145.385 ;
        RECT 110.185 144.755 110.435 145.555 ;
        RECT 110.625 144.905 110.955 145.385 ;
        RECT 111.125 145.095 111.350 145.555 ;
        RECT 111.520 144.905 111.850 145.385 ;
        RECT 109.675 144.705 109.905 144.755 ;
        RECT 110.625 144.735 111.850 144.905 ;
        RECT 112.480 144.775 112.980 145.385 ;
        RECT 114.275 144.830 114.565 145.555 ;
        RECT 109.675 144.145 109.850 144.705 ;
        RECT 110.020 144.395 110.715 144.565 ;
        RECT 110.545 144.145 110.715 144.395 ;
        RECT 110.890 144.365 111.310 144.565 ;
        RECT 111.480 144.365 111.810 144.565 ;
        RECT 111.980 144.365 112.310 144.565 ;
        RECT 112.480 144.145 112.650 144.775 ;
        RECT 115.470 144.745 115.715 145.350 ;
        RECT 115.935 145.020 116.445 145.555 ;
        RECT 115.195 144.575 116.425 144.745 ;
        RECT 112.835 144.315 113.185 144.565 ;
        RECT 109.675 143.175 110.015 144.145 ;
        RECT 110.185 143.005 110.355 144.145 ;
        RECT 110.545 143.975 112.980 144.145 ;
        RECT 110.625 143.005 110.875 143.805 ;
        RECT 111.520 143.175 111.850 143.975 ;
        RECT 112.150 143.005 112.480 143.805 ;
        RECT 112.650 143.175 112.980 143.975 ;
        RECT 114.275 143.005 114.565 144.170 ;
        RECT 115.195 143.765 115.535 144.575 ;
        RECT 115.705 144.010 116.455 144.200 ;
        RECT 115.195 143.355 115.710 143.765 ;
        RECT 115.945 143.005 116.115 143.765 ;
        RECT 116.285 143.345 116.455 144.010 ;
        RECT 116.625 144.025 116.815 145.385 ;
        RECT 116.985 145.215 117.260 145.385 ;
        RECT 116.985 145.045 117.265 145.215 ;
        RECT 116.985 144.225 117.260 145.045 ;
        RECT 117.450 145.020 117.980 145.385 ;
        RECT 118.405 145.155 118.735 145.555 ;
        RECT 117.805 144.985 117.980 145.020 ;
        RECT 117.465 144.025 117.635 144.825 ;
        RECT 116.625 143.855 117.635 144.025 ;
        RECT 117.805 144.815 118.735 144.985 ;
        RECT 118.905 144.815 119.160 145.385 ;
        RECT 117.805 143.685 117.975 144.815 ;
        RECT 118.565 144.645 118.735 144.815 ;
        RECT 116.850 143.515 117.975 143.685 ;
        RECT 118.145 144.315 118.340 144.645 ;
        RECT 118.565 144.315 118.820 144.645 ;
        RECT 118.145 143.345 118.315 144.315 ;
        RECT 118.990 144.145 119.160 144.815 ;
        RECT 119.375 144.735 119.605 145.555 ;
        RECT 119.775 144.755 120.105 145.385 ;
        RECT 119.355 144.315 119.685 144.565 ;
        RECT 119.855 144.155 120.105 144.755 ;
        RECT 120.275 144.735 120.485 145.555 ;
        RECT 121.265 145.005 121.435 145.385 ;
        RECT 121.615 145.175 121.945 145.555 ;
        RECT 121.265 144.835 121.930 145.005 ;
        RECT 122.125 144.880 122.385 145.385 ;
        RECT 121.195 144.285 121.525 144.655 ;
        RECT 121.760 144.580 121.930 144.835 ;
        RECT 116.285 143.175 118.315 143.345 ;
        RECT 118.485 143.005 118.655 144.145 ;
        RECT 118.825 143.175 119.160 144.145 ;
        RECT 119.375 143.005 119.605 144.145 ;
        RECT 119.775 143.175 120.105 144.155 ;
        RECT 121.760 144.250 122.045 144.580 ;
        RECT 120.275 143.005 120.485 144.145 ;
        RECT 121.760 144.105 121.930 144.250 ;
        RECT 121.265 143.935 121.930 144.105 ;
        RECT 122.215 144.080 122.385 144.880 ;
        RECT 122.555 144.785 126.065 145.555 ;
        RECT 126.235 144.805 127.445 145.555 ;
        RECT 121.265 143.175 121.435 143.935 ;
        RECT 121.615 143.005 121.945 143.765 ;
        RECT 122.115 143.175 122.385 144.080 ;
        RECT 122.555 144.095 124.245 144.615 ;
        RECT 124.415 144.265 126.065 144.785 ;
        RECT 126.235 144.095 126.755 144.635 ;
        RECT 126.925 144.265 127.445 144.805 ;
        RECT 122.555 143.005 126.065 144.095 ;
        RECT 126.235 143.005 127.445 144.095 ;
        RECT 14.370 142.835 127.530 143.005 ;
        RECT 14.455 141.745 15.665 142.835 ;
        RECT 14.455 141.035 14.975 141.575 ;
        RECT 15.145 141.205 15.665 141.745 ;
        RECT 15.835 141.745 18.425 142.835 ;
        RECT 18.600 142.400 23.945 142.835 ;
        RECT 15.835 141.225 17.045 141.745 ;
        RECT 17.215 141.055 18.425 141.575 ;
        RECT 20.190 141.150 20.540 142.400 ;
        RECT 24.115 141.670 24.405 142.835 ;
        RECT 25.035 141.745 28.545 142.835 ;
        RECT 28.720 142.400 34.065 142.835 ;
        RECT 14.455 140.285 15.665 141.035 ;
        RECT 15.835 140.285 18.425 141.055 ;
        RECT 22.020 140.830 22.360 141.660 ;
        RECT 25.035 141.225 26.725 141.745 ;
        RECT 26.895 141.055 28.545 141.575 ;
        RECT 30.310 141.150 30.660 142.400 ;
        RECT 34.235 141.695 34.505 142.665 ;
        RECT 34.715 142.035 34.995 142.835 ;
        RECT 35.165 142.325 36.820 142.615 ;
        RECT 35.230 141.985 36.820 142.155 ;
        RECT 35.230 141.865 35.400 141.985 ;
        RECT 34.675 141.695 35.400 141.865 ;
        RECT 18.600 140.285 23.945 140.830 ;
        RECT 24.115 140.285 24.405 141.010 ;
        RECT 25.035 140.285 28.545 141.055 ;
        RECT 32.140 140.830 32.480 141.660 ;
        RECT 34.235 140.960 34.405 141.695 ;
        RECT 34.675 141.525 34.845 141.695 ;
        RECT 34.575 141.195 34.845 141.525 ;
        RECT 35.015 141.195 35.420 141.525 ;
        RECT 35.590 141.195 36.300 141.815 ;
        RECT 36.500 141.695 36.820 141.985 ;
        RECT 37.915 141.745 41.425 142.835 ;
        RECT 41.600 142.400 46.945 142.835 ;
        RECT 34.675 141.025 34.845 141.195 ;
        RECT 28.720 140.285 34.065 140.830 ;
        RECT 34.235 140.615 34.505 140.960 ;
        RECT 34.675 140.855 36.285 141.025 ;
        RECT 36.470 140.955 36.820 141.525 ;
        RECT 37.915 141.225 39.605 141.745 ;
        RECT 39.775 141.055 41.425 141.575 ;
        RECT 43.190 141.150 43.540 142.400 ;
        RECT 47.115 141.695 47.385 142.665 ;
        RECT 47.595 142.035 47.875 142.835 ;
        RECT 48.045 142.325 49.700 142.615 ;
        RECT 48.110 141.985 49.700 142.155 ;
        RECT 48.110 141.865 48.280 141.985 ;
        RECT 47.555 141.695 48.280 141.865 ;
        RECT 34.695 140.285 35.075 140.685 ;
        RECT 35.245 140.505 35.415 140.855 ;
        RECT 35.585 140.285 35.915 140.685 ;
        RECT 36.115 140.505 36.285 140.855 ;
        RECT 36.485 140.285 36.815 140.785 ;
        RECT 37.915 140.285 41.425 141.055 ;
        RECT 45.020 140.830 45.360 141.660 ;
        RECT 47.115 140.960 47.285 141.695 ;
        RECT 47.555 141.525 47.725 141.695 ;
        RECT 47.455 141.195 47.725 141.525 ;
        RECT 47.895 141.195 48.300 141.525 ;
        RECT 48.470 141.195 49.180 141.815 ;
        RECT 49.380 141.695 49.700 141.985 ;
        RECT 49.875 141.670 50.165 142.835 ;
        RECT 50.335 141.745 52.005 142.835 ;
        RECT 47.555 141.025 47.725 141.195 ;
        RECT 41.600 140.285 46.945 140.830 ;
        RECT 47.115 140.615 47.385 140.960 ;
        RECT 47.555 140.855 49.165 141.025 ;
        RECT 49.350 140.955 49.700 141.525 ;
        RECT 50.335 141.225 51.085 141.745 ;
        RECT 52.175 141.695 52.515 142.665 ;
        RECT 52.685 141.695 52.855 142.835 ;
        RECT 53.125 142.035 53.375 142.835 ;
        RECT 54.020 141.865 54.350 142.665 ;
        RECT 54.650 142.035 54.980 142.835 ;
        RECT 55.150 141.865 55.480 142.665 ;
        RECT 55.970 142.205 56.255 142.665 ;
        RECT 56.425 142.375 56.695 142.835 ;
        RECT 55.970 141.985 56.925 142.205 ;
        RECT 53.045 141.695 55.480 141.865 ;
        RECT 51.255 141.055 52.005 141.575 ;
        RECT 47.575 140.285 47.955 140.685 ;
        RECT 48.125 140.505 48.295 140.855 ;
        RECT 48.465 140.285 48.795 140.685 ;
        RECT 48.995 140.505 49.165 140.855 ;
        RECT 49.365 140.285 49.695 140.785 ;
        RECT 49.875 140.285 50.165 141.010 ;
        RECT 50.335 140.285 52.005 141.055 ;
        RECT 52.175 141.135 52.350 141.695 ;
        RECT 53.045 141.445 53.215 141.695 ;
        RECT 52.520 141.275 53.215 141.445 ;
        RECT 53.390 141.275 53.810 141.475 ;
        RECT 53.980 141.275 54.310 141.475 ;
        RECT 54.480 141.275 54.810 141.475 ;
        RECT 52.175 141.085 52.405 141.135 ;
        RECT 52.175 140.455 52.515 141.085 ;
        RECT 52.685 140.285 52.935 141.085 ;
        RECT 53.125 140.935 54.350 141.105 ;
        RECT 53.125 140.455 53.455 140.935 ;
        RECT 53.625 140.285 53.850 140.745 ;
        RECT 54.020 140.455 54.350 140.935 ;
        RECT 54.980 141.065 55.150 141.695 ;
        RECT 55.335 141.275 55.685 141.525 ;
        RECT 55.855 141.255 56.545 141.815 ;
        RECT 56.715 141.085 56.925 141.985 ;
        RECT 54.980 140.455 55.480 141.065 ;
        RECT 55.970 140.915 56.925 141.085 ;
        RECT 57.095 141.815 57.495 142.665 ;
        RECT 57.685 142.205 57.965 142.665 ;
        RECT 58.485 142.375 58.810 142.835 ;
        RECT 57.685 141.985 58.810 142.205 ;
        RECT 57.095 141.255 58.190 141.815 ;
        RECT 58.360 141.525 58.810 141.985 ;
        RECT 58.980 141.695 59.365 142.665 ;
        RECT 55.970 140.455 56.255 140.915 ;
        RECT 56.425 140.285 56.695 140.745 ;
        RECT 57.095 140.455 57.495 141.255 ;
        RECT 58.360 141.195 58.915 141.525 ;
        RECT 58.360 141.085 58.810 141.195 ;
        RECT 57.685 140.915 58.810 141.085 ;
        RECT 59.085 141.025 59.365 141.695 ;
        RECT 57.685 140.455 57.965 140.915 ;
        RECT 58.485 140.285 58.810 140.745 ;
        RECT 58.980 140.455 59.365 141.025 ;
        RECT 59.540 141.645 59.795 142.525 ;
        RECT 59.965 141.695 60.270 142.835 ;
        RECT 60.610 142.455 60.940 142.835 ;
        RECT 61.120 142.285 61.290 142.575 ;
        RECT 61.460 142.375 61.710 142.835 ;
        RECT 60.490 142.115 61.290 142.285 ;
        RECT 61.880 142.325 62.750 142.665 ;
        RECT 59.540 140.995 59.750 141.645 ;
        RECT 60.490 141.525 60.660 142.115 ;
        RECT 61.880 141.945 62.050 142.325 ;
        RECT 62.985 142.205 63.155 142.665 ;
        RECT 63.325 142.375 63.695 142.835 ;
        RECT 63.990 142.235 64.160 142.575 ;
        RECT 64.330 142.405 64.660 142.835 ;
        RECT 64.895 142.235 65.065 142.575 ;
        RECT 60.830 141.775 62.050 141.945 ;
        RECT 62.220 141.865 62.680 142.155 ;
        RECT 62.985 142.035 63.545 142.205 ;
        RECT 63.990 142.065 65.065 142.235 ;
        RECT 65.235 142.335 65.915 142.665 ;
        RECT 66.130 142.335 66.380 142.665 ;
        RECT 66.550 142.375 66.800 142.835 ;
        RECT 63.375 141.895 63.545 142.035 ;
        RECT 62.220 141.855 63.185 141.865 ;
        RECT 61.880 141.685 62.050 141.775 ;
        RECT 62.510 141.695 63.185 141.855 ;
        RECT 59.920 141.495 60.660 141.525 ;
        RECT 59.920 141.195 60.835 141.495 ;
        RECT 60.510 141.020 60.835 141.195 ;
        RECT 59.540 140.465 59.795 140.995 ;
        RECT 59.965 140.285 60.270 140.745 ;
        RECT 60.515 140.665 60.835 141.020 ;
        RECT 61.005 141.235 61.545 141.605 ;
        RECT 61.880 141.515 62.285 141.685 ;
        RECT 61.005 140.835 61.245 141.235 ;
        RECT 61.725 141.065 61.945 141.345 ;
        RECT 61.415 140.895 61.945 141.065 ;
        RECT 61.415 140.665 61.585 140.895 ;
        RECT 62.115 140.735 62.285 141.515 ;
        RECT 62.455 140.905 62.805 141.525 ;
        RECT 62.975 140.905 63.185 141.695 ;
        RECT 63.375 141.725 64.875 141.895 ;
        RECT 63.375 141.035 63.545 141.725 ;
        RECT 65.235 141.555 65.405 142.335 ;
        RECT 66.210 142.205 66.380 142.335 ;
        RECT 63.715 141.385 65.405 141.555 ;
        RECT 65.575 141.775 66.040 142.165 ;
        RECT 66.210 142.035 66.605 142.205 ;
        RECT 63.715 141.205 63.885 141.385 ;
        RECT 60.515 140.495 61.585 140.665 ;
        RECT 61.755 140.285 61.945 140.725 ;
        RECT 62.115 140.455 63.065 140.735 ;
        RECT 63.375 140.645 63.635 141.035 ;
        RECT 64.055 140.965 64.845 141.215 ;
        RECT 63.285 140.475 63.635 140.645 ;
        RECT 63.845 140.285 64.175 140.745 ;
        RECT 65.050 140.675 65.220 141.385 ;
        RECT 65.575 141.185 65.745 141.775 ;
        RECT 65.390 140.965 65.745 141.185 ;
        RECT 65.915 140.965 66.265 141.585 ;
        RECT 66.435 140.675 66.605 142.035 ;
        RECT 66.970 141.865 67.295 142.650 ;
        RECT 66.775 140.815 67.235 141.865 ;
        RECT 65.050 140.505 65.905 140.675 ;
        RECT 66.110 140.505 66.605 140.675 ;
        RECT 66.775 140.285 67.105 140.645 ;
        RECT 67.465 140.545 67.635 142.665 ;
        RECT 67.805 142.335 68.135 142.835 ;
        RECT 68.305 142.165 68.560 142.665 ;
        RECT 67.810 141.995 68.560 142.165 ;
        RECT 67.810 141.005 68.040 141.995 ;
        RECT 68.210 141.175 68.560 141.825 ;
        RECT 68.735 141.760 69.005 142.665 ;
        RECT 69.175 142.075 69.505 142.835 ;
        RECT 69.685 141.905 69.855 142.665 ;
        RECT 67.810 140.835 68.560 141.005 ;
        RECT 67.805 140.285 68.135 140.665 ;
        RECT 68.305 140.545 68.560 140.835 ;
        RECT 68.735 140.960 68.905 141.760 ;
        RECT 69.190 141.735 69.855 141.905 ;
        RECT 70.115 141.745 71.325 142.835 ;
        RECT 69.190 141.590 69.360 141.735 ;
        RECT 69.075 141.260 69.360 141.590 ;
        RECT 69.190 141.005 69.360 141.260 ;
        RECT 69.595 141.185 69.925 141.555 ;
        RECT 70.115 141.205 70.635 141.745 ;
        RECT 71.555 141.695 71.765 142.835 ;
        RECT 71.935 141.685 72.265 142.665 ;
        RECT 72.435 141.695 72.665 142.835 ;
        RECT 72.875 141.745 75.465 142.835 ;
        RECT 70.805 141.035 71.325 141.575 ;
        RECT 68.735 140.455 68.995 140.960 ;
        RECT 69.190 140.835 69.855 141.005 ;
        RECT 69.175 140.285 69.505 140.665 ;
        RECT 69.685 140.455 69.855 140.835 ;
        RECT 70.115 140.285 71.325 141.035 ;
        RECT 71.555 140.285 71.765 141.105 ;
        RECT 71.935 141.085 72.185 141.685 ;
        RECT 72.355 141.275 72.685 141.525 ;
        RECT 72.875 141.225 74.085 141.745 ;
        RECT 75.635 141.670 75.925 142.835 ;
        RECT 76.555 141.745 79.145 142.835 ;
        RECT 79.320 142.400 84.665 142.835 ;
        RECT 84.840 142.400 90.185 142.835 ;
        RECT 90.360 142.400 95.705 142.835 ;
        RECT 95.880 142.400 101.225 142.835 ;
        RECT 71.935 140.455 72.265 141.085 ;
        RECT 72.435 140.285 72.665 141.105 ;
        RECT 74.255 141.055 75.465 141.575 ;
        RECT 76.555 141.225 77.765 141.745 ;
        RECT 77.935 141.055 79.145 141.575 ;
        RECT 80.910 141.150 81.260 142.400 ;
        RECT 72.875 140.285 75.465 141.055 ;
        RECT 75.635 140.285 75.925 141.010 ;
        RECT 76.555 140.285 79.145 141.055 ;
        RECT 82.740 140.830 83.080 141.660 ;
        RECT 86.430 141.150 86.780 142.400 ;
        RECT 88.260 140.830 88.600 141.660 ;
        RECT 91.950 141.150 92.300 142.400 ;
        RECT 93.780 140.830 94.120 141.660 ;
        RECT 97.470 141.150 97.820 142.400 ;
        RECT 101.395 141.670 101.685 142.835 ;
        RECT 101.855 141.745 104.445 142.835 ;
        RECT 104.620 142.400 109.965 142.835 ;
        RECT 110.140 142.400 115.485 142.835 ;
        RECT 99.300 140.830 99.640 141.660 ;
        RECT 101.855 141.225 103.065 141.745 ;
        RECT 103.235 141.055 104.445 141.575 ;
        RECT 106.210 141.150 106.560 142.400 ;
        RECT 79.320 140.285 84.665 140.830 ;
        RECT 84.840 140.285 90.185 140.830 ;
        RECT 90.360 140.285 95.705 140.830 ;
        RECT 95.880 140.285 101.225 140.830 ;
        RECT 101.395 140.285 101.685 141.010 ;
        RECT 101.855 140.285 104.445 141.055 ;
        RECT 108.040 140.830 108.380 141.660 ;
        RECT 111.730 141.150 112.080 142.400 ;
        RECT 115.655 142.075 116.170 142.485 ;
        RECT 116.405 142.075 116.575 142.835 ;
        RECT 116.745 142.495 118.775 142.665 ;
        RECT 113.560 140.830 113.900 141.660 ;
        RECT 115.655 141.265 115.995 142.075 ;
        RECT 116.745 141.830 116.915 142.495 ;
        RECT 117.310 142.155 118.435 142.325 ;
        RECT 116.165 141.640 116.915 141.830 ;
        RECT 117.085 141.815 118.095 141.985 ;
        RECT 115.655 141.095 116.885 141.265 ;
        RECT 104.620 140.285 109.965 140.830 ;
        RECT 110.140 140.285 115.485 140.830 ;
        RECT 115.930 140.490 116.175 141.095 ;
        RECT 116.395 140.285 116.905 140.820 ;
        RECT 117.085 140.455 117.275 141.815 ;
        RECT 117.445 141.475 117.720 141.615 ;
        RECT 117.445 141.305 117.725 141.475 ;
        RECT 117.445 140.455 117.720 141.305 ;
        RECT 117.925 141.015 118.095 141.815 ;
        RECT 118.265 141.025 118.435 142.155 ;
        RECT 118.605 141.525 118.775 142.495 ;
        RECT 118.945 141.695 119.115 142.835 ;
        RECT 119.285 141.695 119.620 142.665 ;
        RECT 119.835 141.695 120.065 142.835 ;
        RECT 118.605 141.195 118.800 141.525 ;
        RECT 119.025 141.195 119.280 141.525 ;
        RECT 119.025 141.025 119.195 141.195 ;
        RECT 119.450 141.025 119.620 141.695 ;
        RECT 120.235 141.685 120.565 142.665 ;
        RECT 120.735 141.695 120.945 142.835 ;
        RECT 121.175 141.745 122.385 142.835 ;
        RECT 122.555 141.745 126.065 142.835 ;
        RECT 126.235 141.745 127.445 142.835 ;
        RECT 119.815 141.275 120.145 141.525 ;
        RECT 118.265 140.855 119.195 141.025 ;
        RECT 118.265 140.820 118.440 140.855 ;
        RECT 117.910 140.455 118.440 140.820 ;
        RECT 118.865 140.285 119.195 140.685 ;
        RECT 119.365 140.455 119.620 141.025 ;
        RECT 119.835 140.285 120.065 141.105 ;
        RECT 120.315 141.085 120.565 141.685 ;
        RECT 121.175 141.205 121.695 141.745 ;
        RECT 120.235 140.455 120.565 141.085 ;
        RECT 120.735 140.285 120.945 141.105 ;
        RECT 121.865 141.035 122.385 141.575 ;
        RECT 122.555 141.225 124.245 141.745 ;
        RECT 124.415 141.055 126.065 141.575 ;
        RECT 126.235 141.205 126.755 141.745 ;
        RECT 121.175 140.285 122.385 141.035 ;
        RECT 122.555 140.285 126.065 141.055 ;
        RECT 126.925 141.035 127.445 141.575 ;
        RECT 126.235 140.285 127.445 141.035 ;
        RECT 14.370 140.115 127.530 140.285 ;
        RECT 14.455 139.365 15.665 140.115 ;
        RECT 16.210 139.405 16.465 139.935 ;
        RECT 16.645 139.655 16.930 140.115 ;
        RECT 14.455 138.825 14.975 139.365 ;
        RECT 15.145 138.655 15.665 139.195 ;
        RECT 14.455 137.565 15.665 138.655 ;
        RECT 16.210 138.545 16.390 139.405 ;
        RECT 17.110 139.205 17.360 139.855 ;
        RECT 16.560 138.875 17.360 139.205 ;
        RECT 16.210 138.075 16.465 138.545 ;
        RECT 16.125 137.905 16.465 138.075 ;
        RECT 16.210 137.875 16.465 137.905 ;
        RECT 16.645 137.565 16.930 138.365 ;
        RECT 17.110 138.285 17.360 138.875 ;
        RECT 17.560 139.520 17.880 139.850 ;
        RECT 18.060 139.635 18.720 140.115 ;
        RECT 18.920 139.725 19.770 139.895 ;
        RECT 17.560 138.625 17.750 139.520 ;
        RECT 18.070 139.195 18.730 139.465 ;
        RECT 18.400 139.135 18.730 139.195 ;
        RECT 17.920 138.965 18.250 139.025 ;
        RECT 18.920 138.965 19.090 139.725 ;
        RECT 20.330 139.655 20.650 140.115 ;
        RECT 20.850 139.475 21.100 139.905 ;
        RECT 21.390 139.675 21.800 140.115 ;
        RECT 21.970 139.735 22.985 139.935 ;
        RECT 19.260 139.305 20.510 139.475 ;
        RECT 19.260 139.185 19.590 139.305 ;
        RECT 17.920 138.795 19.820 138.965 ;
        RECT 17.560 138.455 19.480 138.625 ;
        RECT 17.560 138.435 17.880 138.455 ;
        RECT 17.110 137.775 17.440 138.285 ;
        RECT 17.710 137.825 17.880 138.435 ;
        RECT 19.650 138.285 19.820 138.795 ;
        RECT 19.990 138.725 20.170 139.135 ;
        RECT 20.340 138.545 20.510 139.305 ;
        RECT 18.050 137.565 18.380 138.255 ;
        RECT 18.610 138.115 19.820 138.285 ;
        RECT 19.990 138.235 20.510 138.545 ;
        RECT 20.680 139.135 21.100 139.475 ;
        RECT 21.390 139.135 21.800 139.465 ;
        RECT 20.680 138.365 20.870 139.135 ;
        RECT 21.970 139.005 22.140 139.735 ;
        RECT 23.285 139.565 23.455 139.895 ;
        RECT 23.625 139.735 23.955 140.115 ;
        RECT 22.310 139.185 22.660 139.555 ;
        RECT 21.970 138.965 22.390 139.005 ;
        RECT 21.040 138.795 22.390 138.965 ;
        RECT 21.040 138.635 21.290 138.795 ;
        RECT 21.800 138.365 22.050 138.625 ;
        RECT 20.680 138.115 22.050 138.365 ;
        RECT 18.610 137.825 18.850 138.115 ;
        RECT 19.650 138.035 19.820 138.115 ;
        RECT 19.050 137.565 19.470 137.945 ;
        RECT 19.650 137.785 20.280 138.035 ;
        RECT 20.750 137.565 21.080 137.945 ;
        RECT 21.250 137.825 21.420 138.115 ;
        RECT 22.220 137.950 22.390 138.795 ;
        RECT 22.840 138.625 23.060 139.495 ;
        RECT 23.285 139.375 23.980 139.565 ;
        RECT 22.560 138.245 23.060 138.625 ;
        RECT 23.230 138.575 23.640 139.195 ;
        RECT 23.810 138.405 23.980 139.375 ;
        RECT 23.285 138.235 23.980 138.405 ;
        RECT 21.600 137.565 21.980 137.945 ;
        RECT 22.220 137.780 23.050 137.950 ;
        RECT 23.285 137.735 23.455 138.235 ;
        RECT 23.625 137.565 23.955 138.065 ;
        RECT 24.170 137.735 24.395 139.855 ;
        RECT 24.565 139.735 24.895 140.115 ;
        RECT 25.065 139.565 25.235 139.855 ;
        RECT 24.570 139.395 25.235 139.565 ;
        RECT 24.570 138.405 24.800 139.395 ;
        RECT 25.495 139.345 28.085 140.115 ;
        RECT 28.260 139.570 33.605 140.115 ;
        RECT 24.970 138.575 25.320 139.225 ;
        RECT 25.495 138.655 26.705 139.175 ;
        RECT 26.875 138.825 28.085 139.345 ;
        RECT 24.570 138.235 25.235 138.405 ;
        RECT 24.565 137.565 24.895 138.065 ;
        RECT 25.065 137.735 25.235 138.235 ;
        RECT 25.495 137.565 28.085 138.655 ;
        RECT 29.850 138.000 30.200 139.250 ;
        RECT 31.680 138.740 32.020 139.570 ;
        RECT 33.975 139.485 34.305 139.845 ;
        RECT 34.925 139.655 35.175 140.115 ;
        RECT 35.345 139.655 35.905 139.945 ;
        RECT 33.975 139.295 35.365 139.485 ;
        RECT 35.195 139.205 35.365 139.295 ;
        RECT 33.790 138.875 34.465 139.125 ;
        RECT 34.685 138.875 35.025 139.125 ;
        RECT 35.195 138.875 35.485 139.205 ;
        RECT 33.790 138.515 34.055 138.875 ;
        RECT 35.195 138.625 35.365 138.875 ;
        RECT 34.425 138.455 35.365 138.625 ;
        RECT 28.260 137.565 33.605 138.000 ;
        RECT 33.975 137.565 34.255 138.235 ;
        RECT 34.425 137.905 34.725 138.455 ;
        RECT 35.655 138.285 35.905 139.655 ;
        RECT 36.995 139.390 37.285 140.115 ;
        RECT 38.375 139.440 38.645 139.785 ;
        RECT 38.835 139.715 39.215 140.115 ;
        RECT 39.385 139.545 39.555 139.895 ;
        RECT 39.725 139.715 40.055 140.115 ;
        RECT 40.255 139.545 40.425 139.895 ;
        RECT 40.625 139.615 40.955 140.115 ;
        RECT 34.925 137.565 35.255 138.285 ;
        RECT 35.445 137.735 35.905 138.285 ;
        RECT 36.995 137.565 37.285 138.730 ;
        RECT 38.375 138.705 38.545 139.440 ;
        RECT 38.815 139.375 40.425 139.545 ;
        RECT 38.815 139.205 38.985 139.375 ;
        RECT 38.715 138.875 38.985 139.205 ;
        RECT 39.155 138.875 39.560 139.205 ;
        RECT 38.815 138.705 38.985 138.875 ;
        RECT 38.375 137.735 38.645 138.705 ;
        RECT 38.815 138.535 39.540 138.705 ;
        RECT 39.730 138.585 40.440 139.205 ;
        RECT 40.610 138.875 40.960 139.445 ;
        RECT 41.595 139.345 44.185 140.115 ;
        RECT 44.360 139.570 49.705 140.115 ;
        RECT 49.880 139.570 55.225 140.115 ;
        RECT 39.370 138.415 39.540 138.535 ;
        RECT 40.640 138.415 40.960 138.705 ;
        RECT 38.855 137.565 39.135 138.365 ;
        RECT 39.370 138.245 40.960 138.415 ;
        RECT 41.595 138.655 42.805 139.175 ;
        RECT 42.975 138.825 44.185 139.345 ;
        RECT 39.305 137.785 40.960 138.075 ;
        RECT 41.595 137.565 44.185 138.655 ;
        RECT 45.950 138.000 46.300 139.250 ;
        RECT 47.780 138.740 48.120 139.570 ;
        RECT 51.470 138.000 51.820 139.250 ;
        RECT 53.300 138.740 53.640 139.570 ;
        RECT 55.435 139.295 55.665 140.115 ;
        RECT 55.835 139.315 56.165 139.945 ;
        RECT 55.415 138.875 55.745 139.125 ;
        RECT 55.915 138.715 56.165 139.315 ;
        RECT 56.335 139.295 56.545 140.115 ;
        RECT 57.235 139.345 58.905 140.115 ;
        RECT 44.360 137.565 49.705 138.000 ;
        RECT 49.880 137.565 55.225 138.000 ;
        RECT 55.435 137.565 55.665 138.705 ;
        RECT 55.835 137.735 56.165 138.715 ;
        RECT 56.335 137.565 56.545 138.705 ;
        RECT 57.235 138.655 57.985 139.175 ;
        RECT 58.155 138.825 58.905 139.345 ;
        RECT 59.075 139.315 59.415 139.945 ;
        RECT 59.585 139.315 59.835 140.115 ;
        RECT 60.025 139.465 60.355 139.945 ;
        RECT 60.525 139.655 60.750 140.115 ;
        RECT 60.920 139.465 61.250 139.945 ;
        RECT 59.075 138.705 59.250 139.315 ;
        RECT 60.025 139.295 61.250 139.465 ;
        RECT 61.880 139.335 62.380 139.945 ;
        RECT 62.755 139.390 63.045 140.115 ;
        RECT 59.420 138.955 60.115 139.125 ;
        RECT 59.945 138.705 60.115 138.955 ;
        RECT 60.290 138.925 60.710 139.125 ;
        RECT 60.880 138.925 61.210 139.125 ;
        RECT 61.380 138.925 61.710 139.125 ;
        RECT 61.880 138.705 62.050 139.335 ;
        RECT 63.675 139.315 64.015 139.945 ;
        RECT 64.185 139.315 64.435 140.115 ;
        RECT 64.625 139.465 64.955 139.945 ;
        RECT 65.125 139.655 65.350 140.115 ;
        RECT 65.520 139.465 65.850 139.945 ;
        RECT 62.235 138.875 62.585 139.125 ;
        RECT 57.235 137.565 58.905 138.655 ;
        RECT 59.075 137.735 59.415 138.705 ;
        RECT 59.585 137.565 59.755 138.705 ;
        RECT 59.945 138.535 62.380 138.705 ;
        RECT 60.025 137.565 60.275 138.365 ;
        RECT 60.920 137.735 61.250 138.535 ;
        RECT 61.550 137.565 61.880 138.365 ;
        RECT 62.050 137.735 62.380 138.535 ;
        RECT 62.755 137.565 63.045 138.730 ;
        RECT 63.675 138.705 63.850 139.315 ;
        RECT 64.625 139.295 65.850 139.465 ;
        RECT 66.480 139.335 66.980 139.945 ;
        RECT 67.730 139.775 67.985 139.935 ;
        RECT 67.645 139.605 67.985 139.775 ;
        RECT 68.165 139.655 68.450 140.115 ;
        RECT 67.730 139.405 67.985 139.605 ;
        RECT 64.020 138.955 64.715 139.125 ;
        RECT 64.545 138.705 64.715 138.955 ;
        RECT 64.890 138.925 65.310 139.125 ;
        RECT 65.480 138.925 65.810 139.125 ;
        RECT 65.980 138.925 66.310 139.125 ;
        RECT 66.480 138.705 66.650 139.335 ;
        RECT 66.835 138.875 67.185 139.125 ;
        RECT 63.675 137.735 64.015 138.705 ;
        RECT 64.185 137.565 64.355 138.705 ;
        RECT 64.545 138.535 66.980 138.705 ;
        RECT 64.625 137.565 64.875 138.365 ;
        RECT 65.520 137.735 65.850 138.535 ;
        RECT 66.150 137.565 66.480 138.365 ;
        RECT 66.650 137.735 66.980 138.535 ;
        RECT 67.730 138.545 67.910 139.405 ;
        RECT 68.630 139.205 68.880 139.855 ;
        RECT 68.080 138.875 68.880 139.205 ;
        RECT 67.730 137.875 67.985 138.545 ;
        RECT 68.165 137.565 68.450 138.365 ;
        RECT 68.630 138.285 68.880 138.875 ;
        RECT 69.080 139.520 69.400 139.850 ;
        RECT 69.580 139.635 70.240 140.115 ;
        RECT 70.440 139.725 71.290 139.895 ;
        RECT 69.080 138.625 69.270 139.520 ;
        RECT 69.590 139.195 70.250 139.465 ;
        RECT 69.920 139.135 70.250 139.195 ;
        RECT 69.440 138.965 69.770 139.025 ;
        RECT 70.440 138.965 70.610 139.725 ;
        RECT 71.850 139.655 72.170 140.115 ;
        RECT 72.370 139.475 72.620 139.905 ;
        RECT 72.910 139.675 73.320 140.115 ;
        RECT 73.490 139.735 74.505 139.935 ;
        RECT 70.780 139.305 72.030 139.475 ;
        RECT 70.780 139.185 71.110 139.305 ;
        RECT 69.440 138.795 71.340 138.965 ;
        RECT 69.080 138.455 71.000 138.625 ;
        RECT 69.080 138.435 69.400 138.455 ;
        RECT 68.630 137.775 68.960 138.285 ;
        RECT 69.230 137.825 69.400 138.435 ;
        RECT 71.170 138.285 71.340 138.795 ;
        RECT 71.510 138.725 71.690 139.135 ;
        RECT 71.860 138.545 72.030 139.305 ;
        RECT 69.570 137.565 69.900 138.255 ;
        RECT 70.130 138.115 71.340 138.285 ;
        RECT 71.510 138.235 72.030 138.545 ;
        RECT 72.200 139.135 72.620 139.475 ;
        RECT 72.910 139.135 73.320 139.465 ;
        RECT 72.200 138.365 72.390 139.135 ;
        RECT 73.490 139.005 73.660 139.735 ;
        RECT 74.805 139.565 74.975 139.895 ;
        RECT 75.145 139.735 75.475 140.115 ;
        RECT 73.830 139.185 74.180 139.555 ;
        RECT 73.490 138.965 73.910 139.005 ;
        RECT 72.560 138.795 73.910 138.965 ;
        RECT 72.560 138.635 72.810 138.795 ;
        RECT 73.320 138.365 73.570 138.625 ;
        RECT 72.200 138.115 73.570 138.365 ;
        RECT 70.130 137.825 70.370 138.115 ;
        RECT 71.170 138.035 71.340 138.115 ;
        RECT 70.570 137.565 70.990 137.945 ;
        RECT 71.170 137.785 71.800 138.035 ;
        RECT 72.270 137.565 72.600 137.945 ;
        RECT 72.770 137.825 72.940 138.115 ;
        RECT 73.740 137.950 73.910 138.795 ;
        RECT 74.360 138.625 74.580 139.495 ;
        RECT 74.805 139.375 75.500 139.565 ;
        RECT 74.080 138.245 74.580 138.625 ;
        RECT 74.750 138.575 75.160 139.195 ;
        RECT 75.330 138.405 75.500 139.375 ;
        RECT 74.805 138.235 75.500 138.405 ;
        RECT 73.120 137.565 73.500 137.945 ;
        RECT 73.740 137.780 74.570 137.950 ;
        RECT 74.805 137.735 74.975 138.235 ;
        RECT 75.145 137.565 75.475 138.065 ;
        RECT 75.690 137.735 75.915 139.855 ;
        RECT 76.085 139.735 76.415 140.115 ;
        RECT 76.585 139.565 76.755 139.855 ;
        RECT 76.090 139.395 76.755 139.565 ;
        RECT 76.090 138.405 76.320 139.395 ;
        RECT 77.475 139.345 79.145 140.115 ;
        RECT 76.490 138.575 76.840 139.225 ;
        RECT 77.475 138.655 78.225 139.175 ;
        RECT 78.395 138.825 79.145 139.345 ;
        RECT 79.315 139.315 79.655 139.945 ;
        RECT 79.825 139.315 80.075 140.115 ;
        RECT 80.265 139.465 80.595 139.945 ;
        RECT 80.765 139.655 80.990 140.115 ;
        RECT 81.160 139.465 81.490 139.945 ;
        RECT 79.315 138.705 79.490 139.315 ;
        RECT 80.265 139.295 81.490 139.465 ;
        RECT 82.120 139.335 82.620 139.945 ;
        RECT 82.995 139.365 84.205 140.115 ;
        RECT 79.660 138.955 80.355 139.125 ;
        RECT 80.185 138.705 80.355 138.955 ;
        RECT 80.530 138.925 80.950 139.125 ;
        RECT 81.120 138.925 81.450 139.125 ;
        RECT 81.620 138.925 81.950 139.125 ;
        RECT 82.120 138.705 82.290 139.335 ;
        RECT 82.475 138.875 82.825 139.125 ;
        RECT 76.090 138.235 76.755 138.405 ;
        RECT 76.085 137.565 76.415 138.065 ;
        RECT 76.585 137.735 76.755 138.235 ;
        RECT 77.475 137.565 79.145 138.655 ;
        RECT 79.315 137.735 79.655 138.705 ;
        RECT 79.825 137.565 79.995 138.705 ;
        RECT 80.185 138.535 82.620 138.705 ;
        RECT 80.265 137.565 80.515 138.365 ;
        RECT 81.160 137.735 81.490 138.535 ;
        RECT 81.790 137.565 82.120 138.365 ;
        RECT 82.290 137.735 82.620 138.535 ;
        RECT 82.995 138.655 83.515 139.195 ;
        RECT 83.685 138.825 84.205 139.365 ;
        RECT 84.650 139.305 84.895 139.910 ;
        RECT 85.115 139.580 85.625 140.115 ;
        RECT 84.375 139.135 85.605 139.305 ;
        RECT 82.995 137.565 84.205 138.655 ;
        RECT 84.375 138.325 84.715 139.135 ;
        RECT 84.885 138.570 85.635 138.760 ;
        RECT 84.375 137.915 84.890 138.325 ;
        RECT 85.125 137.565 85.295 138.325 ;
        RECT 85.465 137.905 85.635 138.570 ;
        RECT 85.805 138.585 85.995 139.945 ;
        RECT 86.165 139.095 86.440 139.945 ;
        RECT 86.630 139.580 87.160 139.945 ;
        RECT 87.585 139.715 87.915 140.115 ;
        RECT 86.985 139.545 87.160 139.580 ;
        RECT 86.165 138.925 86.445 139.095 ;
        RECT 86.165 138.785 86.440 138.925 ;
        RECT 86.645 138.585 86.815 139.385 ;
        RECT 85.805 138.415 86.815 138.585 ;
        RECT 86.985 139.375 87.915 139.545 ;
        RECT 88.085 139.375 88.340 139.945 ;
        RECT 88.515 139.390 88.805 140.115 ;
        RECT 89.065 139.565 89.235 139.945 ;
        RECT 89.415 139.735 89.745 140.115 ;
        RECT 89.065 139.395 89.730 139.565 ;
        RECT 89.925 139.440 90.185 139.945 ;
        RECT 86.985 138.245 87.155 139.375 ;
        RECT 87.745 139.205 87.915 139.375 ;
        RECT 86.030 138.075 87.155 138.245 ;
        RECT 87.325 138.875 87.520 139.205 ;
        RECT 87.745 138.875 88.000 139.205 ;
        RECT 87.325 137.905 87.495 138.875 ;
        RECT 88.170 138.705 88.340 139.375 ;
        RECT 88.995 138.845 89.325 139.215 ;
        RECT 89.560 139.140 89.730 139.395 ;
        RECT 89.560 138.810 89.845 139.140 ;
        RECT 85.465 137.735 87.495 137.905 ;
        RECT 87.665 137.565 87.835 138.705 ;
        RECT 88.005 137.735 88.340 138.705 ;
        RECT 88.515 137.565 88.805 138.730 ;
        RECT 89.560 138.665 89.730 138.810 ;
        RECT 89.065 138.495 89.730 138.665 ;
        RECT 90.015 138.640 90.185 139.440 ;
        RECT 90.355 139.345 92.025 140.115 ;
        RECT 92.200 139.570 97.545 140.115 ;
        RECT 89.065 137.735 89.235 138.495 ;
        RECT 89.415 137.565 89.745 138.325 ;
        RECT 89.915 137.735 90.185 138.640 ;
        RECT 90.355 138.655 91.105 139.175 ;
        RECT 91.275 138.825 92.025 139.345 ;
        RECT 90.355 137.565 92.025 138.655 ;
        RECT 93.790 138.000 94.140 139.250 ;
        RECT 95.620 138.740 95.960 139.570 ;
        RECT 98.090 139.405 98.345 139.935 ;
        RECT 98.525 139.655 98.810 140.115 ;
        RECT 98.090 138.755 98.270 139.405 ;
        RECT 98.990 139.205 99.240 139.855 ;
        RECT 98.440 138.875 99.240 139.205 ;
        RECT 98.005 138.585 98.270 138.755 ;
        RECT 98.090 138.545 98.270 138.585 ;
        RECT 92.200 137.565 97.545 138.000 ;
        RECT 98.090 137.875 98.345 138.545 ;
        RECT 98.525 137.565 98.810 138.365 ;
        RECT 98.990 138.285 99.240 138.875 ;
        RECT 99.440 139.520 99.760 139.850 ;
        RECT 99.940 139.635 100.600 140.115 ;
        RECT 100.800 139.725 101.650 139.895 ;
        RECT 99.440 138.625 99.630 139.520 ;
        RECT 99.950 139.195 100.610 139.465 ;
        RECT 100.280 139.135 100.610 139.195 ;
        RECT 99.800 138.965 100.130 139.025 ;
        RECT 100.800 138.965 100.970 139.725 ;
        RECT 102.210 139.655 102.530 140.115 ;
        RECT 102.730 139.475 102.980 139.905 ;
        RECT 103.270 139.675 103.680 140.115 ;
        RECT 103.850 139.735 104.865 139.935 ;
        RECT 101.140 139.305 102.390 139.475 ;
        RECT 101.140 139.185 101.470 139.305 ;
        RECT 99.800 138.795 101.700 138.965 ;
        RECT 99.440 138.455 101.360 138.625 ;
        RECT 99.440 138.435 99.760 138.455 ;
        RECT 98.990 137.775 99.320 138.285 ;
        RECT 99.590 137.825 99.760 138.435 ;
        RECT 101.530 138.285 101.700 138.795 ;
        RECT 101.870 138.725 102.050 139.135 ;
        RECT 102.220 138.545 102.390 139.305 ;
        RECT 99.930 137.565 100.260 138.255 ;
        RECT 100.490 138.115 101.700 138.285 ;
        RECT 101.870 138.235 102.390 138.545 ;
        RECT 102.560 139.135 102.980 139.475 ;
        RECT 103.270 139.135 103.680 139.465 ;
        RECT 102.560 138.365 102.750 139.135 ;
        RECT 103.850 139.005 104.020 139.735 ;
        RECT 105.165 139.565 105.335 139.895 ;
        RECT 105.505 139.735 105.835 140.115 ;
        RECT 104.190 139.185 104.540 139.555 ;
        RECT 103.850 138.965 104.270 139.005 ;
        RECT 102.920 138.795 104.270 138.965 ;
        RECT 102.920 138.635 103.170 138.795 ;
        RECT 103.680 138.365 103.930 138.625 ;
        RECT 102.560 138.115 103.930 138.365 ;
        RECT 100.490 137.825 100.730 138.115 ;
        RECT 101.530 138.035 101.700 138.115 ;
        RECT 100.930 137.565 101.350 137.945 ;
        RECT 101.530 137.785 102.160 138.035 ;
        RECT 102.630 137.565 102.960 137.945 ;
        RECT 103.130 137.825 103.300 138.115 ;
        RECT 104.100 137.950 104.270 138.795 ;
        RECT 104.720 138.625 104.940 139.495 ;
        RECT 105.165 139.375 105.860 139.565 ;
        RECT 104.440 138.245 104.940 138.625 ;
        RECT 105.110 138.575 105.520 139.195 ;
        RECT 105.690 138.405 105.860 139.375 ;
        RECT 105.165 138.235 105.860 138.405 ;
        RECT 103.480 137.565 103.860 137.945 ;
        RECT 104.100 137.780 104.930 137.950 ;
        RECT 105.165 137.735 105.335 138.235 ;
        RECT 105.505 137.565 105.835 138.065 ;
        RECT 106.050 137.735 106.275 139.855 ;
        RECT 106.445 139.735 106.775 140.115 ;
        RECT 106.945 139.565 107.115 139.855 ;
        RECT 106.450 139.395 107.115 139.565 ;
        RECT 106.450 138.405 106.680 139.395 ;
        RECT 107.835 139.345 109.505 140.115 ;
        RECT 106.850 138.575 107.200 139.225 ;
        RECT 107.835 138.655 108.585 139.175 ;
        RECT 108.755 138.825 109.505 139.345 ;
        RECT 109.880 139.335 110.380 139.945 ;
        RECT 109.675 138.875 110.025 139.125 ;
        RECT 110.210 138.705 110.380 139.335 ;
        RECT 111.010 139.465 111.340 139.945 ;
        RECT 111.510 139.655 111.735 140.115 ;
        RECT 111.905 139.465 112.235 139.945 ;
        RECT 111.010 139.295 112.235 139.465 ;
        RECT 112.425 139.315 112.675 140.115 ;
        RECT 112.845 139.315 113.185 139.945 ;
        RECT 114.275 139.390 114.565 140.115 ;
        RECT 112.955 139.265 113.185 139.315 ;
        RECT 115.235 139.295 115.465 140.115 ;
        RECT 115.635 139.315 115.965 139.945 ;
        RECT 110.550 138.925 110.880 139.125 ;
        RECT 111.050 138.925 111.380 139.125 ;
        RECT 111.550 138.925 111.970 139.125 ;
        RECT 112.145 138.955 112.840 139.125 ;
        RECT 112.145 138.705 112.315 138.955 ;
        RECT 113.010 138.705 113.185 139.265 ;
        RECT 115.215 138.875 115.545 139.125 ;
        RECT 106.450 138.235 107.115 138.405 ;
        RECT 106.445 137.565 106.775 138.065 ;
        RECT 106.945 137.735 107.115 138.235 ;
        RECT 107.835 137.565 109.505 138.655 ;
        RECT 109.880 138.535 112.315 138.705 ;
        RECT 109.880 137.735 110.210 138.535 ;
        RECT 110.380 137.565 110.710 138.365 ;
        RECT 111.010 137.735 111.340 138.535 ;
        RECT 111.985 137.565 112.235 138.365 ;
        RECT 112.505 137.565 112.675 138.705 ;
        RECT 112.845 137.735 113.185 138.705 ;
        RECT 114.275 137.565 114.565 138.730 ;
        RECT 115.715 138.715 115.965 139.315 ;
        RECT 116.135 139.295 116.345 140.115 ;
        RECT 116.950 139.435 117.205 139.935 ;
        RECT 117.385 139.655 117.670 140.115 ;
        RECT 116.865 139.405 117.205 139.435 ;
        RECT 116.865 139.265 117.130 139.405 ;
        RECT 115.235 137.565 115.465 138.705 ;
        RECT 115.635 137.735 115.965 138.715 ;
        RECT 116.135 137.565 116.345 138.705 ;
        RECT 116.950 138.545 117.130 139.265 ;
        RECT 117.850 139.205 118.100 139.855 ;
        RECT 117.300 138.875 118.100 139.205 ;
        RECT 116.950 137.875 117.205 138.545 ;
        RECT 117.385 137.565 117.670 138.365 ;
        RECT 117.850 138.285 118.100 138.875 ;
        RECT 118.300 139.520 118.620 139.850 ;
        RECT 118.800 139.635 119.460 140.115 ;
        RECT 119.660 139.725 120.510 139.895 ;
        RECT 118.300 138.625 118.490 139.520 ;
        RECT 118.810 139.195 119.470 139.465 ;
        RECT 119.140 139.135 119.470 139.195 ;
        RECT 118.660 138.965 118.990 139.025 ;
        RECT 119.660 138.965 119.830 139.725 ;
        RECT 121.070 139.655 121.390 140.115 ;
        RECT 121.590 139.475 121.840 139.905 ;
        RECT 122.130 139.675 122.540 140.115 ;
        RECT 122.710 139.735 123.725 139.935 ;
        RECT 120.000 139.305 121.250 139.475 ;
        RECT 120.000 139.185 120.330 139.305 ;
        RECT 118.660 138.795 120.560 138.965 ;
        RECT 118.300 138.455 120.220 138.625 ;
        RECT 118.300 138.435 118.620 138.455 ;
        RECT 117.850 137.775 118.180 138.285 ;
        RECT 118.450 137.825 118.620 138.435 ;
        RECT 120.390 138.285 120.560 138.795 ;
        RECT 120.730 138.725 120.910 139.135 ;
        RECT 121.080 138.545 121.250 139.305 ;
        RECT 118.790 137.565 119.120 138.255 ;
        RECT 119.350 138.115 120.560 138.285 ;
        RECT 120.730 138.235 121.250 138.545 ;
        RECT 121.420 139.135 121.840 139.475 ;
        RECT 122.130 139.135 122.540 139.465 ;
        RECT 121.420 138.365 121.610 139.135 ;
        RECT 122.710 139.005 122.880 139.735 ;
        RECT 124.025 139.565 124.195 139.895 ;
        RECT 124.365 139.735 124.695 140.115 ;
        RECT 123.050 139.185 123.400 139.555 ;
        RECT 122.710 138.965 123.130 139.005 ;
        RECT 121.780 138.795 123.130 138.965 ;
        RECT 121.780 138.635 122.030 138.795 ;
        RECT 122.540 138.365 122.790 138.625 ;
        RECT 121.420 138.115 122.790 138.365 ;
        RECT 119.350 137.825 119.590 138.115 ;
        RECT 120.390 138.035 120.560 138.115 ;
        RECT 119.790 137.565 120.210 137.945 ;
        RECT 120.390 137.785 121.020 138.035 ;
        RECT 121.490 137.565 121.820 137.945 ;
        RECT 121.990 137.825 122.160 138.115 ;
        RECT 122.960 137.950 123.130 138.795 ;
        RECT 123.580 138.625 123.800 139.495 ;
        RECT 124.025 139.375 124.720 139.565 ;
        RECT 123.300 138.245 123.800 138.625 ;
        RECT 123.970 138.575 124.380 139.195 ;
        RECT 124.550 138.405 124.720 139.375 ;
        RECT 124.025 138.235 124.720 138.405 ;
        RECT 122.340 137.565 122.720 137.945 ;
        RECT 122.960 137.780 123.790 137.950 ;
        RECT 124.025 137.735 124.195 138.235 ;
        RECT 124.365 137.565 124.695 138.065 ;
        RECT 124.910 137.735 125.135 139.855 ;
        RECT 125.305 139.735 125.635 140.115 ;
        RECT 125.805 139.565 125.975 139.855 ;
        RECT 125.310 139.395 125.975 139.565 ;
        RECT 125.310 138.405 125.540 139.395 ;
        RECT 126.235 139.365 127.445 140.115 ;
        RECT 125.710 138.575 126.060 139.225 ;
        RECT 126.235 138.655 126.755 139.195 ;
        RECT 126.925 138.825 127.445 139.365 ;
        RECT 125.310 138.235 125.975 138.405 ;
        RECT 125.305 137.565 125.635 138.065 ;
        RECT 125.805 137.735 125.975 138.235 ;
        RECT 126.235 137.565 127.445 138.655 ;
        RECT 14.370 137.395 127.530 137.565 ;
        RECT 14.455 136.305 15.665 137.395 ;
        RECT 14.455 135.595 14.975 136.135 ;
        RECT 15.145 135.765 15.665 136.305 ;
        RECT 16.295 136.305 19.805 137.395 ;
        RECT 16.295 135.785 17.985 136.305 ;
        RECT 19.980 136.255 20.315 137.225 ;
        RECT 20.485 136.255 20.655 137.395 ;
        RECT 20.825 137.055 22.855 137.225 ;
        RECT 18.155 135.615 19.805 136.135 ;
        RECT 14.455 134.845 15.665 135.595 ;
        RECT 16.295 134.845 19.805 135.615 ;
        RECT 19.980 135.585 20.150 136.255 ;
        RECT 20.825 136.085 20.995 137.055 ;
        RECT 20.320 135.755 20.575 136.085 ;
        RECT 20.800 135.755 20.995 136.085 ;
        RECT 21.165 136.715 22.290 136.885 ;
        RECT 20.405 135.585 20.575 135.755 ;
        RECT 21.165 135.585 21.335 136.715 ;
        RECT 19.980 135.015 20.235 135.585 ;
        RECT 20.405 135.415 21.335 135.585 ;
        RECT 21.505 136.375 22.515 136.545 ;
        RECT 21.505 135.575 21.675 136.375 ;
        RECT 21.880 136.035 22.155 136.175 ;
        RECT 21.875 135.865 22.155 136.035 ;
        RECT 21.160 135.380 21.335 135.415 ;
        RECT 20.405 134.845 20.735 135.245 ;
        RECT 21.160 135.015 21.690 135.380 ;
        RECT 21.880 135.015 22.155 135.865 ;
        RECT 22.325 135.015 22.515 136.375 ;
        RECT 22.685 136.390 22.855 137.055 ;
        RECT 23.025 136.635 23.195 137.395 ;
        RECT 23.430 136.635 23.945 137.045 ;
        RECT 22.685 136.200 23.435 136.390 ;
        RECT 23.605 135.825 23.945 136.635 ;
        RECT 24.115 136.230 24.405 137.395 ;
        RECT 24.575 136.305 28.085 137.395 ;
        RECT 22.715 135.655 23.945 135.825 ;
        RECT 24.575 135.785 26.265 136.305 ;
        RECT 28.260 136.255 28.595 137.225 ;
        RECT 28.765 136.255 28.935 137.395 ;
        RECT 29.105 137.055 31.135 137.225 ;
        RECT 22.695 134.845 23.205 135.380 ;
        RECT 23.425 135.050 23.670 135.655 ;
        RECT 26.435 135.615 28.085 136.135 ;
        RECT 24.115 134.845 24.405 135.570 ;
        RECT 24.575 134.845 28.085 135.615 ;
        RECT 28.260 135.585 28.430 136.255 ;
        RECT 29.105 136.085 29.275 137.055 ;
        RECT 28.600 135.755 28.855 136.085 ;
        RECT 29.080 135.755 29.275 136.085 ;
        RECT 29.445 136.715 30.570 136.885 ;
        RECT 28.685 135.585 28.855 135.755 ;
        RECT 29.445 135.585 29.615 136.715 ;
        RECT 28.260 135.015 28.515 135.585 ;
        RECT 28.685 135.415 29.615 135.585 ;
        RECT 29.785 136.375 30.795 136.545 ;
        RECT 29.785 135.575 29.955 136.375 ;
        RECT 30.160 135.695 30.435 136.175 ;
        RECT 30.155 135.525 30.435 135.695 ;
        RECT 29.440 135.380 29.615 135.415 ;
        RECT 28.685 134.845 29.015 135.245 ;
        RECT 29.440 135.015 29.970 135.380 ;
        RECT 30.160 135.015 30.435 135.525 ;
        RECT 30.605 135.015 30.795 136.375 ;
        RECT 30.965 136.390 31.135 137.055 ;
        RECT 31.305 136.635 31.475 137.395 ;
        RECT 31.710 136.635 32.225 137.045 ;
        RECT 32.595 136.725 32.875 137.395 ;
        RECT 30.965 136.200 31.715 136.390 ;
        RECT 31.885 135.825 32.225 136.635 ;
        RECT 33.045 136.505 33.345 137.055 ;
        RECT 33.545 136.675 33.875 137.395 ;
        RECT 34.065 136.675 34.525 137.225 ;
        RECT 32.410 136.085 32.675 136.445 ;
        RECT 33.045 136.335 33.985 136.505 ;
        RECT 33.815 136.085 33.985 136.335 ;
        RECT 32.410 135.835 33.085 136.085 ;
        RECT 33.305 135.835 33.645 136.085 ;
        RECT 30.995 135.655 32.225 135.825 ;
        RECT 33.815 135.755 34.105 136.085 ;
        RECT 33.815 135.665 33.985 135.755 ;
        RECT 30.975 134.845 31.485 135.380 ;
        RECT 31.705 135.050 31.950 135.655 ;
        RECT 32.595 135.475 33.985 135.665 ;
        RECT 32.595 135.115 32.925 135.475 ;
        RECT 34.275 135.305 34.525 136.675 ;
        RECT 33.545 134.845 33.795 135.305 ;
        RECT 33.965 135.015 34.525 135.305 ;
        RECT 34.695 136.255 34.965 137.225 ;
        RECT 35.175 136.595 35.455 137.395 ;
        RECT 35.625 136.885 37.280 137.175 ;
        RECT 35.690 136.545 37.280 136.715 ;
        RECT 35.690 136.425 35.860 136.545 ;
        RECT 35.135 136.255 35.860 136.425 ;
        RECT 34.695 135.520 34.865 136.255 ;
        RECT 35.135 136.085 35.305 136.255 ;
        RECT 35.035 135.755 35.305 136.085 ;
        RECT 35.475 135.755 35.880 136.085 ;
        RECT 36.050 135.755 36.760 136.375 ;
        RECT 36.960 136.255 37.280 136.545 ;
        RECT 37.455 136.255 37.725 137.225 ;
        RECT 37.935 136.595 38.215 137.395 ;
        RECT 38.385 136.885 40.040 137.175 ;
        RECT 38.450 136.545 40.040 136.715 ;
        RECT 38.450 136.425 38.620 136.545 ;
        RECT 37.895 136.255 38.620 136.425 ;
        RECT 35.135 135.585 35.305 135.755 ;
        RECT 34.695 135.175 34.965 135.520 ;
        RECT 35.135 135.415 36.745 135.585 ;
        RECT 36.930 135.515 37.280 136.085 ;
        RECT 37.455 135.520 37.625 136.255 ;
        RECT 37.895 136.085 38.065 136.255 ;
        RECT 37.795 135.755 38.065 136.085 ;
        RECT 38.235 135.755 38.640 136.085 ;
        RECT 38.810 135.755 39.520 136.375 ;
        RECT 39.720 136.255 40.040 136.545 ;
        RECT 40.675 136.305 43.265 137.395 ;
        RECT 37.895 135.585 38.065 135.755 ;
        RECT 35.155 134.845 35.535 135.245 ;
        RECT 35.705 135.065 35.875 135.415 ;
        RECT 36.045 134.845 36.375 135.245 ;
        RECT 36.575 135.065 36.745 135.415 ;
        RECT 36.945 134.845 37.275 135.345 ;
        RECT 37.455 135.175 37.725 135.520 ;
        RECT 37.895 135.415 39.505 135.585 ;
        RECT 39.690 135.515 40.040 136.085 ;
        RECT 40.675 135.785 41.885 136.305 ;
        RECT 43.435 136.255 43.705 137.225 ;
        RECT 43.915 136.595 44.195 137.395 ;
        RECT 44.365 136.885 46.020 137.175 ;
        RECT 44.430 136.545 46.020 136.715 ;
        RECT 44.430 136.425 44.600 136.545 ;
        RECT 43.875 136.255 44.600 136.425 ;
        RECT 42.055 135.615 43.265 136.135 ;
        RECT 37.915 134.845 38.295 135.245 ;
        RECT 38.465 135.065 38.635 135.415 ;
        RECT 38.805 134.845 39.135 135.245 ;
        RECT 39.335 135.065 39.505 135.415 ;
        RECT 39.705 134.845 40.035 135.345 ;
        RECT 40.675 134.845 43.265 135.615 ;
        RECT 43.435 135.520 43.605 136.255 ;
        RECT 43.875 136.085 44.045 136.255 ;
        RECT 44.790 136.205 45.505 136.375 ;
        RECT 45.700 136.255 46.020 136.545 ;
        RECT 46.195 136.255 46.535 137.225 ;
        RECT 46.705 136.255 46.875 137.395 ;
        RECT 47.145 136.595 47.395 137.395 ;
        RECT 48.040 136.425 48.370 137.225 ;
        RECT 48.670 136.595 49.000 137.395 ;
        RECT 49.170 136.425 49.500 137.225 ;
        RECT 47.065 136.255 49.500 136.425 ;
        RECT 43.775 135.755 44.045 136.085 ;
        RECT 44.215 135.755 44.620 136.085 ;
        RECT 44.790 135.755 45.500 136.205 ;
        RECT 43.875 135.585 44.045 135.755 ;
        RECT 43.435 135.175 43.705 135.520 ;
        RECT 43.875 135.415 45.485 135.585 ;
        RECT 45.670 135.515 46.020 136.085 ;
        RECT 46.195 135.695 46.370 136.255 ;
        RECT 47.065 136.005 47.235 136.255 ;
        RECT 46.540 135.835 47.235 136.005 ;
        RECT 47.410 135.835 47.830 136.035 ;
        RECT 48.000 135.835 48.330 136.035 ;
        RECT 48.500 135.835 48.830 136.035 ;
        RECT 46.195 135.645 46.425 135.695 ;
        RECT 43.895 134.845 44.275 135.245 ;
        RECT 44.445 135.065 44.615 135.415 ;
        RECT 44.785 134.845 45.115 135.245 ;
        RECT 45.315 135.065 45.485 135.415 ;
        RECT 45.685 134.845 46.015 135.345 ;
        RECT 46.195 135.015 46.535 135.645 ;
        RECT 46.705 134.845 46.955 135.645 ;
        RECT 47.145 135.495 48.370 135.665 ;
        RECT 47.145 135.015 47.475 135.495 ;
        RECT 47.645 134.845 47.870 135.305 ;
        RECT 48.040 135.015 48.370 135.495 ;
        RECT 49.000 135.625 49.170 136.255 ;
        RECT 49.875 136.230 50.165 137.395 ;
        RECT 50.335 136.305 52.925 137.395 ;
        RECT 53.095 136.635 53.610 137.045 ;
        RECT 53.845 136.635 54.015 137.395 ;
        RECT 54.185 137.055 56.215 137.225 ;
        RECT 49.355 135.835 49.705 136.085 ;
        RECT 50.335 135.785 51.545 136.305 ;
        RECT 49.000 135.015 49.500 135.625 ;
        RECT 51.715 135.615 52.925 136.135 ;
        RECT 53.095 135.825 53.435 136.635 ;
        RECT 54.185 136.390 54.355 137.055 ;
        RECT 54.750 136.715 55.875 136.885 ;
        RECT 53.605 136.200 54.355 136.390 ;
        RECT 54.525 136.375 55.535 136.545 ;
        RECT 53.095 135.655 54.325 135.825 ;
        RECT 49.875 134.845 50.165 135.570 ;
        RECT 50.335 134.845 52.925 135.615 ;
        RECT 53.370 135.050 53.615 135.655 ;
        RECT 53.835 134.845 54.345 135.380 ;
        RECT 54.525 135.015 54.715 136.375 ;
        RECT 54.885 136.035 55.160 136.175 ;
        RECT 54.885 135.865 55.165 136.035 ;
        RECT 54.885 135.015 55.160 135.865 ;
        RECT 55.365 135.575 55.535 136.375 ;
        RECT 55.705 135.585 55.875 136.715 ;
        RECT 56.045 136.085 56.215 137.055 ;
        RECT 56.385 136.255 56.555 137.395 ;
        RECT 56.725 136.255 57.060 137.225 ;
        RECT 57.785 136.465 57.955 137.225 ;
        RECT 58.135 136.635 58.465 137.395 ;
        RECT 57.785 136.295 58.450 136.465 ;
        RECT 58.635 136.320 58.905 137.225 ;
        RECT 56.045 135.755 56.240 136.085 ;
        RECT 56.465 135.755 56.720 136.085 ;
        RECT 56.465 135.585 56.635 135.755 ;
        RECT 56.890 135.585 57.060 136.255 ;
        RECT 58.280 136.150 58.450 136.295 ;
        RECT 57.715 135.745 58.045 136.115 ;
        RECT 58.280 135.820 58.565 136.150 ;
        RECT 55.705 135.415 56.635 135.585 ;
        RECT 55.705 135.380 55.880 135.415 ;
        RECT 55.350 135.015 55.880 135.380 ;
        RECT 56.305 134.845 56.635 135.245 ;
        RECT 56.805 135.015 57.060 135.585 ;
        RECT 58.280 135.565 58.450 135.820 ;
        RECT 57.785 135.395 58.450 135.565 ;
        RECT 58.735 135.520 58.905 136.320 ;
        RECT 59.075 136.305 60.745 137.395 ;
        RECT 59.075 135.785 59.825 136.305 ;
        RECT 60.915 136.255 61.255 137.225 ;
        RECT 61.425 136.255 61.595 137.395 ;
        RECT 61.865 136.595 62.115 137.395 ;
        RECT 62.760 136.425 63.090 137.225 ;
        RECT 63.390 136.595 63.720 137.395 ;
        RECT 63.890 136.425 64.220 137.225 ;
        RECT 64.710 136.765 64.995 137.225 ;
        RECT 65.165 136.935 65.435 137.395 ;
        RECT 64.710 136.545 65.665 136.765 ;
        RECT 61.785 136.255 64.220 136.425 ;
        RECT 59.995 135.615 60.745 136.135 ;
        RECT 57.785 135.015 57.955 135.395 ;
        RECT 58.135 134.845 58.465 135.225 ;
        RECT 58.645 135.015 58.905 135.520 ;
        RECT 59.075 134.845 60.745 135.615 ;
        RECT 60.915 135.645 61.090 136.255 ;
        RECT 61.785 136.005 61.955 136.255 ;
        RECT 61.260 135.835 61.955 136.005 ;
        RECT 62.130 135.835 62.550 136.035 ;
        RECT 62.720 135.835 63.050 136.035 ;
        RECT 63.220 135.835 63.550 136.035 ;
        RECT 60.915 135.015 61.255 135.645 ;
        RECT 61.425 134.845 61.675 135.645 ;
        RECT 61.865 135.495 63.090 135.665 ;
        RECT 61.865 135.015 62.195 135.495 ;
        RECT 62.365 134.845 62.590 135.305 ;
        RECT 62.760 135.015 63.090 135.495 ;
        RECT 63.720 135.625 63.890 136.255 ;
        RECT 64.075 135.835 64.425 136.085 ;
        RECT 64.595 135.815 65.285 136.375 ;
        RECT 65.455 135.645 65.665 136.545 ;
        RECT 63.720 135.015 64.220 135.625 ;
        RECT 64.710 135.475 65.665 135.645 ;
        RECT 65.835 136.375 66.235 137.225 ;
        RECT 66.425 136.765 66.705 137.225 ;
        RECT 67.225 136.935 67.550 137.395 ;
        RECT 66.425 136.545 67.550 136.765 ;
        RECT 65.835 135.815 66.930 136.375 ;
        RECT 67.100 136.085 67.550 136.545 ;
        RECT 67.720 136.255 68.105 137.225 ;
        RECT 64.710 135.015 64.995 135.475 ;
        RECT 65.165 134.845 65.435 135.305 ;
        RECT 65.835 135.015 66.235 135.815 ;
        RECT 67.100 135.755 67.655 136.085 ;
        RECT 67.100 135.645 67.550 135.755 ;
        RECT 66.425 135.475 67.550 135.645 ;
        RECT 67.825 135.585 68.105 136.255 ;
        RECT 68.280 137.005 68.615 137.225 ;
        RECT 69.620 137.015 69.975 137.395 ;
        RECT 68.280 136.385 68.535 137.005 ;
        RECT 68.785 136.845 69.015 136.885 ;
        RECT 70.145 136.845 70.395 137.225 ;
        RECT 68.785 136.645 70.395 136.845 ;
        RECT 68.785 136.555 68.970 136.645 ;
        RECT 69.560 136.635 70.395 136.645 ;
        RECT 70.645 136.615 70.895 137.395 ;
        RECT 71.065 136.545 71.325 137.225 ;
        RECT 69.125 136.445 69.455 136.475 ;
        RECT 69.125 136.385 70.925 136.445 ;
        RECT 68.280 136.275 70.985 136.385 ;
        RECT 68.280 136.215 69.455 136.275 ;
        RECT 70.785 136.240 70.985 136.275 ;
        RECT 68.275 135.835 68.765 136.035 ;
        RECT 68.955 135.835 69.430 136.045 ;
        RECT 66.425 135.015 66.705 135.475 ;
        RECT 67.225 134.845 67.550 135.305 ;
        RECT 67.720 135.015 68.105 135.585 ;
        RECT 68.280 134.845 68.735 135.610 ;
        RECT 69.210 135.435 69.430 135.835 ;
        RECT 69.675 135.835 70.005 136.045 ;
        RECT 69.675 135.435 69.885 135.835 ;
        RECT 70.175 135.800 70.585 136.105 ;
        RECT 70.815 135.665 70.985 136.240 ;
        RECT 70.715 135.545 70.985 135.665 ;
        RECT 70.140 135.500 70.985 135.545 ;
        RECT 70.140 135.375 70.895 135.500 ;
        RECT 70.140 135.225 70.310 135.375 ;
        RECT 71.155 135.345 71.325 136.545 ;
        RECT 71.955 136.305 75.465 137.395 ;
        RECT 71.955 135.785 73.645 136.305 ;
        RECT 75.635 136.230 75.925 137.395 ;
        RECT 77.015 136.255 77.285 137.225 ;
        RECT 77.495 136.595 77.775 137.395 ;
        RECT 77.945 136.885 79.600 137.175 ;
        RECT 78.010 136.545 79.600 136.715 ;
        RECT 78.010 136.425 78.180 136.545 ;
        RECT 77.455 136.255 78.180 136.425 ;
        RECT 73.815 135.615 75.465 136.135 ;
        RECT 69.010 135.015 70.310 135.225 ;
        RECT 70.565 134.845 70.895 135.205 ;
        RECT 71.065 135.015 71.325 135.345 ;
        RECT 71.955 134.845 75.465 135.615 ;
        RECT 75.635 134.845 75.925 135.570 ;
        RECT 77.015 135.520 77.185 136.255 ;
        RECT 77.455 136.085 77.625 136.255 ;
        RECT 77.355 135.755 77.625 136.085 ;
        RECT 77.795 135.755 78.200 136.085 ;
        RECT 78.370 135.755 79.080 136.375 ;
        RECT 79.280 136.255 79.600 136.545 ;
        RECT 79.775 136.255 80.115 137.225 ;
        RECT 80.285 136.255 80.455 137.395 ;
        RECT 80.725 136.595 80.975 137.395 ;
        RECT 81.620 136.425 81.950 137.225 ;
        RECT 82.250 136.595 82.580 137.395 ;
        RECT 82.750 136.425 83.080 137.225 ;
        RECT 83.830 137.055 84.085 137.085 ;
        RECT 83.745 136.885 84.085 137.055 ;
        RECT 80.645 136.255 83.080 136.425 ;
        RECT 83.830 136.415 84.085 136.885 ;
        RECT 84.265 136.595 84.550 137.395 ;
        RECT 84.730 136.675 85.060 137.185 ;
        RECT 77.455 135.585 77.625 135.755 ;
        RECT 77.015 135.175 77.285 135.520 ;
        RECT 77.455 135.415 79.065 135.585 ;
        RECT 79.250 135.515 79.600 136.085 ;
        RECT 79.775 135.645 79.950 136.255 ;
        RECT 80.645 136.005 80.815 136.255 ;
        RECT 80.120 135.835 80.815 136.005 ;
        RECT 80.990 135.835 81.410 136.035 ;
        RECT 81.580 135.835 81.910 136.035 ;
        RECT 82.080 135.835 82.410 136.035 ;
        RECT 77.475 134.845 77.855 135.245 ;
        RECT 78.025 135.065 78.195 135.415 ;
        RECT 78.365 134.845 78.695 135.245 ;
        RECT 78.895 135.065 79.065 135.415 ;
        RECT 79.265 134.845 79.595 135.345 ;
        RECT 79.775 135.015 80.115 135.645 ;
        RECT 80.285 134.845 80.535 135.645 ;
        RECT 80.725 135.495 81.950 135.665 ;
        RECT 80.725 135.015 81.055 135.495 ;
        RECT 81.225 134.845 81.450 135.305 ;
        RECT 81.620 135.015 81.950 135.495 ;
        RECT 82.580 135.625 82.750 136.255 ;
        RECT 82.935 135.835 83.285 136.085 ;
        RECT 82.580 135.015 83.080 135.625 ;
        RECT 83.830 135.555 84.010 136.415 ;
        RECT 84.730 136.085 84.980 136.675 ;
        RECT 85.330 136.525 85.500 137.135 ;
        RECT 85.670 136.705 86.000 137.395 ;
        RECT 86.230 136.845 86.470 137.135 ;
        RECT 86.670 137.015 87.090 137.395 ;
        RECT 87.270 136.925 87.900 137.175 ;
        RECT 88.370 137.015 88.700 137.395 ;
        RECT 87.270 136.845 87.440 136.925 ;
        RECT 88.870 136.845 89.040 137.135 ;
        RECT 89.220 137.015 89.600 137.395 ;
        RECT 89.840 137.010 90.670 137.180 ;
        RECT 86.230 136.675 87.440 136.845 ;
        RECT 84.180 135.755 84.980 136.085 ;
        RECT 83.830 135.025 84.085 135.555 ;
        RECT 84.265 134.845 84.550 135.305 ;
        RECT 84.730 135.105 84.980 135.755 ;
        RECT 85.180 136.505 85.500 136.525 ;
        RECT 85.180 136.335 87.100 136.505 ;
        RECT 85.180 135.440 85.370 136.335 ;
        RECT 87.270 136.165 87.440 136.675 ;
        RECT 87.610 136.415 88.130 136.725 ;
        RECT 85.540 135.995 87.440 136.165 ;
        RECT 85.540 135.935 85.870 135.995 ;
        RECT 86.020 135.765 86.350 135.825 ;
        RECT 85.690 135.495 86.350 135.765 ;
        RECT 85.180 135.110 85.500 135.440 ;
        RECT 85.680 134.845 86.340 135.325 ;
        RECT 86.540 135.235 86.710 135.995 ;
        RECT 87.610 135.825 87.790 136.235 ;
        RECT 86.880 135.655 87.210 135.775 ;
        RECT 87.960 135.655 88.130 136.415 ;
        RECT 86.880 135.485 88.130 135.655 ;
        RECT 88.300 136.595 89.670 136.845 ;
        RECT 88.300 135.825 88.490 136.595 ;
        RECT 89.420 136.335 89.670 136.595 ;
        RECT 88.660 136.165 88.910 136.325 ;
        RECT 89.840 136.165 90.010 137.010 ;
        RECT 90.905 136.725 91.075 137.225 ;
        RECT 91.245 136.895 91.575 137.395 ;
        RECT 90.180 136.335 90.680 136.715 ;
        RECT 90.905 136.555 91.600 136.725 ;
        RECT 88.660 135.995 90.010 136.165 ;
        RECT 89.590 135.955 90.010 135.995 ;
        RECT 88.300 135.485 88.720 135.825 ;
        RECT 89.010 135.495 89.420 135.825 ;
        RECT 86.540 135.065 87.390 135.235 ;
        RECT 87.950 134.845 88.270 135.305 ;
        RECT 88.470 135.055 88.720 135.485 ;
        RECT 89.010 134.845 89.420 135.285 ;
        RECT 89.590 135.225 89.760 135.955 ;
        RECT 89.930 135.405 90.280 135.775 ;
        RECT 90.460 135.465 90.680 136.335 ;
        RECT 90.850 135.765 91.260 136.385 ;
        RECT 91.430 135.585 91.600 136.555 ;
        RECT 90.905 135.395 91.600 135.585 ;
        RECT 89.590 135.025 90.605 135.225 ;
        RECT 90.905 135.065 91.075 135.395 ;
        RECT 91.245 134.845 91.575 135.225 ;
        RECT 91.790 135.105 92.015 137.225 ;
        RECT 92.185 136.895 92.515 137.395 ;
        RECT 92.685 136.725 92.855 137.225 ;
        RECT 92.190 136.555 92.855 136.725 ;
        RECT 92.190 135.565 92.420 136.555 ;
        RECT 92.590 135.735 92.940 136.385 ;
        RECT 93.120 136.255 93.455 137.225 ;
        RECT 93.625 136.255 93.795 137.395 ;
        RECT 93.965 137.055 95.995 137.225 ;
        RECT 93.120 135.585 93.290 136.255 ;
        RECT 93.965 136.085 94.135 137.055 ;
        RECT 93.460 135.755 93.715 136.085 ;
        RECT 93.940 135.755 94.135 136.085 ;
        RECT 94.305 136.715 95.430 136.885 ;
        RECT 93.545 135.585 93.715 135.755 ;
        RECT 94.305 135.585 94.475 136.715 ;
        RECT 92.190 135.395 92.855 135.565 ;
        RECT 92.185 134.845 92.515 135.225 ;
        RECT 92.685 135.105 92.855 135.395 ;
        RECT 93.120 135.015 93.375 135.585 ;
        RECT 93.545 135.415 94.475 135.585 ;
        RECT 94.645 136.375 95.655 136.545 ;
        RECT 94.645 135.575 94.815 136.375 ;
        RECT 94.300 135.380 94.475 135.415 ;
        RECT 93.545 134.845 93.875 135.245 ;
        RECT 94.300 135.015 94.830 135.380 ;
        RECT 95.020 135.355 95.295 136.175 ;
        RECT 95.015 135.185 95.295 135.355 ;
        RECT 95.020 135.015 95.295 135.185 ;
        RECT 95.465 135.015 95.655 136.375 ;
        RECT 95.825 136.390 95.995 137.055 ;
        RECT 96.165 136.635 96.335 137.395 ;
        RECT 96.570 136.635 97.085 137.045 ;
        RECT 95.825 136.200 96.575 136.390 ;
        RECT 96.745 135.825 97.085 136.635 ;
        RECT 97.920 136.425 98.250 137.225 ;
        RECT 98.420 136.595 98.750 137.395 ;
        RECT 99.050 136.425 99.380 137.225 ;
        RECT 100.025 136.595 100.275 137.395 ;
        RECT 97.920 136.255 100.355 136.425 ;
        RECT 100.545 136.255 100.715 137.395 ;
        RECT 100.885 136.255 101.225 137.225 ;
        RECT 97.715 135.835 98.065 136.085 ;
        RECT 95.855 135.655 97.085 135.825 ;
        RECT 95.835 134.845 96.345 135.380 ;
        RECT 96.565 135.050 96.810 135.655 ;
        RECT 98.250 135.625 98.420 136.255 ;
        RECT 98.590 135.835 98.920 136.035 ;
        RECT 99.090 135.835 99.420 136.035 ;
        RECT 99.590 135.835 100.010 136.035 ;
        RECT 100.185 136.005 100.355 136.255 ;
        RECT 100.185 135.835 100.880 136.005 ;
        RECT 97.920 135.015 98.420 135.625 ;
        RECT 99.050 135.495 100.275 135.665 ;
        RECT 101.050 135.645 101.225 136.255 ;
        RECT 101.395 136.230 101.685 137.395 ;
        RECT 102.775 136.635 103.290 137.045 ;
        RECT 103.525 136.635 103.695 137.395 ;
        RECT 103.865 137.055 105.895 137.225 ;
        RECT 102.775 135.825 103.115 136.635 ;
        RECT 103.865 136.390 104.035 137.055 ;
        RECT 104.430 136.715 105.555 136.885 ;
        RECT 103.285 136.200 104.035 136.390 ;
        RECT 104.205 136.375 105.215 136.545 ;
        RECT 102.775 135.655 104.005 135.825 ;
        RECT 99.050 135.015 99.380 135.495 ;
        RECT 99.550 134.845 99.775 135.305 ;
        RECT 99.945 135.015 100.275 135.495 ;
        RECT 100.465 134.845 100.715 135.645 ;
        RECT 100.885 135.015 101.225 135.645 ;
        RECT 101.395 134.845 101.685 135.570 ;
        RECT 103.050 135.050 103.295 135.655 ;
        RECT 103.515 134.845 104.025 135.380 ;
        RECT 104.205 135.015 104.395 136.375 ;
        RECT 104.565 136.035 104.840 136.175 ;
        RECT 104.565 135.865 104.845 136.035 ;
        RECT 104.565 135.015 104.840 135.865 ;
        RECT 105.045 135.575 105.215 136.375 ;
        RECT 105.385 135.585 105.555 136.715 ;
        RECT 105.725 136.085 105.895 137.055 ;
        RECT 106.065 136.255 106.235 137.395 ;
        RECT 106.405 136.255 106.740 137.225 ;
        RECT 105.725 135.755 105.920 136.085 ;
        RECT 106.145 135.755 106.400 136.085 ;
        RECT 106.145 135.585 106.315 135.755 ;
        RECT 106.570 135.585 106.740 136.255 ;
        RECT 105.385 135.415 106.315 135.585 ;
        RECT 105.385 135.380 105.560 135.415 ;
        RECT 105.030 135.015 105.560 135.380 ;
        RECT 105.985 134.845 106.315 135.245 ;
        RECT 106.485 135.015 106.740 135.585 ;
        RECT 106.915 136.320 107.185 137.225 ;
        RECT 107.355 136.635 107.685 137.395 ;
        RECT 107.865 136.465 108.035 137.225 ;
        RECT 106.915 135.520 107.085 136.320 ;
        RECT 107.370 136.295 108.035 136.465 ;
        RECT 109.215 136.635 109.730 137.045 ;
        RECT 109.965 136.635 110.135 137.395 ;
        RECT 110.305 137.055 112.335 137.225 ;
        RECT 107.370 136.150 107.540 136.295 ;
        RECT 107.255 135.820 107.540 136.150 ;
        RECT 107.370 135.565 107.540 135.820 ;
        RECT 107.775 135.745 108.105 136.115 ;
        RECT 109.215 135.825 109.555 136.635 ;
        RECT 110.305 136.390 110.475 137.055 ;
        RECT 110.870 136.715 111.995 136.885 ;
        RECT 109.725 136.200 110.475 136.390 ;
        RECT 110.645 136.375 111.655 136.545 ;
        RECT 109.215 135.655 110.445 135.825 ;
        RECT 106.915 135.015 107.175 135.520 ;
        RECT 107.370 135.395 108.035 135.565 ;
        RECT 107.355 134.845 107.685 135.225 ;
        RECT 107.865 135.015 108.035 135.395 ;
        RECT 109.490 135.050 109.735 135.655 ;
        RECT 109.955 134.845 110.465 135.380 ;
        RECT 110.645 135.015 110.835 136.375 ;
        RECT 111.005 136.035 111.280 136.175 ;
        RECT 111.005 135.865 111.285 136.035 ;
        RECT 111.005 135.015 111.280 135.865 ;
        RECT 111.485 135.575 111.655 136.375 ;
        RECT 111.825 135.585 111.995 136.715 ;
        RECT 112.165 136.085 112.335 137.055 ;
        RECT 112.505 136.255 112.675 137.395 ;
        RECT 112.845 136.255 113.180 137.225 ;
        RECT 112.165 135.755 112.360 136.085 ;
        RECT 112.585 135.755 112.840 136.085 ;
        RECT 112.585 135.585 112.755 135.755 ;
        RECT 113.010 135.585 113.180 136.255 ;
        RECT 113.730 136.415 113.985 137.085 ;
        RECT 114.165 136.595 114.450 137.395 ;
        RECT 114.630 136.675 114.960 137.185 ;
        RECT 113.730 135.695 113.910 136.415 ;
        RECT 114.630 136.085 114.880 136.675 ;
        RECT 115.230 136.525 115.400 137.135 ;
        RECT 115.570 136.705 115.900 137.395 ;
        RECT 116.130 136.845 116.370 137.135 ;
        RECT 116.570 137.015 116.990 137.395 ;
        RECT 117.170 136.925 117.800 137.175 ;
        RECT 118.270 137.015 118.600 137.395 ;
        RECT 117.170 136.845 117.340 136.925 ;
        RECT 118.770 136.845 118.940 137.135 ;
        RECT 119.120 137.015 119.500 137.395 ;
        RECT 119.740 137.010 120.570 137.180 ;
        RECT 116.130 136.675 117.340 136.845 ;
        RECT 114.080 135.755 114.880 136.085 ;
        RECT 111.825 135.415 112.755 135.585 ;
        RECT 111.825 135.380 112.000 135.415 ;
        RECT 111.470 135.015 112.000 135.380 ;
        RECT 112.425 134.845 112.755 135.245 ;
        RECT 112.925 135.015 113.180 135.585 ;
        RECT 113.645 135.555 113.910 135.695 ;
        RECT 113.645 135.525 113.985 135.555 ;
        RECT 113.730 135.025 113.985 135.525 ;
        RECT 114.165 134.845 114.450 135.305 ;
        RECT 114.630 135.105 114.880 135.755 ;
        RECT 115.080 136.505 115.400 136.525 ;
        RECT 115.080 136.335 117.000 136.505 ;
        RECT 115.080 135.440 115.270 136.335 ;
        RECT 117.170 136.165 117.340 136.675 ;
        RECT 117.510 136.415 118.030 136.725 ;
        RECT 115.440 135.995 117.340 136.165 ;
        RECT 115.440 135.935 115.770 135.995 ;
        RECT 115.920 135.765 116.250 135.825 ;
        RECT 115.590 135.495 116.250 135.765 ;
        RECT 115.080 135.110 115.400 135.440 ;
        RECT 115.580 134.845 116.240 135.325 ;
        RECT 116.440 135.235 116.610 135.995 ;
        RECT 117.510 135.825 117.690 136.235 ;
        RECT 116.780 135.655 117.110 135.775 ;
        RECT 117.860 135.655 118.030 136.415 ;
        RECT 116.780 135.485 118.030 135.655 ;
        RECT 118.200 136.595 119.570 136.845 ;
        RECT 118.200 135.825 118.390 136.595 ;
        RECT 119.320 136.335 119.570 136.595 ;
        RECT 118.560 136.165 118.810 136.325 ;
        RECT 119.740 136.165 119.910 137.010 ;
        RECT 120.805 136.725 120.975 137.225 ;
        RECT 121.145 136.895 121.475 137.395 ;
        RECT 120.080 136.335 120.580 136.715 ;
        RECT 120.805 136.555 121.500 136.725 ;
        RECT 118.560 135.995 119.910 136.165 ;
        RECT 119.490 135.955 119.910 135.995 ;
        RECT 118.200 135.485 118.620 135.825 ;
        RECT 118.910 135.495 119.320 135.825 ;
        RECT 116.440 135.065 117.290 135.235 ;
        RECT 117.850 134.845 118.170 135.305 ;
        RECT 118.370 135.055 118.620 135.485 ;
        RECT 118.910 134.845 119.320 135.285 ;
        RECT 119.490 135.225 119.660 135.955 ;
        RECT 119.830 135.405 120.180 135.775 ;
        RECT 120.360 135.465 120.580 136.335 ;
        RECT 120.750 135.765 121.160 136.385 ;
        RECT 121.330 135.585 121.500 136.555 ;
        RECT 120.805 135.395 121.500 135.585 ;
        RECT 119.490 135.025 120.505 135.225 ;
        RECT 120.805 135.065 120.975 135.395 ;
        RECT 121.145 134.845 121.475 135.225 ;
        RECT 121.690 135.105 121.915 137.225 ;
        RECT 122.085 136.895 122.415 137.395 ;
        RECT 122.585 136.725 122.755 137.225 ;
        RECT 122.090 136.555 122.755 136.725 ;
        RECT 122.090 135.565 122.320 136.555 ;
        RECT 123.105 136.465 123.275 137.225 ;
        RECT 123.455 136.635 123.785 137.395 ;
        RECT 122.490 135.735 122.840 136.385 ;
        RECT 123.105 136.295 123.770 136.465 ;
        RECT 123.955 136.320 124.225 137.225 ;
        RECT 123.600 136.150 123.770 136.295 ;
        RECT 123.035 135.745 123.365 136.115 ;
        RECT 123.600 135.820 123.885 136.150 ;
        RECT 123.600 135.565 123.770 135.820 ;
        RECT 122.090 135.395 122.755 135.565 ;
        RECT 122.085 134.845 122.415 135.225 ;
        RECT 122.585 135.105 122.755 135.395 ;
        RECT 123.105 135.395 123.770 135.565 ;
        RECT 124.055 135.520 124.225 136.320 ;
        RECT 124.395 136.305 126.065 137.395 ;
        RECT 126.235 136.305 127.445 137.395 ;
        RECT 124.395 135.785 125.145 136.305 ;
        RECT 125.315 135.615 126.065 136.135 ;
        RECT 126.235 135.765 126.755 136.305 ;
        RECT 123.105 135.015 123.275 135.395 ;
        RECT 123.455 134.845 123.785 135.225 ;
        RECT 123.965 135.015 124.225 135.520 ;
        RECT 124.395 134.845 126.065 135.615 ;
        RECT 126.925 135.595 127.445 136.135 ;
        RECT 126.235 134.845 127.445 135.595 ;
        RECT 14.370 134.675 127.530 134.845 ;
        RECT 14.455 133.925 15.665 134.675 ;
        RECT 14.455 133.385 14.975 133.925 ;
        RECT 16.355 133.855 16.565 134.675 ;
        RECT 16.735 133.875 17.065 134.505 ;
        RECT 15.145 133.215 15.665 133.755 ;
        RECT 16.735 133.275 16.985 133.875 ;
        RECT 17.235 133.855 17.465 134.675 ;
        RECT 17.765 134.125 17.935 134.505 ;
        RECT 18.115 134.295 18.445 134.675 ;
        RECT 17.765 133.955 18.430 134.125 ;
        RECT 18.625 134.000 18.885 134.505 ;
        RECT 17.155 133.435 17.485 133.685 ;
        RECT 17.695 133.405 18.025 133.775 ;
        RECT 18.260 133.700 18.430 133.955 ;
        RECT 18.260 133.370 18.545 133.700 ;
        RECT 14.455 132.125 15.665 133.215 ;
        RECT 16.355 132.125 16.565 133.265 ;
        RECT 16.735 132.295 17.065 133.275 ;
        RECT 17.235 132.125 17.465 133.265 ;
        RECT 18.260 133.225 18.430 133.370 ;
        RECT 17.765 133.055 18.430 133.225 ;
        RECT 18.715 133.200 18.885 134.000 ;
        RECT 19.095 133.855 19.325 134.675 ;
        RECT 19.495 133.875 19.825 134.505 ;
        RECT 19.075 133.435 19.405 133.685 ;
        RECT 19.575 133.275 19.825 133.875 ;
        RECT 19.995 133.855 20.205 134.675 ;
        RECT 20.810 134.335 21.065 134.495 ;
        RECT 20.725 134.165 21.065 134.335 ;
        RECT 21.245 134.215 21.530 134.675 ;
        RECT 20.810 133.965 21.065 134.165 ;
        RECT 17.765 132.295 17.935 133.055 ;
        RECT 18.115 132.125 18.445 132.885 ;
        RECT 18.615 132.295 18.885 133.200 ;
        RECT 19.095 132.125 19.325 133.265 ;
        RECT 19.495 132.295 19.825 133.275 ;
        RECT 19.995 132.125 20.205 133.265 ;
        RECT 20.810 133.105 20.990 133.965 ;
        RECT 21.710 133.765 21.960 134.415 ;
        RECT 21.160 133.435 21.960 133.765 ;
        RECT 20.810 132.435 21.065 133.105 ;
        RECT 21.245 132.125 21.530 132.925 ;
        RECT 21.710 132.845 21.960 133.435 ;
        RECT 22.160 134.080 22.480 134.410 ;
        RECT 22.660 134.195 23.320 134.675 ;
        RECT 23.520 134.285 24.370 134.455 ;
        RECT 22.160 133.185 22.350 134.080 ;
        RECT 22.670 133.755 23.330 134.025 ;
        RECT 23.000 133.695 23.330 133.755 ;
        RECT 22.520 133.525 22.850 133.585 ;
        RECT 23.520 133.525 23.690 134.285 ;
        RECT 24.930 134.215 25.250 134.675 ;
        RECT 25.450 134.035 25.700 134.465 ;
        RECT 25.990 134.235 26.400 134.675 ;
        RECT 26.570 134.295 27.585 134.495 ;
        RECT 23.860 133.865 25.110 134.035 ;
        RECT 23.860 133.745 24.190 133.865 ;
        RECT 22.520 133.355 24.420 133.525 ;
        RECT 22.160 133.015 24.080 133.185 ;
        RECT 22.160 132.995 22.480 133.015 ;
        RECT 21.710 132.335 22.040 132.845 ;
        RECT 22.310 132.385 22.480 132.995 ;
        RECT 24.250 132.845 24.420 133.355 ;
        RECT 24.590 133.285 24.770 133.695 ;
        RECT 24.940 133.105 25.110 133.865 ;
        RECT 22.650 132.125 22.980 132.815 ;
        RECT 23.210 132.675 24.420 132.845 ;
        RECT 24.590 132.795 25.110 133.105 ;
        RECT 25.280 133.695 25.700 134.035 ;
        RECT 25.990 133.695 26.400 134.025 ;
        RECT 25.280 132.925 25.470 133.695 ;
        RECT 26.570 133.565 26.740 134.295 ;
        RECT 27.885 134.125 28.055 134.455 ;
        RECT 28.225 134.295 28.555 134.675 ;
        RECT 26.910 133.745 27.260 134.115 ;
        RECT 26.570 133.525 26.990 133.565 ;
        RECT 25.640 133.355 26.990 133.525 ;
        RECT 25.640 133.195 25.890 133.355 ;
        RECT 26.400 132.925 26.650 133.185 ;
        RECT 25.280 132.675 26.650 132.925 ;
        RECT 23.210 132.385 23.450 132.675 ;
        RECT 24.250 132.595 24.420 132.675 ;
        RECT 23.650 132.125 24.070 132.505 ;
        RECT 24.250 132.345 24.880 132.595 ;
        RECT 25.350 132.125 25.680 132.505 ;
        RECT 25.850 132.385 26.020 132.675 ;
        RECT 26.820 132.510 26.990 133.355 ;
        RECT 27.440 133.185 27.660 134.055 ;
        RECT 27.885 133.935 28.580 134.125 ;
        RECT 27.160 132.805 27.660 133.185 ;
        RECT 27.830 133.135 28.240 133.755 ;
        RECT 28.410 132.965 28.580 133.935 ;
        RECT 27.885 132.795 28.580 132.965 ;
        RECT 26.200 132.125 26.580 132.505 ;
        RECT 26.820 132.340 27.650 132.510 ;
        RECT 27.885 132.295 28.055 132.795 ;
        RECT 28.225 132.125 28.555 132.625 ;
        RECT 28.770 132.295 28.995 134.415 ;
        RECT 29.165 134.295 29.495 134.675 ;
        RECT 29.665 134.125 29.835 134.415 ;
        RECT 29.170 133.955 29.835 134.125 ;
        RECT 30.755 134.045 31.085 134.405 ;
        RECT 31.705 134.215 31.955 134.675 ;
        RECT 32.125 134.215 32.685 134.505 ;
        RECT 29.170 132.965 29.400 133.955 ;
        RECT 30.755 133.855 32.145 134.045 ;
        RECT 29.570 133.135 29.920 133.785 ;
        RECT 31.975 133.765 32.145 133.855 ;
        RECT 30.570 133.435 31.245 133.685 ;
        RECT 31.465 133.435 31.805 133.685 ;
        RECT 31.975 133.435 32.265 133.765 ;
        RECT 30.570 133.075 30.835 133.435 ;
        RECT 31.975 133.185 32.145 133.435 ;
        RECT 31.205 133.015 32.145 133.185 ;
        RECT 29.170 132.795 29.835 132.965 ;
        RECT 29.165 132.125 29.495 132.625 ;
        RECT 29.665 132.295 29.835 132.795 ;
        RECT 30.755 132.125 31.035 132.795 ;
        RECT 31.205 132.465 31.505 133.015 ;
        RECT 32.435 132.845 32.685 134.215 ;
        RECT 33.130 133.865 33.375 134.470 ;
        RECT 33.595 134.140 34.105 134.675 ;
        RECT 31.705 132.125 32.035 132.845 ;
        RECT 32.225 132.295 32.685 132.845 ;
        RECT 32.855 133.695 34.085 133.865 ;
        RECT 32.855 132.885 33.195 133.695 ;
        RECT 33.365 133.130 34.115 133.320 ;
        RECT 32.855 132.475 33.370 132.885 ;
        RECT 33.605 132.125 33.775 132.885 ;
        RECT 33.945 132.465 34.115 133.130 ;
        RECT 34.285 133.145 34.475 134.505 ;
        RECT 34.645 133.655 34.920 134.505 ;
        RECT 35.110 134.140 35.640 134.505 ;
        RECT 36.065 134.275 36.395 134.675 ;
        RECT 35.465 134.105 35.640 134.140 ;
        RECT 34.645 133.485 34.925 133.655 ;
        RECT 34.645 133.345 34.920 133.485 ;
        RECT 35.125 133.145 35.295 133.945 ;
        RECT 34.285 132.975 35.295 133.145 ;
        RECT 35.465 133.935 36.395 134.105 ;
        RECT 36.565 133.935 36.820 134.505 ;
        RECT 36.995 133.950 37.285 134.675 ;
        RECT 35.465 132.805 35.635 133.935 ;
        RECT 36.225 133.765 36.395 133.935 ;
        RECT 34.510 132.635 35.635 132.805 ;
        RECT 35.805 133.435 36.000 133.765 ;
        RECT 36.225 133.435 36.480 133.765 ;
        RECT 35.805 132.465 35.975 133.435 ;
        RECT 36.650 133.265 36.820 133.935 ;
        RECT 37.455 133.905 39.125 134.675 ;
        RECT 39.305 134.175 39.635 134.675 ;
        RECT 39.835 134.105 40.005 134.455 ;
        RECT 40.205 134.275 40.535 134.675 ;
        RECT 40.705 134.105 40.875 134.455 ;
        RECT 41.045 134.275 41.425 134.675 ;
        RECT 33.945 132.295 35.975 132.465 ;
        RECT 36.145 132.125 36.315 133.265 ;
        RECT 36.485 132.295 36.820 133.265 ;
        RECT 36.995 132.125 37.285 133.290 ;
        RECT 37.455 133.215 38.205 133.735 ;
        RECT 38.375 133.385 39.125 133.905 ;
        RECT 39.300 133.435 39.650 134.005 ;
        RECT 39.835 133.935 41.445 134.105 ;
        RECT 41.615 134.000 41.885 134.345 ;
        RECT 42.065 134.175 42.395 134.675 ;
        RECT 42.595 134.105 42.765 134.455 ;
        RECT 42.965 134.275 43.295 134.675 ;
        RECT 43.465 134.105 43.635 134.455 ;
        RECT 43.805 134.275 44.185 134.675 ;
        RECT 41.275 133.765 41.445 133.935 ;
        RECT 37.455 132.125 39.125 133.215 ;
        RECT 39.300 132.975 39.620 133.265 ;
        RECT 39.820 133.145 40.530 133.765 ;
        RECT 40.700 133.435 41.105 133.765 ;
        RECT 41.275 133.435 41.545 133.765 ;
        RECT 41.275 133.265 41.445 133.435 ;
        RECT 41.715 133.265 41.885 134.000 ;
        RECT 42.060 133.435 42.410 134.005 ;
        RECT 42.595 133.935 44.205 134.105 ;
        RECT 44.375 134.000 44.645 134.345 ;
        RECT 44.035 133.765 44.205 133.935 ;
        RECT 40.720 133.095 41.445 133.265 ;
        RECT 40.720 132.975 40.890 133.095 ;
        RECT 39.300 132.805 40.890 132.975 ;
        RECT 39.300 132.345 40.955 132.635 ;
        RECT 41.125 132.125 41.405 132.925 ;
        RECT 41.615 132.295 41.885 133.265 ;
        RECT 42.060 132.975 42.380 133.265 ;
        RECT 42.580 133.145 43.290 133.765 ;
        RECT 43.460 133.435 43.865 133.765 ;
        RECT 44.035 133.435 44.305 133.765 ;
        RECT 44.035 133.265 44.205 133.435 ;
        RECT 44.475 133.265 44.645 134.000 ;
        RECT 43.480 133.095 44.205 133.265 ;
        RECT 43.480 132.975 43.650 133.095 ;
        RECT 42.060 132.805 43.650 132.975 ;
        RECT 42.060 132.345 43.715 132.635 ;
        RECT 43.885 132.125 44.165 132.925 ;
        RECT 44.375 132.295 44.645 133.265 ;
        RECT 44.815 133.875 45.155 134.505 ;
        RECT 45.325 133.875 45.575 134.675 ;
        RECT 45.765 134.025 46.095 134.505 ;
        RECT 46.265 134.215 46.490 134.675 ;
        RECT 46.660 134.025 46.990 134.505 ;
        RECT 44.815 133.315 44.990 133.875 ;
        RECT 45.765 133.855 46.990 134.025 ;
        RECT 47.620 133.895 48.120 134.505 ;
        RECT 45.160 133.515 45.855 133.685 ;
        RECT 44.815 133.265 45.045 133.315 ;
        RECT 45.685 133.265 45.855 133.515 ;
        RECT 46.030 133.485 46.450 133.685 ;
        RECT 46.620 133.485 46.950 133.685 ;
        RECT 47.120 133.485 47.450 133.685 ;
        RECT 47.620 133.265 47.790 133.895 ;
        RECT 48.495 133.875 48.835 134.505 ;
        RECT 49.005 133.875 49.255 134.675 ;
        RECT 49.445 134.025 49.775 134.505 ;
        RECT 49.945 134.215 50.170 134.675 ;
        RECT 50.340 134.025 50.670 134.505 ;
        RECT 48.495 133.825 48.725 133.875 ;
        RECT 49.445 133.855 50.670 134.025 ;
        RECT 51.300 133.895 51.800 134.505 ;
        RECT 52.550 134.335 52.805 134.495 ;
        RECT 52.465 134.165 52.805 134.335 ;
        RECT 52.985 134.215 53.270 134.675 ;
        RECT 52.550 133.965 52.805 134.165 ;
        RECT 47.975 133.435 48.325 133.685 ;
        RECT 48.495 133.265 48.670 133.825 ;
        RECT 48.840 133.515 49.535 133.685 ;
        RECT 49.365 133.265 49.535 133.515 ;
        RECT 49.710 133.485 50.130 133.685 ;
        RECT 50.300 133.485 50.630 133.685 ;
        RECT 50.800 133.485 51.130 133.685 ;
        RECT 51.300 133.265 51.470 133.895 ;
        RECT 51.655 133.435 52.005 133.685 ;
        RECT 44.815 132.295 45.155 133.265 ;
        RECT 45.325 132.125 45.495 133.265 ;
        RECT 45.685 133.095 48.120 133.265 ;
        RECT 45.765 132.125 46.015 132.925 ;
        RECT 46.660 132.295 46.990 133.095 ;
        RECT 47.290 132.125 47.620 132.925 ;
        RECT 47.790 132.295 48.120 133.095 ;
        RECT 48.495 132.295 48.835 133.265 ;
        RECT 49.005 132.125 49.175 133.265 ;
        RECT 49.365 133.095 51.800 133.265 ;
        RECT 49.445 132.125 49.695 132.925 ;
        RECT 50.340 132.295 50.670 133.095 ;
        RECT 50.970 132.125 51.300 132.925 ;
        RECT 51.470 132.295 51.800 133.095 ;
        RECT 52.550 133.105 52.730 133.965 ;
        RECT 53.450 133.765 53.700 134.415 ;
        RECT 52.900 133.435 53.700 133.765 ;
        RECT 52.550 132.435 52.805 133.105 ;
        RECT 52.985 132.125 53.270 132.925 ;
        RECT 53.450 132.845 53.700 133.435 ;
        RECT 53.900 134.080 54.220 134.410 ;
        RECT 54.400 134.195 55.060 134.675 ;
        RECT 55.260 134.285 56.110 134.455 ;
        RECT 53.900 133.185 54.090 134.080 ;
        RECT 54.410 133.755 55.070 134.025 ;
        RECT 54.740 133.695 55.070 133.755 ;
        RECT 54.260 133.525 54.590 133.585 ;
        RECT 55.260 133.525 55.430 134.285 ;
        RECT 56.670 134.215 56.990 134.675 ;
        RECT 57.190 134.035 57.440 134.465 ;
        RECT 57.730 134.235 58.140 134.675 ;
        RECT 58.310 134.295 59.325 134.495 ;
        RECT 55.600 133.865 56.850 134.035 ;
        RECT 55.600 133.745 55.930 133.865 ;
        RECT 54.260 133.355 56.160 133.525 ;
        RECT 53.900 133.015 55.820 133.185 ;
        RECT 53.900 132.995 54.220 133.015 ;
        RECT 53.450 132.335 53.780 132.845 ;
        RECT 54.050 132.385 54.220 132.995 ;
        RECT 55.990 132.845 56.160 133.355 ;
        RECT 56.330 133.285 56.510 133.695 ;
        RECT 56.680 133.105 56.850 133.865 ;
        RECT 54.390 132.125 54.720 132.815 ;
        RECT 54.950 132.675 56.160 132.845 ;
        RECT 56.330 132.795 56.850 133.105 ;
        RECT 57.020 133.695 57.440 134.035 ;
        RECT 57.730 133.695 58.140 134.025 ;
        RECT 57.020 132.925 57.210 133.695 ;
        RECT 58.310 133.565 58.480 134.295 ;
        RECT 59.625 134.125 59.795 134.455 ;
        RECT 59.965 134.295 60.295 134.675 ;
        RECT 58.650 133.745 59.000 134.115 ;
        RECT 58.310 133.525 58.730 133.565 ;
        RECT 57.380 133.355 58.730 133.525 ;
        RECT 57.380 133.195 57.630 133.355 ;
        RECT 58.140 132.925 58.390 133.185 ;
        RECT 57.020 132.675 58.390 132.925 ;
        RECT 54.950 132.385 55.190 132.675 ;
        RECT 55.990 132.595 56.160 132.675 ;
        RECT 55.390 132.125 55.810 132.505 ;
        RECT 55.990 132.345 56.620 132.595 ;
        RECT 57.090 132.125 57.420 132.505 ;
        RECT 57.590 132.385 57.760 132.675 ;
        RECT 58.560 132.510 58.730 133.355 ;
        RECT 59.180 133.185 59.400 134.055 ;
        RECT 59.625 133.935 60.320 134.125 ;
        RECT 58.900 132.805 59.400 133.185 ;
        RECT 59.570 133.135 59.980 133.755 ;
        RECT 60.150 132.965 60.320 133.935 ;
        RECT 59.625 132.795 60.320 132.965 ;
        RECT 57.940 132.125 58.320 132.505 ;
        RECT 58.560 132.340 59.390 132.510 ;
        RECT 59.625 132.295 59.795 132.795 ;
        RECT 59.965 132.125 60.295 132.625 ;
        RECT 60.510 132.295 60.735 134.415 ;
        RECT 60.905 134.295 61.235 134.675 ;
        RECT 61.405 134.125 61.575 134.415 ;
        RECT 60.910 133.955 61.575 134.125 ;
        RECT 60.910 132.965 61.140 133.955 ;
        RECT 62.755 133.950 63.045 134.675 ;
        RECT 63.215 133.875 63.555 134.505 ;
        RECT 63.725 133.875 63.975 134.675 ;
        RECT 64.165 134.025 64.495 134.505 ;
        RECT 64.665 134.215 64.890 134.675 ;
        RECT 65.060 134.025 65.390 134.505 ;
        RECT 61.310 133.135 61.660 133.785 ;
        RECT 63.215 133.315 63.390 133.875 ;
        RECT 64.165 133.855 65.390 134.025 ;
        RECT 66.020 133.895 66.520 134.505 ;
        RECT 67.820 134.130 73.165 134.675 ;
        RECT 73.340 134.130 78.685 134.675 ;
        RECT 78.865 134.175 79.195 134.675 ;
        RECT 63.560 133.515 64.255 133.685 ;
        RECT 60.910 132.795 61.575 132.965 ;
        RECT 60.905 132.125 61.235 132.625 ;
        RECT 61.405 132.295 61.575 132.795 ;
        RECT 62.755 132.125 63.045 133.290 ;
        RECT 63.215 133.265 63.445 133.315 ;
        RECT 64.085 133.265 64.255 133.515 ;
        RECT 64.430 133.485 64.850 133.685 ;
        RECT 65.020 133.485 65.350 133.685 ;
        RECT 65.520 133.485 65.850 133.685 ;
        RECT 66.020 133.265 66.190 133.895 ;
        RECT 66.375 133.435 66.725 133.685 ;
        RECT 63.215 132.295 63.555 133.265 ;
        RECT 63.725 132.125 63.895 133.265 ;
        RECT 64.085 133.095 66.520 133.265 ;
        RECT 64.165 132.125 64.415 132.925 ;
        RECT 65.060 132.295 65.390 133.095 ;
        RECT 65.690 132.125 66.020 132.925 ;
        RECT 66.190 132.295 66.520 133.095 ;
        RECT 69.410 132.560 69.760 133.810 ;
        RECT 71.240 133.300 71.580 134.130 ;
        RECT 74.930 132.560 75.280 133.810 ;
        RECT 76.760 133.300 77.100 134.130 ;
        RECT 79.395 134.105 79.565 134.455 ;
        RECT 79.765 134.275 80.095 134.675 ;
        RECT 80.265 134.105 80.435 134.455 ;
        RECT 80.605 134.275 80.985 134.675 ;
        RECT 78.860 133.435 79.210 134.005 ;
        RECT 79.395 133.935 81.005 134.105 ;
        RECT 81.175 134.000 81.445 134.345 ;
        RECT 81.620 134.130 86.965 134.675 ;
        RECT 80.835 133.765 81.005 133.935 ;
        RECT 78.860 132.975 79.180 133.265 ;
        RECT 79.380 133.145 80.090 133.765 ;
        RECT 80.260 133.435 80.665 133.765 ;
        RECT 80.835 133.435 81.105 133.765 ;
        RECT 80.835 133.265 81.005 133.435 ;
        RECT 81.275 133.265 81.445 134.000 ;
        RECT 80.280 133.095 81.005 133.265 ;
        RECT 80.280 132.975 80.450 133.095 ;
        RECT 78.860 132.805 80.450 132.975 ;
        RECT 67.820 132.125 73.165 132.560 ;
        RECT 73.340 132.125 78.685 132.560 ;
        RECT 78.860 132.345 80.515 132.635 ;
        RECT 80.685 132.125 80.965 132.925 ;
        RECT 81.175 132.295 81.445 133.265 ;
        RECT 83.210 132.560 83.560 133.810 ;
        RECT 85.040 133.300 85.380 134.130 ;
        RECT 87.195 133.855 87.405 134.675 ;
        RECT 87.575 133.875 87.905 134.505 ;
        RECT 87.575 133.275 87.825 133.875 ;
        RECT 88.075 133.855 88.305 134.675 ;
        RECT 88.515 133.950 88.805 134.675 ;
        RECT 89.350 133.965 89.605 134.495 ;
        RECT 89.785 134.215 90.070 134.675 ;
        RECT 87.995 133.435 88.325 133.685 ;
        RECT 89.350 133.315 89.530 133.965 ;
        RECT 90.250 133.765 90.500 134.415 ;
        RECT 89.700 133.435 90.500 133.765 ;
        RECT 81.620 132.125 86.965 132.560 ;
        RECT 87.195 132.125 87.405 133.265 ;
        RECT 87.575 132.295 87.905 133.275 ;
        RECT 88.075 132.125 88.305 133.265 ;
        RECT 88.515 132.125 88.805 133.290 ;
        RECT 89.265 133.145 89.530 133.315 ;
        RECT 89.350 133.105 89.530 133.145 ;
        RECT 89.350 132.435 89.605 133.105 ;
        RECT 89.785 132.125 90.070 132.925 ;
        RECT 90.250 132.845 90.500 133.435 ;
        RECT 90.700 134.080 91.020 134.410 ;
        RECT 91.200 134.195 91.860 134.675 ;
        RECT 92.060 134.285 92.910 134.455 ;
        RECT 90.700 133.185 90.890 134.080 ;
        RECT 91.210 133.755 91.870 134.025 ;
        RECT 91.540 133.695 91.870 133.755 ;
        RECT 91.060 133.525 91.390 133.585 ;
        RECT 92.060 133.525 92.230 134.285 ;
        RECT 93.470 134.215 93.790 134.675 ;
        RECT 93.990 134.035 94.240 134.465 ;
        RECT 94.530 134.235 94.940 134.675 ;
        RECT 95.110 134.295 96.125 134.495 ;
        RECT 92.400 133.865 93.650 134.035 ;
        RECT 92.400 133.745 92.730 133.865 ;
        RECT 91.060 133.355 92.960 133.525 ;
        RECT 90.700 133.015 92.620 133.185 ;
        RECT 90.700 132.995 91.020 133.015 ;
        RECT 90.250 132.335 90.580 132.845 ;
        RECT 90.850 132.385 91.020 132.995 ;
        RECT 92.790 132.845 92.960 133.355 ;
        RECT 93.130 133.285 93.310 133.695 ;
        RECT 93.480 133.105 93.650 133.865 ;
        RECT 91.190 132.125 91.520 132.815 ;
        RECT 91.750 132.675 92.960 132.845 ;
        RECT 93.130 132.795 93.650 133.105 ;
        RECT 93.820 133.695 94.240 134.035 ;
        RECT 94.530 133.695 94.940 134.025 ;
        RECT 93.820 132.925 94.010 133.695 ;
        RECT 95.110 133.565 95.280 134.295 ;
        RECT 96.425 134.125 96.595 134.455 ;
        RECT 96.765 134.295 97.095 134.675 ;
        RECT 95.450 133.745 95.800 134.115 ;
        RECT 95.110 133.525 95.530 133.565 ;
        RECT 94.180 133.355 95.530 133.525 ;
        RECT 94.180 133.195 94.430 133.355 ;
        RECT 94.940 132.925 95.190 133.185 ;
        RECT 93.820 132.675 95.190 132.925 ;
        RECT 91.750 132.385 91.990 132.675 ;
        RECT 92.790 132.595 92.960 132.675 ;
        RECT 92.190 132.125 92.610 132.505 ;
        RECT 92.790 132.345 93.420 132.595 ;
        RECT 93.890 132.125 94.220 132.505 ;
        RECT 94.390 132.385 94.560 132.675 ;
        RECT 95.360 132.510 95.530 133.355 ;
        RECT 95.980 133.185 96.200 134.055 ;
        RECT 96.425 133.935 97.120 134.125 ;
        RECT 95.700 132.805 96.200 133.185 ;
        RECT 96.370 133.135 96.780 133.755 ;
        RECT 96.950 132.965 97.120 133.935 ;
        RECT 96.425 132.795 97.120 132.965 ;
        RECT 94.740 132.125 95.120 132.505 ;
        RECT 95.360 132.340 96.190 132.510 ;
        RECT 96.425 132.295 96.595 132.795 ;
        RECT 96.765 132.125 97.095 132.625 ;
        RECT 97.310 132.295 97.535 134.415 ;
        RECT 97.705 134.295 98.035 134.675 ;
        RECT 98.205 134.125 98.375 134.415 ;
        RECT 97.710 133.955 98.375 134.125 ;
        RECT 98.635 134.000 98.905 134.345 ;
        RECT 99.095 134.275 99.475 134.675 ;
        RECT 99.645 134.105 99.815 134.455 ;
        RECT 99.985 134.275 100.315 134.675 ;
        RECT 100.515 134.105 100.685 134.455 ;
        RECT 100.885 134.175 101.215 134.675 ;
        RECT 97.710 132.965 97.940 133.955 ;
        RECT 98.110 133.135 98.460 133.785 ;
        RECT 98.635 133.265 98.805 134.000 ;
        RECT 99.075 133.935 100.685 134.105 ;
        RECT 99.075 133.765 99.245 133.935 ;
        RECT 98.975 133.435 99.245 133.765 ;
        RECT 99.415 133.435 99.820 133.765 ;
        RECT 99.075 133.265 99.245 133.435 ;
        RECT 99.990 133.315 100.700 133.765 ;
        RECT 100.870 133.435 101.220 134.005 ;
        RECT 101.455 133.855 101.665 134.675 ;
        RECT 101.835 133.875 102.165 134.505 ;
        RECT 97.710 132.795 98.375 132.965 ;
        RECT 97.705 132.125 98.035 132.625 ;
        RECT 98.205 132.295 98.375 132.795 ;
        RECT 98.635 132.295 98.905 133.265 ;
        RECT 99.075 133.095 99.800 133.265 ;
        RECT 99.990 133.145 100.705 133.315 ;
        RECT 101.835 133.275 102.085 133.875 ;
        RECT 102.335 133.855 102.565 134.675 ;
        RECT 103.235 134.000 103.505 134.345 ;
        RECT 103.695 134.275 104.075 134.675 ;
        RECT 104.245 134.105 104.415 134.455 ;
        RECT 104.585 134.275 104.915 134.675 ;
        RECT 105.115 134.105 105.285 134.455 ;
        RECT 105.485 134.175 105.815 134.675 ;
        RECT 102.255 133.435 102.585 133.685 ;
        RECT 99.630 132.975 99.800 133.095 ;
        RECT 100.900 132.975 101.220 133.265 ;
        RECT 99.115 132.125 99.395 132.925 ;
        RECT 99.630 132.805 101.220 132.975 ;
        RECT 99.565 132.345 101.220 132.635 ;
        RECT 101.455 132.125 101.665 133.265 ;
        RECT 101.835 132.295 102.165 133.275 ;
        RECT 103.235 133.265 103.405 134.000 ;
        RECT 103.675 133.935 105.285 134.105 ;
        RECT 103.675 133.765 103.845 133.935 ;
        RECT 103.575 133.435 103.845 133.765 ;
        RECT 104.015 133.435 104.420 133.765 ;
        RECT 103.675 133.265 103.845 133.435 ;
        RECT 102.335 132.125 102.565 133.265 ;
        RECT 103.235 132.295 103.505 133.265 ;
        RECT 103.675 133.095 104.400 133.265 ;
        RECT 104.590 133.145 105.300 133.765 ;
        RECT 105.470 133.435 105.820 134.005 ;
        RECT 105.995 133.875 106.335 134.505 ;
        RECT 106.505 133.875 106.755 134.675 ;
        RECT 106.945 134.025 107.275 134.505 ;
        RECT 107.445 134.215 107.670 134.675 ;
        RECT 107.840 134.025 108.170 134.505 ;
        RECT 105.995 133.825 106.225 133.875 ;
        RECT 106.945 133.855 108.170 134.025 ;
        RECT 108.800 133.895 109.300 134.505 ;
        RECT 109.675 134.000 109.945 134.345 ;
        RECT 110.135 134.275 110.515 134.675 ;
        RECT 110.685 134.105 110.855 134.455 ;
        RECT 111.025 134.275 111.355 134.675 ;
        RECT 111.555 134.105 111.725 134.455 ;
        RECT 111.925 134.175 112.255 134.675 ;
        RECT 105.995 133.265 106.170 133.825 ;
        RECT 106.340 133.515 107.035 133.685 ;
        RECT 106.865 133.265 107.035 133.515 ;
        RECT 107.210 133.485 107.630 133.685 ;
        RECT 107.800 133.485 108.130 133.685 ;
        RECT 108.300 133.485 108.630 133.685 ;
        RECT 108.800 133.265 108.970 133.895 ;
        RECT 109.155 133.435 109.505 133.685 ;
        RECT 109.675 133.265 109.845 134.000 ;
        RECT 110.115 133.935 111.725 134.105 ;
        RECT 110.115 133.765 110.285 133.935 ;
        RECT 110.015 133.435 110.285 133.765 ;
        RECT 110.455 133.435 110.860 133.765 ;
        RECT 110.115 133.265 110.285 133.435 ;
        RECT 104.230 132.975 104.400 133.095 ;
        RECT 105.500 132.975 105.820 133.265 ;
        RECT 103.715 132.125 103.995 132.925 ;
        RECT 104.230 132.805 105.820 132.975 ;
        RECT 104.165 132.345 105.820 132.635 ;
        RECT 105.995 132.295 106.335 133.265 ;
        RECT 106.505 132.125 106.675 133.265 ;
        RECT 106.865 133.095 109.300 133.265 ;
        RECT 106.945 132.125 107.195 132.925 ;
        RECT 107.840 132.295 108.170 133.095 ;
        RECT 108.470 132.125 108.800 132.925 ;
        RECT 108.970 132.295 109.300 133.095 ;
        RECT 109.675 132.295 109.945 133.265 ;
        RECT 110.115 133.095 110.840 133.265 ;
        RECT 111.030 133.145 111.740 133.765 ;
        RECT 111.910 133.435 112.260 134.005 ;
        RECT 112.435 133.905 114.105 134.675 ;
        RECT 114.275 133.950 114.565 134.675 ;
        RECT 115.195 133.905 118.705 134.675 ;
        RECT 118.965 134.125 119.135 134.505 ;
        RECT 119.315 134.295 119.645 134.675 ;
        RECT 118.965 133.955 119.630 134.125 ;
        RECT 119.825 134.000 120.085 134.505 ;
        RECT 120.720 134.130 126.065 134.675 ;
        RECT 110.670 132.975 110.840 133.095 ;
        RECT 111.940 132.975 112.260 133.265 ;
        RECT 110.155 132.125 110.435 132.925 ;
        RECT 110.670 132.805 112.260 132.975 ;
        RECT 112.435 133.215 113.185 133.735 ;
        RECT 113.355 133.385 114.105 133.905 ;
        RECT 110.605 132.345 112.260 132.635 ;
        RECT 112.435 132.125 114.105 133.215 ;
        RECT 114.275 132.125 114.565 133.290 ;
        RECT 115.195 133.215 116.885 133.735 ;
        RECT 117.055 133.385 118.705 133.905 ;
        RECT 118.895 133.405 119.225 133.775 ;
        RECT 119.460 133.700 119.630 133.955 ;
        RECT 119.460 133.370 119.745 133.700 ;
        RECT 119.460 133.225 119.630 133.370 ;
        RECT 115.195 132.125 118.705 133.215 ;
        RECT 118.965 133.055 119.630 133.225 ;
        RECT 119.915 133.200 120.085 134.000 ;
        RECT 118.965 132.295 119.135 133.055 ;
        RECT 119.315 132.125 119.645 132.885 ;
        RECT 119.815 132.295 120.085 133.200 ;
        RECT 122.310 132.560 122.660 133.810 ;
        RECT 124.140 133.300 124.480 134.130 ;
        RECT 126.235 133.925 127.445 134.675 ;
        RECT 126.235 133.215 126.755 133.755 ;
        RECT 126.925 133.385 127.445 133.925 ;
        RECT 120.720 132.125 126.065 132.560 ;
        RECT 126.235 132.125 127.445 133.215 ;
        RECT 14.370 131.955 127.530 132.125 ;
        RECT 14.455 130.865 15.665 131.955 ;
        RECT 14.455 130.155 14.975 130.695 ;
        RECT 15.145 130.325 15.665 130.865 ;
        RECT 16.295 130.865 19.805 131.955 ;
        RECT 19.975 131.195 20.490 131.605 ;
        RECT 20.725 131.195 20.895 131.955 ;
        RECT 21.065 131.615 23.095 131.785 ;
        RECT 16.295 130.345 17.985 130.865 ;
        RECT 18.155 130.175 19.805 130.695 ;
        RECT 19.975 130.385 20.315 131.195 ;
        RECT 21.065 130.950 21.235 131.615 ;
        RECT 21.630 131.275 22.755 131.445 ;
        RECT 20.485 130.760 21.235 130.950 ;
        RECT 21.405 130.935 22.415 131.105 ;
        RECT 19.975 130.215 21.205 130.385 ;
        RECT 14.455 129.405 15.665 130.155 ;
        RECT 16.295 129.405 19.805 130.175 ;
        RECT 20.250 129.610 20.495 130.215 ;
        RECT 20.715 129.405 21.225 129.940 ;
        RECT 21.405 129.575 21.595 130.935 ;
        RECT 21.765 130.255 22.040 130.735 ;
        RECT 21.765 130.085 22.045 130.255 ;
        RECT 22.245 130.135 22.415 130.935 ;
        RECT 22.585 130.145 22.755 131.275 ;
        RECT 22.925 130.645 23.095 131.615 ;
        RECT 23.265 130.815 23.435 131.955 ;
        RECT 23.605 130.815 23.940 131.785 ;
        RECT 22.925 130.315 23.120 130.645 ;
        RECT 23.345 130.315 23.600 130.645 ;
        RECT 23.345 130.145 23.515 130.315 ;
        RECT 23.770 130.145 23.940 130.815 ;
        RECT 24.115 130.790 24.405 131.955 ;
        RECT 25.035 130.865 28.545 131.955 ;
        RECT 28.715 130.880 28.985 131.785 ;
        RECT 29.155 131.195 29.485 131.955 ;
        RECT 29.665 131.025 29.835 131.785 ;
        RECT 30.470 131.615 30.725 131.645 ;
        RECT 30.385 131.445 30.725 131.615 ;
        RECT 25.035 130.345 26.725 130.865 ;
        RECT 26.895 130.175 28.545 130.695 ;
        RECT 21.765 129.575 22.040 130.085 ;
        RECT 22.585 129.975 23.515 130.145 ;
        RECT 22.585 129.940 22.760 129.975 ;
        RECT 22.230 129.575 22.760 129.940 ;
        RECT 23.185 129.405 23.515 129.805 ;
        RECT 23.685 129.575 23.940 130.145 ;
        RECT 24.115 129.405 24.405 130.130 ;
        RECT 25.035 129.405 28.545 130.175 ;
        RECT 28.715 130.080 28.885 130.880 ;
        RECT 29.170 130.855 29.835 131.025 ;
        RECT 30.470 130.975 30.725 131.445 ;
        RECT 30.905 131.155 31.190 131.955 ;
        RECT 31.370 131.235 31.700 131.745 ;
        RECT 29.170 130.710 29.340 130.855 ;
        RECT 29.055 130.380 29.340 130.710 ;
        RECT 29.170 130.125 29.340 130.380 ;
        RECT 29.575 130.305 29.905 130.675 ;
        RECT 28.715 129.575 28.975 130.080 ;
        RECT 29.170 129.955 29.835 130.125 ;
        RECT 29.155 129.405 29.485 129.785 ;
        RECT 29.665 129.575 29.835 129.955 ;
        RECT 30.470 130.115 30.650 130.975 ;
        RECT 31.370 130.645 31.620 131.235 ;
        RECT 31.970 131.085 32.140 131.695 ;
        RECT 32.310 131.265 32.640 131.955 ;
        RECT 32.870 131.405 33.110 131.695 ;
        RECT 33.310 131.575 33.730 131.955 ;
        RECT 33.910 131.485 34.540 131.735 ;
        RECT 35.010 131.575 35.340 131.955 ;
        RECT 33.910 131.405 34.080 131.485 ;
        RECT 35.510 131.405 35.680 131.695 ;
        RECT 35.860 131.575 36.240 131.955 ;
        RECT 36.480 131.570 37.310 131.740 ;
        RECT 32.870 131.235 34.080 131.405 ;
        RECT 30.820 130.315 31.620 130.645 ;
        RECT 30.470 129.585 30.725 130.115 ;
        RECT 30.905 129.405 31.190 129.865 ;
        RECT 31.370 129.665 31.620 130.315 ;
        RECT 31.820 131.065 32.140 131.085 ;
        RECT 31.820 130.895 33.740 131.065 ;
        RECT 31.820 130.000 32.010 130.895 ;
        RECT 33.910 130.725 34.080 131.235 ;
        RECT 34.250 130.975 34.770 131.285 ;
        RECT 32.180 130.555 34.080 130.725 ;
        RECT 32.180 130.495 32.510 130.555 ;
        RECT 32.660 130.325 32.990 130.385 ;
        RECT 32.330 130.055 32.990 130.325 ;
        RECT 31.820 129.670 32.140 130.000 ;
        RECT 32.320 129.405 32.980 129.885 ;
        RECT 33.180 129.795 33.350 130.555 ;
        RECT 34.250 130.385 34.430 130.795 ;
        RECT 33.520 130.215 33.850 130.335 ;
        RECT 34.600 130.215 34.770 130.975 ;
        RECT 33.520 130.045 34.770 130.215 ;
        RECT 34.940 131.155 36.310 131.405 ;
        RECT 34.940 130.385 35.130 131.155 ;
        RECT 36.060 130.895 36.310 131.155 ;
        RECT 35.300 130.725 35.550 130.885 ;
        RECT 36.480 130.725 36.650 131.570 ;
        RECT 37.545 131.285 37.715 131.785 ;
        RECT 37.885 131.455 38.215 131.955 ;
        RECT 36.820 130.895 37.320 131.275 ;
        RECT 37.545 131.115 38.240 131.285 ;
        RECT 35.300 130.555 36.650 130.725 ;
        RECT 36.230 130.515 36.650 130.555 ;
        RECT 34.940 130.045 35.360 130.385 ;
        RECT 35.650 130.055 36.060 130.385 ;
        RECT 33.180 129.625 34.030 129.795 ;
        RECT 34.590 129.405 34.910 129.865 ;
        RECT 35.110 129.615 35.360 130.045 ;
        RECT 35.650 129.405 36.060 129.845 ;
        RECT 36.230 129.785 36.400 130.515 ;
        RECT 36.570 129.965 36.920 130.335 ;
        RECT 37.100 130.025 37.320 130.895 ;
        RECT 37.490 130.325 37.900 130.945 ;
        RECT 38.070 130.145 38.240 131.115 ;
        RECT 37.545 129.955 38.240 130.145 ;
        RECT 36.230 129.585 37.245 129.785 ;
        RECT 37.545 129.625 37.715 129.955 ;
        RECT 37.885 129.405 38.215 129.785 ;
        RECT 38.430 129.665 38.655 131.785 ;
        RECT 38.825 131.455 39.155 131.955 ;
        RECT 39.325 131.285 39.495 131.785 ;
        RECT 38.830 131.115 39.495 131.285 ;
        RECT 39.845 131.210 40.115 131.955 ;
        RECT 40.745 131.950 47.020 131.955 ;
        RECT 38.830 130.125 39.060 131.115 ;
        RECT 40.285 131.040 40.575 131.780 ;
        RECT 40.745 131.225 41.000 131.950 ;
        RECT 41.185 131.055 41.445 131.780 ;
        RECT 41.615 131.225 41.860 131.950 ;
        RECT 42.045 131.055 42.305 131.780 ;
        RECT 42.475 131.225 42.720 131.950 ;
        RECT 42.905 131.055 43.165 131.780 ;
        RECT 43.335 131.225 43.580 131.950 ;
        RECT 43.750 131.055 44.010 131.780 ;
        RECT 44.180 131.225 44.440 131.950 ;
        RECT 44.610 131.055 44.870 131.780 ;
        RECT 45.040 131.225 45.300 131.950 ;
        RECT 45.470 131.055 45.730 131.780 ;
        RECT 45.900 131.225 46.160 131.950 ;
        RECT 46.330 131.055 46.590 131.780 ;
        RECT 46.760 131.155 47.020 131.950 ;
        RECT 41.185 131.040 46.590 131.055 ;
        RECT 39.230 130.295 39.580 130.945 ;
        RECT 39.845 130.815 46.590 131.040 ;
        RECT 39.845 130.225 41.010 130.815 ;
        RECT 47.190 130.645 47.440 131.780 ;
        RECT 47.620 131.145 47.880 131.955 ;
        RECT 48.055 130.645 48.300 131.785 ;
        RECT 48.480 131.145 48.775 131.955 ;
        RECT 49.875 130.790 50.165 131.955 ;
        RECT 50.795 130.865 54.305 131.955 ;
        RECT 54.480 131.520 59.825 131.955 ;
        RECT 60.000 131.520 65.345 131.955 ;
        RECT 41.180 130.395 48.300 130.645 ;
        RECT 38.830 129.955 39.495 130.125 ;
        RECT 39.845 130.055 46.590 130.225 ;
        RECT 38.825 129.405 39.155 129.785 ;
        RECT 39.325 129.665 39.495 129.955 ;
        RECT 39.845 129.405 40.145 129.885 ;
        RECT 40.315 129.600 40.575 130.055 ;
        RECT 40.745 129.405 41.005 129.885 ;
        RECT 41.185 129.600 41.445 130.055 ;
        RECT 41.615 129.405 41.865 129.885 ;
        RECT 42.045 129.600 42.305 130.055 ;
        RECT 42.475 129.405 42.725 129.885 ;
        RECT 42.905 129.600 43.165 130.055 ;
        RECT 43.335 129.405 43.580 129.885 ;
        RECT 43.750 129.600 44.025 130.055 ;
        RECT 44.195 129.405 44.440 129.885 ;
        RECT 44.610 129.600 44.870 130.055 ;
        RECT 45.040 129.405 45.300 129.885 ;
        RECT 45.470 129.600 45.730 130.055 ;
        RECT 45.900 129.405 46.160 129.885 ;
        RECT 46.330 129.600 46.590 130.055 ;
        RECT 46.760 129.405 47.020 129.965 ;
        RECT 47.190 129.585 47.440 130.395 ;
        RECT 47.620 129.405 47.880 129.930 ;
        RECT 48.050 129.585 48.300 130.395 ;
        RECT 48.470 130.085 48.785 130.645 ;
        RECT 50.795 130.345 52.485 130.865 ;
        RECT 52.655 130.175 54.305 130.695 ;
        RECT 56.070 130.270 56.420 131.520 ;
        RECT 48.480 129.405 48.785 129.915 ;
        RECT 49.875 129.405 50.165 130.130 ;
        RECT 50.795 129.405 54.305 130.175 ;
        RECT 57.900 129.950 58.240 130.780 ;
        RECT 61.590 130.270 61.940 131.520 ;
        RECT 65.515 131.195 66.030 131.605 ;
        RECT 66.265 131.195 66.435 131.955 ;
        RECT 66.605 131.615 68.635 131.785 ;
        RECT 63.420 129.950 63.760 130.780 ;
        RECT 65.515 130.385 65.855 131.195 ;
        RECT 66.605 130.950 66.775 131.615 ;
        RECT 67.170 131.275 68.295 131.445 ;
        RECT 66.025 130.760 66.775 130.950 ;
        RECT 66.945 130.935 67.955 131.105 ;
        RECT 65.515 130.215 66.745 130.385 ;
        RECT 54.480 129.405 59.825 129.950 ;
        RECT 60.000 129.405 65.345 129.950 ;
        RECT 65.790 129.610 66.035 130.215 ;
        RECT 66.255 129.405 66.765 129.940 ;
        RECT 66.945 129.575 67.135 130.935 ;
        RECT 67.305 130.255 67.580 130.735 ;
        RECT 67.305 130.085 67.585 130.255 ;
        RECT 67.785 130.135 67.955 130.935 ;
        RECT 68.125 130.145 68.295 131.275 ;
        RECT 68.465 130.645 68.635 131.615 ;
        RECT 68.805 130.815 68.975 131.955 ;
        RECT 69.145 130.815 69.480 131.785 ;
        RECT 69.660 131.530 69.995 131.955 ;
        RECT 70.165 131.350 70.350 131.755 ;
        RECT 68.465 130.315 68.660 130.645 ;
        RECT 68.885 130.315 69.140 130.645 ;
        RECT 68.885 130.145 69.055 130.315 ;
        RECT 69.310 130.145 69.480 130.815 ;
        RECT 67.305 129.575 67.580 130.085 ;
        RECT 68.125 129.975 69.055 130.145 ;
        RECT 68.125 129.940 68.300 129.975 ;
        RECT 67.770 129.575 68.300 129.940 ;
        RECT 68.725 129.405 69.055 129.805 ;
        RECT 69.225 129.575 69.480 130.145 ;
        RECT 69.685 131.175 70.350 131.350 ;
        RECT 70.555 131.175 70.885 131.955 ;
        RECT 69.685 130.145 70.025 131.175 ;
        RECT 71.055 130.985 71.325 131.755 ;
        RECT 70.195 130.815 71.325 130.985 ;
        RECT 70.195 130.315 70.445 130.815 ;
        RECT 69.685 129.975 70.370 130.145 ;
        RECT 70.625 130.065 70.985 130.645 ;
        RECT 69.660 129.405 69.995 129.805 ;
        RECT 70.165 129.575 70.370 129.975 ;
        RECT 71.155 129.905 71.325 130.815 ;
        RECT 70.580 129.405 70.855 129.885 ;
        RECT 71.065 129.575 71.325 129.905 ;
        RECT 71.495 131.235 71.955 131.785 ;
        RECT 72.145 131.235 72.475 131.955 ;
        RECT 71.495 129.865 71.745 131.235 ;
        RECT 72.675 131.065 72.975 131.615 ;
        RECT 73.145 131.285 73.425 131.955 ;
        RECT 72.035 130.895 72.975 131.065 ;
        RECT 72.035 130.645 72.205 130.895 ;
        RECT 73.345 130.645 73.610 131.005 ;
        RECT 71.915 130.315 72.205 130.645 ;
        RECT 72.375 130.395 72.715 130.645 ;
        RECT 72.935 130.395 73.610 130.645 ;
        RECT 73.795 130.985 74.065 131.755 ;
        RECT 74.235 131.175 74.565 131.955 ;
        RECT 74.770 131.350 74.955 131.755 ;
        RECT 75.125 131.530 75.460 131.955 ;
        RECT 74.770 131.175 75.435 131.350 ;
        RECT 73.795 130.815 74.925 130.985 ;
        RECT 72.035 130.225 72.205 130.315 ;
        RECT 72.035 130.035 73.425 130.225 ;
        RECT 71.495 129.575 72.055 129.865 ;
        RECT 72.225 129.405 72.475 129.865 ;
        RECT 73.095 129.675 73.425 130.035 ;
        RECT 73.795 129.905 73.965 130.815 ;
        RECT 74.135 130.065 74.495 130.645 ;
        RECT 74.675 130.315 74.925 130.815 ;
        RECT 75.095 130.145 75.435 131.175 ;
        RECT 75.635 130.790 75.925 131.955 ;
        RECT 76.555 130.865 78.225 131.955 ;
        RECT 78.395 131.235 78.855 131.785 ;
        RECT 79.045 131.235 79.375 131.955 ;
        RECT 76.555 130.345 77.305 130.865 ;
        RECT 77.475 130.175 78.225 130.695 ;
        RECT 74.750 129.975 75.435 130.145 ;
        RECT 73.795 129.575 74.055 129.905 ;
        RECT 74.265 129.405 74.540 129.885 ;
        RECT 74.750 129.575 74.955 129.975 ;
        RECT 75.125 129.405 75.460 129.805 ;
        RECT 75.635 129.405 75.925 130.130 ;
        RECT 76.555 129.405 78.225 130.175 ;
        RECT 78.395 129.865 78.645 131.235 ;
        RECT 79.575 131.065 79.875 131.615 ;
        RECT 80.045 131.285 80.325 131.955 ;
        RECT 78.935 130.895 79.875 131.065 ;
        RECT 78.935 130.645 79.105 130.895 ;
        RECT 80.245 130.645 80.510 131.005 ;
        RECT 78.815 130.315 79.105 130.645 ;
        RECT 79.275 130.395 79.615 130.645 ;
        RECT 79.835 130.395 80.510 130.645 ;
        RECT 80.695 130.865 83.285 131.955 ;
        RECT 83.460 131.520 88.805 131.955 ;
        RECT 80.695 130.345 81.905 130.865 ;
        RECT 78.935 130.225 79.105 130.315 ;
        RECT 78.935 130.035 80.325 130.225 ;
        RECT 82.075 130.175 83.285 130.695 ;
        RECT 85.050 130.270 85.400 131.520 ;
        RECT 89.015 130.815 89.245 131.955 ;
        RECT 89.415 130.805 89.745 131.785 ;
        RECT 89.915 130.815 90.125 131.955 ;
        RECT 90.465 131.155 90.635 131.955 ;
        RECT 90.805 130.935 91.135 131.785 ;
        RECT 91.305 131.155 91.475 131.955 ;
        RECT 91.645 130.935 91.975 131.785 ;
        RECT 92.145 131.155 92.315 131.955 ;
        RECT 92.485 130.935 92.815 131.785 ;
        RECT 92.985 131.155 93.155 131.955 ;
        RECT 93.325 130.935 93.655 131.785 ;
        RECT 93.825 131.155 93.995 131.955 ;
        RECT 94.165 130.935 94.495 131.785 ;
        RECT 94.665 131.155 94.835 131.955 ;
        RECT 95.005 130.935 95.335 131.785 ;
        RECT 95.505 131.155 95.675 131.955 ;
        RECT 95.845 130.935 96.175 131.785 ;
        RECT 96.345 131.155 96.515 131.955 ;
        RECT 96.685 130.935 97.015 131.785 ;
        RECT 97.185 131.155 97.355 131.955 ;
        RECT 97.525 130.935 97.855 131.785 ;
        RECT 98.025 131.155 98.195 131.955 ;
        RECT 98.365 130.935 98.695 131.785 ;
        RECT 98.865 131.155 99.035 131.955 ;
        RECT 99.205 130.935 99.535 131.785 ;
        RECT 99.705 131.105 99.875 131.955 ;
        RECT 100.045 130.935 100.375 131.785 ;
        RECT 100.545 131.105 100.715 131.955 ;
        RECT 100.885 130.935 101.215 131.785 ;
        RECT 78.395 129.575 78.955 129.865 ;
        RECT 79.125 129.405 79.375 129.865 ;
        RECT 79.995 129.675 80.325 130.035 ;
        RECT 80.695 129.405 83.285 130.175 ;
        RECT 86.880 129.950 87.220 130.780 ;
        RECT 88.995 130.395 89.325 130.645 ;
        RECT 83.460 129.405 88.805 129.950 ;
        RECT 89.015 129.405 89.245 130.225 ;
        RECT 89.495 130.205 89.745 130.805 ;
        RECT 90.355 130.765 97.015 130.935 ;
        RECT 97.185 130.765 99.535 130.935 ;
        RECT 99.705 130.765 101.215 130.935 ;
        RECT 101.395 130.790 101.685 131.955 ;
        RECT 102.315 130.865 103.985 131.955 ;
        RECT 104.160 131.520 109.505 131.955 ;
        RECT 90.355 130.225 90.630 130.765 ;
        RECT 97.185 130.595 97.360 130.765 ;
        RECT 99.705 130.595 99.875 130.765 ;
        RECT 90.800 130.395 97.360 130.595 ;
        RECT 97.565 130.395 99.875 130.595 ;
        RECT 100.045 130.395 101.220 130.595 ;
        RECT 97.185 130.225 97.360 130.395 ;
        RECT 99.705 130.225 99.875 130.395 ;
        RECT 102.315 130.345 103.065 130.865 ;
        RECT 89.415 129.575 89.745 130.205 ;
        RECT 89.915 129.405 90.125 130.225 ;
        RECT 90.355 130.055 97.015 130.225 ;
        RECT 97.185 130.055 99.535 130.225 ;
        RECT 99.705 130.055 101.215 130.225 ;
        RECT 103.235 130.175 103.985 130.695 ;
        RECT 105.750 130.270 106.100 131.520 ;
        RECT 109.675 131.235 110.135 131.785 ;
        RECT 110.325 131.235 110.655 131.955 ;
        RECT 90.465 129.405 90.635 129.885 ;
        RECT 90.805 129.580 91.135 130.055 ;
        RECT 91.305 129.405 91.475 129.885 ;
        RECT 91.645 129.580 91.975 130.055 ;
        RECT 92.145 129.405 92.315 129.885 ;
        RECT 92.485 129.580 92.815 130.055 ;
        RECT 92.985 129.405 93.155 129.885 ;
        RECT 93.325 129.580 93.655 130.055 ;
        RECT 93.825 129.405 93.995 129.885 ;
        RECT 94.165 129.580 94.495 130.055 ;
        RECT 94.665 129.405 94.835 129.885 ;
        RECT 95.005 129.580 95.335 130.055 ;
        RECT 95.085 129.575 95.255 129.580 ;
        RECT 95.505 129.405 95.675 129.885 ;
        RECT 95.845 129.580 96.175 130.055 ;
        RECT 95.925 129.575 96.095 129.580 ;
        RECT 96.345 129.405 96.515 129.885 ;
        RECT 96.685 129.580 97.015 130.055 ;
        RECT 96.765 129.575 97.015 129.580 ;
        RECT 97.185 129.405 97.355 129.885 ;
        RECT 97.525 129.580 97.855 130.055 ;
        RECT 98.025 129.405 98.195 129.885 ;
        RECT 98.365 129.580 98.695 130.055 ;
        RECT 98.865 129.405 99.035 129.885 ;
        RECT 99.205 129.580 99.535 130.055 ;
        RECT 99.705 129.405 99.875 129.885 ;
        RECT 100.045 129.580 100.375 130.055 ;
        RECT 100.545 129.405 100.715 129.885 ;
        RECT 100.885 129.580 101.215 130.055 ;
        RECT 101.395 129.405 101.685 130.130 ;
        RECT 102.315 129.405 103.985 130.175 ;
        RECT 107.580 129.950 107.920 130.780 ;
        RECT 104.160 129.405 109.505 129.950 ;
        RECT 109.675 129.865 109.925 131.235 ;
        RECT 110.855 131.065 111.155 131.615 ;
        RECT 111.325 131.285 111.605 131.955 ;
        RECT 110.215 130.895 111.155 131.065 ;
        RECT 110.215 130.645 110.385 130.895 ;
        RECT 111.525 130.645 111.790 131.005 ;
        RECT 110.095 130.315 110.385 130.645 ;
        RECT 110.555 130.395 110.895 130.645 ;
        RECT 111.115 130.395 111.790 130.645 ;
        RECT 112.435 130.865 115.025 131.955 ;
        RECT 115.200 131.520 120.545 131.955 ;
        RECT 120.720 131.520 126.065 131.955 ;
        RECT 112.435 130.345 113.645 130.865 ;
        RECT 110.215 130.225 110.385 130.315 ;
        RECT 110.215 130.035 111.605 130.225 ;
        RECT 113.815 130.175 115.025 130.695 ;
        RECT 116.790 130.270 117.140 131.520 ;
        RECT 109.675 129.575 110.235 129.865 ;
        RECT 110.405 129.405 110.655 129.865 ;
        RECT 111.275 129.675 111.605 130.035 ;
        RECT 112.435 129.405 115.025 130.175 ;
        RECT 118.620 129.950 118.960 130.780 ;
        RECT 122.310 130.270 122.660 131.520 ;
        RECT 126.235 130.865 127.445 131.955 ;
        RECT 124.140 129.950 124.480 130.780 ;
        RECT 126.235 130.325 126.755 130.865 ;
        RECT 126.925 130.155 127.445 130.695 ;
        RECT 115.200 129.405 120.545 129.950 ;
        RECT 120.720 129.405 126.065 129.950 ;
        RECT 126.235 129.405 127.445 130.155 ;
        RECT 14.370 129.235 127.530 129.405 ;
        RECT 14.455 128.485 15.665 129.235 ;
        RECT 15.835 128.485 17.045 129.235 ;
        RECT 17.590 128.895 17.845 129.055 ;
        RECT 17.505 128.725 17.845 128.895 ;
        RECT 18.025 128.775 18.310 129.235 ;
        RECT 14.455 127.945 14.975 128.485 ;
        RECT 15.145 127.775 15.665 128.315 ;
        RECT 14.455 126.685 15.665 127.775 ;
        RECT 15.835 127.775 16.355 128.315 ;
        RECT 16.525 127.945 17.045 128.485 ;
        RECT 17.590 128.525 17.845 128.725 ;
        RECT 15.835 126.685 17.045 127.775 ;
        RECT 17.590 127.665 17.770 128.525 ;
        RECT 18.490 128.325 18.740 128.975 ;
        RECT 17.940 127.995 18.740 128.325 ;
        RECT 17.590 126.995 17.845 127.665 ;
        RECT 18.025 126.685 18.310 127.485 ;
        RECT 18.490 127.405 18.740 127.995 ;
        RECT 18.940 128.640 19.260 128.970 ;
        RECT 19.440 128.755 20.100 129.235 ;
        RECT 20.300 128.845 21.150 129.015 ;
        RECT 18.940 127.745 19.130 128.640 ;
        RECT 19.450 128.315 20.110 128.585 ;
        RECT 19.780 128.255 20.110 128.315 ;
        RECT 19.300 128.085 19.630 128.145 ;
        RECT 20.300 128.085 20.470 128.845 ;
        RECT 21.710 128.775 22.030 129.235 ;
        RECT 22.230 128.595 22.480 129.025 ;
        RECT 22.770 128.795 23.180 129.235 ;
        RECT 23.350 128.855 24.365 129.055 ;
        RECT 20.640 128.425 21.890 128.595 ;
        RECT 20.640 128.305 20.970 128.425 ;
        RECT 19.300 127.915 21.200 128.085 ;
        RECT 18.940 127.575 20.860 127.745 ;
        RECT 18.940 127.555 19.260 127.575 ;
        RECT 18.490 126.895 18.820 127.405 ;
        RECT 19.090 126.945 19.260 127.555 ;
        RECT 21.030 127.405 21.200 127.915 ;
        RECT 21.370 127.845 21.550 128.255 ;
        RECT 21.720 127.665 21.890 128.425 ;
        RECT 19.430 126.685 19.760 127.375 ;
        RECT 19.990 127.235 21.200 127.405 ;
        RECT 21.370 127.355 21.890 127.665 ;
        RECT 22.060 128.255 22.480 128.595 ;
        RECT 22.770 128.255 23.180 128.585 ;
        RECT 22.060 127.485 22.250 128.255 ;
        RECT 23.350 128.125 23.520 128.855 ;
        RECT 24.665 128.685 24.835 129.015 ;
        RECT 25.005 128.855 25.335 129.235 ;
        RECT 23.690 128.305 24.040 128.675 ;
        RECT 23.350 128.085 23.770 128.125 ;
        RECT 22.420 127.915 23.770 128.085 ;
        RECT 22.420 127.755 22.670 127.915 ;
        RECT 23.180 127.485 23.430 127.745 ;
        RECT 22.060 127.235 23.430 127.485 ;
        RECT 19.990 126.945 20.230 127.235 ;
        RECT 21.030 127.155 21.200 127.235 ;
        RECT 20.430 126.685 20.850 127.065 ;
        RECT 21.030 126.905 21.660 127.155 ;
        RECT 22.130 126.685 22.460 127.065 ;
        RECT 22.630 126.945 22.800 127.235 ;
        RECT 23.600 127.070 23.770 127.915 ;
        RECT 24.220 127.745 24.440 128.615 ;
        RECT 24.665 128.495 25.360 128.685 ;
        RECT 23.940 127.365 24.440 127.745 ;
        RECT 24.610 127.695 25.020 128.315 ;
        RECT 25.190 127.525 25.360 128.495 ;
        RECT 24.665 127.355 25.360 127.525 ;
        RECT 22.980 126.685 23.360 127.065 ;
        RECT 23.600 126.900 24.430 127.070 ;
        RECT 24.665 126.855 24.835 127.355 ;
        RECT 25.005 126.685 25.335 127.185 ;
        RECT 25.550 126.855 25.775 128.975 ;
        RECT 25.945 128.855 26.275 129.235 ;
        RECT 26.445 128.685 26.615 128.975 ;
        RECT 27.800 128.690 33.145 129.235 ;
        RECT 25.950 128.515 26.615 128.685 ;
        RECT 25.950 127.525 26.180 128.515 ;
        RECT 26.350 127.695 26.700 128.345 ;
        RECT 25.950 127.355 26.615 127.525 ;
        RECT 25.945 126.685 26.275 127.185 ;
        RECT 26.445 126.855 26.615 127.355 ;
        RECT 29.390 127.120 29.740 128.370 ;
        RECT 31.220 127.860 31.560 128.690 ;
        RECT 33.355 128.415 33.585 129.235 ;
        RECT 33.755 128.435 34.085 129.065 ;
        RECT 33.335 127.995 33.665 128.245 ;
        RECT 33.835 127.835 34.085 128.435 ;
        RECT 34.255 128.415 34.465 129.235 ;
        RECT 35.155 128.465 36.825 129.235 ;
        RECT 36.995 128.510 37.285 129.235 ;
        RECT 38.375 128.560 38.635 129.065 ;
        RECT 38.815 128.855 39.145 129.235 ;
        RECT 39.325 128.685 39.495 129.065 ;
        RECT 27.800 126.685 33.145 127.120 ;
        RECT 33.355 126.685 33.585 127.825 ;
        RECT 33.755 126.855 34.085 127.835 ;
        RECT 34.255 126.685 34.465 127.825 ;
        RECT 35.155 127.775 35.905 128.295 ;
        RECT 36.075 127.945 36.825 128.465 ;
        RECT 35.155 126.685 36.825 127.775 ;
        RECT 36.995 126.685 37.285 127.850 ;
        RECT 38.375 127.760 38.545 128.560 ;
        RECT 38.830 128.515 39.495 128.685 ;
        RECT 39.955 128.605 40.285 128.965 ;
        RECT 40.905 128.775 41.155 129.235 ;
        RECT 41.325 128.775 41.885 129.065 ;
        RECT 38.830 128.260 39.000 128.515 ;
        RECT 39.955 128.415 41.345 128.605 ;
        RECT 38.715 127.930 39.000 128.260 ;
        RECT 39.235 127.965 39.565 128.335 ;
        RECT 41.175 128.325 41.345 128.415 ;
        RECT 39.770 127.995 40.445 128.245 ;
        RECT 40.665 127.995 41.005 128.245 ;
        RECT 41.175 127.995 41.465 128.325 ;
        RECT 38.830 127.785 39.000 127.930 ;
        RECT 38.375 126.855 38.645 127.760 ;
        RECT 38.830 127.615 39.495 127.785 ;
        RECT 39.770 127.635 40.035 127.995 ;
        RECT 41.175 127.745 41.345 127.995 ;
        RECT 38.815 126.685 39.145 127.445 ;
        RECT 39.325 126.855 39.495 127.615 ;
        RECT 40.405 127.575 41.345 127.745 ;
        RECT 39.955 126.685 40.235 127.355 ;
        RECT 40.405 127.025 40.705 127.575 ;
        RECT 41.635 127.405 41.885 128.775 ;
        RECT 42.255 128.605 42.585 128.965 ;
        RECT 43.205 128.775 43.455 129.235 ;
        RECT 43.625 128.775 44.185 129.065 ;
        RECT 42.255 128.415 43.645 128.605 ;
        RECT 43.475 128.325 43.645 128.415 ;
        RECT 42.070 127.995 42.745 128.245 ;
        RECT 42.965 127.995 43.305 128.245 ;
        RECT 43.475 127.995 43.765 128.325 ;
        RECT 42.070 127.635 42.335 127.995 ;
        RECT 43.475 127.745 43.645 127.995 ;
        RECT 40.905 126.685 41.235 127.405 ;
        RECT 41.425 126.855 41.885 127.405 ;
        RECT 42.705 127.575 43.645 127.745 ;
        RECT 42.255 126.685 42.535 127.355 ;
        RECT 42.705 127.025 43.005 127.575 ;
        RECT 43.935 127.405 44.185 128.775 ;
        RECT 45.025 128.545 45.355 129.235 ;
        RECT 45.815 128.640 46.435 129.065 ;
        RECT 46.605 128.745 46.935 129.235 ;
        RECT 46.075 128.305 46.435 128.640 ;
        RECT 47.315 128.605 47.645 128.965 ;
        RECT 48.265 128.775 48.515 129.235 ;
        RECT 48.685 128.775 49.245 129.065 ;
        RECT 45.015 128.025 46.435 128.305 ;
        RECT 43.205 126.685 43.535 127.405 ;
        RECT 43.725 126.855 44.185 127.405 ;
        RECT 44.485 126.685 44.815 127.855 ;
        RECT 45.015 126.855 45.345 128.025 ;
        RECT 45.545 126.685 45.875 127.855 ;
        RECT 46.075 126.855 46.435 128.025 ;
        RECT 46.605 127.995 46.945 128.575 ;
        RECT 47.315 128.415 48.705 128.605 ;
        RECT 48.535 128.325 48.705 128.415 ;
        RECT 47.130 127.995 47.805 128.245 ;
        RECT 48.025 127.995 48.365 128.245 ;
        RECT 48.535 127.995 48.825 128.325 ;
        RECT 46.605 126.685 46.935 127.825 ;
        RECT 47.130 127.635 47.395 127.995 ;
        RECT 48.535 127.745 48.705 127.995 ;
        RECT 47.765 127.575 48.705 127.745 ;
        RECT 47.315 126.685 47.595 127.355 ;
        RECT 47.765 127.025 48.065 127.575 ;
        RECT 48.995 127.405 49.245 128.775 ;
        RECT 49.415 128.485 50.625 129.235 ;
        RECT 48.265 126.685 48.595 127.405 ;
        RECT 48.785 126.855 49.245 127.405 ;
        RECT 49.415 127.775 49.935 128.315 ;
        RECT 50.105 127.945 50.625 128.485 ;
        RECT 50.795 128.465 54.305 129.235 ;
        RECT 50.795 127.775 52.485 128.295 ;
        RECT 52.655 127.945 54.305 128.465 ;
        RECT 54.750 128.425 54.995 129.030 ;
        RECT 55.215 128.700 55.725 129.235 ;
        RECT 54.475 128.255 55.705 128.425 ;
        RECT 49.415 126.685 50.625 127.775 ;
        RECT 50.795 126.685 54.305 127.775 ;
        RECT 54.475 127.445 54.815 128.255 ;
        RECT 54.985 127.690 55.735 127.880 ;
        RECT 54.475 127.035 54.990 127.445 ;
        RECT 55.225 126.685 55.395 127.445 ;
        RECT 55.565 127.025 55.735 127.690 ;
        RECT 55.905 127.705 56.095 129.065 ;
        RECT 56.265 128.895 56.540 129.065 ;
        RECT 56.265 128.725 56.545 128.895 ;
        RECT 56.265 127.905 56.540 128.725 ;
        RECT 56.730 128.700 57.260 129.065 ;
        RECT 57.685 128.835 58.015 129.235 ;
        RECT 57.085 128.665 57.260 128.700 ;
        RECT 56.745 127.705 56.915 128.505 ;
        RECT 55.905 127.535 56.915 127.705 ;
        RECT 57.085 128.495 58.015 128.665 ;
        RECT 58.185 128.495 58.440 129.065 ;
        RECT 57.085 127.365 57.255 128.495 ;
        RECT 57.845 128.325 58.015 128.495 ;
        RECT 56.130 127.195 57.255 127.365 ;
        RECT 57.425 127.995 57.620 128.325 ;
        RECT 57.845 127.995 58.100 128.325 ;
        RECT 57.425 127.025 57.595 127.995 ;
        RECT 58.270 127.825 58.440 128.495 ;
        RECT 59.075 128.465 62.585 129.235 ;
        RECT 62.755 128.510 63.045 129.235 ;
        RECT 63.215 128.485 64.425 129.235 ;
        RECT 64.970 128.895 65.225 129.055 ;
        RECT 64.885 128.725 65.225 128.895 ;
        RECT 65.405 128.775 65.690 129.235 ;
        RECT 55.565 126.855 57.595 127.025 ;
        RECT 57.765 126.685 57.935 127.825 ;
        RECT 58.105 126.855 58.440 127.825 ;
        RECT 59.075 127.775 60.765 128.295 ;
        RECT 60.935 127.945 62.585 128.465 ;
        RECT 59.075 126.685 62.585 127.775 ;
        RECT 62.755 126.685 63.045 127.850 ;
        RECT 63.215 127.775 63.735 128.315 ;
        RECT 63.905 127.945 64.425 128.485 ;
        RECT 64.970 128.525 65.225 128.725 ;
        RECT 63.215 126.685 64.425 127.775 ;
        RECT 64.970 127.665 65.150 128.525 ;
        RECT 65.870 128.325 66.120 128.975 ;
        RECT 65.320 127.995 66.120 128.325 ;
        RECT 64.970 126.995 65.225 127.665 ;
        RECT 65.405 126.685 65.690 127.485 ;
        RECT 65.870 127.405 66.120 127.995 ;
        RECT 66.320 128.640 66.640 128.970 ;
        RECT 66.820 128.755 67.480 129.235 ;
        RECT 67.680 128.845 68.530 129.015 ;
        RECT 66.320 127.745 66.510 128.640 ;
        RECT 66.830 128.315 67.490 128.585 ;
        RECT 67.160 128.255 67.490 128.315 ;
        RECT 66.680 128.085 67.010 128.145 ;
        RECT 67.680 128.085 67.850 128.845 ;
        RECT 69.090 128.775 69.410 129.235 ;
        RECT 69.610 128.595 69.860 129.025 ;
        RECT 70.150 128.795 70.560 129.235 ;
        RECT 70.730 128.855 71.745 129.055 ;
        RECT 68.020 128.425 69.270 128.595 ;
        RECT 68.020 128.305 68.350 128.425 ;
        RECT 66.680 127.915 68.580 128.085 ;
        RECT 66.320 127.575 68.240 127.745 ;
        RECT 66.320 127.555 66.640 127.575 ;
        RECT 65.870 126.895 66.200 127.405 ;
        RECT 66.470 126.945 66.640 127.555 ;
        RECT 68.410 127.405 68.580 127.915 ;
        RECT 68.750 127.845 68.930 128.255 ;
        RECT 69.100 127.665 69.270 128.425 ;
        RECT 66.810 126.685 67.140 127.375 ;
        RECT 67.370 127.235 68.580 127.405 ;
        RECT 68.750 127.355 69.270 127.665 ;
        RECT 69.440 128.255 69.860 128.595 ;
        RECT 70.150 128.255 70.560 128.585 ;
        RECT 69.440 127.485 69.630 128.255 ;
        RECT 70.730 128.125 70.900 128.855 ;
        RECT 72.045 128.685 72.215 129.015 ;
        RECT 72.385 128.855 72.715 129.235 ;
        RECT 71.070 128.305 71.420 128.675 ;
        RECT 70.730 128.085 71.150 128.125 ;
        RECT 69.800 127.915 71.150 128.085 ;
        RECT 69.800 127.755 70.050 127.915 ;
        RECT 70.560 127.485 70.810 127.745 ;
        RECT 69.440 127.235 70.810 127.485 ;
        RECT 67.370 126.945 67.610 127.235 ;
        RECT 68.410 127.155 68.580 127.235 ;
        RECT 67.810 126.685 68.230 127.065 ;
        RECT 68.410 126.905 69.040 127.155 ;
        RECT 69.510 126.685 69.840 127.065 ;
        RECT 70.010 126.945 70.180 127.235 ;
        RECT 70.980 127.070 71.150 127.915 ;
        RECT 71.600 127.745 71.820 128.615 ;
        RECT 72.045 128.495 72.740 128.685 ;
        RECT 71.320 127.365 71.820 127.745 ;
        RECT 71.990 127.695 72.400 128.315 ;
        RECT 72.570 127.525 72.740 128.495 ;
        RECT 72.045 127.355 72.740 127.525 ;
        RECT 70.360 126.685 70.740 127.065 ;
        RECT 70.980 126.900 71.810 127.070 ;
        RECT 72.045 126.855 72.215 127.355 ;
        RECT 72.385 126.685 72.715 127.185 ;
        RECT 72.930 126.855 73.155 128.975 ;
        RECT 73.325 128.855 73.655 129.235 ;
        RECT 73.825 128.685 73.995 128.975 ;
        RECT 73.330 128.515 73.995 128.685 ;
        RECT 74.455 128.605 74.785 128.965 ;
        RECT 75.405 128.775 75.655 129.235 ;
        RECT 75.825 128.775 76.385 129.065 ;
        RECT 73.330 127.525 73.560 128.515 ;
        RECT 74.455 128.415 75.845 128.605 ;
        RECT 73.730 127.695 74.080 128.345 ;
        RECT 75.675 128.325 75.845 128.415 ;
        RECT 74.270 127.995 74.945 128.245 ;
        RECT 75.165 127.995 75.505 128.245 ;
        RECT 75.675 127.995 75.965 128.325 ;
        RECT 74.270 127.635 74.535 127.995 ;
        RECT 75.675 127.745 75.845 127.995 ;
        RECT 74.905 127.575 75.845 127.745 ;
        RECT 73.330 127.355 73.995 127.525 ;
        RECT 73.325 126.685 73.655 127.185 ;
        RECT 73.825 126.855 73.995 127.355 ;
        RECT 74.455 126.685 74.735 127.355 ;
        RECT 74.905 127.025 75.205 127.575 ;
        RECT 76.135 127.405 76.385 128.775 ;
        RECT 76.755 128.605 77.085 128.965 ;
        RECT 77.705 128.775 77.955 129.235 ;
        RECT 78.125 128.775 78.685 129.065 ;
        RECT 76.755 128.415 78.145 128.605 ;
        RECT 77.975 128.325 78.145 128.415 ;
        RECT 76.570 127.995 77.245 128.245 ;
        RECT 77.465 127.995 77.805 128.245 ;
        RECT 77.975 127.995 78.265 128.325 ;
        RECT 76.570 127.635 76.835 127.995 ;
        RECT 77.975 127.745 78.145 127.995 ;
        RECT 75.405 126.685 75.735 127.405 ;
        RECT 75.925 126.855 76.385 127.405 ;
        RECT 77.205 127.575 78.145 127.745 ;
        RECT 76.755 126.685 77.035 127.355 ;
        RECT 77.205 127.025 77.505 127.575 ;
        RECT 78.435 127.405 78.685 128.775 ;
        RECT 79.130 128.425 79.375 129.030 ;
        RECT 79.595 128.700 80.105 129.235 ;
        RECT 77.705 126.685 78.035 127.405 ;
        RECT 78.225 126.855 78.685 127.405 ;
        RECT 78.855 128.255 80.085 128.425 ;
        RECT 78.855 127.445 79.195 128.255 ;
        RECT 79.365 127.690 80.115 127.880 ;
        RECT 78.855 127.035 79.370 127.445 ;
        RECT 79.605 126.685 79.775 127.445 ;
        RECT 79.945 127.025 80.115 127.690 ;
        RECT 80.285 127.705 80.475 129.065 ;
        RECT 80.645 128.215 80.920 129.065 ;
        RECT 81.110 128.700 81.640 129.065 ;
        RECT 82.065 128.835 82.395 129.235 ;
        RECT 81.465 128.665 81.640 128.700 ;
        RECT 80.645 128.045 80.925 128.215 ;
        RECT 80.645 127.905 80.920 128.045 ;
        RECT 81.125 127.705 81.295 128.505 ;
        RECT 80.285 127.535 81.295 127.705 ;
        RECT 81.465 128.495 82.395 128.665 ;
        RECT 82.565 128.495 82.820 129.065 ;
        RECT 81.465 127.365 81.635 128.495 ;
        RECT 82.225 128.325 82.395 128.495 ;
        RECT 80.510 127.195 81.635 127.365 ;
        RECT 81.805 127.995 82.000 128.325 ;
        RECT 82.225 127.995 82.480 128.325 ;
        RECT 81.805 127.025 81.975 127.995 ;
        RECT 82.650 127.825 82.820 128.495 ;
        RECT 79.945 126.855 81.975 127.025 ;
        RECT 82.145 126.685 82.315 127.825 ;
        RECT 82.485 126.855 82.820 127.825 ;
        RECT 82.995 128.775 83.555 129.065 ;
        RECT 83.725 128.775 83.975 129.235 ;
        RECT 82.995 127.405 83.245 128.775 ;
        RECT 84.595 128.605 84.925 128.965 ;
        RECT 83.535 128.415 84.925 128.605 ;
        RECT 85.295 128.465 86.965 129.235 ;
        RECT 87.225 128.685 87.395 129.065 ;
        RECT 87.575 128.855 87.905 129.235 ;
        RECT 87.225 128.515 87.890 128.685 ;
        RECT 88.085 128.560 88.345 129.065 ;
        RECT 83.535 128.325 83.705 128.415 ;
        RECT 83.415 127.995 83.705 128.325 ;
        RECT 83.875 127.995 84.215 128.245 ;
        RECT 84.435 127.995 85.110 128.245 ;
        RECT 83.535 127.745 83.705 127.995 ;
        RECT 83.535 127.575 84.475 127.745 ;
        RECT 84.845 127.635 85.110 127.995 ;
        RECT 85.295 127.775 86.045 128.295 ;
        RECT 86.215 127.945 86.965 128.465 ;
        RECT 87.155 127.965 87.485 128.335 ;
        RECT 87.720 128.260 87.890 128.515 ;
        RECT 87.720 127.930 88.005 128.260 ;
        RECT 87.720 127.785 87.890 127.930 ;
        RECT 82.995 126.855 83.455 127.405 ;
        RECT 83.645 126.685 83.975 127.405 ;
        RECT 84.175 127.025 84.475 127.575 ;
        RECT 84.645 126.685 84.925 127.355 ;
        RECT 85.295 126.685 86.965 127.775 ;
        RECT 87.225 127.615 87.890 127.785 ;
        RECT 88.175 127.760 88.345 128.560 ;
        RECT 88.515 128.510 88.805 129.235 ;
        RECT 89.440 128.495 89.695 129.065 ;
        RECT 89.865 128.835 90.195 129.235 ;
        RECT 90.620 128.700 91.150 129.065 ;
        RECT 90.620 128.665 90.795 128.700 ;
        RECT 89.865 128.495 90.795 128.665 ;
        RECT 87.225 126.855 87.395 127.615 ;
        RECT 87.575 126.685 87.905 127.445 ;
        RECT 88.075 126.855 88.345 127.760 ;
        RECT 88.515 126.685 88.805 127.850 ;
        RECT 89.440 127.825 89.610 128.495 ;
        RECT 89.865 128.325 90.035 128.495 ;
        RECT 89.780 127.995 90.035 128.325 ;
        RECT 90.260 127.995 90.455 128.325 ;
        RECT 89.440 126.855 89.775 127.825 ;
        RECT 89.945 126.685 90.115 127.825 ;
        RECT 90.285 127.025 90.455 127.995 ;
        RECT 90.625 127.365 90.795 128.495 ;
        RECT 90.965 127.705 91.135 128.505 ;
        RECT 91.340 128.215 91.615 129.065 ;
        RECT 91.335 128.045 91.615 128.215 ;
        RECT 91.340 127.905 91.615 128.045 ;
        RECT 91.785 127.705 91.975 129.065 ;
        RECT 92.155 128.700 92.665 129.235 ;
        RECT 92.885 128.425 93.130 129.030 ;
        RECT 94.125 128.685 94.295 129.065 ;
        RECT 94.475 128.855 94.805 129.235 ;
        RECT 94.125 128.515 94.790 128.685 ;
        RECT 94.985 128.560 95.245 129.065 ;
        RECT 95.415 128.725 95.720 129.235 ;
        RECT 92.175 128.255 93.405 128.425 ;
        RECT 90.965 127.535 91.975 127.705 ;
        RECT 92.145 127.690 92.895 127.880 ;
        RECT 90.625 127.195 91.750 127.365 ;
        RECT 92.145 127.025 92.315 127.690 ;
        RECT 93.065 127.445 93.405 128.255 ;
        RECT 94.055 127.965 94.385 128.335 ;
        RECT 94.620 128.260 94.790 128.515 ;
        RECT 94.620 127.930 94.905 128.260 ;
        RECT 94.620 127.785 94.790 127.930 ;
        RECT 90.285 126.855 92.315 127.025 ;
        RECT 92.485 126.685 92.655 127.445 ;
        RECT 92.890 127.035 93.405 127.445 ;
        RECT 94.125 127.615 94.790 127.785 ;
        RECT 95.075 127.760 95.245 128.560 ;
        RECT 95.415 127.995 95.730 128.555 ;
        RECT 95.900 128.245 96.150 129.055 ;
        RECT 96.320 128.710 96.580 129.235 ;
        RECT 96.760 128.245 97.010 129.055 ;
        RECT 97.180 128.675 97.440 129.235 ;
        RECT 97.610 128.585 97.870 129.040 ;
        RECT 98.040 128.755 98.300 129.235 ;
        RECT 98.470 128.585 98.730 129.040 ;
        RECT 98.900 128.755 99.160 129.235 ;
        RECT 99.330 128.585 99.590 129.040 ;
        RECT 99.760 128.755 100.005 129.235 ;
        RECT 100.175 128.585 100.450 129.040 ;
        RECT 100.620 128.755 100.865 129.235 ;
        RECT 101.035 128.585 101.295 129.040 ;
        RECT 101.475 128.755 101.725 129.235 ;
        RECT 101.895 128.585 102.155 129.040 ;
        RECT 102.335 128.755 102.585 129.235 ;
        RECT 102.755 128.585 103.015 129.040 ;
        RECT 103.195 128.755 103.455 129.235 ;
        RECT 103.625 128.585 103.885 129.040 ;
        RECT 104.055 128.755 104.355 129.235 ;
        RECT 104.615 128.775 105.175 129.065 ;
        RECT 105.345 128.775 105.595 129.235 ;
        RECT 97.610 128.415 104.355 128.585 ;
        RECT 95.900 127.995 103.020 128.245 ;
        RECT 94.125 126.855 94.295 127.615 ;
        RECT 94.475 126.685 94.805 127.445 ;
        RECT 94.975 126.855 95.245 127.760 ;
        RECT 95.425 126.685 95.720 127.495 ;
        RECT 95.900 126.855 96.145 127.995 ;
        RECT 96.320 126.685 96.580 127.495 ;
        RECT 96.760 126.860 97.010 127.995 ;
        RECT 103.190 127.825 104.355 128.415 ;
        RECT 97.610 127.600 104.355 127.825 ;
        RECT 97.610 127.585 103.015 127.600 ;
        RECT 97.180 126.690 97.440 127.485 ;
        RECT 97.610 126.860 97.870 127.585 ;
        RECT 98.040 126.690 98.300 127.415 ;
        RECT 98.470 126.860 98.730 127.585 ;
        RECT 98.900 126.690 99.160 127.415 ;
        RECT 99.330 126.860 99.590 127.585 ;
        RECT 99.760 126.690 100.020 127.415 ;
        RECT 100.190 126.860 100.450 127.585 ;
        RECT 100.620 126.690 100.865 127.415 ;
        RECT 101.035 126.860 101.295 127.585 ;
        RECT 101.480 126.690 101.725 127.415 ;
        RECT 101.895 126.860 102.155 127.585 ;
        RECT 102.340 126.690 102.585 127.415 ;
        RECT 102.755 126.860 103.015 127.585 ;
        RECT 103.200 126.690 103.455 127.415 ;
        RECT 103.625 126.860 103.915 127.600 ;
        RECT 97.180 126.685 103.455 126.690 ;
        RECT 104.085 126.685 104.355 127.430 ;
        RECT 104.615 127.405 104.865 128.775 ;
        RECT 106.215 128.605 106.545 128.965 ;
        RECT 105.155 128.415 106.545 128.605 ;
        RECT 106.915 128.775 107.475 129.065 ;
        RECT 107.645 128.775 107.895 129.235 ;
        RECT 105.155 128.325 105.325 128.415 ;
        RECT 105.035 127.995 105.325 128.325 ;
        RECT 105.495 127.995 105.835 128.245 ;
        RECT 106.055 127.995 106.730 128.245 ;
        RECT 105.155 127.745 105.325 127.995 ;
        RECT 105.155 127.575 106.095 127.745 ;
        RECT 106.465 127.635 106.730 127.995 ;
        RECT 104.615 126.855 105.075 127.405 ;
        RECT 105.265 126.685 105.595 127.405 ;
        RECT 105.795 127.025 106.095 127.575 ;
        RECT 106.915 127.405 107.165 128.775 ;
        RECT 108.515 128.605 108.845 128.965 ;
        RECT 107.455 128.415 108.845 128.605 ;
        RECT 109.415 128.605 109.745 128.965 ;
        RECT 110.365 128.775 110.615 129.235 ;
        RECT 110.785 128.775 111.345 129.065 ;
        RECT 109.415 128.415 110.805 128.605 ;
        RECT 107.455 128.325 107.625 128.415 ;
        RECT 107.335 127.995 107.625 128.325 ;
        RECT 110.635 128.325 110.805 128.415 ;
        RECT 107.795 127.995 108.135 128.245 ;
        RECT 108.355 127.995 109.030 128.245 ;
        RECT 107.455 127.745 107.625 127.995 ;
        RECT 107.455 127.575 108.395 127.745 ;
        RECT 108.765 127.635 109.030 127.995 ;
        RECT 109.230 127.995 109.905 128.245 ;
        RECT 110.125 127.995 110.465 128.245 ;
        RECT 110.635 127.995 110.925 128.325 ;
        RECT 109.230 127.635 109.495 127.995 ;
        RECT 110.635 127.745 110.805 127.995 ;
        RECT 106.265 126.685 106.545 127.355 ;
        RECT 106.915 126.855 107.375 127.405 ;
        RECT 107.565 126.685 107.895 127.405 ;
        RECT 108.095 127.025 108.395 127.575 ;
        RECT 109.865 127.575 110.805 127.745 ;
        RECT 108.565 126.685 108.845 127.355 ;
        RECT 109.415 126.685 109.695 127.355 ;
        RECT 109.865 127.025 110.165 127.575 ;
        RECT 111.095 127.405 111.345 128.775 ;
        RECT 110.365 126.685 110.695 127.405 ;
        RECT 110.885 126.855 111.345 127.405 ;
        RECT 111.515 128.775 112.075 129.065 ;
        RECT 112.245 128.775 112.495 129.235 ;
        RECT 111.515 127.405 111.765 128.775 ;
        RECT 113.115 128.605 113.445 128.965 ;
        RECT 112.055 128.415 113.445 128.605 ;
        RECT 114.275 128.510 114.565 129.235 ;
        RECT 115.195 128.465 117.785 129.235 ;
        RECT 112.055 128.325 112.225 128.415 ;
        RECT 111.935 127.995 112.225 128.325 ;
        RECT 112.395 127.995 112.735 128.245 ;
        RECT 112.955 127.995 113.630 128.245 ;
        RECT 112.055 127.745 112.225 127.995 ;
        RECT 112.055 127.575 112.995 127.745 ;
        RECT 113.365 127.635 113.630 127.995 ;
        RECT 111.515 126.855 111.975 127.405 ;
        RECT 112.165 126.685 112.495 127.405 ;
        RECT 112.695 127.025 112.995 127.575 ;
        RECT 113.165 126.685 113.445 127.355 ;
        RECT 114.275 126.685 114.565 127.850 ;
        RECT 115.195 127.775 116.405 128.295 ;
        RECT 116.575 127.945 117.785 128.465 ;
        RECT 117.995 128.415 118.225 129.235 ;
        RECT 118.395 128.435 118.725 129.065 ;
        RECT 117.975 127.995 118.305 128.245 ;
        RECT 118.475 127.835 118.725 128.435 ;
        RECT 118.895 128.415 119.105 129.235 ;
        RECT 119.425 128.685 119.595 129.065 ;
        RECT 119.775 128.855 120.105 129.235 ;
        RECT 119.425 128.515 120.090 128.685 ;
        RECT 120.285 128.560 120.545 129.065 ;
        RECT 120.720 128.690 126.065 129.235 ;
        RECT 119.355 127.965 119.685 128.335 ;
        RECT 119.920 128.260 120.090 128.515 ;
        RECT 115.195 126.685 117.785 127.775 ;
        RECT 117.995 126.685 118.225 127.825 ;
        RECT 118.395 126.855 118.725 127.835 ;
        RECT 119.920 127.930 120.205 128.260 ;
        RECT 118.895 126.685 119.105 127.825 ;
        RECT 119.920 127.785 120.090 127.930 ;
        RECT 119.425 127.615 120.090 127.785 ;
        RECT 120.375 127.760 120.545 128.560 ;
        RECT 119.425 126.855 119.595 127.615 ;
        RECT 119.775 126.685 120.105 127.445 ;
        RECT 120.275 126.855 120.545 127.760 ;
        RECT 122.310 127.120 122.660 128.370 ;
        RECT 124.140 127.860 124.480 128.690 ;
        RECT 126.235 128.485 127.445 129.235 ;
        RECT 126.235 127.775 126.755 128.315 ;
        RECT 126.925 127.945 127.445 128.485 ;
        RECT 120.720 126.685 126.065 127.120 ;
        RECT 126.235 126.685 127.445 127.775 ;
        RECT 14.370 126.515 127.530 126.685 ;
        RECT 14.455 125.425 15.665 126.515 ;
        RECT 14.455 124.715 14.975 125.255 ;
        RECT 15.145 124.885 15.665 125.425 ;
        RECT 15.835 125.425 17.045 126.515 ;
        RECT 17.215 125.425 20.725 126.515 ;
        RECT 15.835 124.885 16.355 125.425 ;
        RECT 16.525 124.715 17.045 125.255 ;
        RECT 17.215 124.905 18.905 125.425 ;
        RECT 20.955 125.375 21.165 126.515 ;
        RECT 21.335 125.365 21.665 126.345 ;
        RECT 21.835 125.375 22.065 126.515 ;
        RECT 22.825 125.585 22.995 126.345 ;
        RECT 23.175 125.755 23.505 126.515 ;
        RECT 22.825 125.415 23.490 125.585 ;
        RECT 23.675 125.440 23.945 126.345 ;
        RECT 19.075 124.735 20.725 125.255 ;
        RECT 14.455 123.965 15.665 124.715 ;
        RECT 15.835 123.965 17.045 124.715 ;
        RECT 17.215 123.965 20.725 124.735 ;
        RECT 20.955 123.965 21.165 124.785 ;
        RECT 21.335 124.765 21.585 125.365 ;
        RECT 23.320 125.270 23.490 125.415 ;
        RECT 21.755 124.955 22.085 125.205 ;
        RECT 22.755 124.865 23.085 125.235 ;
        RECT 23.320 124.940 23.605 125.270 ;
        RECT 21.335 124.135 21.665 124.765 ;
        RECT 21.835 123.965 22.065 124.785 ;
        RECT 23.320 124.685 23.490 124.940 ;
        RECT 22.825 124.515 23.490 124.685 ;
        RECT 23.775 124.640 23.945 125.440 ;
        RECT 24.115 125.350 24.405 126.515 ;
        RECT 25.500 126.080 30.845 126.515 ;
        RECT 31.020 126.080 36.365 126.515 ;
        RECT 27.090 124.830 27.440 126.080 ;
        RECT 22.825 124.135 22.995 124.515 ;
        RECT 23.175 123.965 23.505 124.345 ;
        RECT 23.685 124.135 23.945 124.640 ;
        RECT 24.115 123.965 24.405 124.690 ;
        RECT 28.920 124.510 29.260 125.340 ;
        RECT 32.610 124.830 32.960 126.080 ;
        RECT 36.735 125.845 37.015 126.515 ;
        RECT 37.185 125.625 37.485 126.175 ;
        RECT 37.685 125.795 38.015 126.515 ;
        RECT 38.205 125.795 38.665 126.345 ;
        RECT 34.440 124.510 34.780 125.340 ;
        RECT 36.550 125.205 36.815 125.565 ;
        RECT 37.185 125.455 38.125 125.625 ;
        RECT 37.955 125.205 38.125 125.455 ;
        RECT 36.550 124.955 37.225 125.205 ;
        RECT 37.445 124.955 37.785 125.205 ;
        RECT 37.955 124.875 38.245 125.205 ;
        RECT 37.955 124.785 38.125 124.875 ;
        RECT 36.735 124.595 38.125 124.785 ;
        RECT 25.500 123.965 30.845 124.510 ;
        RECT 31.020 123.965 36.365 124.510 ;
        RECT 36.735 124.235 37.065 124.595 ;
        RECT 38.415 124.425 38.665 125.795 ;
        RECT 38.835 125.425 40.045 126.515 ;
        RECT 40.215 125.795 40.675 126.345 ;
        RECT 40.865 125.795 41.195 126.515 ;
        RECT 38.835 124.885 39.355 125.425 ;
        RECT 39.525 124.715 40.045 125.255 ;
        RECT 37.685 123.965 37.935 124.425 ;
        RECT 38.105 124.135 38.665 124.425 ;
        RECT 38.835 123.965 40.045 124.715 ;
        RECT 40.215 124.425 40.465 125.795 ;
        RECT 41.395 125.625 41.695 126.175 ;
        RECT 41.865 125.845 42.145 126.515 ;
        RECT 42.715 125.845 42.995 126.515 ;
        RECT 40.755 125.455 41.695 125.625 ;
        RECT 43.165 125.625 43.465 126.175 ;
        RECT 43.665 125.795 43.995 126.515 ;
        RECT 44.185 125.795 44.645 126.345 ;
        RECT 40.755 125.205 40.925 125.455 ;
        RECT 42.065 125.205 42.330 125.565 ;
        RECT 40.635 124.875 40.925 125.205 ;
        RECT 41.095 124.955 41.435 125.205 ;
        RECT 41.655 124.955 42.330 125.205 ;
        RECT 42.530 125.205 42.795 125.565 ;
        RECT 43.165 125.455 44.105 125.625 ;
        RECT 43.935 125.205 44.105 125.455 ;
        RECT 42.530 124.955 43.205 125.205 ;
        RECT 43.425 124.955 43.765 125.205 ;
        RECT 40.755 124.785 40.925 124.875 ;
        RECT 43.935 124.875 44.225 125.205 ;
        RECT 43.935 124.785 44.105 124.875 ;
        RECT 40.755 124.595 42.145 124.785 ;
        RECT 40.215 124.135 40.775 124.425 ;
        RECT 40.945 123.965 41.195 124.425 ;
        RECT 41.815 124.235 42.145 124.595 ;
        RECT 42.715 124.595 44.105 124.785 ;
        RECT 42.715 124.235 43.045 124.595 ;
        RECT 44.395 124.425 44.645 125.795 ;
        RECT 43.665 123.965 43.915 124.425 ;
        RECT 44.085 124.135 44.645 124.425 ;
        RECT 44.815 125.795 45.275 126.345 ;
        RECT 45.465 125.795 45.795 126.515 ;
        RECT 44.815 124.425 45.065 125.795 ;
        RECT 45.995 125.625 46.295 126.175 ;
        RECT 46.465 125.845 46.745 126.515 ;
        RECT 47.170 125.645 47.455 126.515 ;
        RECT 47.625 125.885 47.885 126.345 ;
        RECT 48.060 126.055 48.315 126.515 ;
        RECT 48.485 125.885 48.745 126.345 ;
        RECT 47.625 125.715 48.745 125.885 ;
        RECT 48.915 125.715 49.225 126.515 ;
        RECT 45.355 125.455 46.295 125.625 ;
        RECT 45.355 125.205 45.525 125.455 ;
        RECT 46.665 125.205 46.930 125.565 ;
        RECT 47.625 125.465 47.885 125.715 ;
        RECT 49.395 125.545 49.705 126.345 ;
        RECT 45.235 124.875 45.525 125.205 ;
        RECT 45.695 124.955 46.035 125.205 ;
        RECT 46.255 124.955 46.930 125.205 ;
        RECT 47.130 125.295 47.885 125.465 ;
        RECT 48.675 125.375 49.705 125.545 ;
        RECT 45.355 124.785 45.525 124.875 ;
        RECT 47.130 124.785 47.535 125.295 ;
        RECT 48.675 125.125 48.845 125.375 ;
        RECT 47.705 124.955 48.845 125.125 ;
        RECT 45.355 124.595 46.745 124.785 ;
        RECT 47.130 124.615 48.780 124.785 ;
        RECT 49.015 124.635 49.365 125.205 ;
        RECT 44.815 124.135 45.375 124.425 ;
        RECT 45.545 123.965 45.795 124.425 ;
        RECT 46.415 124.235 46.745 124.595 ;
        RECT 47.175 123.965 47.455 124.445 ;
        RECT 47.625 124.225 47.885 124.615 ;
        RECT 48.060 123.965 48.315 124.445 ;
        RECT 48.485 124.225 48.780 124.615 ;
        RECT 49.535 124.465 49.705 125.375 ;
        RECT 49.875 125.350 50.165 126.515 ;
        RECT 50.335 125.425 52.005 126.515 ;
        RECT 52.180 126.080 57.525 126.515 ;
        RECT 50.335 124.905 51.085 125.425 ;
        RECT 51.255 124.735 52.005 125.255 ;
        RECT 53.770 124.830 54.120 126.080 ;
        RECT 57.785 125.585 57.955 126.345 ;
        RECT 58.135 125.755 58.465 126.515 ;
        RECT 57.785 125.415 58.450 125.585 ;
        RECT 58.635 125.440 58.905 126.345 ;
        RECT 48.960 123.965 49.235 124.445 ;
        RECT 49.405 124.135 49.705 124.465 ;
        RECT 49.875 123.965 50.165 124.690 ;
        RECT 50.335 123.965 52.005 124.735 ;
        RECT 55.600 124.510 55.940 125.340 ;
        RECT 58.280 125.270 58.450 125.415 ;
        RECT 57.715 124.865 58.045 125.235 ;
        RECT 58.280 124.940 58.565 125.270 ;
        RECT 58.280 124.685 58.450 124.940 ;
        RECT 57.785 124.515 58.450 124.685 ;
        RECT 58.735 124.640 58.905 125.440 ;
        RECT 59.075 125.755 59.590 126.165 ;
        RECT 59.825 125.755 59.995 126.515 ;
        RECT 60.165 126.175 62.195 126.345 ;
        RECT 59.075 124.945 59.415 125.755 ;
        RECT 60.165 125.510 60.335 126.175 ;
        RECT 60.730 125.835 61.855 126.005 ;
        RECT 59.585 125.320 60.335 125.510 ;
        RECT 60.505 125.495 61.515 125.665 ;
        RECT 59.075 124.775 60.305 124.945 ;
        RECT 52.180 123.965 57.525 124.510 ;
        RECT 57.785 124.135 57.955 124.515 ;
        RECT 58.135 123.965 58.465 124.345 ;
        RECT 58.645 124.135 58.905 124.640 ;
        RECT 59.350 124.170 59.595 124.775 ;
        RECT 59.815 123.965 60.325 124.500 ;
        RECT 60.505 124.135 60.695 125.495 ;
        RECT 60.865 125.155 61.140 125.295 ;
        RECT 60.865 124.985 61.145 125.155 ;
        RECT 60.865 124.135 61.140 124.985 ;
        RECT 61.345 124.695 61.515 125.495 ;
        RECT 61.685 124.705 61.855 125.835 ;
        RECT 62.025 125.205 62.195 126.175 ;
        RECT 62.365 125.375 62.535 126.515 ;
        RECT 62.705 125.375 63.040 126.345 ;
        RECT 62.025 124.875 62.220 125.205 ;
        RECT 62.445 124.875 62.700 125.205 ;
        RECT 62.445 124.705 62.615 124.875 ;
        RECT 62.870 124.705 63.040 125.375 ;
        RECT 63.215 125.425 64.425 126.515 ;
        RECT 64.595 125.425 68.105 126.515 ;
        RECT 63.215 124.885 63.735 125.425 ;
        RECT 63.905 124.715 64.425 125.255 ;
        RECT 64.595 124.905 66.285 125.425 ;
        RECT 68.335 125.375 68.545 126.515 ;
        RECT 68.715 125.365 69.045 126.345 ;
        RECT 69.215 125.375 69.445 126.515 ;
        RECT 70.205 125.585 70.375 126.345 ;
        RECT 70.555 125.755 70.885 126.515 ;
        RECT 70.205 125.415 70.870 125.585 ;
        RECT 71.055 125.440 71.325 126.345 ;
        RECT 66.455 124.735 68.105 125.255 ;
        RECT 61.685 124.535 62.615 124.705 ;
        RECT 61.685 124.500 61.860 124.535 ;
        RECT 61.330 124.135 61.860 124.500 ;
        RECT 62.285 123.965 62.615 124.365 ;
        RECT 62.785 124.135 63.040 124.705 ;
        RECT 63.215 123.965 64.425 124.715 ;
        RECT 64.595 123.965 68.105 124.735 ;
        RECT 68.335 123.965 68.545 124.785 ;
        RECT 68.715 124.765 68.965 125.365 ;
        RECT 70.700 125.270 70.870 125.415 ;
        RECT 69.135 124.955 69.465 125.205 ;
        RECT 70.135 124.865 70.465 125.235 ;
        RECT 70.700 124.940 70.985 125.270 ;
        RECT 68.715 124.135 69.045 124.765 ;
        RECT 69.215 123.965 69.445 124.785 ;
        RECT 70.700 124.685 70.870 124.940 ;
        RECT 70.205 124.515 70.870 124.685 ;
        RECT 71.155 124.640 71.325 125.440 ;
        RECT 70.205 124.135 70.375 124.515 ;
        RECT 70.555 123.965 70.885 124.345 ;
        RECT 71.065 124.135 71.325 124.640 ;
        RECT 72.415 125.545 72.725 126.345 ;
        RECT 72.895 125.715 73.205 126.515 ;
        RECT 73.375 125.885 73.635 126.345 ;
        RECT 73.805 126.055 74.060 126.515 ;
        RECT 74.235 125.885 74.495 126.345 ;
        RECT 73.375 125.715 74.495 125.885 ;
        RECT 72.415 125.375 73.445 125.545 ;
        RECT 72.415 124.465 72.585 125.375 ;
        RECT 72.755 124.635 73.105 125.205 ;
        RECT 73.275 125.125 73.445 125.375 ;
        RECT 74.235 125.465 74.495 125.715 ;
        RECT 74.665 125.645 74.950 126.515 ;
        RECT 74.235 125.295 74.990 125.465 ;
        RECT 75.635 125.350 75.925 126.515 ;
        RECT 76.095 125.425 77.765 126.515 ;
        RECT 78.310 126.175 78.565 126.205 ;
        RECT 78.225 126.005 78.565 126.175 ;
        RECT 78.310 125.535 78.565 126.005 ;
        RECT 78.745 125.715 79.030 126.515 ;
        RECT 79.210 125.795 79.540 126.305 ;
        RECT 73.275 124.955 74.415 125.125 ;
        RECT 74.585 124.785 74.990 125.295 ;
        RECT 76.095 124.905 76.845 125.425 ;
        RECT 73.340 124.615 74.990 124.785 ;
        RECT 77.015 124.735 77.765 125.255 ;
        RECT 72.415 124.135 72.715 124.465 ;
        RECT 72.885 123.965 73.160 124.445 ;
        RECT 73.340 124.225 73.635 124.615 ;
        RECT 73.805 123.965 74.060 124.445 ;
        RECT 74.235 124.225 74.495 124.615 ;
        RECT 74.665 123.965 74.945 124.445 ;
        RECT 75.635 123.965 75.925 124.690 ;
        RECT 76.095 123.965 77.765 124.735 ;
        RECT 78.310 124.675 78.490 125.535 ;
        RECT 79.210 125.205 79.460 125.795 ;
        RECT 79.810 125.645 79.980 126.255 ;
        RECT 80.150 125.825 80.480 126.515 ;
        RECT 80.710 125.965 80.950 126.255 ;
        RECT 81.150 126.135 81.570 126.515 ;
        RECT 81.750 126.045 82.380 126.295 ;
        RECT 82.850 126.135 83.180 126.515 ;
        RECT 81.750 125.965 81.920 126.045 ;
        RECT 83.350 125.965 83.520 126.255 ;
        RECT 83.700 126.135 84.080 126.515 ;
        RECT 84.320 126.130 85.150 126.300 ;
        RECT 80.710 125.795 81.920 125.965 ;
        RECT 78.660 124.875 79.460 125.205 ;
        RECT 78.310 124.145 78.565 124.675 ;
        RECT 78.745 123.965 79.030 124.425 ;
        RECT 79.210 124.225 79.460 124.875 ;
        RECT 79.660 125.625 79.980 125.645 ;
        RECT 79.660 125.455 81.580 125.625 ;
        RECT 79.660 124.560 79.850 125.455 ;
        RECT 81.750 125.285 81.920 125.795 ;
        RECT 82.090 125.535 82.610 125.845 ;
        RECT 80.020 125.115 81.920 125.285 ;
        RECT 80.020 125.055 80.350 125.115 ;
        RECT 80.500 124.885 80.830 124.945 ;
        RECT 80.170 124.615 80.830 124.885 ;
        RECT 79.660 124.230 79.980 124.560 ;
        RECT 80.160 123.965 80.820 124.445 ;
        RECT 81.020 124.355 81.190 125.115 ;
        RECT 82.090 124.945 82.270 125.355 ;
        RECT 81.360 124.775 81.690 124.895 ;
        RECT 82.440 124.775 82.610 125.535 ;
        RECT 81.360 124.605 82.610 124.775 ;
        RECT 82.780 125.715 84.150 125.965 ;
        RECT 82.780 124.945 82.970 125.715 ;
        RECT 83.900 125.455 84.150 125.715 ;
        RECT 83.140 125.285 83.390 125.445 ;
        RECT 84.320 125.285 84.490 126.130 ;
        RECT 85.385 125.845 85.555 126.345 ;
        RECT 85.725 126.015 86.055 126.515 ;
        RECT 84.660 125.455 85.160 125.835 ;
        RECT 85.385 125.675 86.080 125.845 ;
        RECT 83.140 125.115 84.490 125.285 ;
        RECT 84.070 125.075 84.490 125.115 ;
        RECT 82.780 124.605 83.200 124.945 ;
        RECT 83.490 124.615 83.900 124.945 ;
        RECT 81.020 124.185 81.870 124.355 ;
        RECT 82.430 123.965 82.750 124.425 ;
        RECT 82.950 124.175 83.200 124.605 ;
        RECT 83.490 123.965 83.900 124.405 ;
        RECT 84.070 124.345 84.240 125.075 ;
        RECT 84.410 124.525 84.760 124.895 ;
        RECT 84.940 124.585 85.160 125.455 ;
        RECT 85.330 124.885 85.740 125.505 ;
        RECT 85.910 124.705 86.080 125.675 ;
        RECT 85.385 124.515 86.080 124.705 ;
        RECT 84.070 124.145 85.085 124.345 ;
        RECT 85.385 124.185 85.555 124.515 ;
        RECT 85.725 123.965 86.055 124.345 ;
        RECT 86.270 124.225 86.495 126.345 ;
        RECT 86.665 126.015 86.995 126.515 ;
        RECT 87.165 125.845 87.335 126.345 ;
        RECT 86.670 125.675 87.335 125.845 ;
        RECT 86.670 124.685 86.900 125.675 ;
        RECT 87.070 124.855 87.420 125.505 ;
        RECT 87.595 125.425 89.265 126.515 ;
        RECT 89.525 125.845 89.695 126.345 ;
        RECT 89.865 126.015 90.195 126.515 ;
        RECT 89.525 125.675 90.190 125.845 ;
        RECT 87.595 124.905 88.345 125.425 ;
        RECT 88.515 124.735 89.265 125.255 ;
        RECT 89.440 124.855 89.790 125.505 ;
        RECT 86.670 124.515 87.335 124.685 ;
        RECT 86.665 123.965 86.995 124.345 ;
        RECT 87.165 124.225 87.335 124.515 ;
        RECT 87.595 123.965 89.265 124.735 ;
        RECT 89.960 124.685 90.190 125.675 ;
        RECT 89.525 124.515 90.190 124.685 ;
        RECT 89.525 124.225 89.695 124.515 ;
        RECT 89.865 123.965 90.195 124.345 ;
        RECT 90.365 124.225 90.590 126.345 ;
        RECT 90.805 126.015 91.135 126.515 ;
        RECT 91.305 125.845 91.475 126.345 ;
        RECT 91.710 126.130 92.540 126.300 ;
        RECT 92.780 126.135 93.160 126.515 ;
        RECT 90.780 125.675 91.475 125.845 ;
        RECT 90.780 124.705 90.950 125.675 ;
        RECT 91.120 124.885 91.530 125.505 ;
        RECT 91.700 125.455 92.200 125.835 ;
        RECT 90.780 124.515 91.475 124.705 ;
        RECT 91.700 124.585 91.920 125.455 ;
        RECT 92.370 125.285 92.540 126.130 ;
        RECT 93.340 125.965 93.510 126.255 ;
        RECT 93.680 126.135 94.010 126.515 ;
        RECT 94.480 126.045 95.110 126.295 ;
        RECT 95.290 126.135 95.710 126.515 ;
        RECT 94.940 125.965 95.110 126.045 ;
        RECT 95.910 125.965 96.150 126.255 ;
        RECT 92.710 125.715 94.080 125.965 ;
        RECT 92.710 125.455 92.960 125.715 ;
        RECT 93.470 125.285 93.720 125.445 ;
        RECT 92.370 125.115 93.720 125.285 ;
        RECT 92.370 125.075 92.790 125.115 ;
        RECT 92.100 124.525 92.450 124.895 ;
        RECT 90.805 123.965 91.135 124.345 ;
        RECT 91.305 124.185 91.475 124.515 ;
        RECT 92.620 124.345 92.790 125.075 ;
        RECT 93.890 124.945 94.080 125.715 ;
        RECT 92.960 124.615 93.370 124.945 ;
        RECT 93.660 124.605 94.080 124.945 ;
        RECT 94.250 125.535 94.770 125.845 ;
        RECT 94.940 125.795 96.150 125.965 ;
        RECT 96.380 125.825 96.710 126.515 ;
        RECT 94.250 124.775 94.420 125.535 ;
        RECT 94.590 124.945 94.770 125.355 ;
        RECT 94.940 125.285 95.110 125.795 ;
        RECT 96.880 125.645 97.050 126.255 ;
        RECT 97.320 125.795 97.650 126.305 ;
        RECT 96.880 125.625 97.200 125.645 ;
        RECT 95.280 125.455 97.200 125.625 ;
        RECT 94.940 125.115 96.840 125.285 ;
        RECT 95.170 124.775 95.500 124.895 ;
        RECT 94.250 124.605 95.500 124.775 ;
        RECT 91.775 124.145 92.790 124.345 ;
        RECT 92.960 123.965 93.370 124.405 ;
        RECT 93.660 124.175 93.910 124.605 ;
        RECT 94.110 123.965 94.430 124.425 ;
        RECT 95.670 124.355 95.840 125.115 ;
        RECT 96.510 125.055 96.840 125.115 ;
        RECT 96.030 124.885 96.360 124.945 ;
        RECT 96.030 124.615 96.690 124.885 ;
        RECT 97.010 124.560 97.200 125.455 ;
        RECT 94.990 124.185 95.840 124.355 ;
        RECT 96.040 123.965 96.700 124.445 ;
        RECT 96.880 124.230 97.200 124.560 ;
        RECT 97.400 125.205 97.650 125.795 ;
        RECT 97.830 125.715 98.115 126.515 ;
        RECT 98.295 126.175 98.550 126.205 ;
        RECT 98.295 126.005 98.635 126.175 ;
        RECT 98.295 125.535 98.550 126.005 ;
        RECT 99.295 125.845 99.575 126.515 ;
        RECT 99.745 125.625 100.045 126.175 ;
        RECT 100.245 125.795 100.575 126.515 ;
        RECT 100.765 125.795 101.225 126.345 ;
        RECT 97.400 124.875 98.200 125.205 ;
        RECT 97.400 124.225 97.650 124.875 ;
        RECT 98.370 124.675 98.550 125.535 ;
        RECT 99.110 125.205 99.375 125.565 ;
        RECT 99.745 125.455 100.685 125.625 ;
        RECT 100.515 125.205 100.685 125.455 ;
        RECT 99.110 124.955 99.785 125.205 ;
        RECT 100.005 124.955 100.345 125.205 ;
        RECT 100.515 124.875 100.805 125.205 ;
        RECT 100.515 124.785 100.685 124.875 ;
        RECT 97.830 123.965 98.115 124.425 ;
        RECT 98.295 124.145 98.550 124.675 ;
        RECT 99.295 124.595 100.685 124.785 ;
        RECT 99.295 124.235 99.625 124.595 ;
        RECT 100.975 124.425 101.225 125.795 ;
        RECT 101.395 125.350 101.685 126.515 ;
        RECT 101.855 125.425 105.365 126.515 ;
        RECT 105.540 126.080 110.885 126.515 ;
        RECT 101.855 124.905 103.545 125.425 ;
        RECT 103.715 124.735 105.365 125.255 ;
        RECT 107.130 124.830 107.480 126.080 ;
        RECT 111.055 125.755 111.570 126.165 ;
        RECT 111.805 125.755 111.975 126.515 ;
        RECT 112.145 126.175 114.175 126.345 ;
        RECT 100.245 123.965 100.495 124.425 ;
        RECT 100.665 124.135 101.225 124.425 ;
        RECT 101.395 123.965 101.685 124.690 ;
        RECT 101.855 123.965 105.365 124.735 ;
        RECT 108.960 124.510 109.300 125.340 ;
        RECT 111.055 124.945 111.395 125.755 ;
        RECT 112.145 125.510 112.315 126.175 ;
        RECT 112.710 125.835 113.835 126.005 ;
        RECT 111.565 125.320 112.315 125.510 ;
        RECT 112.485 125.495 113.495 125.665 ;
        RECT 111.055 124.775 112.285 124.945 ;
        RECT 105.540 123.965 110.885 124.510 ;
        RECT 111.330 124.170 111.575 124.775 ;
        RECT 111.795 123.965 112.305 124.500 ;
        RECT 112.485 124.135 112.675 125.495 ;
        RECT 112.845 124.475 113.120 125.295 ;
        RECT 113.325 124.695 113.495 125.495 ;
        RECT 113.665 124.705 113.835 125.835 ;
        RECT 114.005 125.205 114.175 126.175 ;
        RECT 114.345 125.375 114.515 126.515 ;
        RECT 114.685 125.375 115.020 126.345 ;
        RECT 114.005 124.875 114.200 125.205 ;
        RECT 114.425 124.875 114.680 125.205 ;
        RECT 114.425 124.705 114.595 124.875 ;
        RECT 114.850 124.705 115.020 125.375 ;
        RECT 113.665 124.535 114.595 124.705 ;
        RECT 113.665 124.500 113.840 124.535 ;
        RECT 112.845 124.305 113.125 124.475 ;
        RECT 112.845 124.135 113.120 124.305 ;
        RECT 113.310 124.135 113.840 124.500 ;
        RECT 114.265 123.965 114.595 124.365 ;
        RECT 114.765 124.135 115.020 124.705 ;
        RECT 115.570 125.535 115.825 126.205 ;
        RECT 116.005 125.715 116.290 126.515 ;
        RECT 116.470 125.795 116.800 126.305 ;
        RECT 115.570 124.675 115.750 125.535 ;
        RECT 116.470 125.205 116.720 125.795 ;
        RECT 117.070 125.645 117.240 126.255 ;
        RECT 117.410 125.825 117.740 126.515 ;
        RECT 117.970 125.965 118.210 126.255 ;
        RECT 118.410 126.135 118.830 126.515 ;
        RECT 119.010 126.045 119.640 126.295 ;
        RECT 120.110 126.135 120.440 126.515 ;
        RECT 119.010 125.965 119.180 126.045 ;
        RECT 120.610 125.965 120.780 126.255 ;
        RECT 120.960 126.135 121.340 126.515 ;
        RECT 121.580 126.130 122.410 126.300 ;
        RECT 117.970 125.795 119.180 125.965 ;
        RECT 115.920 124.875 116.720 125.205 ;
        RECT 115.570 124.475 115.825 124.675 ;
        RECT 115.485 124.305 115.825 124.475 ;
        RECT 115.570 124.145 115.825 124.305 ;
        RECT 116.005 123.965 116.290 124.425 ;
        RECT 116.470 124.225 116.720 124.875 ;
        RECT 116.920 125.625 117.240 125.645 ;
        RECT 116.920 125.455 118.840 125.625 ;
        RECT 116.920 124.560 117.110 125.455 ;
        RECT 119.010 125.285 119.180 125.795 ;
        RECT 119.350 125.535 119.870 125.845 ;
        RECT 117.280 125.115 119.180 125.285 ;
        RECT 117.280 125.055 117.610 125.115 ;
        RECT 117.760 124.885 118.090 124.945 ;
        RECT 117.430 124.615 118.090 124.885 ;
        RECT 116.920 124.230 117.240 124.560 ;
        RECT 117.420 123.965 118.080 124.445 ;
        RECT 118.280 124.355 118.450 125.115 ;
        RECT 119.350 124.945 119.530 125.355 ;
        RECT 118.620 124.775 118.950 124.895 ;
        RECT 119.700 124.775 119.870 125.535 ;
        RECT 118.620 124.605 119.870 124.775 ;
        RECT 120.040 125.715 121.410 125.965 ;
        RECT 120.040 124.945 120.230 125.715 ;
        RECT 121.160 125.455 121.410 125.715 ;
        RECT 120.400 125.285 120.650 125.445 ;
        RECT 121.580 125.285 121.750 126.130 ;
        RECT 122.645 125.845 122.815 126.345 ;
        RECT 122.985 126.015 123.315 126.515 ;
        RECT 121.920 125.455 122.420 125.835 ;
        RECT 122.645 125.675 123.340 125.845 ;
        RECT 120.400 125.115 121.750 125.285 ;
        RECT 121.330 125.075 121.750 125.115 ;
        RECT 120.040 124.605 120.460 124.945 ;
        RECT 120.750 124.615 121.160 124.945 ;
        RECT 118.280 124.185 119.130 124.355 ;
        RECT 119.690 123.965 120.010 124.425 ;
        RECT 120.210 124.175 120.460 124.605 ;
        RECT 120.750 123.965 121.160 124.405 ;
        RECT 121.330 124.345 121.500 125.075 ;
        RECT 121.670 124.525 122.020 124.895 ;
        RECT 122.200 124.585 122.420 125.455 ;
        RECT 122.590 124.885 123.000 125.505 ;
        RECT 123.170 124.705 123.340 125.675 ;
        RECT 122.645 124.515 123.340 124.705 ;
        RECT 121.330 124.145 122.345 124.345 ;
        RECT 122.645 124.185 122.815 124.515 ;
        RECT 122.985 123.965 123.315 124.345 ;
        RECT 123.530 124.225 123.755 126.345 ;
        RECT 123.925 126.015 124.255 126.515 ;
        RECT 124.425 125.845 124.595 126.345 ;
        RECT 123.930 125.675 124.595 125.845 ;
        RECT 123.930 124.685 124.160 125.675 ;
        RECT 124.330 124.855 124.680 125.505 ;
        RECT 124.855 125.425 126.065 126.515 ;
        RECT 126.235 125.425 127.445 126.515 ;
        RECT 124.855 124.885 125.375 125.425 ;
        RECT 125.545 124.715 126.065 125.255 ;
        RECT 126.235 124.885 126.755 125.425 ;
        RECT 126.925 124.715 127.445 125.255 ;
        RECT 123.930 124.515 124.595 124.685 ;
        RECT 123.925 123.965 124.255 124.345 ;
        RECT 124.425 124.225 124.595 124.515 ;
        RECT 124.855 123.965 126.065 124.715 ;
        RECT 126.235 123.965 127.445 124.715 ;
        RECT 14.370 123.795 127.530 123.965 ;
        RECT 14.455 123.045 15.665 123.795 ;
        RECT 15.835 123.045 17.045 123.795 ;
        RECT 17.220 123.250 22.565 123.795 ;
        RECT 14.455 122.505 14.975 123.045 ;
        RECT 15.145 122.335 15.665 122.875 ;
        RECT 14.455 121.245 15.665 122.335 ;
        RECT 15.835 122.335 16.355 122.875 ;
        RECT 16.525 122.505 17.045 123.045 ;
        RECT 15.835 121.245 17.045 122.335 ;
        RECT 18.810 121.680 19.160 122.930 ;
        RECT 20.640 122.420 20.980 123.250 ;
        RECT 23.010 122.985 23.255 123.590 ;
        RECT 23.475 123.260 23.985 123.795 ;
        RECT 22.735 122.815 23.965 122.985 ;
        RECT 22.735 122.005 23.075 122.815 ;
        RECT 23.245 122.250 23.995 122.440 ;
        RECT 17.220 121.245 22.565 121.680 ;
        RECT 22.735 121.595 23.250 122.005 ;
        RECT 23.485 121.245 23.655 122.005 ;
        RECT 23.825 121.585 23.995 122.250 ;
        RECT 24.165 122.265 24.355 123.625 ;
        RECT 24.525 123.455 24.800 123.625 ;
        RECT 24.525 123.285 24.805 123.455 ;
        RECT 24.525 122.465 24.800 123.285 ;
        RECT 24.990 123.260 25.520 123.625 ;
        RECT 25.945 123.395 26.275 123.795 ;
        RECT 25.345 123.225 25.520 123.260 ;
        RECT 25.005 122.265 25.175 123.065 ;
        RECT 24.165 122.095 25.175 122.265 ;
        RECT 25.345 123.055 26.275 123.225 ;
        RECT 26.445 123.055 26.700 123.625 ;
        RECT 27.340 123.250 32.685 123.795 ;
        RECT 25.345 121.925 25.515 123.055 ;
        RECT 26.105 122.885 26.275 123.055 ;
        RECT 24.390 121.755 25.515 121.925 ;
        RECT 25.685 122.555 25.880 122.885 ;
        RECT 26.105 122.555 26.360 122.885 ;
        RECT 25.685 121.585 25.855 122.555 ;
        RECT 26.530 122.385 26.700 123.055 ;
        RECT 23.825 121.415 25.855 121.585 ;
        RECT 26.025 121.245 26.195 122.385 ;
        RECT 26.365 121.415 26.700 122.385 ;
        RECT 28.930 121.680 29.280 122.930 ;
        RECT 30.760 122.420 31.100 123.250 ;
        RECT 33.130 122.985 33.375 123.590 ;
        RECT 33.595 123.260 34.105 123.795 ;
        RECT 32.855 122.815 34.085 122.985 ;
        RECT 32.855 122.005 33.195 122.815 ;
        RECT 33.365 122.250 34.115 122.440 ;
        RECT 27.340 121.245 32.685 121.680 ;
        RECT 32.855 121.595 33.370 122.005 ;
        RECT 33.605 121.245 33.775 122.005 ;
        RECT 33.945 121.585 34.115 122.250 ;
        RECT 34.285 122.265 34.475 123.625 ;
        RECT 34.645 122.775 34.920 123.625 ;
        RECT 35.110 123.260 35.640 123.625 ;
        RECT 36.065 123.395 36.395 123.795 ;
        RECT 35.465 123.225 35.640 123.260 ;
        RECT 34.645 122.605 34.925 122.775 ;
        RECT 34.645 122.465 34.920 122.605 ;
        RECT 35.125 122.265 35.295 123.065 ;
        RECT 34.285 122.095 35.295 122.265 ;
        RECT 35.465 123.055 36.395 123.225 ;
        RECT 36.565 123.055 36.820 123.625 ;
        RECT 36.995 123.070 37.285 123.795 ;
        RECT 35.465 121.925 35.635 123.055 ;
        RECT 36.225 122.885 36.395 123.055 ;
        RECT 34.510 121.755 35.635 121.925 ;
        RECT 35.805 122.555 36.000 122.885 ;
        RECT 36.225 122.555 36.480 122.885 ;
        RECT 35.805 121.585 35.975 122.555 ;
        RECT 36.650 122.385 36.820 123.055 ;
        RECT 37.915 123.025 41.425 123.795 ;
        RECT 41.600 123.250 46.945 123.795 ;
        RECT 47.120 123.250 52.465 123.795 ;
        RECT 53.010 123.455 53.265 123.615 ;
        RECT 52.925 123.285 53.265 123.455 ;
        RECT 53.445 123.335 53.730 123.795 ;
        RECT 33.945 121.415 35.975 121.585 ;
        RECT 36.145 121.245 36.315 122.385 ;
        RECT 36.485 121.415 36.820 122.385 ;
        RECT 36.995 121.245 37.285 122.410 ;
        RECT 37.915 122.335 39.605 122.855 ;
        RECT 39.775 122.505 41.425 123.025 ;
        RECT 37.915 121.245 41.425 122.335 ;
        RECT 43.190 121.680 43.540 122.930 ;
        RECT 45.020 122.420 45.360 123.250 ;
        RECT 48.710 121.680 49.060 122.930 ;
        RECT 50.540 122.420 50.880 123.250 ;
        RECT 53.010 123.085 53.265 123.285 ;
        RECT 53.010 122.225 53.190 123.085 ;
        RECT 53.910 122.885 54.160 123.535 ;
        RECT 53.360 122.555 54.160 122.885 ;
        RECT 41.600 121.245 46.945 121.680 ;
        RECT 47.120 121.245 52.465 121.680 ;
        RECT 53.010 121.555 53.265 122.225 ;
        RECT 53.445 121.245 53.730 122.045 ;
        RECT 53.910 121.965 54.160 122.555 ;
        RECT 54.360 123.200 54.680 123.530 ;
        RECT 54.860 123.315 55.520 123.795 ;
        RECT 55.720 123.405 56.570 123.575 ;
        RECT 54.360 122.305 54.550 123.200 ;
        RECT 54.870 122.875 55.530 123.145 ;
        RECT 55.200 122.815 55.530 122.875 ;
        RECT 54.720 122.645 55.050 122.705 ;
        RECT 55.720 122.645 55.890 123.405 ;
        RECT 57.130 123.335 57.450 123.795 ;
        RECT 57.650 123.155 57.900 123.585 ;
        RECT 58.190 123.355 58.600 123.795 ;
        RECT 58.770 123.415 59.785 123.615 ;
        RECT 56.060 122.985 57.310 123.155 ;
        RECT 56.060 122.865 56.390 122.985 ;
        RECT 54.720 122.475 56.620 122.645 ;
        RECT 54.360 122.135 56.280 122.305 ;
        RECT 54.360 122.115 54.680 122.135 ;
        RECT 53.910 121.455 54.240 121.965 ;
        RECT 54.510 121.505 54.680 122.115 ;
        RECT 56.450 121.965 56.620 122.475 ;
        RECT 56.790 122.405 56.970 122.815 ;
        RECT 57.140 122.225 57.310 122.985 ;
        RECT 54.850 121.245 55.180 121.935 ;
        RECT 55.410 121.795 56.620 121.965 ;
        RECT 56.790 121.915 57.310 122.225 ;
        RECT 57.480 122.815 57.900 123.155 ;
        RECT 58.190 122.815 58.600 123.145 ;
        RECT 57.480 122.045 57.670 122.815 ;
        RECT 58.770 122.685 58.940 123.415 ;
        RECT 60.085 123.245 60.255 123.575 ;
        RECT 60.425 123.415 60.755 123.795 ;
        RECT 59.110 122.865 59.460 123.235 ;
        RECT 58.770 122.645 59.190 122.685 ;
        RECT 57.840 122.475 59.190 122.645 ;
        RECT 57.840 122.315 58.090 122.475 ;
        RECT 58.600 122.045 58.850 122.305 ;
        RECT 57.480 121.795 58.850 122.045 ;
        RECT 55.410 121.505 55.650 121.795 ;
        RECT 56.450 121.715 56.620 121.795 ;
        RECT 55.850 121.245 56.270 121.625 ;
        RECT 56.450 121.465 57.080 121.715 ;
        RECT 57.550 121.245 57.880 121.625 ;
        RECT 58.050 121.505 58.220 121.795 ;
        RECT 59.020 121.630 59.190 122.475 ;
        RECT 59.640 122.305 59.860 123.175 ;
        RECT 60.085 123.055 60.780 123.245 ;
        RECT 59.360 121.925 59.860 122.305 ;
        RECT 60.030 122.255 60.440 122.875 ;
        RECT 60.610 122.085 60.780 123.055 ;
        RECT 60.085 121.915 60.780 122.085 ;
        RECT 58.400 121.245 58.780 121.625 ;
        RECT 59.020 121.460 59.850 121.630 ;
        RECT 60.085 121.415 60.255 121.915 ;
        RECT 60.425 121.245 60.755 121.745 ;
        RECT 60.970 121.415 61.195 123.535 ;
        RECT 61.365 123.415 61.695 123.795 ;
        RECT 61.865 123.245 62.035 123.535 ;
        RECT 61.370 123.075 62.035 123.245 ;
        RECT 61.370 122.085 61.600 123.075 ;
        RECT 62.755 123.070 63.045 123.795 ;
        RECT 63.950 122.985 64.195 123.590 ;
        RECT 64.415 123.260 64.925 123.795 ;
        RECT 61.770 122.255 62.120 122.905 ;
        RECT 63.675 122.815 64.905 122.985 ;
        RECT 61.370 121.915 62.035 122.085 ;
        RECT 61.365 121.245 61.695 121.745 ;
        RECT 61.865 121.415 62.035 121.915 ;
        RECT 62.755 121.245 63.045 122.410 ;
        RECT 63.675 122.005 64.015 122.815 ;
        RECT 64.185 122.250 64.935 122.440 ;
        RECT 63.675 121.595 64.190 122.005 ;
        RECT 64.425 121.245 64.595 122.005 ;
        RECT 64.765 121.585 64.935 122.250 ;
        RECT 65.105 122.265 65.295 123.625 ;
        RECT 65.465 123.455 65.740 123.625 ;
        RECT 65.465 123.285 65.745 123.455 ;
        RECT 65.465 122.465 65.740 123.285 ;
        RECT 65.930 123.260 66.460 123.625 ;
        RECT 66.885 123.395 67.215 123.795 ;
        RECT 66.285 123.225 66.460 123.260 ;
        RECT 65.945 122.265 66.115 123.065 ;
        RECT 65.105 122.095 66.115 122.265 ;
        RECT 66.285 123.055 67.215 123.225 ;
        RECT 67.385 123.055 67.640 123.625 ;
        RECT 66.285 121.925 66.455 123.055 ;
        RECT 67.045 122.885 67.215 123.055 ;
        RECT 65.330 121.755 66.455 121.925 ;
        RECT 66.625 122.555 66.820 122.885 ;
        RECT 67.045 122.555 67.300 122.885 ;
        RECT 66.625 121.585 66.795 122.555 ;
        RECT 67.470 122.385 67.640 123.055 ;
        RECT 67.815 123.025 70.405 123.795 ;
        RECT 70.580 123.250 75.925 123.795 ;
        RECT 76.100 123.250 81.445 123.795 ;
        RECT 64.765 121.415 66.795 121.585 ;
        RECT 66.965 121.245 67.135 122.385 ;
        RECT 67.305 121.415 67.640 122.385 ;
        RECT 67.815 122.335 69.025 122.855 ;
        RECT 69.195 122.505 70.405 123.025 ;
        RECT 67.815 121.245 70.405 122.335 ;
        RECT 72.170 121.680 72.520 122.930 ;
        RECT 74.000 122.420 74.340 123.250 ;
        RECT 77.690 121.680 78.040 122.930 ;
        RECT 79.520 122.420 79.860 123.250 ;
        RECT 81.675 122.975 81.885 123.795 ;
        RECT 82.055 122.995 82.385 123.625 ;
        RECT 82.055 122.395 82.305 122.995 ;
        RECT 82.555 122.975 82.785 123.795 ;
        RECT 83.545 123.245 83.715 123.625 ;
        RECT 83.895 123.415 84.225 123.795 ;
        RECT 83.545 123.075 84.210 123.245 ;
        RECT 84.405 123.120 84.665 123.625 ;
        RECT 82.475 122.555 82.805 122.805 ;
        RECT 83.475 122.525 83.805 122.895 ;
        RECT 84.040 122.820 84.210 123.075 ;
        RECT 84.040 122.490 84.325 122.820 ;
        RECT 70.580 121.245 75.925 121.680 ;
        RECT 76.100 121.245 81.445 121.680 ;
        RECT 81.675 121.245 81.885 122.385 ;
        RECT 82.055 121.415 82.385 122.395 ;
        RECT 82.555 121.245 82.785 122.385 ;
        RECT 84.040 122.345 84.210 122.490 ;
        RECT 83.545 122.175 84.210 122.345 ;
        RECT 84.495 122.320 84.665 123.120 ;
        RECT 84.835 123.025 88.345 123.795 ;
        RECT 88.515 123.070 88.805 123.795 ;
        RECT 88.975 123.025 92.485 123.795 ;
        RECT 83.545 121.415 83.715 122.175 ;
        RECT 83.895 121.245 84.225 122.005 ;
        RECT 84.395 121.415 84.665 122.320 ;
        RECT 84.835 122.335 86.525 122.855 ;
        RECT 86.695 122.505 88.345 123.025 ;
        RECT 84.835 121.245 88.345 122.335 ;
        RECT 88.515 121.245 88.805 122.410 ;
        RECT 88.975 122.335 90.665 122.855 ;
        RECT 90.835 122.505 92.485 123.025 ;
        RECT 92.695 122.975 92.925 123.795 ;
        RECT 93.095 122.995 93.425 123.625 ;
        RECT 92.675 122.555 93.005 122.805 ;
        RECT 93.175 122.395 93.425 122.995 ;
        RECT 93.595 122.975 93.805 123.795 ;
        RECT 94.035 123.045 95.245 123.795 ;
        RECT 88.975 121.245 92.485 122.335 ;
        RECT 92.695 121.245 92.925 122.385 ;
        RECT 93.095 121.415 93.425 122.395 ;
        RECT 93.595 121.245 93.805 122.385 ;
        RECT 94.035 122.335 94.555 122.875 ;
        RECT 94.725 122.505 95.245 123.045 ;
        RECT 95.415 123.025 98.925 123.795 ;
        RECT 99.100 123.250 104.445 123.795 ;
        RECT 104.620 123.250 109.965 123.795 ;
        RECT 95.415 122.335 97.105 122.855 ;
        RECT 97.275 122.505 98.925 123.025 ;
        RECT 94.035 121.245 95.245 122.335 ;
        RECT 95.415 121.245 98.925 122.335 ;
        RECT 100.690 121.680 101.040 122.930 ;
        RECT 102.520 122.420 102.860 123.250 ;
        RECT 106.210 121.680 106.560 122.930 ;
        RECT 108.040 122.420 108.380 123.250 ;
        RECT 110.410 122.985 110.655 123.590 ;
        RECT 110.875 123.260 111.385 123.795 ;
        RECT 110.135 122.815 111.365 122.985 ;
        RECT 110.135 122.005 110.475 122.815 ;
        RECT 110.645 122.250 111.395 122.440 ;
        RECT 99.100 121.245 104.445 121.680 ;
        RECT 104.620 121.245 109.965 121.680 ;
        RECT 110.135 121.595 110.650 122.005 ;
        RECT 110.885 121.245 111.055 122.005 ;
        RECT 111.225 121.585 111.395 122.250 ;
        RECT 111.565 122.265 111.755 123.625 ;
        RECT 111.925 122.775 112.200 123.625 ;
        RECT 112.390 123.260 112.920 123.625 ;
        RECT 113.345 123.395 113.675 123.795 ;
        RECT 112.745 123.225 112.920 123.260 ;
        RECT 111.925 122.605 112.205 122.775 ;
        RECT 111.925 122.465 112.200 122.605 ;
        RECT 112.405 122.265 112.575 123.065 ;
        RECT 111.565 122.095 112.575 122.265 ;
        RECT 112.745 123.055 113.675 123.225 ;
        RECT 113.845 123.055 114.100 123.625 ;
        RECT 114.275 123.070 114.565 123.795 ;
        RECT 115.570 123.085 115.825 123.615 ;
        RECT 116.005 123.335 116.290 123.795 ;
        RECT 112.745 121.925 112.915 123.055 ;
        RECT 113.505 122.885 113.675 123.055 ;
        RECT 111.790 121.755 112.915 121.925 ;
        RECT 113.085 122.555 113.280 122.885 ;
        RECT 113.505 122.555 113.760 122.885 ;
        RECT 113.085 121.585 113.255 122.555 ;
        RECT 113.930 122.385 114.100 123.055 ;
        RECT 115.570 122.775 115.750 123.085 ;
        RECT 116.470 122.885 116.720 123.535 ;
        RECT 115.485 122.605 115.750 122.775 ;
        RECT 111.225 121.415 113.255 121.585 ;
        RECT 113.425 121.245 113.595 122.385 ;
        RECT 113.765 121.415 114.100 122.385 ;
        RECT 114.275 121.245 114.565 122.410 ;
        RECT 115.570 122.225 115.750 122.605 ;
        RECT 115.920 122.555 116.720 122.885 ;
        RECT 115.570 121.555 115.825 122.225 ;
        RECT 116.005 121.245 116.290 122.045 ;
        RECT 116.470 121.965 116.720 122.555 ;
        RECT 116.920 123.200 117.240 123.530 ;
        RECT 117.420 123.315 118.080 123.795 ;
        RECT 118.280 123.405 119.130 123.575 ;
        RECT 116.920 122.305 117.110 123.200 ;
        RECT 117.430 122.875 118.090 123.145 ;
        RECT 117.760 122.815 118.090 122.875 ;
        RECT 117.280 122.645 117.610 122.705 ;
        RECT 118.280 122.645 118.450 123.405 ;
        RECT 119.690 123.335 120.010 123.795 ;
        RECT 120.210 123.155 120.460 123.585 ;
        RECT 120.750 123.355 121.160 123.795 ;
        RECT 121.330 123.415 122.345 123.615 ;
        RECT 118.620 122.985 119.870 123.155 ;
        RECT 118.620 122.865 118.950 122.985 ;
        RECT 117.280 122.475 119.180 122.645 ;
        RECT 116.920 122.135 118.840 122.305 ;
        RECT 116.920 122.115 117.240 122.135 ;
        RECT 116.470 121.455 116.800 121.965 ;
        RECT 117.070 121.505 117.240 122.115 ;
        RECT 119.010 121.965 119.180 122.475 ;
        RECT 119.350 122.405 119.530 122.815 ;
        RECT 119.700 122.225 119.870 122.985 ;
        RECT 117.410 121.245 117.740 121.935 ;
        RECT 117.970 121.795 119.180 121.965 ;
        RECT 119.350 121.915 119.870 122.225 ;
        RECT 120.040 122.815 120.460 123.155 ;
        RECT 120.750 122.815 121.160 123.145 ;
        RECT 120.040 122.045 120.230 122.815 ;
        RECT 121.330 122.685 121.500 123.415 ;
        RECT 122.645 123.245 122.815 123.575 ;
        RECT 122.985 123.415 123.315 123.795 ;
        RECT 121.670 122.865 122.020 123.235 ;
        RECT 121.330 122.645 121.750 122.685 ;
        RECT 120.400 122.475 121.750 122.645 ;
        RECT 120.400 122.315 120.650 122.475 ;
        RECT 121.160 122.045 121.410 122.305 ;
        RECT 120.040 121.795 121.410 122.045 ;
        RECT 117.970 121.505 118.210 121.795 ;
        RECT 119.010 121.715 119.180 121.795 ;
        RECT 118.410 121.245 118.830 121.625 ;
        RECT 119.010 121.465 119.640 121.715 ;
        RECT 120.110 121.245 120.440 121.625 ;
        RECT 120.610 121.505 120.780 121.795 ;
        RECT 121.580 121.630 121.750 122.475 ;
        RECT 122.200 122.305 122.420 123.175 ;
        RECT 122.645 123.055 123.340 123.245 ;
        RECT 121.920 121.925 122.420 122.305 ;
        RECT 122.590 122.255 123.000 122.875 ;
        RECT 123.170 122.085 123.340 123.055 ;
        RECT 122.645 121.915 123.340 122.085 ;
        RECT 120.960 121.245 121.340 121.625 ;
        RECT 121.580 121.460 122.410 121.630 ;
        RECT 122.645 121.415 122.815 121.915 ;
        RECT 122.985 121.245 123.315 121.745 ;
        RECT 123.530 121.415 123.755 123.535 ;
        RECT 123.925 123.415 124.255 123.795 ;
        RECT 124.425 123.245 124.595 123.535 ;
        RECT 123.930 123.075 124.595 123.245 ;
        RECT 123.930 122.085 124.160 123.075 ;
        RECT 124.855 123.045 126.065 123.795 ;
        RECT 126.235 123.045 127.445 123.795 ;
        RECT 124.330 122.255 124.680 122.905 ;
        RECT 124.855 122.335 125.375 122.875 ;
        RECT 125.545 122.505 126.065 123.045 ;
        RECT 126.235 122.335 126.755 122.875 ;
        RECT 126.925 122.505 127.445 123.045 ;
        RECT 123.930 121.915 124.595 122.085 ;
        RECT 123.925 121.245 124.255 121.745 ;
        RECT 124.425 121.415 124.595 121.915 ;
        RECT 124.855 121.245 126.065 122.335 ;
        RECT 126.235 121.245 127.445 122.335 ;
        RECT 14.370 121.075 127.530 121.245 ;
        RECT 14.455 119.985 15.665 121.075 ;
        RECT 14.455 119.275 14.975 119.815 ;
        RECT 15.145 119.445 15.665 119.985 ;
        RECT 16.295 119.985 19.805 121.075 ;
        RECT 16.295 119.465 17.985 119.985 ;
        RECT 19.980 119.935 20.315 120.905 ;
        RECT 20.485 119.935 20.655 121.075 ;
        RECT 20.825 120.735 22.855 120.905 ;
        RECT 18.155 119.295 19.805 119.815 ;
        RECT 14.455 118.525 15.665 119.275 ;
        RECT 16.295 118.525 19.805 119.295 ;
        RECT 19.980 119.265 20.150 119.935 ;
        RECT 20.825 119.765 20.995 120.735 ;
        RECT 20.320 119.435 20.575 119.765 ;
        RECT 20.800 119.435 20.995 119.765 ;
        RECT 21.165 120.395 22.290 120.565 ;
        RECT 20.405 119.265 20.575 119.435 ;
        RECT 21.165 119.265 21.335 120.395 ;
        RECT 19.980 118.695 20.235 119.265 ;
        RECT 20.405 119.095 21.335 119.265 ;
        RECT 21.505 120.055 22.515 120.225 ;
        RECT 21.505 119.255 21.675 120.055 ;
        RECT 21.880 119.375 22.155 119.855 ;
        RECT 21.875 119.205 22.155 119.375 ;
        RECT 21.160 119.060 21.335 119.095 ;
        RECT 20.405 118.525 20.735 118.925 ;
        RECT 21.160 118.695 21.690 119.060 ;
        RECT 21.880 118.695 22.155 119.205 ;
        RECT 22.325 118.695 22.515 120.055 ;
        RECT 22.685 120.070 22.855 120.735 ;
        RECT 23.025 120.315 23.195 121.075 ;
        RECT 23.430 120.315 23.945 120.725 ;
        RECT 22.685 119.880 23.435 120.070 ;
        RECT 23.605 119.505 23.945 120.315 ;
        RECT 24.115 119.910 24.405 121.075 ;
        RECT 24.575 119.985 25.785 121.075 ;
        RECT 25.955 120.000 26.225 120.905 ;
        RECT 26.395 120.315 26.725 121.075 ;
        RECT 26.905 120.145 27.075 120.905 ;
        RECT 22.715 119.335 23.945 119.505 ;
        RECT 24.575 119.445 25.095 119.985 ;
        RECT 22.695 118.525 23.205 119.060 ;
        RECT 23.425 118.730 23.670 119.335 ;
        RECT 25.265 119.275 25.785 119.815 ;
        RECT 24.115 118.525 24.405 119.250 ;
        RECT 24.575 118.525 25.785 119.275 ;
        RECT 25.955 119.200 26.125 120.000 ;
        RECT 26.410 119.975 27.075 120.145 ;
        RECT 27.335 119.985 29.925 121.075 ;
        RECT 30.470 120.735 30.725 120.765 ;
        RECT 30.385 120.565 30.725 120.735 ;
        RECT 30.470 120.095 30.725 120.565 ;
        RECT 30.905 120.275 31.190 121.075 ;
        RECT 31.370 120.355 31.700 120.865 ;
        RECT 26.410 119.830 26.580 119.975 ;
        RECT 26.295 119.500 26.580 119.830 ;
        RECT 26.410 119.245 26.580 119.500 ;
        RECT 26.815 119.425 27.145 119.795 ;
        RECT 27.335 119.465 28.545 119.985 ;
        RECT 28.715 119.295 29.925 119.815 ;
        RECT 25.955 118.695 26.215 119.200 ;
        RECT 26.410 119.075 27.075 119.245 ;
        RECT 26.395 118.525 26.725 118.905 ;
        RECT 26.905 118.695 27.075 119.075 ;
        RECT 27.335 118.525 29.925 119.295 ;
        RECT 30.470 119.235 30.650 120.095 ;
        RECT 31.370 119.765 31.620 120.355 ;
        RECT 31.970 120.205 32.140 120.815 ;
        RECT 32.310 120.385 32.640 121.075 ;
        RECT 32.870 120.525 33.110 120.815 ;
        RECT 33.310 120.695 33.730 121.075 ;
        RECT 33.910 120.605 34.540 120.855 ;
        RECT 35.010 120.695 35.340 121.075 ;
        RECT 33.910 120.525 34.080 120.605 ;
        RECT 35.510 120.525 35.680 120.815 ;
        RECT 35.860 120.695 36.240 121.075 ;
        RECT 36.480 120.690 37.310 120.860 ;
        RECT 32.870 120.355 34.080 120.525 ;
        RECT 30.820 119.435 31.620 119.765 ;
        RECT 30.470 118.705 30.725 119.235 ;
        RECT 30.905 118.525 31.190 118.985 ;
        RECT 31.370 118.785 31.620 119.435 ;
        RECT 31.820 120.185 32.140 120.205 ;
        RECT 31.820 120.015 33.740 120.185 ;
        RECT 31.820 119.120 32.010 120.015 ;
        RECT 33.910 119.845 34.080 120.355 ;
        RECT 34.250 120.095 34.770 120.405 ;
        RECT 32.180 119.675 34.080 119.845 ;
        RECT 32.180 119.615 32.510 119.675 ;
        RECT 32.660 119.445 32.990 119.505 ;
        RECT 32.330 119.175 32.990 119.445 ;
        RECT 31.820 118.790 32.140 119.120 ;
        RECT 32.320 118.525 32.980 119.005 ;
        RECT 33.180 118.915 33.350 119.675 ;
        RECT 34.250 119.505 34.430 119.915 ;
        RECT 33.520 119.335 33.850 119.455 ;
        RECT 34.600 119.335 34.770 120.095 ;
        RECT 33.520 119.165 34.770 119.335 ;
        RECT 34.940 120.275 36.310 120.525 ;
        RECT 34.940 119.505 35.130 120.275 ;
        RECT 36.060 120.015 36.310 120.275 ;
        RECT 35.300 119.845 35.550 120.005 ;
        RECT 36.480 119.845 36.650 120.690 ;
        RECT 37.545 120.405 37.715 120.905 ;
        RECT 37.885 120.575 38.215 121.075 ;
        RECT 36.820 120.015 37.320 120.395 ;
        RECT 37.545 120.235 38.240 120.405 ;
        RECT 35.300 119.675 36.650 119.845 ;
        RECT 36.230 119.635 36.650 119.675 ;
        RECT 34.940 119.165 35.360 119.505 ;
        RECT 35.650 119.175 36.060 119.505 ;
        RECT 33.180 118.745 34.030 118.915 ;
        RECT 34.590 118.525 34.910 118.985 ;
        RECT 35.110 118.735 35.360 119.165 ;
        RECT 35.650 118.525 36.060 118.965 ;
        RECT 36.230 118.905 36.400 119.635 ;
        RECT 36.570 119.085 36.920 119.455 ;
        RECT 37.100 119.145 37.320 120.015 ;
        RECT 37.490 119.445 37.900 120.065 ;
        RECT 38.070 119.265 38.240 120.235 ;
        RECT 37.545 119.075 38.240 119.265 ;
        RECT 36.230 118.705 37.245 118.905 ;
        RECT 37.545 118.745 37.715 119.075 ;
        RECT 37.885 118.525 38.215 118.905 ;
        RECT 38.430 118.785 38.655 120.905 ;
        RECT 38.825 120.575 39.155 121.075 ;
        RECT 39.325 120.405 39.495 120.905 ;
        RECT 38.830 120.235 39.495 120.405 ;
        RECT 38.830 119.245 39.060 120.235 ;
        RECT 39.230 119.415 39.580 120.065 ;
        RECT 39.760 119.935 40.095 120.905 ;
        RECT 40.265 119.935 40.435 121.075 ;
        RECT 40.605 120.735 42.635 120.905 ;
        RECT 39.760 119.265 39.930 119.935 ;
        RECT 40.605 119.765 40.775 120.735 ;
        RECT 40.100 119.435 40.355 119.765 ;
        RECT 40.580 119.435 40.775 119.765 ;
        RECT 40.945 120.395 42.070 120.565 ;
        RECT 40.185 119.265 40.355 119.435 ;
        RECT 40.945 119.265 41.115 120.395 ;
        RECT 38.830 119.075 39.495 119.245 ;
        RECT 38.825 118.525 39.155 118.905 ;
        RECT 39.325 118.785 39.495 119.075 ;
        RECT 39.760 118.695 40.015 119.265 ;
        RECT 40.185 119.095 41.115 119.265 ;
        RECT 41.285 120.055 42.295 120.225 ;
        RECT 41.285 119.255 41.455 120.055 ;
        RECT 41.660 119.715 41.935 119.855 ;
        RECT 41.655 119.545 41.935 119.715 ;
        RECT 40.940 119.060 41.115 119.095 ;
        RECT 40.185 118.525 40.515 118.925 ;
        RECT 40.940 118.695 41.470 119.060 ;
        RECT 41.660 118.695 41.935 119.545 ;
        RECT 42.105 118.695 42.295 120.055 ;
        RECT 42.465 120.070 42.635 120.735 ;
        RECT 42.805 120.315 42.975 121.075 ;
        RECT 43.210 120.315 43.725 120.725 ;
        RECT 42.465 119.880 43.215 120.070 ;
        RECT 43.385 119.505 43.725 120.315 ;
        RECT 42.495 119.335 43.725 119.505 ;
        RECT 44.355 120.000 44.625 120.905 ;
        RECT 44.795 120.315 45.125 121.075 ;
        RECT 45.305 120.145 45.475 120.905 ;
        RECT 42.475 118.525 42.985 119.060 ;
        RECT 43.205 118.730 43.450 119.335 ;
        RECT 44.355 119.200 44.525 120.000 ;
        RECT 44.810 119.975 45.475 120.145 ;
        RECT 45.735 120.315 46.250 120.725 ;
        RECT 46.485 120.315 46.655 121.075 ;
        RECT 46.825 120.735 48.855 120.905 ;
        RECT 44.810 119.830 44.980 119.975 ;
        RECT 44.695 119.500 44.980 119.830 ;
        RECT 44.810 119.245 44.980 119.500 ;
        RECT 45.215 119.425 45.545 119.795 ;
        RECT 45.735 119.505 46.075 120.315 ;
        RECT 46.825 120.070 46.995 120.735 ;
        RECT 47.390 120.395 48.515 120.565 ;
        RECT 46.245 119.880 46.995 120.070 ;
        RECT 47.165 120.055 48.175 120.225 ;
        RECT 45.735 119.335 46.965 119.505 ;
        RECT 44.355 118.695 44.615 119.200 ;
        RECT 44.810 119.075 45.475 119.245 ;
        RECT 44.795 118.525 45.125 118.905 ;
        RECT 45.305 118.695 45.475 119.075 ;
        RECT 46.010 118.730 46.255 119.335 ;
        RECT 46.475 118.525 46.985 119.060 ;
        RECT 47.165 118.695 47.355 120.055 ;
        RECT 47.525 119.715 47.800 119.855 ;
        RECT 47.525 119.545 47.805 119.715 ;
        RECT 47.525 118.695 47.800 119.545 ;
        RECT 48.005 119.255 48.175 120.055 ;
        RECT 48.345 119.265 48.515 120.395 ;
        RECT 48.685 119.765 48.855 120.735 ;
        RECT 49.025 119.935 49.195 121.075 ;
        RECT 49.365 119.935 49.700 120.905 ;
        RECT 48.685 119.435 48.880 119.765 ;
        RECT 49.105 119.435 49.360 119.765 ;
        RECT 49.105 119.265 49.275 119.435 ;
        RECT 49.530 119.265 49.700 119.935 ;
        RECT 49.875 119.910 50.165 121.075 ;
        RECT 50.375 119.935 50.605 121.075 ;
        RECT 50.775 119.925 51.105 120.905 ;
        RECT 51.275 119.935 51.485 121.075 ;
        RECT 51.715 119.985 52.925 121.075 ;
        RECT 50.355 119.515 50.685 119.765 ;
        RECT 48.345 119.095 49.275 119.265 ;
        RECT 48.345 119.060 48.520 119.095 ;
        RECT 47.990 118.695 48.520 119.060 ;
        RECT 48.945 118.525 49.275 118.925 ;
        RECT 49.445 118.695 49.700 119.265 ;
        RECT 49.875 118.525 50.165 119.250 ;
        RECT 50.375 118.525 50.605 119.345 ;
        RECT 50.855 119.325 51.105 119.925 ;
        RECT 51.715 119.445 52.235 119.985 ;
        RECT 53.245 119.925 53.575 121.075 ;
        RECT 53.745 120.055 53.915 120.905 ;
        RECT 54.085 120.275 54.415 121.075 ;
        RECT 54.585 120.055 54.755 120.905 ;
        RECT 54.935 120.275 55.175 121.075 ;
        RECT 55.345 120.095 55.675 120.905 ;
        RECT 53.745 119.885 54.755 120.055 ;
        RECT 54.960 119.925 55.675 120.095 ;
        RECT 56.835 119.935 57.045 121.075 ;
        RECT 57.215 119.925 57.545 120.905 ;
        RECT 57.715 119.935 57.945 121.075 ;
        RECT 59.450 120.735 59.705 120.765 ;
        RECT 59.365 120.565 59.705 120.735 ;
        RECT 59.450 120.095 59.705 120.565 ;
        RECT 59.885 120.275 60.170 121.075 ;
        RECT 60.350 120.355 60.680 120.865 ;
        RECT 50.775 118.695 51.105 119.325 ;
        RECT 51.275 118.525 51.485 119.345 ;
        RECT 52.405 119.275 52.925 119.815 ;
        RECT 53.745 119.715 54.240 119.885 ;
        RECT 53.745 119.545 54.245 119.715 ;
        RECT 54.960 119.685 55.130 119.925 ;
        RECT 53.745 119.345 54.240 119.545 ;
        RECT 54.630 119.515 55.130 119.685 ;
        RECT 55.300 119.515 55.680 119.755 ;
        RECT 54.960 119.345 55.130 119.515 ;
        RECT 51.715 118.525 52.925 119.275 ;
        RECT 53.245 118.525 53.575 119.325 ;
        RECT 53.745 119.175 54.755 119.345 ;
        RECT 54.960 119.175 55.595 119.345 ;
        RECT 53.745 118.695 53.915 119.175 ;
        RECT 54.085 118.525 54.415 119.005 ;
        RECT 54.585 118.695 54.755 119.175 ;
        RECT 55.005 118.525 55.245 119.005 ;
        RECT 55.425 118.695 55.595 119.175 ;
        RECT 56.835 118.525 57.045 119.345 ;
        RECT 57.215 119.325 57.465 119.925 ;
        RECT 57.635 119.515 57.965 119.765 ;
        RECT 57.215 118.695 57.545 119.325 ;
        RECT 57.715 118.525 57.945 119.345 ;
        RECT 59.450 119.235 59.630 120.095 ;
        RECT 60.350 119.765 60.600 120.355 ;
        RECT 60.950 120.205 61.120 120.815 ;
        RECT 61.290 120.385 61.620 121.075 ;
        RECT 61.850 120.525 62.090 120.815 ;
        RECT 62.290 120.695 62.710 121.075 ;
        RECT 62.890 120.605 63.520 120.855 ;
        RECT 63.990 120.695 64.320 121.075 ;
        RECT 62.890 120.525 63.060 120.605 ;
        RECT 64.490 120.525 64.660 120.815 ;
        RECT 64.840 120.695 65.220 121.075 ;
        RECT 65.460 120.690 66.290 120.860 ;
        RECT 61.850 120.355 63.060 120.525 ;
        RECT 59.800 119.435 60.600 119.765 ;
        RECT 59.450 118.705 59.705 119.235 ;
        RECT 59.885 118.525 60.170 118.985 ;
        RECT 60.350 118.785 60.600 119.435 ;
        RECT 60.800 120.185 61.120 120.205 ;
        RECT 60.800 120.015 62.720 120.185 ;
        RECT 60.800 119.120 60.990 120.015 ;
        RECT 62.890 119.845 63.060 120.355 ;
        RECT 63.230 120.095 63.750 120.405 ;
        RECT 61.160 119.675 63.060 119.845 ;
        RECT 61.160 119.615 61.490 119.675 ;
        RECT 61.640 119.445 61.970 119.505 ;
        RECT 61.310 119.175 61.970 119.445 ;
        RECT 60.800 118.790 61.120 119.120 ;
        RECT 61.300 118.525 61.960 119.005 ;
        RECT 62.160 118.915 62.330 119.675 ;
        RECT 63.230 119.505 63.410 119.915 ;
        RECT 62.500 119.335 62.830 119.455 ;
        RECT 63.580 119.335 63.750 120.095 ;
        RECT 62.500 119.165 63.750 119.335 ;
        RECT 63.920 120.275 65.290 120.525 ;
        RECT 63.920 119.505 64.110 120.275 ;
        RECT 65.040 120.015 65.290 120.275 ;
        RECT 64.280 119.845 64.530 120.005 ;
        RECT 65.460 119.845 65.630 120.690 ;
        RECT 66.525 120.405 66.695 120.905 ;
        RECT 66.865 120.575 67.195 121.075 ;
        RECT 65.800 120.015 66.300 120.395 ;
        RECT 66.525 120.235 67.220 120.405 ;
        RECT 64.280 119.675 65.630 119.845 ;
        RECT 65.210 119.635 65.630 119.675 ;
        RECT 63.920 119.165 64.340 119.505 ;
        RECT 64.630 119.175 65.040 119.505 ;
        RECT 62.160 118.745 63.010 118.915 ;
        RECT 63.570 118.525 63.890 118.985 ;
        RECT 64.090 118.735 64.340 119.165 ;
        RECT 64.630 118.525 65.040 118.965 ;
        RECT 65.210 118.905 65.380 119.635 ;
        RECT 65.550 119.085 65.900 119.455 ;
        RECT 66.080 119.145 66.300 120.015 ;
        RECT 66.470 119.445 66.880 120.065 ;
        RECT 67.050 119.265 67.220 120.235 ;
        RECT 66.525 119.075 67.220 119.265 ;
        RECT 65.210 118.705 66.225 118.905 ;
        RECT 66.525 118.745 66.695 119.075 ;
        RECT 66.865 118.525 67.195 118.905 ;
        RECT 67.410 118.785 67.635 120.905 ;
        RECT 67.805 120.575 68.135 121.075 ;
        RECT 68.305 120.405 68.475 120.905 ;
        RECT 67.810 120.235 68.475 120.405 ;
        RECT 67.810 119.245 68.040 120.235 ;
        RECT 68.210 119.415 68.560 120.065 ;
        RECT 68.735 120.000 69.005 120.905 ;
        RECT 69.175 120.315 69.505 121.075 ;
        RECT 69.685 120.145 69.855 120.905 ;
        RECT 67.810 119.075 68.475 119.245 ;
        RECT 67.805 118.525 68.135 118.905 ;
        RECT 68.305 118.785 68.475 119.075 ;
        RECT 68.735 119.200 68.905 120.000 ;
        RECT 69.190 119.975 69.855 120.145 ;
        RECT 70.575 119.985 74.085 121.075 ;
        RECT 69.190 119.830 69.360 119.975 ;
        RECT 69.075 119.500 69.360 119.830 ;
        RECT 69.190 119.245 69.360 119.500 ;
        RECT 69.595 119.425 69.925 119.795 ;
        RECT 70.575 119.465 72.265 119.985 ;
        RECT 74.295 119.935 74.525 121.075 ;
        RECT 74.695 119.925 75.025 120.905 ;
        RECT 75.195 119.935 75.405 121.075 ;
        RECT 72.435 119.295 74.085 119.815 ;
        RECT 74.275 119.515 74.605 119.765 ;
        RECT 68.735 118.695 68.995 119.200 ;
        RECT 69.190 119.075 69.855 119.245 ;
        RECT 69.175 118.525 69.505 118.905 ;
        RECT 69.685 118.695 69.855 119.075 ;
        RECT 70.575 118.525 74.085 119.295 ;
        RECT 74.295 118.525 74.525 119.345 ;
        RECT 74.775 119.325 75.025 119.925 ;
        RECT 75.635 119.910 75.925 121.075 ;
        RECT 76.555 120.315 77.070 120.725 ;
        RECT 77.305 120.315 77.475 121.075 ;
        RECT 77.645 120.735 79.675 120.905 ;
        RECT 76.555 119.505 76.895 120.315 ;
        RECT 77.645 120.070 77.815 120.735 ;
        RECT 78.210 120.395 79.335 120.565 ;
        RECT 77.065 119.880 77.815 120.070 ;
        RECT 77.985 120.055 78.995 120.225 ;
        RECT 74.695 118.695 75.025 119.325 ;
        RECT 75.195 118.525 75.405 119.345 ;
        RECT 76.555 119.335 77.785 119.505 ;
        RECT 75.635 118.525 75.925 119.250 ;
        RECT 76.830 118.730 77.075 119.335 ;
        RECT 77.295 118.525 77.805 119.060 ;
        RECT 77.985 118.695 78.175 120.055 ;
        RECT 78.345 119.035 78.620 119.855 ;
        RECT 78.825 119.255 78.995 120.055 ;
        RECT 79.165 119.265 79.335 120.395 ;
        RECT 79.505 119.765 79.675 120.735 ;
        RECT 79.845 119.935 80.015 121.075 ;
        RECT 80.185 119.935 80.520 120.905 ;
        RECT 79.505 119.435 79.700 119.765 ;
        RECT 79.925 119.435 80.180 119.765 ;
        RECT 79.925 119.265 80.095 119.435 ;
        RECT 80.350 119.265 80.520 119.935 ;
        RECT 79.165 119.095 80.095 119.265 ;
        RECT 79.165 119.060 79.340 119.095 ;
        RECT 78.345 118.865 78.625 119.035 ;
        RECT 78.345 118.695 78.620 118.865 ;
        RECT 78.810 118.695 79.340 119.060 ;
        RECT 79.765 118.525 80.095 118.925 ;
        RECT 80.265 118.695 80.520 119.265 ;
        RECT 80.695 120.000 80.965 120.905 ;
        RECT 81.135 120.315 81.465 121.075 ;
        RECT 81.645 120.145 81.815 120.905 ;
        RECT 80.695 119.200 80.865 120.000 ;
        RECT 81.150 119.975 81.815 120.145 ;
        RECT 81.150 119.830 81.320 119.975 ;
        RECT 82.135 119.935 82.345 121.075 ;
        RECT 81.035 119.500 81.320 119.830 ;
        RECT 82.515 119.925 82.845 120.905 ;
        RECT 83.015 119.935 83.245 121.075 ;
        RECT 84.005 120.145 84.175 120.905 ;
        RECT 84.355 120.315 84.685 121.075 ;
        RECT 84.005 119.975 84.670 120.145 ;
        RECT 84.855 120.000 85.125 120.905 ;
        RECT 85.300 120.640 90.645 121.075 ;
        RECT 81.150 119.245 81.320 119.500 ;
        RECT 81.555 119.425 81.885 119.795 ;
        RECT 80.695 118.695 80.955 119.200 ;
        RECT 81.150 119.075 81.815 119.245 ;
        RECT 81.135 118.525 81.465 118.905 ;
        RECT 81.645 118.695 81.815 119.075 ;
        RECT 82.135 118.525 82.345 119.345 ;
        RECT 82.515 119.325 82.765 119.925 ;
        RECT 84.500 119.830 84.670 119.975 ;
        RECT 82.935 119.515 83.265 119.765 ;
        RECT 83.935 119.425 84.265 119.795 ;
        RECT 84.500 119.500 84.785 119.830 ;
        RECT 82.515 118.695 82.845 119.325 ;
        RECT 83.015 118.525 83.245 119.345 ;
        RECT 84.500 119.245 84.670 119.500 ;
        RECT 84.005 119.075 84.670 119.245 ;
        RECT 84.955 119.200 85.125 120.000 ;
        RECT 86.890 119.390 87.240 120.640 ;
        RECT 90.820 119.935 91.155 120.905 ;
        RECT 91.325 119.935 91.495 121.075 ;
        RECT 91.665 120.735 93.695 120.905 ;
        RECT 84.005 118.695 84.175 119.075 ;
        RECT 84.355 118.525 84.685 118.905 ;
        RECT 84.865 118.695 85.125 119.200 ;
        RECT 88.720 119.070 89.060 119.900 ;
        RECT 90.820 119.265 90.990 119.935 ;
        RECT 91.665 119.765 91.835 120.735 ;
        RECT 91.160 119.435 91.415 119.765 ;
        RECT 91.640 119.435 91.835 119.765 ;
        RECT 92.005 120.395 93.130 120.565 ;
        RECT 91.245 119.265 91.415 119.435 ;
        RECT 92.005 119.265 92.175 120.395 ;
        RECT 85.300 118.525 90.645 119.070 ;
        RECT 90.820 118.695 91.075 119.265 ;
        RECT 91.245 119.095 92.175 119.265 ;
        RECT 92.345 120.055 93.355 120.225 ;
        RECT 92.345 119.255 92.515 120.055 ;
        RECT 92.000 119.060 92.175 119.095 ;
        RECT 91.245 118.525 91.575 118.925 ;
        RECT 92.000 118.695 92.530 119.060 ;
        RECT 92.720 119.035 92.995 119.855 ;
        RECT 92.715 118.865 92.995 119.035 ;
        RECT 92.720 118.695 92.995 118.865 ;
        RECT 93.165 118.695 93.355 120.055 ;
        RECT 93.525 120.070 93.695 120.735 ;
        RECT 93.865 120.315 94.035 121.075 ;
        RECT 94.270 120.315 94.785 120.725 ;
        RECT 93.525 119.880 94.275 120.070 ;
        RECT 94.445 119.505 94.785 120.315 ;
        RECT 93.555 119.335 94.785 119.505 ;
        RECT 95.415 119.985 97.085 121.075 ;
        RECT 97.255 120.315 97.770 120.725 ;
        RECT 98.005 120.315 98.175 121.075 ;
        RECT 98.345 120.735 100.375 120.905 ;
        RECT 95.415 119.465 96.165 119.985 ;
        RECT 93.535 118.525 94.045 119.060 ;
        RECT 94.265 118.730 94.510 119.335 ;
        RECT 96.335 119.295 97.085 119.815 ;
        RECT 97.255 119.505 97.595 120.315 ;
        RECT 98.345 120.070 98.515 120.735 ;
        RECT 98.910 120.395 100.035 120.565 ;
        RECT 97.765 119.880 98.515 120.070 ;
        RECT 98.685 120.055 99.695 120.225 ;
        RECT 97.255 119.335 98.485 119.505 ;
        RECT 95.415 118.525 97.085 119.295 ;
        RECT 97.530 118.730 97.775 119.335 ;
        RECT 97.995 118.525 98.505 119.060 ;
        RECT 98.685 118.695 98.875 120.055 ;
        RECT 99.045 119.715 99.320 119.855 ;
        RECT 99.045 119.545 99.325 119.715 ;
        RECT 99.045 118.695 99.320 119.545 ;
        RECT 99.525 119.255 99.695 120.055 ;
        RECT 99.865 119.265 100.035 120.395 ;
        RECT 100.205 119.765 100.375 120.735 ;
        RECT 100.545 119.935 100.715 121.075 ;
        RECT 100.885 119.935 101.220 120.905 ;
        RECT 100.205 119.435 100.400 119.765 ;
        RECT 100.625 119.435 100.880 119.765 ;
        RECT 100.625 119.265 100.795 119.435 ;
        RECT 101.050 119.265 101.220 119.935 ;
        RECT 101.395 119.910 101.685 121.075 ;
        RECT 101.855 119.985 103.065 121.075 ;
        RECT 101.855 119.445 102.375 119.985 ;
        RECT 103.275 119.935 103.505 121.075 ;
        RECT 103.675 119.925 104.005 120.905 ;
        RECT 104.175 119.935 104.385 121.075 ;
        RECT 104.615 120.315 105.130 120.725 ;
        RECT 105.365 120.315 105.535 121.075 ;
        RECT 105.705 120.735 107.735 120.905 ;
        RECT 102.545 119.275 103.065 119.815 ;
        RECT 103.255 119.515 103.585 119.765 ;
        RECT 99.865 119.095 100.795 119.265 ;
        RECT 99.865 119.060 100.040 119.095 ;
        RECT 99.510 118.695 100.040 119.060 ;
        RECT 100.465 118.525 100.795 118.925 ;
        RECT 100.965 118.695 101.220 119.265 ;
        RECT 101.395 118.525 101.685 119.250 ;
        RECT 101.855 118.525 103.065 119.275 ;
        RECT 103.275 118.525 103.505 119.345 ;
        RECT 103.755 119.325 104.005 119.925 ;
        RECT 104.615 119.505 104.955 120.315 ;
        RECT 105.705 120.070 105.875 120.735 ;
        RECT 106.270 120.395 107.395 120.565 ;
        RECT 105.125 119.880 105.875 120.070 ;
        RECT 106.045 120.055 107.055 120.225 ;
        RECT 103.675 118.695 104.005 119.325 ;
        RECT 104.175 118.525 104.385 119.345 ;
        RECT 104.615 119.335 105.845 119.505 ;
        RECT 104.890 118.730 105.135 119.335 ;
        RECT 105.355 118.525 105.865 119.060 ;
        RECT 106.045 118.695 106.235 120.055 ;
        RECT 106.405 119.375 106.680 119.855 ;
        RECT 106.405 119.205 106.685 119.375 ;
        RECT 106.885 119.255 107.055 120.055 ;
        RECT 107.225 119.265 107.395 120.395 ;
        RECT 107.565 119.765 107.735 120.735 ;
        RECT 107.905 119.935 108.075 121.075 ;
        RECT 108.245 119.935 108.580 120.905 ;
        RECT 109.130 120.095 109.385 120.765 ;
        RECT 109.565 120.275 109.850 121.075 ;
        RECT 110.030 120.355 110.360 120.865 ;
        RECT 109.130 120.055 109.310 120.095 ;
        RECT 107.565 119.435 107.760 119.765 ;
        RECT 107.985 119.435 108.240 119.765 ;
        RECT 107.985 119.265 108.155 119.435 ;
        RECT 108.410 119.265 108.580 119.935 ;
        RECT 109.045 119.885 109.310 120.055 ;
        RECT 106.405 118.695 106.680 119.205 ;
        RECT 107.225 119.095 108.155 119.265 ;
        RECT 107.225 119.060 107.400 119.095 ;
        RECT 106.870 118.695 107.400 119.060 ;
        RECT 107.825 118.525 108.155 118.925 ;
        RECT 108.325 118.695 108.580 119.265 ;
        RECT 109.130 119.235 109.310 119.885 ;
        RECT 110.030 119.765 110.280 120.355 ;
        RECT 110.630 120.205 110.800 120.815 ;
        RECT 110.970 120.385 111.300 121.075 ;
        RECT 111.530 120.525 111.770 120.815 ;
        RECT 111.970 120.695 112.390 121.075 ;
        RECT 112.570 120.605 113.200 120.855 ;
        RECT 113.670 120.695 114.000 121.075 ;
        RECT 112.570 120.525 112.740 120.605 ;
        RECT 114.170 120.525 114.340 120.815 ;
        RECT 114.520 120.695 114.900 121.075 ;
        RECT 115.140 120.690 115.970 120.860 ;
        RECT 111.530 120.355 112.740 120.525 ;
        RECT 109.480 119.435 110.280 119.765 ;
        RECT 109.130 118.705 109.385 119.235 ;
        RECT 109.565 118.525 109.850 118.985 ;
        RECT 110.030 118.785 110.280 119.435 ;
        RECT 110.480 120.185 110.800 120.205 ;
        RECT 110.480 120.015 112.400 120.185 ;
        RECT 110.480 119.120 110.670 120.015 ;
        RECT 112.570 119.845 112.740 120.355 ;
        RECT 112.910 120.095 113.430 120.405 ;
        RECT 110.840 119.675 112.740 119.845 ;
        RECT 110.840 119.615 111.170 119.675 ;
        RECT 111.320 119.445 111.650 119.505 ;
        RECT 110.990 119.175 111.650 119.445 ;
        RECT 110.480 118.790 110.800 119.120 ;
        RECT 110.980 118.525 111.640 119.005 ;
        RECT 111.840 118.915 112.010 119.675 ;
        RECT 112.910 119.505 113.090 119.915 ;
        RECT 112.180 119.335 112.510 119.455 ;
        RECT 113.260 119.335 113.430 120.095 ;
        RECT 112.180 119.165 113.430 119.335 ;
        RECT 113.600 120.275 114.970 120.525 ;
        RECT 113.600 119.505 113.790 120.275 ;
        RECT 114.720 120.015 114.970 120.275 ;
        RECT 113.960 119.845 114.210 120.005 ;
        RECT 115.140 119.845 115.310 120.690 ;
        RECT 116.205 120.405 116.375 120.905 ;
        RECT 116.545 120.575 116.875 121.075 ;
        RECT 115.480 120.015 115.980 120.395 ;
        RECT 116.205 120.235 116.900 120.405 ;
        RECT 113.960 119.675 115.310 119.845 ;
        RECT 114.890 119.635 115.310 119.675 ;
        RECT 113.600 119.165 114.020 119.505 ;
        RECT 114.310 119.175 114.720 119.505 ;
        RECT 111.840 118.745 112.690 118.915 ;
        RECT 113.250 118.525 113.570 118.985 ;
        RECT 113.770 118.735 114.020 119.165 ;
        RECT 114.310 118.525 114.720 118.965 ;
        RECT 114.890 118.905 115.060 119.635 ;
        RECT 115.230 119.085 115.580 119.455 ;
        RECT 115.760 119.145 115.980 120.015 ;
        RECT 116.150 119.445 116.560 120.065 ;
        RECT 116.730 119.265 116.900 120.235 ;
        RECT 116.205 119.075 116.900 119.265 ;
        RECT 114.890 118.705 115.905 118.905 ;
        RECT 116.205 118.745 116.375 119.075 ;
        RECT 116.545 118.525 116.875 118.905 ;
        RECT 117.090 118.785 117.315 120.905 ;
        RECT 117.485 120.575 117.815 121.075 ;
        RECT 117.985 120.405 118.155 120.905 ;
        RECT 117.490 120.235 118.155 120.405 ;
        RECT 117.490 119.245 117.720 120.235 ;
        RECT 117.890 119.415 118.240 120.065 ;
        RECT 118.455 119.935 118.685 121.075 ;
        RECT 118.855 119.925 119.185 120.905 ;
        RECT 119.355 119.935 119.565 121.075 ;
        RECT 120.345 120.145 120.515 120.905 ;
        RECT 120.695 120.315 121.025 121.075 ;
        RECT 120.345 119.975 121.010 120.145 ;
        RECT 121.195 120.000 121.465 120.905 ;
        RECT 118.435 119.515 118.765 119.765 ;
        RECT 117.490 119.075 118.155 119.245 ;
        RECT 117.485 118.525 117.815 118.905 ;
        RECT 117.985 118.785 118.155 119.075 ;
        RECT 118.455 118.525 118.685 119.345 ;
        RECT 118.935 119.325 119.185 119.925 ;
        RECT 120.840 119.830 121.010 119.975 ;
        RECT 120.275 119.425 120.605 119.795 ;
        RECT 120.840 119.500 121.125 119.830 ;
        RECT 118.855 118.695 119.185 119.325 ;
        RECT 119.355 118.525 119.565 119.345 ;
        RECT 120.840 119.245 121.010 119.500 ;
        RECT 120.345 119.075 121.010 119.245 ;
        RECT 121.295 119.200 121.465 120.000 ;
        RECT 122.555 119.985 126.065 121.075 ;
        RECT 126.235 119.985 127.445 121.075 ;
        RECT 122.555 119.465 124.245 119.985 ;
        RECT 124.415 119.295 126.065 119.815 ;
        RECT 126.235 119.445 126.755 119.985 ;
        RECT 120.345 118.695 120.515 119.075 ;
        RECT 120.695 118.525 121.025 118.905 ;
        RECT 121.205 118.695 121.465 119.200 ;
        RECT 122.555 118.525 126.065 119.295 ;
        RECT 126.925 119.275 127.445 119.815 ;
        RECT 126.235 118.525 127.445 119.275 ;
        RECT 14.370 118.355 127.530 118.525 ;
        RECT 14.455 117.605 15.665 118.355 ;
        RECT 14.455 117.065 14.975 117.605 ;
        RECT 16.355 117.535 16.565 118.355 ;
        RECT 16.735 117.555 17.065 118.185 ;
        RECT 15.145 116.895 15.665 117.435 ;
        RECT 16.735 116.955 16.985 117.555 ;
        RECT 17.235 117.535 17.465 118.355 ;
        RECT 18.050 118.015 18.305 118.175 ;
        RECT 17.965 117.845 18.305 118.015 ;
        RECT 18.485 117.895 18.770 118.355 ;
        RECT 18.050 117.645 18.305 117.845 ;
        RECT 17.155 117.115 17.485 117.365 ;
        RECT 14.455 115.805 15.665 116.895 ;
        RECT 16.355 115.805 16.565 116.945 ;
        RECT 16.735 115.975 17.065 116.955 ;
        RECT 17.235 115.805 17.465 116.945 ;
        RECT 18.050 116.785 18.230 117.645 ;
        RECT 18.950 117.445 19.200 118.095 ;
        RECT 18.400 117.115 19.200 117.445 ;
        RECT 18.050 116.115 18.305 116.785 ;
        RECT 18.485 115.805 18.770 116.605 ;
        RECT 18.950 116.525 19.200 117.115 ;
        RECT 19.400 117.760 19.720 118.090 ;
        RECT 19.900 117.875 20.560 118.355 ;
        RECT 20.760 117.965 21.610 118.135 ;
        RECT 19.400 116.865 19.590 117.760 ;
        RECT 19.910 117.435 20.570 117.705 ;
        RECT 20.240 117.375 20.570 117.435 ;
        RECT 19.760 117.205 20.090 117.265 ;
        RECT 20.760 117.205 20.930 117.965 ;
        RECT 22.170 117.895 22.490 118.355 ;
        RECT 22.690 117.715 22.940 118.145 ;
        RECT 23.230 117.915 23.640 118.355 ;
        RECT 23.810 117.975 24.825 118.175 ;
        RECT 21.100 117.545 22.350 117.715 ;
        RECT 21.100 117.425 21.430 117.545 ;
        RECT 19.760 117.035 21.660 117.205 ;
        RECT 19.400 116.695 21.320 116.865 ;
        RECT 19.400 116.675 19.720 116.695 ;
        RECT 18.950 116.015 19.280 116.525 ;
        RECT 19.550 116.065 19.720 116.675 ;
        RECT 21.490 116.525 21.660 117.035 ;
        RECT 21.830 116.965 22.010 117.375 ;
        RECT 22.180 116.785 22.350 117.545 ;
        RECT 19.890 115.805 20.220 116.495 ;
        RECT 20.450 116.355 21.660 116.525 ;
        RECT 21.830 116.475 22.350 116.785 ;
        RECT 22.520 117.375 22.940 117.715 ;
        RECT 23.230 117.375 23.640 117.705 ;
        RECT 22.520 116.605 22.710 117.375 ;
        RECT 23.810 117.245 23.980 117.975 ;
        RECT 25.125 117.805 25.295 118.135 ;
        RECT 25.465 117.975 25.795 118.355 ;
        RECT 24.150 117.425 24.500 117.795 ;
        RECT 23.810 117.205 24.230 117.245 ;
        RECT 22.880 117.035 24.230 117.205 ;
        RECT 22.880 116.875 23.130 117.035 ;
        RECT 23.640 116.605 23.890 116.865 ;
        RECT 22.520 116.355 23.890 116.605 ;
        RECT 20.450 116.065 20.690 116.355 ;
        RECT 21.490 116.275 21.660 116.355 ;
        RECT 20.890 115.805 21.310 116.185 ;
        RECT 21.490 116.025 22.120 116.275 ;
        RECT 22.590 115.805 22.920 116.185 ;
        RECT 23.090 116.065 23.260 116.355 ;
        RECT 24.060 116.190 24.230 117.035 ;
        RECT 24.680 116.865 24.900 117.735 ;
        RECT 25.125 117.615 25.820 117.805 ;
        RECT 24.400 116.485 24.900 116.865 ;
        RECT 25.070 116.815 25.480 117.435 ;
        RECT 25.650 116.645 25.820 117.615 ;
        RECT 25.125 116.475 25.820 116.645 ;
        RECT 23.440 115.805 23.820 116.185 ;
        RECT 24.060 116.020 24.890 116.190 ;
        RECT 25.125 115.975 25.295 116.475 ;
        RECT 25.465 115.805 25.795 116.305 ;
        RECT 26.010 115.975 26.235 118.095 ;
        RECT 26.405 117.975 26.735 118.355 ;
        RECT 26.905 117.805 27.075 118.095 ;
        RECT 26.410 117.635 27.075 117.805 ;
        RECT 27.425 117.805 27.595 118.095 ;
        RECT 27.765 117.975 28.095 118.355 ;
        RECT 27.425 117.635 28.090 117.805 ;
        RECT 26.410 116.645 26.640 117.635 ;
        RECT 26.810 116.815 27.160 117.465 ;
        RECT 27.340 116.815 27.690 117.465 ;
        RECT 27.860 116.645 28.090 117.635 ;
        RECT 26.410 116.475 27.075 116.645 ;
        RECT 26.405 115.805 26.735 116.305 ;
        RECT 26.905 115.975 27.075 116.475 ;
        RECT 27.425 116.475 28.090 116.645 ;
        RECT 27.425 115.975 27.595 116.475 ;
        RECT 27.765 115.805 28.095 116.305 ;
        RECT 28.265 115.975 28.490 118.095 ;
        RECT 28.705 117.975 29.035 118.355 ;
        RECT 29.205 117.805 29.375 118.135 ;
        RECT 29.675 117.975 30.690 118.175 ;
        RECT 28.680 117.615 29.375 117.805 ;
        RECT 28.680 116.645 28.850 117.615 ;
        RECT 29.020 116.815 29.430 117.435 ;
        RECT 29.600 116.865 29.820 117.735 ;
        RECT 30.000 117.425 30.350 117.795 ;
        RECT 30.520 117.245 30.690 117.975 ;
        RECT 30.860 117.915 31.270 118.355 ;
        RECT 31.560 117.715 31.810 118.145 ;
        RECT 32.010 117.895 32.330 118.355 ;
        RECT 32.890 117.965 33.740 118.135 ;
        RECT 30.860 117.375 31.270 117.705 ;
        RECT 31.560 117.375 31.980 117.715 ;
        RECT 30.270 117.205 30.690 117.245 ;
        RECT 30.270 117.035 31.620 117.205 ;
        RECT 28.680 116.475 29.375 116.645 ;
        RECT 29.600 116.485 30.100 116.865 ;
        RECT 28.705 115.805 29.035 116.305 ;
        RECT 29.205 115.975 29.375 116.475 ;
        RECT 30.270 116.190 30.440 117.035 ;
        RECT 31.370 116.875 31.620 117.035 ;
        RECT 30.610 116.605 30.860 116.865 ;
        RECT 31.790 116.605 31.980 117.375 ;
        RECT 30.610 116.355 31.980 116.605 ;
        RECT 32.150 117.545 33.400 117.715 ;
        RECT 32.150 116.785 32.320 117.545 ;
        RECT 33.070 117.425 33.400 117.545 ;
        RECT 32.490 116.965 32.670 117.375 ;
        RECT 33.570 117.205 33.740 117.965 ;
        RECT 33.940 117.875 34.600 118.355 ;
        RECT 34.780 117.760 35.100 118.090 ;
        RECT 33.930 117.435 34.590 117.705 ;
        RECT 33.930 117.375 34.260 117.435 ;
        RECT 34.410 117.205 34.740 117.265 ;
        RECT 32.840 117.035 34.740 117.205 ;
        RECT 32.150 116.475 32.670 116.785 ;
        RECT 32.840 116.525 33.010 117.035 ;
        RECT 34.910 116.865 35.100 117.760 ;
        RECT 33.180 116.695 35.100 116.865 ;
        RECT 34.780 116.675 35.100 116.695 ;
        RECT 35.300 117.445 35.550 118.095 ;
        RECT 35.730 117.895 36.015 118.355 ;
        RECT 36.195 118.015 36.450 118.175 ;
        RECT 36.195 117.845 36.535 118.015 ;
        RECT 36.195 117.645 36.450 117.845 ;
        RECT 35.300 117.115 36.100 117.445 ;
        RECT 32.840 116.355 34.050 116.525 ;
        RECT 29.610 116.020 30.440 116.190 ;
        RECT 30.680 115.805 31.060 116.185 ;
        RECT 31.240 116.065 31.410 116.355 ;
        RECT 32.840 116.275 33.010 116.355 ;
        RECT 31.580 115.805 31.910 116.185 ;
        RECT 32.380 116.025 33.010 116.275 ;
        RECT 33.190 115.805 33.610 116.185 ;
        RECT 33.810 116.065 34.050 116.355 ;
        RECT 34.280 115.805 34.610 116.495 ;
        RECT 34.780 116.065 34.950 116.675 ;
        RECT 35.300 116.525 35.550 117.115 ;
        RECT 36.270 116.785 36.450 117.645 ;
        RECT 36.995 117.630 37.285 118.355 ;
        RECT 37.830 118.015 38.085 118.175 ;
        RECT 37.745 117.845 38.085 118.015 ;
        RECT 38.265 117.895 38.550 118.355 ;
        RECT 37.830 117.645 38.085 117.845 ;
        RECT 35.220 116.015 35.550 116.525 ;
        RECT 35.730 115.805 36.015 116.605 ;
        RECT 36.195 116.115 36.450 116.785 ;
        RECT 36.995 115.805 37.285 116.970 ;
        RECT 37.830 116.785 38.010 117.645 ;
        RECT 38.730 117.445 38.980 118.095 ;
        RECT 38.180 117.115 38.980 117.445 ;
        RECT 37.830 116.115 38.085 116.785 ;
        RECT 38.265 115.805 38.550 116.605 ;
        RECT 38.730 116.525 38.980 117.115 ;
        RECT 39.180 117.760 39.500 118.090 ;
        RECT 39.680 117.875 40.340 118.355 ;
        RECT 40.540 117.965 41.390 118.135 ;
        RECT 39.180 116.865 39.370 117.760 ;
        RECT 39.690 117.435 40.350 117.705 ;
        RECT 40.020 117.375 40.350 117.435 ;
        RECT 39.540 117.205 39.870 117.265 ;
        RECT 40.540 117.205 40.710 117.965 ;
        RECT 41.950 117.895 42.270 118.355 ;
        RECT 42.470 117.715 42.720 118.145 ;
        RECT 43.010 117.915 43.420 118.355 ;
        RECT 43.590 117.975 44.605 118.175 ;
        RECT 40.880 117.545 42.130 117.715 ;
        RECT 40.880 117.425 41.210 117.545 ;
        RECT 39.540 117.035 41.440 117.205 ;
        RECT 39.180 116.695 41.100 116.865 ;
        RECT 39.180 116.675 39.500 116.695 ;
        RECT 38.730 116.015 39.060 116.525 ;
        RECT 39.330 116.065 39.500 116.675 ;
        RECT 41.270 116.525 41.440 117.035 ;
        RECT 41.610 116.965 41.790 117.375 ;
        RECT 41.960 116.785 42.130 117.545 ;
        RECT 39.670 115.805 40.000 116.495 ;
        RECT 40.230 116.355 41.440 116.525 ;
        RECT 41.610 116.475 42.130 116.785 ;
        RECT 42.300 117.375 42.720 117.715 ;
        RECT 43.010 117.375 43.420 117.705 ;
        RECT 42.300 116.605 42.490 117.375 ;
        RECT 43.590 117.245 43.760 117.975 ;
        RECT 44.905 117.805 45.075 118.135 ;
        RECT 45.245 117.975 45.575 118.355 ;
        RECT 43.930 117.425 44.280 117.795 ;
        RECT 43.590 117.205 44.010 117.245 ;
        RECT 42.660 117.035 44.010 117.205 ;
        RECT 42.660 116.875 42.910 117.035 ;
        RECT 43.420 116.605 43.670 116.865 ;
        RECT 42.300 116.355 43.670 116.605 ;
        RECT 40.230 116.065 40.470 116.355 ;
        RECT 41.270 116.275 41.440 116.355 ;
        RECT 40.670 115.805 41.090 116.185 ;
        RECT 41.270 116.025 41.900 116.275 ;
        RECT 42.370 115.805 42.700 116.185 ;
        RECT 42.870 116.065 43.040 116.355 ;
        RECT 43.840 116.190 44.010 117.035 ;
        RECT 44.460 116.865 44.680 117.735 ;
        RECT 44.905 117.615 45.600 117.805 ;
        RECT 44.180 116.485 44.680 116.865 ;
        RECT 44.850 116.815 45.260 117.435 ;
        RECT 45.430 116.645 45.600 117.615 ;
        RECT 44.905 116.475 45.600 116.645 ;
        RECT 43.220 115.805 43.600 116.185 ;
        RECT 43.840 116.020 44.670 116.190 ;
        RECT 44.905 115.975 45.075 116.475 ;
        RECT 45.245 115.805 45.575 116.305 ;
        RECT 45.790 115.975 46.015 118.095 ;
        RECT 46.185 117.975 46.515 118.355 ;
        RECT 46.685 117.805 46.855 118.095 ;
        RECT 46.190 117.635 46.855 117.805 ;
        RECT 47.490 117.645 47.745 118.175 ;
        RECT 47.925 117.895 48.210 118.355 ;
        RECT 46.190 116.645 46.420 117.635 ;
        RECT 46.590 116.815 46.940 117.465 ;
        RECT 47.490 116.785 47.670 117.645 ;
        RECT 48.390 117.445 48.640 118.095 ;
        RECT 47.840 117.115 48.640 117.445 ;
        RECT 46.190 116.475 46.855 116.645 ;
        RECT 46.185 115.805 46.515 116.305 ;
        RECT 46.685 115.975 46.855 116.475 ;
        RECT 47.490 116.315 47.745 116.785 ;
        RECT 47.405 116.145 47.745 116.315 ;
        RECT 47.490 116.115 47.745 116.145 ;
        RECT 47.925 115.805 48.210 116.605 ;
        RECT 48.390 116.525 48.640 117.115 ;
        RECT 48.840 117.760 49.160 118.090 ;
        RECT 49.340 117.875 50.000 118.355 ;
        RECT 50.200 117.965 51.050 118.135 ;
        RECT 48.840 116.865 49.030 117.760 ;
        RECT 49.350 117.435 50.010 117.705 ;
        RECT 49.680 117.375 50.010 117.435 ;
        RECT 49.200 117.205 49.530 117.265 ;
        RECT 50.200 117.205 50.370 117.965 ;
        RECT 51.610 117.895 51.930 118.355 ;
        RECT 52.130 117.715 52.380 118.145 ;
        RECT 52.670 117.915 53.080 118.355 ;
        RECT 53.250 117.975 54.265 118.175 ;
        RECT 50.540 117.545 51.790 117.715 ;
        RECT 50.540 117.425 50.870 117.545 ;
        RECT 49.200 117.035 51.100 117.205 ;
        RECT 48.840 116.695 50.760 116.865 ;
        RECT 48.840 116.675 49.160 116.695 ;
        RECT 48.390 116.015 48.720 116.525 ;
        RECT 48.990 116.065 49.160 116.675 ;
        RECT 50.930 116.525 51.100 117.035 ;
        RECT 51.270 116.965 51.450 117.375 ;
        RECT 51.620 116.785 51.790 117.545 ;
        RECT 49.330 115.805 49.660 116.495 ;
        RECT 49.890 116.355 51.100 116.525 ;
        RECT 51.270 116.475 51.790 116.785 ;
        RECT 51.960 117.375 52.380 117.715 ;
        RECT 52.670 117.375 53.080 117.705 ;
        RECT 51.960 116.605 52.150 117.375 ;
        RECT 53.250 117.245 53.420 117.975 ;
        RECT 54.565 117.805 54.735 118.135 ;
        RECT 54.905 117.975 55.235 118.355 ;
        RECT 53.590 117.425 53.940 117.795 ;
        RECT 53.250 117.205 53.670 117.245 ;
        RECT 52.320 117.035 53.670 117.205 ;
        RECT 52.320 116.875 52.570 117.035 ;
        RECT 53.080 116.605 53.330 116.865 ;
        RECT 51.960 116.355 53.330 116.605 ;
        RECT 49.890 116.065 50.130 116.355 ;
        RECT 50.930 116.275 51.100 116.355 ;
        RECT 50.330 115.805 50.750 116.185 ;
        RECT 50.930 116.025 51.560 116.275 ;
        RECT 52.030 115.805 52.360 116.185 ;
        RECT 52.530 116.065 52.700 116.355 ;
        RECT 53.500 116.190 53.670 117.035 ;
        RECT 54.120 116.865 54.340 117.735 ;
        RECT 54.565 117.615 55.260 117.805 ;
        RECT 53.840 116.485 54.340 116.865 ;
        RECT 54.510 116.815 54.920 117.435 ;
        RECT 55.090 116.645 55.260 117.615 ;
        RECT 54.565 116.475 55.260 116.645 ;
        RECT 52.880 115.805 53.260 116.185 ;
        RECT 53.500 116.020 54.330 116.190 ;
        RECT 54.565 115.975 54.735 116.475 ;
        RECT 54.905 115.805 55.235 116.305 ;
        RECT 55.450 115.975 55.675 118.095 ;
        RECT 55.845 117.975 56.175 118.355 ;
        RECT 56.345 117.805 56.515 118.095 ;
        RECT 55.850 117.635 56.515 117.805 ;
        RECT 55.850 116.645 56.080 117.635 ;
        RECT 57.695 117.585 61.205 118.355 ;
        RECT 56.250 116.815 56.600 117.465 ;
        RECT 57.695 116.895 59.385 117.415 ;
        RECT 59.555 117.065 61.205 117.585 ;
        RECT 61.415 117.535 61.645 118.355 ;
        RECT 61.815 117.555 62.145 118.185 ;
        RECT 61.395 117.115 61.725 117.365 ;
        RECT 61.895 116.955 62.145 117.555 ;
        RECT 62.315 117.535 62.525 118.355 ;
        RECT 62.755 117.630 63.045 118.355 ;
        RECT 63.590 118.015 63.845 118.175 ;
        RECT 63.505 117.845 63.845 118.015 ;
        RECT 64.025 117.895 64.310 118.355 ;
        RECT 63.590 117.645 63.845 117.845 ;
        RECT 55.850 116.475 56.515 116.645 ;
        RECT 55.845 115.805 56.175 116.305 ;
        RECT 56.345 115.975 56.515 116.475 ;
        RECT 57.695 115.805 61.205 116.895 ;
        RECT 61.415 115.805 61.645 116.945 ;
        RECT 61.815 115.975 62.145 116.955 ;
        RECT 62.315 115.805 62.525 116.945 ;
        RECT 62.755 115.805 63.045 116.970 ;
        RECT 63.590 116.785 63.770 117.645 ;
        RECT 64.490 117.445 64.740 118.095 ;
        RECT 63.940 117.115 64.740 117.445 ;
        RECT 63.590 116.115 63.845 116.785 ;
        RECT 64.025 115.805 64.310 116.605 ;
        RECT 64.490 116.525 64.740 117.115 ;
        RECT 64.940 117.760 65.260 118.090 ;
        RECT 65.440 117.875 66.100 118.355 ;
        RECT 66.300 117.965 67.150 118.135 ;
        RECT 64.940 116.865 65.130 117.760 ;
        RECT 65.450 117.435 66.110 117.705 ;
        RECT 65.780 117.375 66.110 117.435 ;
        RECT 65.300 117.205 65.630 117.265 ;
        RECT 66.300 117.205 66.470 117.965 ;
        RECT 67.710 117.895 68.030 118.355 ;
        RECT 68.230 117.715 68.480 118.145 ;
        RECT 68.770 117.915 69.180 118.355 ;
        RECT 69.350 117.975 70.365 118.175 ;
        RECT 66.640 117.545 67.890 117.715 ;
        RECT 66.640 117.425 66.970 117.545 ;
        RECT 65.300 117.035 67.200 117.205 ;
        RECT 64.940 116.695 66.860 116.865 ;
        RECT 64.940 116.675 65.260 116.695 ;
        RECT 64.490 116.015 64.820 116.525 ;
        RECT 65.090 116.065 65.260 116.675 ;
        RECT 67.030 116.525 67.200 117.035 ;
        RECT 67.370 116.965 67.550 117.375 ;
        RECT 67.720 116.785 67.890 117.545 ;
        RECT 65.430 115.805 65.760 116.495 ;
        RECT 65.990 116.355 67.200 116.525 ;
        RECT 67.370 116.475 67.890 116.785 ;
        RECT 68.060 117.375 68.480 117.715 ;
        RECT 68.770 117.375 69.180 117.705 ;
        RECT 68.060 116.605 68.250 117.375 ;
        RECT 69.350 117.245 69.520 117.975 ;
        RECT 70.665 117.805 70.835 118.135 ;
        RECT 71.005 117.975 71.335 118.355 ;
        RECT 69.690 117.425 70.040 117.795 ;
        RECT 69.350 117.205 69.770 117.245 ;
        RECT 68.420 117.035 69.770 117.205 ;
        RECT 68.420 116.875 68.670 117.035 ;
        RECT 69.180 116.605 69.430 116.865 ;
        RECT 68.060 116.355 69.430 116.605 ;
        RECT 65.990 116.065 66.230 116.355 ;
        RECT 67.030 116.275 67.200 116.355 ;
        RECT 66.430 115.805 66.850 116.185 ;
        RECT 67.030 116.025 67.660 116.275 ;
        RECT 68.130 115.805 68.460 116.185 ;
        RECT 68.630 116.065 68.800 116.355 ;
        RECT 69.600 116.190 69.770 117.035 ;
        RECT 70.220 116.865 70.440 117.735 ;
        RECT 70.665 117.615 71.360 117.805 ;
        RECT 69.940 116.485 70.440 116.865 ;
        RECT 70.610 116.815 71.020 117.435 ;
        RECT 71.190 116.645 71.360 117.615 ;
        RECT 70.665 116.475 71.360 116.645 ;
        RECT 68.980 115.805 69.360 116.185 ;
        RECT 69.600 116.020 70.430 116.190 ;
        RECT 70.665 115.975 70.835 116.475 ;
        RECT 71.005 115.805 71.335 116.305 ;
        RECT 71.550 115.975 71.775 118.095 ;
        RECT 71.945 117.975 72.275 118.355 ;
        RECT 72.445 117.805 72.615 118.095 ;
        RECT 73.250 118.015 73.505 118.175 ;
        RECT 73.165 117.845 73.505 118.015 ;
        RECT 73.685 117.895 73.970 118.355 ;
        RECT 71.950 117.635 72.615 117.805 ;
        RECT 73.250 117.645 73.505 117.845 ;
        RECT 71.950 116.645 72.180 117.635 ;
        RECT 72.350 116.815 72.700 117.465 ;
        RECT 73.250 116.785 73.430 117.645 ;
        RECT 74.150 117.445 74.400 118.095 ;
        RECT 73.600 117.115 74.400 117.445 ;
        RECT 71.950 116.475 72.615 116.645 ;
        RECT 71.945 115.805 72.275 116.305 ;
        RECT 72.445 115.975 72.615 116.475 ;
        RECT 73.250 116.115 73.505 116.785 ;
        RECT 73.685 115.805 73.970 116.605 ;
        RECT 74.150 116.525 74.400 117.115 ;
        RECT 74.600 117.760 74.920 118.090 ;
        RECT 75.100 117.875 75.760 118.355 ;
        RECT 75.960 117.965 76.810 118.135 ;
        RECT 74.600 116.865 74.790 117.760 ;
        RECT 75.110 117.435 75.770 117.705 ;
        RECT 75.440 117.375 75.770 117.435 ;
        RECT 74.960 117.205 75.290 117.265 ;
        RECT 75.960 117.205 76.130 117.965 ;
        RECT 77.370 117.895 77.690 118.355 ;
        RECT 77.890 117.715 78.140 118.145 ;
        RECT 78.430 117.915 78.840 118.355 ;
        RECT 79.010 117.975 80.025 118.175 ;
        RECT 76.300 117.545 77.550 117.715 ;
        RECT 76.300 117.425 76.630 117.545 ;
        RECT 74.960 117.035 76.860 117.205 ;
        RECT 74.600 116.695 76.520 116.865 ;
        RECT 74.600 116.675 74.920 116.695 ;
        RECT 74.150 116.015 74.480 116.525 ;
        RECT 74.750 116.065 74.920 116.675 ;
        RECT 76.690 116.525 76.860 117.035 ;
        RECT 77.030 116.965 77.210 117.375 ;
        RECT 77.380 116.785 77.550 117.545 ;
        RECT 75.090 115.805 75.420 116.495 ;
        RECT 75.650 116.355 76.860 116.525 ;
        RECT 77.030 116.475 77.550 116.785 ;
        RECT 77.720 117.375 78.140 117.715 ;
        RECT 78.430 117.375 78.840 117.705 ;
        RECT 77.720 116.605 77.910 117.375 ;
        RECT 79.010 117.245 79.180 117.975 ;
        RECT 80.325 117.805 80.495 118.135 ;
        RECT 80.665 117.975 80.995 118.355 ;
        RECT 79.350 117.425 79.700 117.795 ;
        RECT 79.010 117.205 79.430 117.245 ;
        RECT 78.080 117.035 79.430 117.205 ;
        RECT 78.080 116.875 78.330 117.035 ;
        RECT 78.840 116.605 79.090 116.865 ;
        RECT 77.720 116.355 79.090 116.605 ;
        RECT 75.650 116.065 75.890 116.355 ;
        RECT 76.690 116.275 76.860 116.355 ;
        RECT 76.090 115.805 76.510 116.185 ;
        RECT 76.690 116.025 77.320 116.275 ;
        RECT 77.790 115.805 78.120 116.185 ;
        RECT 78.290 116.065 78.460 116.355 ;
        RECT 79.260 116.190 79.430 117.035 ;
        RECT 79.880 116.865 80.100 117.735 ;
        RECT 80.325 117.615 81.020 117.805 ;
        RECT 79.600 116.485 80.100 116.865 ;
        RECT 80.270 116.815 80.680 117.435 ;
        RECT 80.850 116.645 81.020 117.615 ;
        RECT 80.325 116.475 81.020 116.645 ;
        RECT 78.640 115.805 79.020 116.185 ;
        RECT 79.260 116.020 80.090 116.190 ;
        RECT 80.325 115.975 80.495 116.475 ;
        RECT 80.665 115.805 80.995 116.305 ;
        RECT 81.210 115.975 81.435 118.095 ;
        RECT 81.605 117.975 81.935 118.355 ;
        RECT 82.105 117.805 82.275 118.095 ;
        RECT 81.610 117.635 82.275 117.805 ;
        RECT 81.610 116.645 81.840 117.635 ;
        RECT 82.540 117.615 82.795 118.185 ;
        RECT 82.965 117.955 83.295 118.355 ;
        RECT 83.720 117.820 84.250 118.185 ;
        RECT 83.720 117.785 83.895 117.820 ;
        RECT 82.965 117.615 83.895 117.785 ;
        RECT 82.010 116.815 82.360 117.465 ;
        RECT 82.540 116.945 82.710 117.615 ;
        RECT 82.965 117.445 83.135 117.615 ;
        RECT 82.880 117.115 83.135 117.445 ;
        RECT 83.360 117.115 83.555 117.445 ;
        RECT 81.610 116.475 82.275 116.645 ;
        RECT 81.605 115.805 81.935 116.305 ;
        RECT 82.105 115.975 82.275 116.475 ;
        RECT 82.540 115.975 82.875 116.945 ;
        RECT 83.045 115.805 83.215 116.945 ;
        RECT 83.385 116.145 83.555 117.115 ;
        RECT 83.725 116.485 83.895 117.615 ;
        RECT 84.065 116.825 84.235 117.625 ;
        RECT 84.440 117.335 84.715 118.185 ;
        RECT 84.435 117.165 84.715 117.335 ;
        RECT 84.440 117.025 84.715 117.165 ;
        RECT 84.885 116.825 85.075 118.185 ;
        RECT 85.255 117.820 85.765 118.355 ;
        RECT 85.985 117.545 86.230 118.150 ;
        RECT 87.225 117.805 87.395 118.185 ;
        RECT 87.575 117.975 87.905 118.355 ;
        RECT 87.225 117.635 87.890 117.805 ;
        RECT 88.085 117.680 88.345 118.185 ;
        RECT 85.275 117.375 86.505 117.545 ;
        RECT 84.065 116.655 85.075 116.825 ;
        RECT 85.245 116.810 85.995 117.000 ;
        RECT 83.725 116.315 84.850 116.485 ;
        RECT 85.245 116.145 85.415 116.810 ;
        RECT 86.165 116.565 86.505 117.375 ;
        RECT 87.155 117.085 87.485 117.455 ;
        RECT 87.720 117.380 87.890 117.635 ;
        RECT 87.720 117.050 88.005 117.380 ;
        RECT 87.720 116.905 87.890 117.050 ;
        RECT 83.385 115.975 85.415 116.145 ;
        RECT 85.585 115.805 85.755 116.565 ;
        RECT 85.990 116.155 86.505 116.565 ;
        RECT 87.225 116.735 87.890 116.905 ;
        RECT 88.175 116.880 88.345 117.680 ;
        RECT 88.515 117.630 88.805 118.355 ;
        RECT 89.015 117.535 89.245 118.355 ;
        RECT 89.415 117.555 89.745 118.185 ;
        RECT 88.995 117.115 89.325 117.365 ;
        RECT 87.225 115.975 87.395 116.735 ;
        RECT 87.575 115.805 87.905 116.565 ;
        RECT 88.075 115.975 88.345 116.880 ;
        RECT 88.515 115.805 88.805 116.970 ;
        RECT 89.495 116.955 89.745 117.555 ;
        RECT 89.915 117.535 90.125 118.355 ;
        RECT 90.395 117.535 90.625 118.355 ;
        RECT 90.795 117.555 91.125 118.185 ;
        RECT 90.375 117.115 90.705 117.365 ;
        RECT 90.875 116.955 91.125 117.555 ;
        RECT 91.295 117.535 91.505 118.355 ;
        RECT 93.030 118.015 93.285 118.175 ;
        RECT 92.945 117.845 93.285 118.015 ;
        RECT 93.465 117.895 93.750 118.355 ;
        RECT 93.030 117.645 93.285 117.845 ;
        RECT 89.015 115.805 89.245 116.945 ;
        RECT 89.415 115.975 89.745 116.955 ;
        RECT 89.915 115.805 90.125 116.945 ;
        RECT 90.395 115.805 90.625 116.945 ;
        RECT 90.795 115.975 91.125 116.955 ;
        RECT 91.295 115.805 91.505 116.945 ;
        RECT 93.030 116.785 93.210 117.645 ;
        RECT 93.930 117.445 94.180 118.095 ;
        RECT 93.380 117.115 94.180 117.445 ;
        RECT 93.030 116.115 93.285 116.785 ;
        RECT 93.465 115.805 93.750 116.605 ;
        RECT 93.930 116.525 94.180 117.115 ;
        RECT 94.380 117.760 94.700 118.090 ;
        RECT 94.880 117.875 95.540 118.355 ;
        RECT 95.740 117.965 96.590 118.135 ;
        RECT 94.380 116.865 94.570 117.760 ;
        RECT 94.890 117.435 95.550 117.705 ;
        RECT 95.220 117.375 95.550 117.435 ;
        RECT 94.740 117.205 95.070 117.265 ;
        RECT 95.740 117.205 95.910 117.965 ;
        RECT 97.150 117.895 97.470 118.355 ;
        RECT 97.670 117.715 97.920 118.145 ;
        RECT 98.210 117.915 98.620 118.355 ;
        RECT 98.790 117.975 99.805 118.175 ;
        RECT 96.080 117.545 97.330 117.715 ;
        RECT 96.080 117.425 96.410 117.545 ;
        RECT 94.740 117.035 96.640 117.205 ;
        RECT 94.380 116.695 96.300 116.865 ;
        RECT 94.380 116.675 94.700 116.695 ;
        RECT 93.930 116.015 94.260 116.525 ;
        RECT 94.530 116.065 94.700 116.675 ;
        RECT 96.470 116.525 96.640 117.035 ;
        RECT 96.810 116.965 96.990 117.375 ;
        RECT 97.160 116.785 97.330 117.545 ;
        RECT 94.870 115.805 95.200 116.495 ;
        RECT 95.430 116.355 96.640 116.525 ;
        RECT 96.810 116.475 97.330 116.785 ;
        RECT 97.500 117.375 97.920 117.715 ;
        RECT 98.210 117.375 98.620 117.705 ;
        RECT 97.500 116.605 97.690 117.375 ;
        RECT 98.790 117.245 98.960 117.975 ;
        RECT 100.105 117.805 100.275 118.135 ;
        RECT 100.445 117.975 100.775 118.355 ;
        RECT 99.130 117.425 99.480 117.795 ;
        RECT 98.790 117.205 99.210 117.245 ;
        RECT 97.860 117.035 99.210 117.205 ;
        RECT 97.860 116.875 98.110 117.035 ;
        RECT 98.620 116.605 98.870 116.865 ;
        RECT 97.500 116.355 98.870 116.605 ;
        RECT 95.430 116.065 95.670 116.355 ;
        RECT 96.470 116.275 96.640 116.355 ;
        RECT 95.870 115.805 96.290 116.185 ;
        RECT 96.470 116.025 97.100 116.275 ;
        RECT 97.570 115.805 97.900 116.185 ;
        RECT 98.070 116.065 98.240 116.355 ;
        RECT 99.040 116.190 99.210 117.035 ;
        RECT 99.660 116.865 99.880 117.735 ;
        RECT 100.105 117.615 100.800 117.805 ;
        RECT 99.380 116.485 99.880 116.865 ;
        RECT 100.050 116.815 100.460 117.435 ;
        RECT 100.630 116.645 100.800 117.615 ;
        RECT 100.105 116.475 100.800 116.645 ;
        RECT 98.420 115.805 98.800 116.185 ;
        RECT 99.040 116.020 99.870 116.190 ;
        RECT 100.105 115.975 100.275 116.475 ;
        RECT 100.445 115.805 100.775 116.305 ;
        RECT 100.990 115.975 101.215 118.095 ;
        RECT 101.385 117.975 101.715 118.355 ;
        RECT 101.885 117.805 102.055 118.095 ;
        RECT 102.690 118.015 102.945 118.175 ;
        RECT 102.605 117.845 102.945 118.015 ;
        RECT 103.125 117.895 103.410 118.355 ;
        RECT 101.390 117.635 102.055 117.805 ;
        RECT 102.690 117.645 102.945 117.845 ;
        RECT 101.390 116.645 101.620 117.635 ;
        RECT 101.790 116.815 102.140 117.465 ;
        RECT 102.690 116.785 102.870 117.645 ;
        RECT 103.590 117.445 103.840 118.095 ;
        RECT 103.040 117.115 103.840 117.445 ;
        RECT 101.390 116.475 102.055 116.645 ;
        RECT 101.385 115.805 101.715 116.305 ;
        RECT 101.885 115.975 102.055 116.475 ;
        RECT 102.690 116.115 102.945 116.785 ;
        RECT 103.125 115.805 103.410 116.605 ;
        RECT 103.590 116.525 103.840 117.115 ;
        RECT 104.040 117.760 104.360 118.090 ;
        RECT 104.540 117.875 105.200 118.355 ;
        RECT 105.400 117.965 106.250 118.135 ;
        RECT 104.040 116.865 104.230 117.760 ;
        RECT 104.550 117.435 105.210 117.705 ;
        RECT 104.880 117.375 105.210 117.435 ;
        RECT 104.400 117.205 104.730 117.265 ;
        RECT 105.400 117.205 105.570 117.965 ;
        RECT 106.810 117.895 107.130 118.355 ;
        RECT 107.330 117.715 107.580 118.145 ;
        RECT 107.870 117.915 108.280 118.355 ;
        RECT 108.450 117.975 109.465 118.175 ;
        RECT 105.740 117.545 106.990 117.715 ;
        RECT 105.740 117.425 106.070 117.545 ;
        RECT 104.400 117.035 106.300 117.205 ;
        RECT 104.040 116.695 105.960 116.865 ;
        RECT 104.040 116.675 104.360 116.695 ;
        RECT 103.590 116.015 103.920 116.525 ;
        RECT 104.190 116.065 104.360 116.675 ;
        RECT 106.130 116.525 106.300 117.035 ;
        RECT 106.470 116.965 106.650 117.375 ;
        RECT 106.820 116.785 106.990 117.545 ;
        RECT 104.530 115.805 104.860 116.495 ;
        RECT 105.090 116.355 106.300 116.525 ;
        RECT 106.470 116.475 106.990 116.785 ;
        RECT 107.160 117.375 107.580 117.715 ;
        RECT 107.870 117.375 108.280 117.705 ;
        RECT 107.160 116.605 107.350 117.375 ;
        RECT 108.450 117.245 108.620 117.975 ;
        RECT 109.765 117.805 109.935 118.135 ;
        RECT 110.105 117.975 110.435 118.355 ;
        RECT 108.790 117.425 109.140 117.795 ;
        RECT 108.450 117.205 108.870 117.245 ;
        RECT 107.520 117.035 108.870 117.205 ;
        RECT 107.520 116.875 107.770 117.035 ;
        RECT 108.280 116.605 108.530 116.865 ;
        RECT 107.160 116.355 108.530 116.605 ;
        RECT 105.090 116.065 105.330 116.355 ;
        RECT 106.130 116.275 106.300 116.355 ;
        RECT 105.530 115.805 105.950 116.185 ;
        RECT 106.130 116.025 106.760 116.275 ;
        RECT 107.230 115.805 107.560 116.185 ;
        RECT 107.730 116.065 107.900 116.355 ;
        RECT 108.700 116.190 108.870 117.035 ;
        RECT 109.320 116.865 109.540 117.735 ;
        RECT 109.765 117.615 110.460 117.805 ;
        RECT 109.040 116.485 109.540 116.865 ;
        RECT 109.710 116.815 110.120 117.435 ;
        RECT 110.290 116.645 110.460 117.615 ;
        RECT 109.765 116.475 110.460 116.645 ;
        RECT 108.080 115.805 108.460 116.185 ;
        RECT 108.700 116.020 109.530 116.190 ;
        RECT 109.765 115.975 109.935 116.475 ;
        RECT 110.105 115.805 110.435 116.305 ;
        RECT 110.650 115.975 110.875 118.095 ;
        RECT 111.045 117.975 111.375 118.355 ;
        RECT 111.545 117.805 111.715 118.095 ;
        RECT 111.050 117.635 111.715 117.805 ;
        RECT 111.050 116.645 111.280 117.635 ;
        RECT 112.955 117.535 113.165 118.355 ;
        RECT 113.335 117.555 113.665 118.185 ;
        RECT 111.450 116.815 111.800 117.465 ;
        RECT 113.335 116.955 113.585 117.555 ;
        RECT 113.835 117.535 114.065 118.355 ;
        RECT 114.275 117.630 114.565 118.355 ;
        RECT 115.285 117.805 115.455 118.185 ;
        RECT 115.635 117.975 115.965 118.355 ;
        RECT 115.285 117.635 115.950 117.805 ;
        RECT 116.145 117.680 116.405 118.185 ;
        RECT 113.755 117.115 114.085 117.365 ;
        RECT 115.215 117.085 115.545 117.455 ;
        RECT 115.780 117.380 115.950 117.635 ;
        RECT 115.780 117.050 116.065 117.380 ;
        RECT 111.050 116.475 111.715 116.645 ;
        RECT 111.045 115.805 111.375 116.305 ;
        RECT 111.545 115.975 111.715 116.475 ;
        RECT 112.955 115.805 113.165 116.945 ;
        RECT 113.335 115.975 113.665 116.955 ;
        RECT 113.835 115.805 114.065 116.945 ;
        RECT 114.275 115.805 114.565 116.970 ;
        RECT 115.780 116.905 115.950 117.050 ;
        RECT 115.285 116.735 115.950 116.905 ;
        RECT 116.235 116.880 116.405 117.680 ;
        RECT 117.035 117.585 120.545 118.355 ;
        RECT 120.720 117.810 126.065 118.355 ;
        RECT 115.285 115.975 115.455 116.735 ;
        RECT 115.635 115.805 115.965 116.565 ;
        RECT 116.135 115.975 116.405 116.880 ;
        RECT 117.035 116.895 118.725 117.415 ;
        RECT 118.895 117.065 120.545 117.585 ;
        RECT 117.035 115.805 120.545 116.895 ;
        RECT 122.310 116.240 122.660 117.490 ;
        RECT 124.140 116.980 124.480 117.810 ;
        RECT 126.235 117.605 127.445 118.355 ;
        RECT 126.235 116.895 126.755 117.435 ;
        RECT 126.925 117.065 127.445 117.605 ;
        RECT 120.720 115.805 126.065 116.240 ;
        RECT 126.235 115.805 127.445 116.895 ;
        RECT 14.370 115.635 127.530 115.805 ;
        RECT 14.455 114.545 15.665 115.635 ;
        RECT 14.455 113.835 14.975 114.375 ;
        RECT 15.145 114.005 15.665 114.545 ;
        RECT 15.835 114.545 17.045 115.635 ;
        RECT 17.215 114.545 20.725 115.635 ;
        RECT 20.985 114.705 21.155 115.465 ;
        RECT 21.335 114.875 21.665 115.635 ;
        RECT 15.835 114.005 16.355 114.545 ;
        RECT 16.525 113.835 17.045 114.375 ;
        RECT 17.215 114.025 18.905 114.545 ;
        RECT 20.985 114.535 21.650 114.705 ;
        RECT 21.835 114.560 22.105 115.465 ;
        RECT 21.480 114.390 21.650 114.535 ;
        RECT 19.075 113.855 20.725 114.375 ;
        RECT 20.915 113.985 21.245 114.355 ;
        RECT 21.480 114.060 21.765 114.390 ;
        RECT 14.455 113.085 15.665 113.835 ;
        RECT 15.835 113.085 17.045 113.835 ;
        RECT 17.215 113.085 20.725 113.855 ;
        RECT 21.480 113.805 21.650 114.060 ;
        RECT 20.985 113.635 21.650 113.805 ;
        RECT 21.935 113.760 22.105 114.560 ;
        RECT 22.335 114.495 22.545 115.635 ;
        RECT 22.715 114.485 23.045 115.465 ;
        RECT 23.215 114.495 23.445 115.635 ;
        RECT 20.985 113.255 21.155 113.635 ;
        RECT 21.335 113.085 21.665 113.465 ;
        RECT 21.845 113.255 22.105 113.760 ;
        RECT 22.335 113.085 22.545 113.905 ;
        RECT 22.715 113.885 22.965 114.485 ;
        RECT 24.115 114.470 24.405 115.635 ;
        RECT 24.665 114.965 24.835 115.465 ;
        RECT 25.005 115.135 25.335 115.635 ;
        RECT 24.665 114.795 25.330 114.965 ;
        RECT 23.135 114.075 23.465 114.325 ;
        RECT 24.580 113.975 24.930 114.625 ;
        RECT 22.715 113.255 23.045 113.885 ;
        RECT 23.215 113.085 23.445 113.905 ;
        RECT 24.115 113.085 24.405 113.810 ;
        RECT 25.100 113.805 25.330 114.795 ;
        RECT 24.665 113.635 25.330 113.805 ;
        RECT 24.665 113.345 24.835 113.635 ;
        RECT 25.005 113.085 25.335 113.465 ;
        RECT 25.505 113.345 25.730 115.465 ;
        RECT 25.945 115.135 26.275 115.635 ;
        RECT 26.445 114.965 26.615 115.465 ;
        RECT 26.850 115.250 27.680 115.420 ;
        RECT 27.920 115.255 28.300 115.635 ;
        RECT 25.920 114.795 26.615 114.965 ;
        RECT 25.920 113.825 26.090 114.795 ;
        RECT 26.260 114.005 26.670 114.625 ;
        RECT 26.840 114.575 27.340 114.955 ;
        RECT 25.920 113.635 26.615 113.825 ;
        RECT 26.840 113.705 27.060 114.575 ;
        RECT 27.510 114.405 27.680 115.250 ;
        RECT 28.480 115.085 28.650 115.375 ;
        RECT 28.820 115.255 29.150 115.635 ;
        RECT 29.620 115.165 30.250 115.415 ;
        RECT 30.430 115.255 30.850 115.635 ;
        RECT 30.080 115.085 30.250 115.165 ;
        RECT 31.050 115.085 31.290 115.375 ;
        RECT 27.850 114.835 29.220 115.085 ;
        RECT 27.850 114.575 28.100 114.835 ;
        RECT 28.610 114.405 28.860 114.565 ;
        RECT 27.510 114.235 28.860 114.405 ;
        RECT 27.510 114.195 27.930 114.235 ;
        RECT 27.240 113.645 27.590 114.015 ;
        RECT 25.945 113.085 26.275 113.465 ;
        RECT 26.445 113.305 26.615 113.635 ;
        RECT 27.760 113.465 27.930 114.195 ;
        RECT 29.030 114.065 29.220 114.835 ;
        RECT 28.100 113.735 28.510 114.065 ;
        RECT 28.800 113.725 29.220 114.065 ;
        RECT 29.390 114.655 29.910 114.965 ;
        RECT 30.080 114.915 31.290 115.085 ;
        RECT 31.520 114.945 31.850 115.635 ;
        RECT 29.390 113.895 29.560 114.655 ;
        RECT 29.730 114.065 29.910 114.475 ;
        RECT 30.080 114.405 30.250 114.915 ;
        RECT 32.020 114.765 32.190 115.375 ;
        RECT 32.460 114.915 32.790 115.425 ;
        RECT 32.020 114.745 32.340 114.765 ;
        RECT 30.420 114.575 32.340 114.745 ;
        RECT 30.080 114.235 31.980 114.405 ;
        RECT 30.310 113.895 30.640 114.015 ;
        RECT 29.390 113.725 30.640 113.895 ;
        RECT 26.915 113.265 27.930 113.465 ;
        RECT 28.100 113.085 28.510 113.525 ;
        RECT 28.800 113.295 29.050 113.725 ;
        RECT 29.250 113.085 29.570 113.545 ;
        RECT 30.810 113.475 30.980 114.235 ;
        RECT 31.650 114.175 31.980 114.235 ;
        RECT 31.170 114.005 31.500 114.065 ;
        RECT 31.170 113.735 31.830 114.005 ;
        RECT 32.150 113.680 32.340 114.575 ;
        RECT 30.130 113.305 30.980 113.475 ;
        RECT 31.180 113.085 31.840 113.565 ;
        RECT 32.020 113.350 32.340 113.680 ;
        RECT 32.540 114.325 32.790 114.915 ;
        RECT 32.970 114.835 33.255 115.635 ;
        RECT 33.435 115.295 33.690 115.325 ;
        RECT 33.435 115.125 33.775 115.295 ;
        RECT 33.435 114.655 33.690 115.125 ;
        RECT 32.540 113.995 33.340 114.325 ;
        RECT 32.540 113.345 32.790 113.995 ;
        RECT 33.510 113.795 33.690 114.655 ;
        RECT 34.755 114.495 34.965 115.635 ;
        RECT 35.135 114.485 35.465 115.465 ;
        RECT 35.635 114.495 35.865 115.635 ;
        RECT 36.625 114.705 36.795 115.465 ;
        RECT 36.975 114.875 37.305 115.635 ;
        RECT 36.625 114.535 37.290 114.705 ;
        RECT 37.475 114.560 37.745 115.465 ;
        RECT 32.970 113.085 33.255 113.545 ;
        RECT 33.435 113.265 33.690 113.795 ;
        RECT 34.755 113.085 34.965 113.905 ;
        RECT 35.135 113.885 35.385 114.485 ;
        RECT 37.120 114.390 37.290 114.535 ;
        RECT 35.555 114.075 35.885 114.325 ;
        RECT 36.555 113.985 36.885 114.355 ;
        RECT 37.120 114.060 37.405 114.390 ;
        RECT 35.135 113.255 35.465 113.885 ;
        RECT 35.635 113.085 35.865 113.905 ;
        RECT 37.120 113.805 37.290 114.060 ;
        RECT 36.625 113.635 37.290 113.805 ;
        RECT 37.575 113.760 37.745 114.560 ;
        RECT 36.625 113.255 36.795 113.635 ;
        RECT 36.975 113.085 37.305 113.465 ;
        RECT 37.485 113.255 37.745 113.760 ;
        RECT 38.835 114.560 39.105 115.465 ;
        RECT 39.275 114.875 39.605 115.635 ;
        RECT 39.785 114.705 39.955 115.465 ;
        RECT 38.835 113.760 39.005 114.560 ;
        RECT 39.290 114.535 39.955 114.705 ;
        RECT 40.215 114.545 43.725 115.635 ;
        RECT 39.290 114.390 39.460 114.535 ;
        RECT 39.175 114.060 39.460 114.390 ;
        RECT 39.290 113.805 39.460 114.060 ;
        RECT 39.695 113.985 40.025 114.355 ;
        RECT 40.215 114.025 41.905 114.545 ;
        RECT 43.955 114.495 44.165 115.635 ;
        RECT 44.335 114.485 44.665 115.465 ;
        RECT 44.835 114.495 45.065 115.635 ;
        RECT 45.280 114.495 45.615 115.465 ;
        RECT 45.785 114.495 45.955 115.635 ;
        RECT 46.125 115.295 48.155 115.465 ;
        RECT 42.075 113.855 43.725 114.375 ;
        RECT 38.835 113.255 39.095 113.760 ;
        RECT 39.290 113.635 39.955 113.805 ;
        RECT 39.275 113.085 39.605 113.465 ;
        RECT 39.785 113.255 39.955 113.635 ;
        RECT 40.215 113.085 43.725 113.855 ;
        RECT 43.955 113.085 44.165 113.905 ;
        RECT 44.335 113.885 44.585 114.485 ;
        RECT 44.755 114.075 45.085 114.325 ;
        RECT 44.335 113.255 44.665 113.885 ;
        RECT 44.835 113.085 45.065 113.905 ;
        RECT 45.280 113.825 45.450 114.495 ;
        RECT 46.125 114.325 46.295 115.295 ;
        RECT 45.620 113.995 45.875 114.325 ;
        RECT 46.100 113.995 46.295 114.325 ;
        RECT 46.465 114.955 47.590 115.125 ;
        RECT 45.705 113.825 45.875 113.995 ;
        RECT 46.465 113.825 46.635 114.955 ;
        RECT 45.280 113.255 45.535 113.825 ;
        RECT 45.705 113.655 46.635 113.825 ;
        RECT 46.805 114.615 47.815 114.785 ;
        RECT 46.805 113.815 46.975 114.615 ;
        RECT 47.180 113.935 47.455 114.415 ;
        RECT 47.175 113.765 47.455 113.935 ;
        RECT 46.460 113.620 46.635 113.655 ;
        RECT 45.705 113.085 46.035 113.485 ;
        RECT 46.460 113.255 46.990 113.620 ;
        RECT 47.180 113.255 47.455 113.765 ;
        RECT 47.625 113.255 47.815 114.615 ;
        RECT 47.985 114.630 48.155 115.295 ;
        RECT 48.325 114.875 48.495 115.635 ;
        RECT 48.730 114.875 49.245 115.285 ;
        RECT 47.985 114.440 48.735 114.630 ;
        RECT 48.905 114.065 49.245 114.875 ;
        RECT 49.875 114.470 50.165 115.635 ;
        RECT 50.335 114.545 52.005 115.635 ;
        RECT 52.265 114.705 52.435 115.465 ;
        RECT 52.615 114.875 52.945 115.635 ;
        RECT 48.015 113.895 49.245 114.065 ;
        RECT 50.335 114.025 51.085 114.545 ;
        RECT 52.265 114.535 52.930 114.705 ;
        RECT 53.115 114.560 53.385 115.465 ;
        RECT 52.760 114.390 52.930 114.535 ;
        RECT 47.995 113.085 48.505 113.620 ;
        RECT 48.725 113.290 48.970 113.895 ;
        RECT 51.255 113.855 52.005 114.375 ;
        RECT 52.195 113.985 52.525 114.355 ;
        RECT 52.760 114.060 53.045 114.390 ;
        RECT 49.875 113.085 50.165 113.810 ;
        RECT 50.335 113.085 52.005 113.855 ;
        RECT 52.760 113.805 52.930 114.060 ;
        RECT 52.265 113.635 52.930 113.805 ;
        RECT 53.215 113.760 53.385 114.560 ;
        RECT 53.555 114.545 54.765 115.635 ;
        RECT 54.940 115.200 60.285 115.635 ;
        RECT 60.460 115.200 65.805 115.635 ;
        RECT 53.555 114.005 54.075 114.545 ;
        RECT 54.245 113.835 54.765 114.375 ;
        RECT 56.530 113.950 56.880 115.200 ;
        RECT 52.265 113.255 52.435 113.635 ;
        RECT 52.615 113.085 52.945 113.465 ;
        RECT 53.125 113.255 53.385 113.760 ;
        RECT 53.555 113.085 54.765 113.835 ;
        RECT 58.360 113.630 58.700 114.460 ;
        RECT 62.050 113.950 62.400 115.200 ;
        RECT 66.015 114.495 66.245 115.635 ;
        RECT 66.415 114.485 66.745 115.465 ;
        RECT 66.915 114.495 67.125 115.635 ;
        RECT 67.905 114.705 68.075 115.465 ;
        RECT 68.255 114.875 68.585 115.635 ;
        RECT 67.905 114.535 68.570 114.705 ;
        RECT 68.755 114.560 69.025 115.465 ;
        RECT 70.120 115.200 75.465 115.635 ;
        RECT 63.880 113.630 64.220 114.460 ;
        RECT 65.995 114.075 66.325 114.325 ;
        RECT 54.940 113.085 60.285 113.630 ;
        RECT 60.460 113.085 65.805 113.630 ;
        RECT 66.015 113.085 66.245 113.905 ;
        RECT 66.495 113.885 66.745 114.485 ;
        RECT 68.400 114.390 68.570 114.535 ;
        RECT 67.835 113.985 68.165 114.355 ;
        RECT 68.400 114.060 68.685 114.390 ;
        RECT 66.415 113.255 66.745 113.885 ;
        RECT 66.915 113.085 67.125 113.905 ;
        RECT 68.400 113.805 68.570 114.060 ;
        RECT 67.905 113.635 68.570 113.805 ;
        RECT 68.855 113.760 69.025 114.560 ;
        RECT 71.710 113.950 72.060 115.200 ;
        RECT 75.635 114.470 75.925 115.635 ;
        RECT 77.390 115.295 77.645 115.325 ;
        RECT 77.305 115.125 77.645 115.295 ;
        RECT 77.390 114.655 77.645 115.125 ;
        RECT 77.825 114.835 78.110 115.635 ;
        RECT 78.290 114.915 78.620 115.425 ;
        RECT 67.905 113.255 68.075 113.635 ;
        RECT 68.255 113.085 68.585 113.465 ;
        RECT 68.765 113.255 69.025 113.760 ;
        RECT 73.540 113.630 73.880 114.460 ;
        RECT 70.120 113.085 75.465 113.630 ;
        RECT 75.635 113.085 75.925 113.810 ;
        RECT 77.390 113.795 77.570 114.655 ;
        RECT 78.290 114.325 78.540 114.915 ;
        RECT 78.890 114.765 79.060 115.375 ;
        RECT 79.230 114.945 79.560 115.635 ;
        RECT 79.790 115.085 80.030 115.375 ;
        RECT 80.230 115.255 80.650 115.635 ;
        RECT 80.830 115.165 81.460 115.415 ;
        RECT 81.930 115.255 82.260 115.635 ;
        RECT 80.830 115.085 81.000 115.165 ;
        RECT 82.430 115.085 82.600 115.375 ;
        RECT 82.780 115.255 83.160 115.635 ;
        RECT 83.400 115.250 84.230 115.420 ;
        RECT 79.790 114.915 81.000 115.085 ;
        RECT 77.740 113.995 78.540 114.325 ;
        RECT 77.390 113.265 77.645 113.795 ;
        RECT 77.825 113.085 78.110 113.545 ;
        RECT 78.290 113.345 78.540 113.995 ;
        RECT 78.740 114.745 79.060 114.765 ;
        RECT 78.740 114.575 80.660 114.745 ;
        RECT 78.740 113.680 78.930 114.575 ;
        RECT 80.830 114.405 81.000 114.915 ;
        RECT 81.170 114.655 81.690 114.965 ;
        RECT 79.100 114.235 81.000 114.405 ;
        RECT 79.100 114.175 79.430 114.235 ;
        RECT 79.580 114.005 79.910 114.065 ;
        RECT 79.250 113.735 79.910 114.005 ;
        RECT 78.740 113.350 79.060 113.680 ;
        RECT 79.240 113.085 79.900 113.565 ;
        RECT 80.100 113.475 80.270 114.235 ;
        RECT 81.170 114.065 81.350 114.475 ;
        RECT 80.440 113.895 80.770 114.015 ;
        RECT 81.520 113.895 81.690 114.655 ;
        RECT 80.440 113.725 81.690 113.895 ;
        RECT 81.860 114.835 83.230 115.085 ;
        RECT 81.860 114.065 82.050 114.835 ;
        RECT 82.980 114.575 83.230 114.835 ;
        RECT 82.220 114.405 82.470 114.565 ;
        RECT 83.400 114.405 83.570 115.250 ;
        RECT 84.465 114.965 84.635 115.465 ;
        RECT 84.805 115.135 85.135 115.635 ;
        RECT 83.740 114.575 84.240 114.955 ;
        RECT 84.465 114.795 85.160 114.965 ;
        RECT 82.220 114.235 83.570 114.405 ;
        RECT 83.150 114.195 83.570 114.235 ;
        RECT 81.860 113.725 82.280 114.065 ;
        RECT 82.570 113.735 82.980 114.065 ;
        RECT 80.100 113.305 80.950 113.475 ;
        RECT 81.510 113.085 81.830 113.545 ;
        RECT 82.030 113.295 82.280 113.725 ;
        RECT 82.570 113.085 82.980 113.525 ;
        RECT 83.150 113.465 83.320 114.195 ;
        RECT 83.490 113.645 83.840 114.015 ;
        RECT 84.020 113.705 84.240 114.575 ;
        RECT 84.410 114.005 84.820 114.625 ;
        RECT 84.990 113.825 85.160 114.795 ;
        RECT 84.465 113.635 85.160 113.825 ;
        RECT 83.150 113.265 84.165 113.465 ;
        RECT 84.465 113.305 84.635 113.635 ;
        RECT 84.805 113.085 85.135 113.465 ;
        RECT 85.350 113.345 85.575 115.465 ;
        RECT 85.745 115.135 86.075 115.635 ;
        RECT 86.245 114.965 86.415 115.465 ;
        RECT 85.750 114.795 86.415 114.965 ;
        RECT 87.225 114.965 87.395 115.465 ;
        RECT 87.565 115.135 87.895 115.635 ;
        RECT 87.225 114.795 87.890 114.965 ;
        RECT 85.750 113.805 85.980 114.795 ;
        RECT 86.150 113.975 86.500 114.625 ;
        RECT 87.140 113.975 87.490 114.625 ;
        RECT 87.660 113.805 87.890 114.795 ;
        RECT 85.750 113.635 86.415 113.805 ;
        RECT 85.745 113.085 86.075 113.465 ;
        RECT 86.245 113.345 86.415 113.635 ;
        RECT 87.225 113.635 87.890 113.805 ;
        RECT 87.225 113.345 87.395 113.635 ;
        RECT 87.565 113.085 87.895 113.465 ;
        RECT 88.065 113.345 88.290 115.465 ;
        RECT 88.505 115.135 88.835 115.635 ;
        RECT 89.005 114.965 89.175 115.465 ;
        RECT 89.410 115.250 90.240 115.420 ;
        RECT 90.480 115.255 90.860 115.635 ;
        RECT 88.480 114.795 89.175 114.965 ;
        RECT 88.480 113.825 88.650 114.795 ;
        RECT 88.820 114.005 89.230 114.625 ;
        RECT 89.400 114.575 89.900 114.955 ;
        RECT 88.480 113.635 89.175 113.825 ;
        RECT 89.400 113.705 89.620 114.575 ;
        RECT 90.070 114.405 90.240 115.250 ;
        RECT 91.040 115.085 91.210 115.375 ;
        RECT 91.380 115.255 91.710 115.635 ;
        RECT 92.180 115.165 92.810 115.415 ;
        RECT 92.990 115.255 93.410 115.635 ;
        RECT 92.640 115.085 92.810 115.165 ;
        RECT 93.610 115.085 93.850 115.375 ;
        RECT 90.410 114.835 91.780 115.085 ;
        RECT 90.410 114.575 90.660 114.835 ;
        RECT 91.170 114.405 91.420 114.565 ;
        RECT 90.070 114.235 91.420 114.405 ;
        RECT 90.070 114.195 90.490 114.235 ;
        RECT 89.800 113.645 90.150 114.015 ;
        RECT 88.505 113.085 88.835 113.465 ;
        RECT 89.005 113.305 89.175 113.635 ;
        RECT 90.320 113.465 90.490 114.195 ;
        RECT 91.590 114.065 91.780 114.835 ;
        RECT 90.660 113.735 91.070 114.065 ;
        RECT 91.360 113.725 91.780 114.065 ;
        RECT 91.950 114.655 92.470 114.965 ;
        RECT 92.640 114.915 93.850 115.085 ;
        RECT 94.080 114.945 94.410 115.635 ;
        RECT 91.950 113.895 92.120 114.655 ;
        RECT 92.290 114.065 92.470 114.475 ;
        RECT 92.640 114.405 92.810 114.915 ;
        RECT 94.580 114.765 94.750 115.375 ;
        RECT 95.020 114.915 95.350 115.425 ;
        RECT 94.580 114.745 94.900 114.765 ;
        RECT 92.980 114.575 94.900 114.745 ;
        RECT 92.640 114.235 94.540 114.405 ;
        RECT 92.870 113.895 93.200 114.015 ;
        RECT 91.950 113.725 93.200 113.895 ;
        RECT 89.475 113.265 90.490 113.465 ;
        RECT 90.660 113.085 91.070 113.525 ;
        RECT 91.360 113.295 91.610 113.725 ;
        RECT 91.810 113.085 92.130 113.545 ;
        RECT 93.370 113.475 93.540 114.235 ;
        RECT 94.210 114.175 94.540 114.235 ;
        RECT 93.730 114.005 94.060 114.065 ;
        RECT 93.730 113.735 94.390 114.005 ;
        RECT 94.710 113.680 94.900 114.575 ;
        RECT 92.690 113.305 93.540 113.475 ;
        RECT 93.740 113.085 94.400 113.565 ;
        RECT 94.580 113.350 94.900 113.680 ;
        RECT 95.100 114.325 95.350 114.915 ;
        RECT 95.530 114.835 95.815 115.635 ;
        RECT 95.995 115.295 96.250 115.325 ;
        RECT 95.995 115.125 96.335 115.295 ;
        RECT 95.995 114.655 96.250 115.125 ;
        RECT 95.100 113.995 95.900 114.325 ;
        RECT 95.100 113.345 95.350 113.995 ;
        RECT 96.070 113.795 96.250 114.655 ;
        RECT 97.255 114.545 99.845 115.635 ;
        RECT 100.015 114.560 100.285 115.465 ;
        RECT 100.455 114.875 100.785 115.635 ;
        RECT 100.965 114.705 101.135 115.465 ;
        RECT 97.255 114.025 98.465 114.545 ;
        RECT 98.635 113.855 99.845 114.375 ;
        RECT 95.530 113.085 95.815 113.545 ;
        RECT 95.995 113.265 96.250 113.795 ;
        RECT 97.255 113.085 99.845 113.855 ;
        RECT 100.015 113.760 100.185 114.560 ;
        RECT 100.470 114.535 101.135 114.705 ;
        RECT 100.470 114.390 100.640 114.535 ;
        RECT 101.395 114.470 101.685 115.635 ;
        RECT 102.320 115.200 107.665 115.635 ;
        RECT 100.355 114.060 100.640 114.390 ;
        RECT 100.470 113.805 100.640 114.060 ;
        RECT 100.875 113.985 101.205 114.355 ;
        RECT 103.910 113.950 104.260 115.200 ;
        RECT 107.925 114.705 108.095 115.465 ;
        RECT 108.275 114.875 108.605 115.635 ;
        RECT 107.925 114.535 108.590 114.705 ;
        RECT 108.775 114.560 109.045 115.465 ;
        RECT 100.015 113.255 100.275 113.760 ;
        RECT 100.470 113.635 101.135 113.805 ;
        RECT 100.455 113.085 100.785 113.465 ;
        RECT 100.965 113.255 101.135 113.635 ;
        RECT 101.395 113.085 101.685 113.810 ;
        RECT 105.740 113.630 106.080 114.460 ;
        RECT 108.420 114.390 108.590 114.535 ;
        RECT 107.855 113.985 108.185 114.355 ;
        RECT 108.420 114.060 108.705 114.390 ;
        RECT 108.420 113.805 108.590 114.060 ;
        RECT 107.925 113.635 108.590 113.805 ;
        RECT 108.875 113.760 109.045 114.560 ;
        RECT 109.215 114.545 110.885 115.635 ;
        RECT 111.055 114.875 111.570 115.285 ;
        RECT 111.805 114.875 111.975 115.635 ;
        RECT 112.145 115.295 114.175 115.465 ;
        RECT 109.215 114.025 109.965 114.545 ;
        RECT 110.135 113.855 110.885 114.375 ;
        RECT 111.055 114.065 111.395 114.875 ;
        RECT 112.145 114.630 112.315 115.295 ;
        RECT 112.710 114.955 113.835 115.125 ;
        RECT 111.565 114.440 112.315 114.630 ;
        RECT 112.485 114.615 113.495 114.785 ;
        RECT 111.055 113.895 112.285 114.065 ;
        RECT 102.320 113.085 107.665 113.630 ;
        RECT 107.925 113.255 108.095 113.635 ;
        RECT 108.275 113.085 108.605 113.465 ;
        RECT 108.785 113.255 109.045 113.760 ;
        RECT 109.215 113.085 110.885 113.855 ;
        RECT 111.330 113.290 111.575 113.895 ;
        RECT 111.795 113.085 112.305 113.620 ;
        RECT 112.485 113.255 112.675 114.615 ;
        RECT 112.845 114.275 113.120 114.415 ;
        RECT 112.845 114.105 113.125 114.275 ;
        RECT 112.845 113.255 113.120 114.105 ;
        RECT 113.325 113.815 113.495 114.615 ;
        RECT 113.665 113.825 113.835 114.955 ;
        RECT 114.005 114.325 114.175 115.295 ;
        RECT 114.345 114.495 114.515 115.635 ;
        RECT 114.685 114.495 115.020 115.465 ;
        RECT 115.200 115.200 120.545 115.635 ;
        RECT 120.720 115.200 126.065 115.635 ;
        RECT 114.005 113.995 114.200 114.325 ;
        RECT 114.425 113.995 114.680 114.325 ;
        RECT 114.425 113.825 114.595 113.995 ;
        RECT 114.850 113.825 115.020 114.495 ;
        RECT 116.790 113.950 117.140 115.200 ;
        RECT 113.665 113.655 114.595 113.825 ;
        RECT 113.665 113.620 113.840 113.655 ;
        RECT 113.310 113.255 113.840 113.620 ;
        RECT 114.265 113.085 114.595 113.485 ;
        RECT 114.765 113.255 115.020 113.825 ;
        RECT 118.620 113.630 118.960 114.460 ;
        RECT 122.310 113.950 122.660 115.200 ;
        RECT 126.235 114.545 127.445 115.635 ;
        RECT 124.140 113.630 124.480 114.460 ;
        RECT 126.235 114.005 126.755 114.545 ;
        RECT 126.925 113.835 127.445 114.375 ;
        RECT 115.200 113.085 120.545 113.630 ;
        RECT 120.720 113.085 126.065 113.630 ;
        RECT 126.235 113.085 127.445 113.835 ;
        RECT 14.370 112.915 127.530 113.085 ;
        RECT 14.455 112.165 15.665 112.915 ;
        RECT 16.145 112.445 16.315 112.915 ;
        RECT 16.485 112.265 16.815 112.745 ;
        RECT 16.985 112.445 17.155 112.915 ;
        RECT 17.325 112.265 17.655 112.745 ;
        RECT 14.455 111.625 14.975 112.165 ;
        RECT 15.890 112.095 17.655 112.265 ;
        RECT 17.825 112.105 17.995 112.915 ;
        RECT 18.195 112.535 19.265 112.705 ;
        RECT 18.195 112.180 18.515 112.535 ;
        RECT 15.145 111.455 15.665 111.995 ;
        RECT 14.455 110.365 15.665 111.455 ;
        RECT 15.890 111.545 16.300 112.095 ;
        RECT 18.190 111.925 18.515 112.180 ;
        RECT 16.485 111.715 18.515 111.925 ;
        RECT 18.170 111.705 18.515 111.715 ;
        RECT 18.685 111.965 18.925 112.365 ;
        RECT 19.095 112.305 19.265 112.535 ;
        RECT 19.435 112.475 19.625 112.915 ;
        RECT 19.795 112.465 20.745 112.745 ;
        RECT 20.965 112.555 21.315 112.725 ;
        RECT 19.095 112.135 19.625 112.305 ;
        RECT 15.890 111.375 17.615 111.545 ;
        RECT 16.145 110.365 16.315 111.205 ;
        RECT 16.525 110.535 16.775 111.375 ;
        RECT 16.985 110.365 17.155 111.205 ;
        RECT 17.325 110.535 17.615 111.375 ;
        RECT 17.825 110.365 17.995 111.425 ;
        RECT 18.170 111.085 18.340 111.705 ;
        RECT 18.685 111.595 19.225 111.965 ;
        RECT 19.405 111.855 19.625 112.135 ;
        RECT 19.795 111.685 19.965 112.465 ;
        RECT 19.560 111.515 19.965 111.685 ;
        RECT 20.135 111.675 20.485 112.295 ;
        RECT 19.560 111.425 19.730 111.515 ;
        RECT 20.655 111.505 20.865 112.295 ;
        RECT 18.510 111.255 19.730 111.425 ;
        RECT 20.190 111.345 20.865 111.505 ;
        RECT 18.170 110.915 18.970 111.085 ;
        RECT 18.290 110.365 18.620 110.745 ;
        RECT 18.800 110.625 18.970 110.915 ;
        RECT 19.560 110.875 19.730 111.255 ;
        RECT 19.900 111.335 20.865 111.345 ;
        RECT 21.055 112.165 21.315 112.555 ;
        RECT 21.525 112.455 21.855 112.915 ;
        RECT 22.730 112.525 23.585 112.695 ;
        RECT 23.790 112.525 24.285 112.695 ;
        RECT 24.455 112.555 24.785 112.915 ;
        RECT 21.055 111.475 21.225 112.165 ;
        RECT 21.395 111.815 21.565 111.995 ;
        RECT 21.735 111.985 22.525 112.235 ;
        RECT 22.730 111.815 22.900 112.525 ;
        RECT 23.070 112.015 23.425 112.235 ;
        RECT 21.395 111.645 23.085 111.815 ;
        RECT 19.900 111.045 20.360 111.335 ;
        RECT 21.055 111.305 22.555 111.475 ;
        RECT 21.055 111.165 21.225 111.305 ;
        RECT 20.665 110.995 21.225 111.165 ;
        RECT 19.140 110.365 19.390 110.825 ;
        RECT 19.560 110.535 20.430 110.875 ;
        RECT 20.665 110.535 20.835 110.995 ;
        RECT 21.670 110.965 22.745 111.135 ;
        RECT 21.005 110.365 21.375 110.825 ;
        RECT 21.670 110.625 21.840 110.965 ;
        RECT 22.010 110.365 22.340 110.795 ;
        RECT 22.575 110.625 22.745 110.965 ;
        RECT 22.915 110.865 23.085 111.645 ;
        RECT 23.255 111.425 23.425 112.015 ;
        RECT 23.595 111.615 23.945 112.235 ;
        RECT 23.255 111.035 23.720 111.425 ;
        RECT 24.115 111.165 24.285 112.525 ;
        RECT 24.455 111.335 24.915 112.385 ;
        RECT 23.890 110.995 24.285 111.165 ;
        RECT 23.890 110.865 24.060 110.995 ;
        RECT 22.915 110.535 23.595 110.865 ;
        RECT 23.810 110.535 24.060 110.865 ;
        RECT 24.230 110.365 24.480 110.825 ;
        RECT 24.650 110.550 24.975 111.335 ;
        RECT 25.145 110.535 25.315 112.655 ;
        RECT 25.485 112.535 25.815 112.915 ;
        RECT 25.985 112.365 26.240 112.655 ;
        RECT 25.490 112.195 26.240 112.365 ;
        RECT 25.490 111.205 25.720 112.195 ;
        RECT 26.415 112.145 28.085 112.915 ;
        RECT 28.260 112.370 33.605 112.915 ;
        RECT 25.890 111.375 26.240 112.025 ;
        RECT 26.415 111.455 27.165 111.975 ;
        RECT 27.335 111.625 28.085 112.145 ;
        RECT 25.490 111.035 26.240 111.205 ;
        RECT 25.485 110.365 25.815 110.865 ;
        RECT 25.985 110.535 26.240 111.035 ;
        RECT 26.415 110.365 28.085 111.455 ;
        RECT 29.850 110.800 30.200 112.050 ;
        RECT 31.680 111.540 32.020 112.370 ;
        RECT 33.835 112.095 34.045 112.915 ;
        RECT 34.215 112.115 34.545 112.745 ;
        RECT 34.215 111.515 34.465 112.115 ;
        RECT 34.715 112.095 34.945 112.915 ;
        RECT 35.155 112.145 36.825 112.915 ;
        RECT 36.995 112.190 37.285 112.915 ;
        RECT 38.005 112.435 38.305 112.915 ;
        RECT 38.475 112.265 38.735 112.720 ;
        RECT 38.905 112.435 39.165 112.915 ;
        RECT 39.345 112.265 39.605 112.720 ;
        RECT 39.775 112.435 40.025 112.915 ;
        RECT 40.205 112.265 40.465 112.720 ;
        RECT 40.635 112.435 40.885 112.915 ;
        RECT 41.065 112.265 41.325 112.720 ;
        RECT 41.495 112.435 41.740 112.915 ;
        RECT 41.910 112.265 42.185 112.720 ;
        RECT 42.355 112.435 42.600 112.915 ;
        RECT 42.770 112.265 43.030 112.720 ;
        RECT 43.200 112.435 43.460 112.915 ;
        RECT 43.630 112.265 43.890 112.720 ;
        RECT 44.060 112.435 44.320 112.915 ;
        RECT 44.490 112.265 44.750 112.720 ;
        RECT 44.920 112.355 45.180 112.915 ;
        RECT 34.635 111.675 34.965 111.925 ;
        RECT 28.260 110.365 33.605 110.800 ;
        RECT 33.835 110.365 34.045 111.505 ;
        RECT 34.215 110.535 34.545 111.515 ;
        RECT 34.715 110.365 34.945 111.505 ;
        RECT 35.155 111.455 35.905 111.975 ;
        RECT 36.075 111.625 36.825 112.145 ;
        RECT 38.005 112.095 44.750 112.265 ;
        RECT 35.155 110.365 36.825 111.455 ;
        RECT 36.995 110.365 37.285 111.530 ;
        RECT 38.005 111.505 39.170 112.095 ;
        RECT 45.350 111.925 45.600 112.735 ;
        RECT 45.780 112.390 46.040 112.915 ;
        RECT 46.210 111.925 46.460 112.735 ;
        RECT 46.640 112.405 46.945 112.915 ;
        RECT 39.340 111.675 46.460 111.925 ;
        RECT 46.630 111.675 46.945 112.235 ;
        RECT 48.035 112.145 51.545 112.915 ;
        RECT 51.720 112.370 57.065 112.915 ;
        RECT 57.240 112.370 62.585 112.915 ;
        RECT 38.005 111.280 44.750 111.505 ;
        RECT 38.005 110.365 38.275 111.110 ;
        RECT 38.445 110.540 38.735 111.280 ;
        RECT 39.345 111.265 44.750 111.280 ;
        RECT 38.905 110.370 39.160 111.095 ;
        RECT 39.345 110.540 39.605 111.265 ;
        RECT 39.775 110.370 40.020 111.095 ;
        RECT 40.205 110.540 40.465 111.265 ;
        RECT 40.635 110.370 40.880 111.095 ;
        RECT 41.065 110.540 41.325 111.265 ;
        RECT 41.495 110.370 41.740 111.095 ;
        RECT 41.910 110.540 42.170 111.265 ;
        RECT 42.340 110.370 42.600 111.095 ;
        RECT 42.770 110.540 43.030 111.265 ;
        RECT 43.200 110.370 43.460 111.095 ;
        RECT 43.630 110.540 43.890 111.265 ;
        RECT 44.060 110.370 44.320 111.095 ;
        RECT 44.490 110.540 44.750 111.265 ;
        RECT 44.920 110.370 45.180 111.165 ;
        RECT 45.350 110.540 45.600 111.675 ;
        RECT 38.905 110.365 45.180 110.370 ;
        RECT 45.780 110.365 46.040 111.175 ;
        RECT 46.215 110.535 46.460 111.675 ;
        RECT 48.035 111.455 49.725 111.975 ;
        RECT 49.895 111.625 51.545 112.145 ;
        RECT 46.640 110.365 46.935 111.175 ;
        RECT 48.035 110.365 51.545 111.455 ;
        RECT 53.310 110.800 53.660 112.050 ;
        RECT 55.140 111.540 55.480 112.370 ;
        RECT 58.830 110.800 59.180 112.050 ;
        RECT 60.660 111.540 61.000 112.370 ;
        RECT 62.755 112.190 63.045 112.915 ;
        RECT 63.680 112.370 69.025 112.915 ;
        RECT 69.200 112.370 74.545 112.915 ;
        RECT 74.720 112.370 80.065 112.915 ;
        RECT 51.720 110.365 57.065 110.800 ;
        RECT 57.240 110.365 62.585 110.800 ;
        RECT 62.755 110.365 63.045 111.530 ;
        RECT 65.270 110.800 65.620 112.050 ;
        RECT 67.100 111.540 67.440 112.370 ;
        RECT 70.790 110.800 71.140 112.050 ;
        RECT 72.620 111.540 72.960 112.370 ;
        RECT 76.310 110.800 76.660 112.050 ;
        RECT 78.140 111.540 78.480 112.370 ;
        RECT 80.295 112.095 80.505 112.915 ;
        RECT 80.675 112.115 81.005 112.745 ;
        RECT 80.675 111.515 80.925 112.115 ;
        RECT 81.175 112.095 81.405 112.915 ;
        RECT 81.615 112.165 82.825 112.915 ;
        RECT 83.000 112.370 88.345 112.915 ;
        RECT 81.095 111.675 81.425 111.925 ;
        RECT 63.680 110.365 69.025 110.800 ;
        RECT 69.200 110.365 74.545 110.800 ;
        RECT 74.720 110.365 80.065 110.800 ;
        RECT 80.295 110.365 80.505 111.505 ;
        RECT 80.675 110.535 81.005 111.515 ;
        RECT 81.175 110.365 81.405 111.505 ;
        RECT 81.615 111.455 82.135 111.995 ;
        RECT 82.305 111.625 82.825 112.165 ;
        RECT 81.615 110.365 82.825 111.455 ;
        RECT 84.590 110.800 84.940 112.050 ;
        RECT 86.420 111.540 86.760 112.370 ;
        RECT 88.515 112.190 88.805 112.915 ;
        RECT 88.975 112.145 92.485 112.915 ;
        RECT 92.655 112.405 92.960 112.915 ;
        RECT 83.000 110.365 88.345 110.800 ;
        RECT 88.515 110.365 88.805 111.530 ;
        RECT 88.975 111.455 90.665 111.975 ;
        RECT 90.835 111.625 92.485 112.145 ;
        RECT 92.655 111.675 92.970 112.235 ;
        RECT 93.140 111.925 93.390 112.735 ;
        RECT 93.560 112.390 93.820 112.915 ;
        RECT 94.000 111.925 94.250 112.735 ;
        RECT 94.420 112.355 94.680 112.915 ;
        RECT 94.850 112.265 95.110 112.720 ;
        RECT 95.280 112.435 95.540 112.915 ;
        RECT 95.710 112.265 95.970 112.720 ;
        RECT 96.140 112.435 96.400 112.915 ;
        RECT 96.570 112.265 96.830 112.720 ;
        RECT 97.000 112.435 97.245 112.915 ;
        RECT 97.415 112.265 97.690 112.720 ;
        RECT 97.860 112.435 98.105 112.915 ;
        RECT 98.275 112.265 98.535 112.720 ;
        RECT 98.715 112.435 98.965 112.915 ;
        RECT 99.135 112.265 99.395 112.720 ;
        RECT 99.575 112.435 99.825 112.915 ;
        RECT 99.995 112.265 100.255 112.720 ;
        RECT 100.435 112.435 100.695 112.915 ;
        RECT 100.865 112.265 101.125 112.720 ;
        RECT 101.295 112.435 101.595 112.915 ;
        RECT 101.855 112.410 102.140 112.915 ;
        RECT 94.850 112.235 101.595 112.265 ;
        RECT 102.310 112.240 102.635 112.745 ;
        RECT 94.850 112.095 101.625 112.235 ;
        RECT 100.430 112.065 101.625 112.095 ;
        RECT 93.140 111.675 100.260 111.925 ;
        RECT 88.975 110.365 92.485 111.455 ;
        RECT 92.665 110.365 92.960 111.175 ;
        RECT 93.140 110.535 93.385 111.675 ;
        RECT 93.560 110.365 93.820 111.175 ;
        RECT 94.000 110.540 94.250 111.675 ;
        RECT 100.430 111.505 101.595 112.065 ;
        RECT 101.855 111.710 102.635 112.240 ;
        RECT 94.850 111.280 101.595 111.505 ;
        RECT 94.850 111.265 100.255 111.280 ;
        RECT 94.420 110.370 94.680 111.165 ;
        RECT 94.850 110.540 95.110 111.265 ;
        RECT 95.280 110.370 95.540 111.095 ;
        RECT 95.710 110.540 95.970 111.265 ;
        RECT 96.140 110.370 96.400 111.095 ;
        RECT 96.570 110.540 96.830 111.265 ;
        RECT 97.000 110.370 97.260 111.095 ;
        RECT 97.430 110.540 97.690 111.265 ;
        RECT 97.860 110.370 98.105 111.095 ;
        RECT 98.275 110.540 98.535 111.265 ;
        RECT 98.720 110.370 98.965 111.095 ;
        RECT 99.135 110.540 99.395 111.265 ;
        RECT 99.580 110.370 99.825 111.095 ;
        RECT 99.995 110.540 100.255 111.265 ;
        RECT 100.440 110.370 100.695 111.095 ;
        RECT 100.865 110.540 101.155 111.280 ;
        RECT 94.420 110.365 100.695 110.370 ;
        RECT 101.325 110.365 101.595 111.110 ;
        RECT 101.855 110.365 102.135 111.335 ;
        RECT 102.305 110.535 102.635 111.710 ;
        RECT 102.825 111.675 103.065 112.625 ;
        RECT 103.240 112.370 108.585 112.915 ;
        RECT 108.760 112.370 114.105 112.915 ;
        RECT 102.805 110.365 103.065 111.335 ;
        RECT 104.830 110.800 105.180 112.050 ;
        RECT 106.660 111.540 107.000 112.370 ;
        RECT 110.350 110.800 110.700 112.050 ;
        RECT 112.180 111.540 112.520 112.370 ;
        RECT 114.275 112.190 114.565 112.915 ;
        RECT 115.655 112.145 119.165 112.915 ;
        RECT 103.240 110.365 108.585 110.800 ;
        RECT 108.760 110.365 114.105 110.800 ;
        RECT 114.275 110.365 114.565 111.530 ;
        RECT 115.655 111.455 117.345 111.975 ;
        RECT 117.515 111.625 119.165 112.145 ;
        RECT 119.375 112.095 119.605 112.915 ;
        RECT 119.775 112.115 120.105 112.745 ;
        RECT 119.355 111.675 119.685 111.925 ;
        RECT 119.855 111.515 120.105 112.115 ;
        RECT 120.275 112.095 120.485 112.915 ;
        RECT 120.715 112.240 120.975 112.745 ;
        RECT 121.155 112.535 121.485 112.915 ;
        RECT 121.665 112.365 121.835 112.745 ;
        RECT 115.655 110.365 119.165 111.455 ;
        RECT 119.375 110.365 119.605 111.505 ;
        RECT 119.775 110.535 120.105 111.515 ;
        RECT 120.275 110.365 120.485 111.505 ;
        RECT 120.715 111.440 120.885 112.240 ;
        RECT 121.170 112.195 121.835 112.365 ;
        RECT 122.095 112.240 122.355 112.745 ;
        RECT 122.535 112.535 122.865 112.915 ;
        RECT 123.045 112.365 123.215 112.745 ;
        RECT 121.170 111.940 121.340 112.195 ;
        RECT 121.055 111.610 121.340 111.940 ;
        RECT 121.575 111.645 121.905 112.015 ;
        RECT 121.170 111.465 121.340 111.610 ;
        RECT 120.715 110.535 120.985 111.440 ;
        RECT 121.170 111.295 121.835 111.465 ;
        RECT 121.155 110.365 121.485 111.125 ;
        RECT 121.665 110.535 121.835 111.295 ;
        RECT 122.095 111.440 122.265 112.240 ;
        RECT 122.550 112.195 123.215 112.365 ;
        RECT 122.550 111.940 122.720 112.195 ;
        RECT 123.475 112.145 126.065 112.915 ;
        RECT 126.235 112.165 127.445 112.915 ;
        RECT 122.435 111.610 122.720 111.940 ;
        RECT 122.955 111.645 123.285 112.015 ;
        RECT 122.550 111.465 122.720 111.610 ;
        RECT 122.095 110.535 122.365 111.440 ;
        RECT 122.550 111.295 123.215 111.465 ;
        RECT 122.535 110.365 122.865 111.125 ;
        RECT 123.045 110.535 123.215 111.295 ;
        RECT 123.475 111.455 124.685 111.975 ;
        RECT 124.855 111.625 126.065 112.145 ;
        RECT 126.235 111.455 126.755 111.995 ;
        RECT 126.925 111.625 127.445 112.165 ;
        RECT 123.475 110.365 126.065 111.455 ;
        RECT 126.235 110.365 127.445 111.455 ;
        RECT 14.370 110.195 127.530 110.365 ;
        RECT 14.455 109.105 15.665 110.195 ;
        RECT 14.455 108.395 14.975 108.935 ;
        RECT 15.145 108.565 15.665 109.105 ;
        RECT 16.755 109.105 20.265 110.195 ;
        RECT 16.755 108.585 18.445 109.105 ;
        RECT 20.495 109.055 20.705 110.195 ;
        RECT 20.875 109.045 21.205 110.025 ;
        RECT 21.375 109.055 21.605 110.195 ;
        RECT 22.795 109.055 23.005 110.195 ;
        RECT 23.175 109.045 23.505 110.025 ;
        RECT 23.675 109.055 23.905 110.195 ;
        RECT 18.615 108.415 20.265 108.935 ;
        RECT 14.455 107.645 15.665 108.395 ;
        RECT 16.755 107.645 20.265 108.415 ;
        RECT 20.495 107.645 20.705 108.465 ;
        RECT 20.875 108.445 21.125 109.045 ;
        RECT 21.295 108.635 21.625 108.885 ;
        RECT 20.875 107.815 21.205 108.445 ;
        RECT 21.375 107.645 21.605 108.465 ;
        RECT 22.795 107.645 23.005 108.465 ;
        RECT 23.175 108.445 23.425 109.045 ;
        RECT 24.115 109.030 24.405 110.195 ;
        RECT 24.575 109.105 27.165 110.195 ;
        RECT 27.335 109.120 27.605 110.025 ;
        RECT 27.775 109.435 28.105 110.195 ;
        RECT 28.285 109.265 28.455 110.025 ;
        RECT 23.595 108.635 23.925 108.885 ;
        RECT 24.575 108.585 25.785 109.105 ;
        RECT 23.175 107.815 23.505 108.445 ;
        RECT 23.675 107.645 23.905 108.465 ;
        RECT 25.955 108.415 27.165 108.935 ;
        RECT 24.115 107.645 24.405 108.370 ;
        RECT 24.575 107.645 27.165 108.415 ;
        RECT 27.335 108.320 27.505 109.120 ;
        RECT 27.790 109.095 28.455 109.265 ;
        RECT 28.715 109.105 30.385 110.195 ;
        RECT 27.790 108.950 27.960 109.095 ;
        RECT 27.675 108.620 27.960 108.950 ;
        RECT 27.790 108.365 27.960 108.620 ;
        RECT 28.195 108.545 28.525 108.915 ;
        RECT 28.715 108.585 29.465 109.105 ;
        RECT 30.615 109.055 30.825 110.195 ;
        RECT 30.995 109.045 31.325 110.025 ;
        RECT 31.495 109.055 31.725 110.195 ;
        RECT 31.935 109.120 32.205 110.025 ;
        RECT 32.375 109.435 32.705 110.195 ;
        RECT 32.885 109.265 33.055 110.025 ;
        RECT 29.635 108.415 30.385 108.935 ;
        RECT 27.335 107.815 27.595 108.320 ;
        RECT 27.790 108.195 28.455 108.365 ;
        RECT 27.775 107.645 28.105 108.025 ;
        RECT 28.285 107.815 28.455 108.195 ;
        RECT 28.715 107.645 30.385 108.415 ;
        RECT 30.615 107.645 30.825 108.465 ;
        RECT 30.995 108.445 31.245 109.045 ;
        RECT 31.415 108.635 31.745 108.885 ;
        RECT 30.995 107.815 31.325 108.445 ;
        RECT 31.495 107.645 31.725 108.465 ;
        RECT 31.935 108.320 32.105 109.120 ;
        RECT 32.390 109.095 33.055 109.265 ;
        RECT 34.235 109.120 34.505 110.025 ;
        RECT 34.675 109.435 35.005 110.195 ;
        RECT 35.185 109.265 35.355 110.025 ;
        RECT 32.390 108.950 32.560 109.095 ;
        RECT 32.275 108.620 32.560 108.950 ;
        RECT 32.390 108.365 32.560 108.620 ;
        RECT 32.795 108.545 33.125 108.915 ;
        RECT 31.935 107.815 32.195 108.320 ;
        RECT 32.390 108.195 33.055 108.365 ;
        RECT 32.375 107.645 32.705 108.025 ;
        RECT 32.885 107.815 33.055 108.195 ;
        RECT 34.235 108.320 34.405 109.120 ;
        RECT 34.690 109.095 35.355 109.265 ;
        RECT 36.075 109.105 38.665 110.195 ;
        RECT 38.840 109.760 44.185 110.195 ;
        RECT 44.360 109.760 49.705 110.195 ;
        RECT 34.690 108.950 34.860 109.095 ;
        RECT 34.575 108.620 34.860 108.950 ;
        RECT 34.690 108.365 34.860 108.620 ;
        RECT 35.095 108.545 35.425 108.915 ;
        RECT 36.075 108.585 37.285 109.105 ;
        RECT 37.455 108.415 38.665 108.935 ;
        RECT 40.430 108.510 40.780 109.760 ;
        RECT 34.235 107.815 34.495 108.320 ;
        RECT 34.690 108.195 35.355 108.365 ;
        RECT 34.675 107.645 35.005 108.025 ;
        RECT 35.185 107.815 35.355 108.195 ;
        RECT 36.075 107.645 38.665 108.415 ;
        RECT 42.260 108.190 42.600 109.020 ;
        RECT 45.950 108.510 46.300 109.760 ;
        RECT 49.875 109.030 50.165 110.195 ;
        RECT 50.885 109.265 51.055 110.025 ;
        RECT 51.235 109.435 51.565 110.195 ;
        RECT 50.885 109.095 51.550 109.265 ;
        RECT 51.735 109.120 52.005 110.025 ;
        RECT 47.780 108.190 48.120 109.020 ;
        RECT 51.380 108.950 51.550 109.095 ;
        RECT 50.815 108.545 51.145 108.915 ;
        RECT 51.380 108.620 51.665 108.950 ;
        RECT 38.840 107.645 44.185 108.190 ;
        RECT 44.360 107.645 49.705 108.190 ;
        RECT 49.875 107.645 50.165 108.370 ;
        RECT 51.380 108.365 51.550 108.620 ;
        RECT 50.885 108.195 51.550 108.365 ;
        RECT 51.835 108.320 52.005 109.120 ;
        RECT 53.095 109.105 56.605 110.195 ;
        RECT 56.865 109.265 57.035 110.025 ;
        RECT 57.215 109.435 57.545 110.195 ;
        RECT 53.095 108.585 54.785 109.105 ;
        RECT 56.865 109.095 57.530 109.265 ;
        RECT 57.715 109.120 57.985 110.025 ;
        RECT 57.360 108.950 57.530 109.095 ;
        RECT 54.955 108.415 56.605 108.935 ;
        RECT 56.795 108.545 57.125 108.915 ;
        RECT 57.360 108.620 57.645 108.950 ;
        RECT 50.885 107.815 51.055 108.195 ;
        RECT 51.235 107.645 51.565 108.025 ;
        RECT 51.745 107.815 52.005 108.320 ;
        RECT 53.095 107.645 56.605 108.415 ;
        RECT 57.360 108.365 57.530 108.620 ;
        RECT 56.865 108.195 57.530 108.365 ;
        RECT 57.815 108.320 57.985 109.120 ;
        RECT 58.155 109.105 59.365 110.195 ;
        RECT 59.545 109.215 59.875 110.025 ;
        RECT 60.045 109.395 60.285 110.195 ;
        RECT 58.155 108.565 58.675 109.105 ;
        RECT 59.545 109.045 60.260 109.215 ;
        RECT 58.845 108.395 59.365 108.935 ;
        RECT 59.540 108.635 59.920 108.875 ;
        RECT 60.090 108.805 60.260 109.045 ;
        RECT 60.465 109.175 60.635 110.025 ;
        RECT 60.805 109.395 61.135 110.195 ;
        RECT 61.305 109.175 61.475 110.025 ;
        RECT 60.465 109.005 61.475 109.175 ;
        RECT 61.645 109.045 61.975 110.195 ;
        RECT 62.755 109.105 64.425 110.195 ;
        RECT 60.980 108.835 61.475 109.005 ;
        RECT 60.090 108.635 60.590 108.805 ;
        RECT 60.975 108.665 61.475 108.835 ;
        RECT 60.090 108.465 60.260 108.635 ;
        RECT 60.980 108.465 61.475 108.665 ;
        RECT 62.755 108.585 63.505 109.105 ;
        RECT 64.635 109.055 64.865 110.195 ;
        RECT 65.035 109.045 65.365 110.025 ;
        RECT 65.535 109.055 65.745 110.195 ;
        RECT 66.435 109.105 68.105 110.195 ;
        RECT 68.365 109.265 68.535 110.025 ;
        RECT 68.715 109.435 69.045 110.195 ;
        RECT 56.865 107.815 57.035 108.195 ;
        RECT 57.215 107.645 57.545 108.025 ;
        RECT 57.725 107.815 57.985 108.320 ;
        RECT 58.155 107.645 59.365 108.395 ;
        RECT 59.625 108.295 60.260 108.465 ;
        RECT 60.465 108.295 61.475 108.465 ;
        RECT 59.625 107.815 59.795 108.295 ;
        RECT 59.975 107.645 60.215 108.125 ;
        RECT 60.465 107.815 60.635 108.295 ;
        RECT 60.805 107.645 61.135 108.125 ;
        RECT 61.305 107.815 61.475 108.295 ;
        RECT 61.645 107.645 61.975 108.445 ;
        RECT 63.675 108.415 64.425 108.935 ;
        RECT 64.615 108.635 64.945 108.885 ;
        RECT 62.755 107.645 64.425 108.415 ;
        RECT 64.635 107.645 64.865 108.465 ;
        RECT 65.115 108.445 65.365 109.045 ;
        RECT 66.435 108.585 67.185 109.105 ;
        RECT 68.365 109.095 69.030 109.265 ;
        RECT 69.215 109.120 69.485 110.025 ;
        RECT 70.120 109.760 75.465 110.195 ;
        RECT 68.860 108.950 69.030 109.095 ;
        RECT 65.035 107.815 65.365 108.445 ;
        RECT 65.535 107.645 65.745 108.465 ;
        RECT 67.355 108.415 68.105 108.935 ;
        RECT 68.295 108.545 68.625 108.915 ;
        RECT 68.860 108.620 69.145 108.950 ;
        RECT 66.435 107.645 68.105 108.415 ;
        RECT 68.860 108.365 69.030 108.620 ;
        RECT 68.365 108.195 69.030 108.365 ;
        RECT 69.315 108.320 69.485 109.120 ;
        RECT 71.710 108.510 72.060 109.760 ;
        RECT 75.635 109.030 75.925 110.195 ;
        RECT 76.155 109.055 76.365 110.195 ;
        RECT 76.535 109.045 76.865 110.025 ;
        RECT 77.035 109.055 77.265 110.195 ;
        RECT 77.535 109.055 77.745 110.195 ;
        RECT 77.915 109.045 78.245 110.025 ;
        RECT 78.415 109.055 78.645 110.195 ;
        RECT 79.785 109.215 80.115 110.025 ;
        RECT 80.285 109.395 80.525 110.195 ;
        RECT 79.785 109.045 80.500 109.215 ;
        RECT 68.365 107.815 68.535 108.195 ;
        RECT 68.715 107.645 69.045 108.025 ;
        RECT 69.225 107.815 69.485 108.320 ;
        RECT 73.540 108.190 73.880 109.020 ;
        RECT 70.120 107.645 75.465 108.190 ;
        RECT 75.635 107.645 75.925 108.370 ;
        RECT 76.155 107.645 76.365 108.465 ;
        RECT 76.535 108.445 76.785 109.045 ;
        RECT 76.955 108.635 77.285 108.885 ;
        RECT 76.535 107.815 76.865 108.445 ;
        RECT 77.035 107.645 77.265 108.465 ;
        RECT 77.535 107.645 77.745 108.465 ;
        RECT 77.915 108.445 78.165 109.045 ;
        RECT 78.335 108.635 78.665 108.885 ;
        RECT 79.780 108.635 80.160 108.875 ;
        RECT 80.330 108.805 80.500 109.045 ;
        RECT 80.705 109.175 80.875 110.025 ;
        RECT 81.045 109.395 81.375 110.195 ;
        RECT 81.545 109.175 81.715 110.025 ;
        RECT 80.705 109.005 81.715 109.175 ;
        RECT 81.885 109.045 82.215 110.195 ;
        RECT 82.625 109.265 82.795 110.025 ;
        RECT 82.975 109.435 83.305 110.195 ;
        RECT 82.625 109.095 83.290 109.265 ;
        RECT 83.475 109.120 83.745 110.025 ;
        RECT 80.330 108.635 80.830 108.805 ;
        RECT 80.330 108.465 80.500 108.635 ;
        RECT 81.220 108.465 81.715 109.005 ;
        RECT 83.120 108.950 83.290 109.095 ;
        RECT 82.555 108.545 82.885 108.915 ;
        RECT 83.120 108.620 83.405 108.950 ;
        RECT 77.915 107.815 78.245 108.445 ;
        RECT 78.415 107.645 78.645 108.465 ;
        RECT 79.865 108.295 80.500 108.465 ;
        RECT 80.705 108.295 81.715 108.465 ;
        RECT 79.865 107.815 80.035 108.295 ;
        RECT 80.215 107.645 80.455 108.125 ;
        RECT 80.705 107.815 80.875 108.295 ;
        RECT 81.045 107.645 81.375 108.125 ;
        RECT 81.545 107.815 81.715 108.295 ;
        RECT 81.885 107.645 82.215 108.445 ;
        RECT 83.120 108.365 83.290 108.620 ;
        RECT 82.625 108.195 83.290 108.365 ;
        RECT 83.575 108.320 83.745 109.120 ;
        RECT 84.375 109.105 86.965 110.195 ;
        RECT 84.375 108.585 85.585 109.105 ;
        RECT 87.175 109.055 87.405 110.195 ;
        RECT 87.575 109.045 87.905 110.025 ;
        RECT 88.075 109.055 88.285 110.195 ;
        RECT 88.515 109.105 92.025 110.195 ;
        RECT 85.755 108.415 86.965 108.935 ;
        RECT 87.155 108.635 87.485 108.885 ;
        RECT 82.625 107.815 82.795 108.195 ;
        RECT 82.975 107.645 83.305 108.025 ;
        RECT 83.485 107.815 83.745 108.320 ;
        RECT 84.375 107.645 86.965 108.415 ;
        RECT 87.175 107.645 87.405 108.465 ;
        RECT 87.655 108.445 87.905 109.045 ;
        RECT 88.515 108.585 90.205 109.105 ;
        RECT 92.235 109.055 92.465 110.195 ;
        RECT 92.635 109.045 92.965 110.025 ;
        RECT 93.135 109.055 93.345 110.195 ;
        RECT 93.665 109.265 93.835 110.025 ;
        RECT 94.015 109.435 94.345 110.195 ;
        RECT 93.665 109.095 94.330 109.265 ;
        RECT 94.515 109.120 94.785 110.025 ;
        RECT 87.575 107.815 87.905 108.445 ;
        RECT 88.075 107.645 88.285 108.465 ;
        RECT 90.375 108.415 92.025 108.935 ;
        RECT 92.215 108.635 92.545 108.885 ;
        RECT 88.515 107.645 92.025 108.415 ;
        RECT 92.235 107.645 92.465 108.465 ;
        RECT 92.715 108.445 92.965 109.045 ;
        RECT 94.160 108.950 94.330 109.095 ;
        RECT 93.595 108.545 93.925 108.915 ;
        RECT 94.160 108.620 94.445 108.950 ;
        RECT 92.635 107.815 92.965 108.445 ;
        RECT 93.135 107.645 93.345 108.465 ;
        RECT 94.160 108.365 94.330 108.620 ;
        RECT 93.665 108.195 94.330 108.365 ;
        RECT 94.615 108.320 94.785 109.120 ;
        RECT 94.955 109.105 96.165 110.195 ;
        RECT 96.335 109.105 99.845 110.195 ;
        RECT 100.015 109.120 100.285 110.025 ;
        RECT 100.455 109.435 100.785 110.195 ;
        RECT 100.965 109.265 101.135 110.025 ;
        RECT 94.955 108.565 95.475 109.105 ;
        RECT 95.645 108.395 96.165 108.935 ;
        RECT 96.335 108.585 98.025 109.105 ;
        RECT 98.195 108.415 99.845 108.935 ;
        RECT 93.665 107.815 93.835 108.195 ;
        RECT 94.015 107.645 94.345 108.025 ;
        RECT 94.525 107.815 94.785 108.320 ;
        RECT 94.955 107.645 96.165 108.395 ;
        RECT 96.335 107.645 99.845 108.415 ;
        RECT 100.015 108.320 100.185 109.120 ;
        RECT 100.470 109.095 101.135 109.265 ;
        RECT 100.470 108.950 100.640 109.095 ;
        RECT 101.395 109.030 101.685 110.195 ;
        RECT 102.315 109.105 105.825 110.195 ;
        RECT 106.085 109.265 106.255 110.025 ;
        RECT 106.435 109.435 106.765 110.195 ;
        RECT 100.355 108.620 100.640 108.950 ;
        RECT 100.470 108.365 100.640 108.620 ;
        RECT 100.875 108.545 101.205 108.915 ;
        RECT 102.315 108.585 104.005 109.105 ;
        RECT 106.085 109.095 106.750 109.265 ;
        RECT 106.935 109.120 107.205 110.025 ;
        RECT 106.580 108.950 106.750 109.095 ;
        RECT 104.175 108.415 105.825 108.935 ;
        RECT 106.015 108.545 106.345 108.915 ;
        RECT 106.580 108.620 106.865 108.950 ;
        RECT 100.015 107.815 100.275 108.320 ;
        RECT 100.470 108.195 101.135 108.365 ;
        RECT 100.455 107.645 100.785 108.025 ;
        RECT 100.965 107.815 101.135 108.195 ;
        RECT 101.395 107.645 101.685 108.370 ;
        RECT 102.315 107.645 105.825 108.415 ;
        RECT 106.580 108.365 106.750 108.620 ;
        RECT 106.085 108.195 106.750 108.365 ;
        RECT 107.035 108.320 107.205 109.120 ;
        RECT 107.375 109.105 108.585 110.195 ;
        RECT 107.375 108.565 107.895 109.105 ;
        RECT 108.815 109.055 109.025 110.195 ;
        RECT 109.195 109.045 109.525 110.025 ;
        RECT 109.695 109.055 109.925 110.195 ;
        RECT 110.225 109.265 110.395 110.025 ;
        RECT 110.575 109.435 110.905 110.195 ;
        RECT 110.225 109.095 110.890 109.265 ;
        RECT 111.075 109.120 111.345 110.025 ;
        RECT 108.065 108.395 108.585 108.935 ;
        RECT 106.085 107.815 106.255 108.195 ;
        RECT 106.435 107.645 106.765 108.025 ;
        RECT 106.945 107.815 107.205 108.320 ;
        RECT 107.375 107.645 108.585 108.395 ;
        RECT 108.815 107.645 109.025 108.465 ;
        RECT 109.195 108.445 109.445 109.045 ;
        RECT 110.720 108.950 110.890 109.095 ;
        RECT 109.615 108.635 109.945 108.885 ;
        RECT 110.155 108.545 110.485 108.915 ;
        RECT 110.720 108.620 111.005 108.950 ;
        RECT 109.195 107.815 109.525 108.445 ;
        RECT 109.695 107.645 109.925 108.465 ;
        RECT 110.720 108.365 110.890 108.620 ;
        RECT 110.225 108.195 110.890 108.365 ;
        RECT 111.175 108.320 111.345 109.120 ;
        RECT 111.605 109.265 111.775 110.025 ;
        RECT 111.955 109.435 112.285 110.195 ;
        RECT 111.605 109.095 112.270 109.265 ;
        RECT 112.455 109.120 112.725 110.025 ;
        RECT 112.100 108.950 112.270 109.095 ;
        RECT 111.535 108.545 111.865 108.915 ;
        RECT 112.100 108.620 112.385 108.950 ;
        RECT 112.100 108.365 112.270 108.620 ;
        RECT 110.225 107.815 110.395 108.195 ;
        RECT 110.575 107.645 110.905 108.025 ;
        RECT 111.085 107.815 111.345 108.320 ;
        RECT 111.605 108.195 112.270 108.365 ;
        RECT 112.555 108.320 112.725 109.120 ;
        RECT 112.895 109.105 114.105 110.195 ;
        RECT 112.895 108.565 113.415 109.105 ;
        RECT 114.315 109.055 114.545 110.195 ;
        RECT 114.715 109.045 115.045 110.025 ;
        RECT 115.215 109.055 115.425 110.195 ;
        RECT 115.660 109.525 115.915 110.025 ;
        RECT 116.085 109.695 116.415 110.195 ;
        RECT 115.660 109.355 116.410 109.525 ;
        RECT 113.585 108.395 114.105 108.935 ;
        RECT 114.295 108.635 114.625 108.885 ;
        RECT 111.605 107.815 111.775 108.195 ;
        RECT 111.955 107.645 112.285 108.025 ;
        RECT 112.465 107.815 112.725 108.320 ;
        RECT 112.895 107.645 114.105 108.395 ;
        RECT 114.315 107.645 114.545 108.465 ;
        RECT 114.795 108.445 115.045 109.045 ;
        RECT 115.660 108.535 116.010 109.185 ;
        RECT 114.715 107.815 115.045 108.445 ;
        RECT 115.215 107.645 115.425 108.465 ;
        RECT 116.180 108.365 116.410 109.355 ;
        RECT 115.660 108.195 116.410 108.365 ;
        RECT 115.660 107.905 115.915 108.195 ;
        RECT 116.085 107.645 116.415 108.025 ;
        RECT 116.585 107.905 116.755 110.025 ;
        RECT 116.925 109.225 117.250 110.010 ;
        RECT 117.420 109.735 117.670 110.195 ;
        RECT 117.840 109.695 118.090 110.025 ;
        RECT 118.305 109.695 118.985 110.025 ;
        RECT 117.840 109.565 118.010 109.695 ;
        RECT 117.615 109.395 118.010 109.565 ;
        RECT 116.985 108.175 117.445 109.225 ;
        RECT 117.615 108.035 117.785 109.395 ;
        RECT 118.180 109.135 118.645 109.525 ;
        RECT 117.955 108.325 118.305 108.945 ;
        RECT 118.475 108.545 118.645 109.135 ;
        RECT 118.815 108.915 118.985 109.695 ;
        RECT 119.155 109.595 119.325 109.935 ;
        RECT 119.560 109.765 119.890 110.195 ;
        RECT 120.060 109.595 120.230 109.935 ;
        RECT 120.525 109.735 120.895 110.195 ;
        RECT 119.155 109.425 120.230 109.595 ;
        RECT 121.065 109.565 121.235 110.025 ;
        RECT 121.470 109.685 122.340 110.025 ;
        RECT 122.510 109.735 122.760 110.195 ;
        RECT 120.675 109.395 121.235 109.565 ;
        RECT 120.675 109.255 120.845 109.395 ;
        RECT 119.345 109.085 120.845 109.255 ;
        RECT 121.540 109.225 122.000 109.515 ;
        RECT 118.815 108.745 120.505 108.915 ;
        RECT 118.475 108.325 118.830 108.545 ;
        RECT 119.000 108.035 119.170 108.745 ;
        RECT 119.375 108.325 120.165 108.575 ;
        RECT 120.335 108.565 120.505 108.745 ;
        RECT 120.675 108.395 120.845 109.085 ;
        RECT 117.115 107.645 117.445 108.005 ;
        RECT 117.615 107.865 118.110 108.035 ;
        RECT 118.315 107.865 119.170 108.035 ;
        RECT 120.045 107.645 120.375 108.105 ;
        RECT 120.585 108.005 120.845 108.395 ;
        RECT 121.035 109.215 122.000 109.225 ;
        RECT 122.170 109.305 122.340 109.685 ;
        RECT 122.930 109.645 123.100 109.935 ;
        RECT 123.280 109.815 123.610 110.195 ;
        RECT 122.930 109.475 123.730 109.645 ;
        RECT 121.035 109.055 121.710 109.215 ;
        RECT 122.170 109.135 123.390 109.305 ;
        RECT 121.035 108.265 121.245 109.055 ;
        RECT 122.170 109.045 122.340 109.135 ;
        RECT 121.415 108.265 121.765 108.885 ;
        RECT 121.935 108.875 122.340 109.045 ;
        RECT 121.935 108.095 122.105 108.875 ;
        RECT 122.275 108.425 122.495 108.705 ;
        RECT 122.675 108.595 123.215 108.965 ;
        RECT 123.560 108.855 123.730 109.475 ;
        RECT 123.905 109.135 124.075 110.195 ;
        RECT 124.285 109.185 124.575 110.025 ;
        RECT 124.745 109.355 124.915 110.195 ;
        RECT 125.125 109.185 125.375 110.025 ;
        RECT 125.585 109.355 125.755 110.195 ;
        RECT 124.285 109.015 126.010 109.185 ;
        RECT 122.275 108.255 122.805 108.425 ;
        RECT 120.585 107.835 120.935 108.005 ;
        RECT 121.155 107.815 122.105 108.095 ;
        RECT 122.275 107.645 122.465 108.085 ;
        RECT 122.635 108.025 122.805 108.255 ;
        RECT 122.975 108.195 123.215 108.595 ;
        RECT 123.385 108.845 123.730 108.855 ;
        RECT 123.385 108.635 125.415 108.845 ;
        RECT 123.385 108.380 123.710 108.635 ;
        RECT 125.600 108.465 126.010 109.015 ;
        RECT 126.235 109.105 127.445 110.195 ;
        RECT 126.235 108.565 126.755 109.105 ;
        RECT 123.385 108.025 123.705 108.380 ;
        RECT 122.635 107.855 123.705 108.025 ;
        RECT 123.905 107.645 124.075 108.455 ;
        RECT 124.245 108.295 126.010 108.465 ;
        RECT 126.925 108.395 127.445 108.935 ;
        RECT 124.245 107.815 124.575 108.295 ;
        RECT 124.745 107.645 124.915 108.115 ;
        RECT 125.085 107.815 125.415 108.295 ;
        RECT 125.585 107.645 125.755 108.115 ;
        RECT 126.235 107.645 127.445 108.395 ;
        RECT 14.370 107.475 127.530 107.645 ;
        RECT 14.455 106.725 15.665 107.475 ;
        RECT 16.145 107.005 16.315 107.475 ;
        RECT 16.485 106.825 16.815 107.305 ;
        RECT 16.985 107.005 17.155 107.475 ;
        RECT 17.325 106.825 17.655 107.305 ;
        RECT 14.455 106.185 14.975 106.725 ;
        RECT 15.890 106.655 17.655 106.825 ;
        RECT 17.825 106.665 17.995 107.475 ;
        RECT 18.195 107.095 19.265 107.265 ;
        RECT 18.195 106.740 18.515 107.095 ;
        RECT 15.145 106.015 15.665 106.555 ;
        RECT 14.455 104.925 15.665 106.015 ;
        RECT 15.890 106.105 16.300 106.655 ;
        RECT 18.190 106.485 18.515 106.740 ;
        RECT 16.485 106.275 18.515 106.485 ;
        RECT 18.170 106.265 18.515 106.275 ;
        RECT 18.685 106.525 18.925 106.925 ;
        RECT 19.095 106.865 19.265 107.095 ;
        RECT 19.435 107.035 19.625 107.475 ;
        RECT 19.795 107.025 20.745 107.305 ;
        RECT 20.965 107.115 21.315 107.285 ;
        RECT 19.095 106.695 19.625 106.865 ;
        RECT 15.890 105.935 17.615 106.105 ;
        RECT 16.145 104.925 16.315 105.765 ;
        RECT 16.525 105.095 16.775 105.935 ;
        RECT 16.985 104.925 17.155 105.765 ;
        RECT 17.325 105.095 17.615 105.935 ;
        RECT 17.825 104.925 17.995 105.985 ;
        RECT 18.170 105.645 18.340 106.265 ;
        RECT 18.685 106.155 19.225 106.525 ;
        RECT 19.405 106.415 19.625 106.695 ;
        RECT 19.795 106.245 19.965 107.025 ;
        RECT 19.560 106.075 19.965 106.245 ;
        RECT 20.135 106.235 20.485 106.855 ;
        RECT 19.560 105.985 19.730 106.075 ;
        RECT 20.655 106.065 20.865 106.855 ;
        RECT 18.510 105.815 19.730 105.985 ;
        RECT 20.190 105.905 20.865 106.065 ;
        RECT 18.170 105.475 18.970 105.645 ;
        RECT 18.290 104.925 18.620 105.305 ;
        RECT 18.800 105.185 18.970 105.475 ;
        RECT 19.560 105.435 19.730 105.815 ;
        RECT 19.900 105.895 20.865 105.905 ;
        RECT 21.055 106.725 21.315 107.115 ;
        RECT 21.525 107.015 21.855 107.475 ;
        RECT 22.730 107.085 23.585 107.255 ;
        RECT 23.790 107.085 24.285 107.255 ;
        RECT 24.455 107.115 24.785 107.475 ;
        RECT 21.055 106.035 21.225 106.725 ;
        RECT 21.395 106.375 21.565 106.555 ;
        RECT 21.735 106.545 22.525 106.795 ;
        RECT 22.730 106.375 22.900 107.085 ;
        RECT 23.070 106.575 23.425 106.795 ;
        RECT 21.395 106.205 23.085 106.375 ;
        RECT 19.900 105.605 20.360 105.895 ;
        RECT 21.055 105.865 22.555 106.035 ;
        RECT 21.055 105.725 21.225 105.865 ;
        RECT 20.665 105.555 21.225 105.725 ;
        RECT 19.140 104.925 19.390 105.385 ;
        RECT 19.560 105.095 20.430 105.435 ;
        RECT 20.665 105.095 20.835 105.555 ;
        RECT 21.670 105.525 22.745 105.695 ;
        RECT 21.005 104.925 21.375 105.385 ;
        RECT 21.670 105.185 21.840 105.525 ;
        RECT 22.010 104.925 22.340 105.355 ;
        RECT 22.575 105.185 22.745 105.525 ;
        RECT 22.915 105.425 23.085 106.205 ;
        RECT 23.255 105.985 23.425 106.575 ;
        RECT 23.595 106.175 23.945 106.795 ;
        RECT 23.255 105.595 23.720 105.985 ;
        RECT 24.115 105.725 24.285 107.085 ;
        RECT 24.455 105.895 24.915 106.945 ;
        RECT 23.890 105.555 24.285 105.725 ;
        RECT 23.890 105.425 24.060 105.555 ;
        RECT 22.915 105.095 23.595 105.425 ;
        RECT 23.810 105.095 24.060 105.425 ;
        RECT 24.230 104.925 24.480 105.385 ;
        RECT 24.650 105.110 24.975 105.895 ;
        RECT 25.145 105.095 25.315 107.215 ;
        RECT 25.485 107.095 25.815 107.475 ;
        RECT 25.985 106.925 26.240 107.215 ;
        RECT 26.725 107.005 26.895 107.475 ;
        RECT 25.490 106.755 26.240 106.925 ;
        RECT 27.065 106.825 27.395 107.305 ;
        RECT 27.565 107.005 27.735 107.475 ;
        RECT 27.905 106.825 28.235 107.305 ;
        RECT 25.490 105.765 25.720 106.755 ;
        RECT 26.470 106.655 28.235 106.825 ;
        RECT 28.405 106.665 28.575 107.475 ;
        RECT 28.775 107.095 29.845 107.265 ;
        RECT 28.775 106.740 29.095 107.095 ;
        RECT 25.890 105.935 26.240 106.585 ;
        RECT 26.470 106.105 26.880 106.655 ;
        RECT 28.770 106.485 29.095 106.740 ;
        RECT 27.065 106.275 29.095 106.485 ;
        RECT 28.750 106.265 29.095 106.275 ;
        RECT 29.265 106.525 29.505 106.925 ;
        RECT 29.675 106.865 29.845 107.095 ;
        RECT 30.015 107.035 30.205 107.475 ;
        RECT 30.375 107.025 31.325 107.305 ;
        RECT 31.545 107.115 31.895 107.285 ;
        RECT 29.675 106.695 30.205 106.865 ;
        RECT 26.470 105.935 28.195 106.105 ;
        RECT 25.490 105.595 26.240 105.765 ;
        RECT 25.485 104.925 25.815 105.425 ;
        RECT 25.985 105.095 26.240 105.595 ;
        RECT 26.725 104.925 26.895 105.765 ;
        RECT 27.105 105.095 27.355 105.935 ;
        RECT 27.565 104.925 27.735 105.765 ;
        RECT 27.905 105.095 28.195 105.935 ;
        RECT 28.405 104.925 28.575 105.985 ;
        RECT 28.750 105.645 28.920 106.265 ;
        RECT 29.265 106.155 29.805 106.525 ;
        RECT 29.985 106.415 30.205 106.695 ;
        RECT 30.375 106.245 30.545 107.025 ;
        RECT 30.140 106.075 30.545 106.245 ;
        RECT 30.715 106.235 31.065 106.855 ;
        RECT 30.140 105.985 30.310 106.075 ;
        RECT 31.235 106.065 31.445 106.855 ;
        RECT 29.090 105.815 30.310 105.985 ;
        RECT 30.770 105.905 31.445 106.065 ;
        RECT 28.750 105.475 29.550 105.645 ;
        RECT 28.870 104.925 29.200 105.305 ;
        RECT 29.380 105.185 29.550 105.475 ;
        RECT 30.140 105.435 30.310 105.815 ;
        RECT 30.480 105.895 31.445 105.905 ;
        RECT 31.635 106.725 31.895 107.115 ;
        RECT 32.105 107.015 32.435 107.475 ;
        RECT 33.310 107.085 34.165 107.255 ;
        RECT 34.370 107.085 34.865 107.255 ;
        RECT 35.035 107.115 35.365 107.475 ;
        RECT 31.635 106.035 31.805 106.725 ;
        RECT 31.975 106.375 32.145 106.555 ;
        RECT 32.315 106.545 33.105 106.795 ;
        RECT 33.310 106.375 33.480 107.085 ;
        RECT 33.650 106.575 34.005 106.795 ;
        RECT 31.975 106.205 33.665 106.375 ;
        RECT 30.480 105.605 30.940 105.895 ;
        RECT 31.635 105.865 33.135 106.035 ;
        RECT 31.635 105.725 31.805 105.865 ;
        RECT 31.245 105.555 31.805 105.725 ;
        RECT 29.720 104.925 29.970 105.385 ;
        RECT 30.140 105.095 31.010 105.435 ;
        RECT 31.245 105.095 31.415 105.555 ;
        RECT 32.250 105.525 33.325 105.695 ;
        RECT 31.585 104.925 31.955 105.385 ;
        RECT 32.250 105.185 32.420 105.525 ;
        RECT 32.590 104.925 32.920 105.355 ;
        RECT 33.155 105.185 33.325 105.525 ;
        RECT 33.495 105.425 33.665 106.205 ;
        RECT 33.835 105.985 34.005 106.575 ;
        RECT 34.175 106.175 34.525 106.795 ;
        RECT 33.835 105.595 34.300 105.985 ;
        RECT 34.695 105.725 34.865 107.085 ;
        RECT 35.035 105.895 35.495 106.945 ;
        RECT 34.470 105.555 34.865 105.725 ;
        RECT 34.470 105.425 34.640 105.555 ;
        RECT 33.495 105.095 34.175 105.425 ;
        RECT 34.390 105.095 34.640 105.425 ;
        RECT 34.810 104.925 35.060 105.385 ;
        RECT 35.230 105.110 35.555 105.895 ;
        RECT 35.725 105.095 35.895 107.215 ;
        RECT 36.065 107.095 36.395 107.475 ;
        RECT 36.565 106.925 36.820 107.215 ;
        RECT 36.070 106.755 36.820 106.925 ;
        RECT 36.070 105.765 36.300 106.755 ;
        RECT 36.995 106.750 37.285 107.475 ;
        RECT 37.455 106.800 37.715 107.305 ;
        RECT 37.895 107.095 38.225 107.475 ;
        RECT 38.405 106.925 38.575 107.305 ;
        RECT 36.470 105.935 36.820 106.585 ;
        RECT 36.070 105.595 36.820 105.765 ;
        RECT 36.065 104.925 36.395 105.425 ;
        RECT 36.565 105.095 36.820 105.595 ;
        RECT 36.995 104.925 37.285 106.090 ;
        RECT 37.455 106.000 37.625 106.800 ;
        RECT 37.910 106.755 38.575 106.925 ;
        RECT 37.910 106.500 38.080 106.755 ;
        RECT 39.355 106.655 39.565 107.475 ;
        RECT 39.735 106.675 40.065 107.305 ;
        RECT 37.795 106.170 38.080 106.500 ;
        RECT 38.315 106.205 38.645 106.575 ;
        RECT 37.910 106.025 38.080 106.170 ;
        RECT 39.735 106.075 39.985 106.675 ;
        RECT 40.235 106.655 40.465 107.475 ;
        RECT 40.675 106.725 41.885 107.475 ;
        RECT 40.155 106.235 40.485 106.485 ;
        RECT 37.455 105.095 37.725 106.000 ;
        RECT 37.910 105.855 38.575 106.025 ;
        RECT 37.895 104.925 38.225 105.685 ;
        RECT 38.405 105.095 38.575 105.855 ;
        RECT 39.355 104.925 39.565 106.065 ;
        RECT 39.735 105.095 40.065 106.075 ;
        RECT 40.235 104.925 40.465 106.065 ;
        RECT 40.675 106.015 41.195 106.555 ;
        RECT 41.365 106.185 41.885 106.725 ;
        RECT 42.055 106.800 42.315 107.305 ;
        RECT 42.495 107.095 42.825 107.475 ;
        RECT 43.005 106.925 43.175 107.305 ;
        RECT 40.675 104.925 41.885 106.015 ;
        RECT 42.055 106.000 42.225 106.800 ;
        RECT 42.510 106.755 43.175 106.925 ;
        RECT 42.510 106.500 42.680 106.755 ;
        RECT 43.955 106.655 44.165 107.475 ;
        RECT 44.335 106.675 44.665 107.305 ;
        RECT 42.395 106.170 42.680 106.500 ;
        RECT 42.915 106.205 43.245 106.575 ;
        RECT 42.510 106.025 42.680 106.170 ;
        RECT 44.335 106.075 44.585 106.675 ;
        RECT 44.835 106.655 45.065 107.475 ;
        RECT 45.365 106.925 45.535 107.305 ;
        RECT 45.715 107.095 46.045 107.475 ;
        RECT 45.365 106.755 46.030 106.925 ;
        RECT 46.225 106.800 46.485 107.305 ;
        RECT 46.965 107.005 47.135 107.475 ;
        RECT 47.305 106.825 47.635 107.305 ;
        RECT 47.805 107.005 47.975 107.475 ;
        RECT 48.145 106.825 48.475 107.305 ;
        RECT 44.755 106.235 45.085 106.485 ;
        RECT 45.295 106.205 45.625 106.575 ;
        RECT 45.860 106.500 46.030 106.755 ;
        RECT 45.860 106.170 46.145 106.500 ;
        RECT 42.055 105.095 42.325 106.000 ;
        RECT 42.510 105.855 43.175 106.025 ;
        RECT 42.495 104.925 42.825 105.685 ;
        RECT 43.005 105.095 43.175 105.855 ;
        RECT 43.955 104.925 44.165 106.065 ;
        RECT 44.335 105.095 44.665 106.075 ;
        RECT 44.835 104.925 45.065 106.065 ;
        RECT 45.860 106.025 46.030 106.170 ;
        RECT 45.365 105.855 46.030 106.025 ;
        RECT 46.315 106.000 46.485 106.800 ;
        RECT 45.365 105.095 45.535 105.855 ;
        RECT 45.715 104.925 46.045 105.685 ;
        RECT 46.215 105.095 46.485 106.000 ;
        RECT 46.710 106.655 48.475 106.825 ;
        RECT 48.645 106.665 48.815 107.475 ;
        RECT 49.015 107.095 50.085 107.265 ;
        RECT 49.015 106.740 49.335 107.095 ;
        RECT 46.710 106.105 47.120 106.655 ;
        RECT 49.010 106.485 49.335 106.740 ;
        RECT 47.305 106.275 49.335 106.485 ;
        RECT 48.990 106.265 49.335 106.275 ;
        RECT 49.505 106.525 49.745 106.925 ;
        RECT 49.915 106.865 50.085 107.095 ;
        RECT 50.255 107.035 50.445 107.475 ;
        RECT 50.615 107.025 51.565 107.305 ;
        RECT 51.785 107.115 52.135 107.285 ;
        RECT 49.915 106.695 50.445 106.865 ;
        RECT 46.710 105.935 48.435 106.105 ;
        RECT 46.965 104.925 47.135 105.765 ;
        RECT 47.345 105.095 47.595 105.935 ;
        RECT 47.805 104.925 47.975 105.765 ;
        RECT 48.145 105.095 48.435 105.935 ;
        RECT 48.645 104.925 48.815 105.985 ;
        RECT 48.990 105.645 49.160 106.265 ;
        RECT 49.505 106.155 50.045 106.525 ;
        RECT 50.225 106.415 50.445 106.695 ;
        RECT 50.615 106.245 50.785 107.025 ;
        RECT 50.380 106.075 50.785 106.245 ;
        RECT 50.955 106.235 51.305 106.855 ;
        RECT 50.380 105.985 50.550 106.075 ;
        RECT 51.475 106.065 51.685 106.855 ;
        RECT 49.330 105.815 50.550 105.985 ;
        RECT 51.010 105.905 51.685 106.065 ;
        RECT 48.990 105.475 49.790 105.645 ;
        RECT 49.110 104.925 49.440 105.305 ;
        RECT 49.620 105.185 49.790 105.475 ;
        RECT 50.380 105.435 50.550 105.815 ;
        RECT 50.720 105.895 51.685 105.905 ;
        RECT 51.875 106.725 52.135 107.115 ;
        RECT 52.345 107.015 52.675 107.475 ;
        RECT 53.550 107.085 54.405 107.255 ;
        RECT 54.610 107.085 55.105 107.255 ;
        RECT 55.275 107.115 55.605 107.475 ;
        RECT 51.875 106.035 52.045 106.725 ;
        RECT 52.215 106.375 52.385 106.555 ;
        RECT 52.555 106.545 53.345 106.795 ;
        RECT 53.550 106.375 53.720 107.085 ;
        RECT 53.890 106.575 54.245 106.795 ;
        RECT 52.215 106.205 53.905 106.375 ;
        RECT 50.720 105.605 51.180 105.895 ;
        RECT 51.875 105.865 53.375 106.035 ;
        RECT 51.875 105.725 52.045 105.865 ;
        RECT 51.485 105.555 52.045 105.725 ;
        RECT 49.960 104.925 50.210 105.385 ;
        RECT 50.380 105.095 51.250 105.435 ;
        RECT 51.485 105.095 51.655 105.555 ;
        RECT 52.490 105.525 53.565 105.695 ;
        RECT 51.825 104.925 52.195 105.385 ;
        RECT 52.490 105.185 52.660 105.525 ;
        RECT 52.830 104.925 53.160 105.355 ;
        RECT 53.395 105.185 53.565 105.525 ;
        RECT 53.735 105.425 53.905 106.205 ;
        RECT 54.075 105.985 54.245 106.575 ;
        RECT 54.415 106.175 54.765 106.795 ;
        RECT 54.075 105.595 54.540 105.985 ;
        RECT 54.935 105.725 55.105 107.085 ;
        RECT 55.275 105.895 55.735 106.945 ;
        RECT 54.710 105.555 55.105 105.725 ;
        RECT 54.710 105.425 54.880 105.555 ;
        RECT 53.735 105.095 54.415 105.425 ;
        RECT 54.630 105.095 54.880 105.425 ;
        RECT 55.050 104.925 55.300 105.385 ;
        RECT 55.470 105.110 55.795 105.895 ;
        RECT 55.965 105.095 56.135 107.215 ;
        RECT 56.305 107.095 56.635 107.475 ;
        RECT 56.805 106.925 57.060 107.215 ;
        RECT 56.310 106.755 57.060 106.925 ;
        RECT 56.310 105.765 56.540 106.755 ;
        RECT 57.295 106.655 57.505 107.475 ;
        RECT 57.675 106.675 58.005 107.305 ;
        RECT 56.710 105.935 57.060 106.585 ;
        RECT 57.675 106.075 57.925 106.675 ;
        RECT 58.175 106.655 58.405 107.475 ;
        RECT 58.615 106.725 59.825 107.475 ;
        RECT 58.095 106.235 58.425 106.485 ;
        RECT 56.310 105.595 57.060 105.765 ;
        RECT 56.305 104.925 56.635 105.425 ;
        RECT 56.805 105.095 57.060 105.595 ;
        RECT 57.295 104.925 57.505 106.065 ;
        RECT 57.675 105.095 58.005 106.075 ;
        RECT 58.175 104.925 58.405 106.065 ;
        RECT 58.615 106.015 59.135 106.555 ;
        RECT 59.305 106.185 59.825 106.725 ;
        RECT 60.035 106.655 60.265 107.475 ;
        RECT 60.435 106.675 60.765 107.305 ;
        RECT 60.015 106.235 60.345 106.485 ;
        RECT 60.515 106.075 60.765 106.675 ;
        RECT 60.935 106.655 61.145 107.475 ;
        RECT 61.465 106.925 61.635 107.305 ;
        RECT 61.815 107.095 62.145 107.475 ;
        RECT 61.465 106.755 62.130 106.925 ;
        RECT 62.325 106.800 62.585 107.305 ;
        RECT 61.395 106.205 61.725 106.575 ;
        RECT 61.960 106.500 62.130 106.755 ;
        RECT 58.615 104.925 59.825 106.015 ;
        RECT 60.035 104.925 60.265 106.065 ;
        RECT 60.435 105.095 60.765 106.075 ;
        RECT 61.960 106.170 62.245 106.500 ;
        RECT 60.935 104.925 61.145 106.065 ;
        RECT 61.960 106.025 62.130 106.170 ;
        RECT 61.465 105.855 62.130 106.025 ;
        RECT 62.415 106.000 62.585 106.800 ;
        RECT 62.755 106.750 63.045 107.475 ;
        RECT 63.525 107.005 63.695 107.475 ;
        RECT 63.865 106.825 64.195 107.305 ;
        RECT 64.365 107.005 64.535 107.475 ;
        RECT 64.705 106.825 65.035 107.305 ;
        RECT 63.270 106.655 65.035 106.825 ;
        RECT 65.205 106.665 65.375 107.475 ;
        RECT 65.575 107.095 66.645 107.265 ;
        RECT 65.575 106.740 65.895 107.095 ;
        RECT 63.270 106.105 63.680 106.655 ;
        RECT 65.570 106.485 65.895 106.740 ;
        RECT 63.865 106.275 65.895 106.485 ;
        RECT 65.550 106.265 65.895 106.275 ;
        RECT 66.065 106.525 66.305 106.925 ;
        RECT 66.475 106.865 66.645 107.095 ;
        RECT 66.815 107.035 67.005 107.475 ;
        RECT 67.175 107.025 68.125 107.305 ;
        RECT 68.345 107.115 68.695 107.285 ;
        RECT 66.475 106.695 67.005 106.865 ;
        RECT 61.465 105.095 61.635 105.855 ;
        RECT 61.815 104.925 62.145 105.685 ;
        RECT 62.315 105.095 62.585 106.000 ;
        RECT 62.755 104.925 63.045 106.090 ;
        RECT 63.270 105.935 64.995 106.105 ;
        RECT 63.525 104.925 63.695 105.765 ;
        RECT 63.905 105.095 64.155 105.935 ;
        RECT 64.365 104.925 64.535 105.765 ;
        RECT 64.705 105.095 64.995 105.935 ;
        RECT 65.205 104.925 65.375 105.985 ;
        RECT 65.550 105.645 65.720 106.265 ;
        RECT 66.065 106.155 66.605 106.525 ;
        RECT 66.785 106.415 67.005 106.695 ;
        RECT 67.175 106.245 67.345 107.025 ;
        RECT 66.940 106.075 67.345 106.245 ;
        RECT 67.515 106.235 67.865 106.855 ;
        RECT 66.940 105.985 67.110 106.075 ;
        RECT 68.035 106.065 68.245 106.855 ;
        RECT 65.890 105.815 67.110 105.985 ;
        RECT 67.570 105.905 68.245 106.065 ;
        RECT 65.550 105.475 66.350 105.645 ;
        RECT 65.670 104.925 66.000 105.305 ;
        RECT 66.180 105.185 66.350 105.475 ;
        RECT 66.940 105.435 67.110 105.815 ;
        RECT 67.280 105.895 68.245 105.905 ;
        RECT 68.435 106.725 68.695 107.115 ;
        RECT 68.905 107.015 69.235 107.475 ;
        RECT 70.110 107.085 70.965 107.255 ;
        RECT 71.170 107.085 71.665 107.255 ;
        RECT 71.835 107.115 72.165 107.475 ;
        RECT 68.435 106.035 68.605 106.725 ;
        RECT 68.775 106.375 68.945 106.555 ;
        RECT 69.115 106.545 69.905 106.795 ;
        RECT 70.110 106.375 70.280 107.085 ;
        RECT 70.450 106.575 70.805 106.795 ;
        RECT 68.775 106.205 70.465 106.375 ;
        RECT 67.280 105.605 67.740 105.895 ;
        RECT 68.435 105.865 69.935 106.035 ;
        RECT 68.435 105.725 68.605 105.865 ;
        RECT 68.045 105.555 68.605 105.725 ;
        RECT 66.520 104.925 66.770 105.385 ;
        RECT 66.940 105.095 67.810 105.435 ;
        RECT 68.045 105.095 68.215 105.555 ;
        RECT 69.050 105.525 70.125 105.695 ;
        RECT 68.385 104.925 68.755 105.385 ;
        RECT 69.050 105.185 69.220 105.525 ;
        RECT 69.390 104.925 69.720 105.355 ;
        RECT 69.955 105.185 70.125 105.525 ;
        RECT 70.295 105.425 70.465 106.205 ;
        RECT 70.635 105.985 70.805 106.575 ;
        RECT 70.975 106.175 71.325 106.795 ;
        RECT 70.635 105.595 71.100 105.985 ;
        RECT 71.495 105.725 71.665 107.085 ;
        RECT 71.835 105.895 72.295 106.945 ;
        RECT 71.270 105.555 71.665 105.725 ;
        RECT 71.270 105.425 71.440 105.555 ;
        RECT 70.295 105.095 70.975 105.425 ;
        RECT 71.190 105.095 71.440 105.425 ;
        RECT 71.610 104.925 71.860 105.385 ;
        RECT 72.030 105.110 72.355 105.895 ;
        RECT 72.525 105.095 72.695 107.215 ;
        RECT 72.865 107.095 73.195 107.475 ;
        RECT 73.365 106.925 73.620 107.215 ;
        RECT 72.870 106.755 73.620 106.925 ;
        RECT 74.805 106.925 74.975 107.305 ;
        RECT 75.155 107.095 75.485 107.475 ;
        RECT 74.805 106.755 75.470 106.925 ;
        RECT 75.665 106.800 75.925 107.305 ;
        RECT 76.405 107.005 76.575 107.475 ;
        RECT 76.745 106.825 77.075 107.305 ;
        RECT 77.245 107.005 77.415 107.475 ;
        RECT 77.585 106.825 77.915 107.305 ;
        RECT 72.870 105.765 73.100 106.755 ;
        RECT 73.270 105.935 73.620 106.585 ;
        RECT 74.735 106.205 75.065 106.575 ;
        RECT 75.300 106.500 75.470 106.755 ;
        RECT 75.300 106.170 75.585 106.500 ;
        RECT 75.300 106.025 75.470 106.170 ;
        RECT 74.805 105.855 75.470 106.025 ;
        RECT 75.755 106.000 75.925 106.800 ;
        RECT 72.870 105.595 73.620 105.765 ;
        RECT 72.865 104.925 73.195 105.425 ;
        RECT 73.365 105.095 73.620 105.595 ;
        RECT 74.805 105.095 74.975 105.855 ;
        RECT 75.155 104.925 75.485 105.685 ;
        RECT 75.655 105.095 75.925 106.000 ;
        RECT 76.150 106.655 77.915 106.825 ;
        RECT 78.085 106.665 78.255 107.475 ;
        RECT 78.455 107.095 79.525 107.265 ;
        RECT 78.455 106.740 78.775 107.095 ;
        RECT 76.150 106.105 76.560 106.655 ;
        RECT 78.450 106.485 78.775 106.740 ;
        RECT 76.745 106.275 78.775 106.485 ;
        RECT 78.430 106.265 78.775 106.275 ;
        RECT 78.945 106.525 79.185 106.925 ;
        RECT 79.355 106.865 79.525 107.095 ;
        RECT 79.695 107.035 79.885 107.475 ;
        RECT 80.055 107.025 81.005 107.305 ;
        RECT 81.225 107.115 81.575 107.285 ;
        RECT 79.355 106.695 79.885 106.865 ;
        RECT 76.150 105.935 77.875 106.105 ;
        RECT 76.405 104.925 76.575 105.765 ;
        RECT 76.785 105.095 77.035 105.935 ;
        RECT 77.245 104.925 77.415 105.765 ;
        RECT 77.585 105.095 77.875 105.935 ;
        RECT 78.085 104.925 78.255 105.985 ;
        RECT 78.430 105.645 78.600 106.265 ;
        RECT 78.945 106.155 79.485 106.525 ;
        RECT 79.665 106.415 79.885 106.695 ;
        RECT 80.055 106.245 80.225 107.025 ;
        RECT 79.820 106.075 80.225 106.245 ;
        RECT 80.395 106.235 80.745 106.855 ;
        RECT 79.820 105.985 79.990 106.075 ;
        RECT 80.915 106.065 81.125 106.855 ;
        RECT 78.770 105.815 79.990 105.985 ;
        RECT 80.450 105.905 81.125 106.065 ;
        RECT 78.430 105.475 79.230 105.645 ;
        RECT 78.550 104.925 78.880 105.305 ;
        RECT 79.060 105.185 79.230 105.475 ;
        RECT 79.820 105.435 79.990 105.815 ;
        RECT 80.160 105.895 81.125 105.905 ;
        RECT 81.315 106.725 81.575 107.115 ;
        RECT 81.785 107.015 82.115 107.475 ;
        RECT 82.990 107.085 83.845 107.255 ;
        RECT 84.050 107.085 84.545 107.255 ;
        RECT 84.715 107.115 85.045 107.475 ;
        RECT 81.315 106.035 81.485 106.725 ;
        RECT 81.655 106.375 81.825 106.555 ;
        RECT 81.995 106.545 82.785 106.795 ;
        RECT 82.990 106.375 83.160 107.085 ;
        RECT 83.330 106.575 83.685 106.795 ;
        RECT 81.655 106.205 83.345 106.375 ;
        RECT 80.160 105.605 80.620 105.895 ;
        RECT 81.315 105.865 82.815 106.035 ;
        RECT 81.315 105.725 81.485 105.865 ;
        RECT 80.925 105.555 81.485 105.725 ;
        RECT 79.400 104.925 79.650 105.385 ;
        RECT 79.820 105.095 80.690 105.435 ;
        RECT 80.925 105.095 81.095 105.555 ;
        RECT 81.930 105.525 83.005 105.695 ;
        RECT 81.265 104.925 81.635 105.385 ;
        RECT 81.930 105.185 82.100 105.525 ;
        RECT 82.270 104.925 82.600 105.355 ;
        RECT 82.835 105.185 83.005 105.525 ;
        RECT 83.175 105.425 83.345 106.205 ;
        RECT 83.515 105.985 83.685 106.575 ;
        RECT 83.855 106.175 84.205 106.795 ;
        RECT 83.515 105.595 83.980 105.985 ;
        RECT 84.375 105.725 84.545 107.085 ;
        RECT 84.715 105.895 85.175 106.945 ;
        RECT 84.150 105.555 84.545 105.725 ;
        RECT 84.150 105.425 84.320 105.555 ;
        RECT 83.175 105.095 83.855 105.425 ;
        RECT 84.070 105.095 84.320 105.425 ;
        RECT 84.490 104.925 84.740 105.385 ;
        RECT 84.910 105.110 85.235 105.895 ;
        RECT 85.405 105.095 85.575 107.215 ;
        RECT 85.745 107.095 86.075 107.475 ;
        RECT 86.245 106.925 86.500 107.215 ;
        RECT 85.750 106.755 86.500 106.925 ;
        RECT 87.225 106.925 87.395 107.305 ;
        RECT 87.575 107.095 87.905 107.475 ;
        RECT 87.225 106.755 87.890 106.925 ;
        RECT 88.085 106.800 88.345 107.305 ;
        RECT 85.750 105.765 85.980 106.755 ;
        RECT 86.150 105.935 86.500 106.585 ;
        RECT 87.155 106.205 87.485 106.575 ;
        RECT 87.720 106.500 87.890 106.755 ;
        RECT 87.720 106.170 88.005 106.500 ;
        RECT 87.720 106.025 87.890 106.170 ;
        RECT 87.225 105.855 87.890 106.025 ;
        RECT 88.175 106.000 88.345 106.800 ;
        RECT 88.515 106.750 88.805 107.475 ;
        RECT 89.285 107.005 89.455 107.475 ;
        RECT 89.625 106.825 89.955 107.305 ;
        RECT 90.125 107.005 90.295 107.475 ;
        RECT 90.465 106.825 90.795 107.305 ;
        RECT 89.030 106.655 90.795 106.825 ;
        RECT 90.965 106.665 91.135 107.475 ;
        RECT 91.335 107.095 92.405 107.265 ;
        RECT 91.335 106.740 91.655 107.095 ;
        RECT 89.030 106.105 89.440 106.655 ;
        RECT 91.330 106.485 91.655 106.740 ;
        RECT 89.625 106.275 91.655 106.485 ;
        RECT 91.310 106.265 91.655 106.275 ;
        RECT 91.825 106.525 92.065 106.925 ;
        RECT 92.235 106.865 92.405 107.095 ;
        RECT 92.575 107.035 92.765 107.475 ;
        RECT 92.935 107.025 93.885 107.305 ;
        RECT 94.105 107.115 94.455 107.285 ;
        RECT 92.235 106.695 92.765 106.865 ;
        RECT 85.750 105.595 86.500 105.765 ;
        RECT 85.745 104.925 86.075 105.425 ;
        RECT 86.245 105.095 86.500 105.595 ;
        RECT 87.225 105.095 87.395 105.855 ;
        RECT 87.575 104.925 87.905 105.685 ;
        RECT 88.075 105.095 88.345 106.000 ;
        RECT 88.515 104.925 88.805 106.090 ;
        RECT 89.030 105.935 90.755 106.105 ;
        RECT 89.285 104.925 89.455 105.765 ;
        RECT 89.665 105.095 89.915 105.935 ;
        RECT 90.125 104.925 90.295 105.765 ;
        RECT 90.465 105.095 90.755 105.935 ;
        RECT 90.965 104.925 91.135 105.985 ;
        RECT 91.310 105.645 91.480 106.265 ;
        RECT 91.825 106.155 92.365 106.525 ;
        RECT 92.545 106.415 92.765 106.695 ;
        RECT 92.935 106.245 93.105 107.025 ;
        RECT 92.700 106.075 93.105 106.245 ;
        RECT 93.275 106.235 93.625 106.855 ;
        RECT 92.700 105.985 92.870 106.075 ;
        RECT 93.795 106.065 94.005 106.855 ;
        RECT 91.650 105.815 92.870 105.985 ;
        RECT 93.330 105.905 94.005 106.065 ;
        RECT 91.310 105.475 92.110 105.645 ;
        RECT 91.430 104.925 91.760 105.305 ;
        RECT 91.940 105.185 92.110 105.475 ;
        RECT 92.700 105.435 92.870 105.815 ;
        RECT 93.040 105.895 94.005 105.905 ;
        RECT 94.195 106.725 94.455 107.115 ;
        RECT 94.665 107.015 94.995 107.475 ;
        RECT 95.870 107.085 96.725 107.255 ;
        RECT 96.930 107.085 97.425 107.255 ;
        RECT 97.595 107.115 97.925 107.475 ;
        RECT 94.195 106.035 94.365 106.725 ;
        RECT 94.535 106.375 94.705 106.555 ;
        RECT 94.875 106.545 95.665 106.795 ;
        RECT 95.870 106.375 96.040 107.085 ;
        RECT 96.210 106.575 96.565 106.795 ;
        RECT 94.535 106.205 96.225 106.375 ;
        RECT 93.040 105.605 93.500 105.895 ;
        RECT 94.195 105.865 95.695 106.035 ;
        RECT 94.195 105.725 94.365 105.865 ;
        RECT 93.805 105.555 94.365 105.725 ;
        RECT 92.280 104.925 92.530 105.385 ;
        RECT 92.700 105.095 93.570 105.435 ;
        RECT 93.805 105.095 93.975 105.555 ;
        RECT 94.810 105.525 95.885 105.695 ;
        RECT 94.145 104.925 94.515 105.385 ;
        RECT 94.810 105.185 94.980 105.525 ;
        RECT 95.150 104.925 95.480 105.355 ;
        RECT 95.715 105.185 95.885 105.525 ;
        RECT 96.055 105.425 96.225 106.205 ;
        RECT 96.395 105.985 96.565 106.575 ;
        RECT 96.735 106.175 97.085 106.795 ;
        RECT 96.395 105.595 96.860 105.985 ;
        RECT 97.255 105.725 97.425 107.085 ;
        RECT 97.595 105.895 98.055 106.945 ;
        RECT 97.030 105.555 97.425 105.725 ;
        RECT 97.030 105.425 97.200 105.555 ;
        RECT 96.055 105.095 96.735 105.425 ;
        RECT 96.950 105.095 97.200 105.425 ;
        RECT 97.370 104.925 97.620 105.385 ;
        RECT 97.790 105.110 98.115 105.895 ;
        RECT 98.285 105.095 98.455 107.215 ;
        RECT 98.625 107.095 98.955 107.475 ;
        RECT 99.125 106.925 99.380 107.215 ;
        RECT 98.630 106.755 99.380 106.925 ;
        RECT 98.630 105.765 98.860 106.755 ;
        RECT 99.615 106.655 99.825 107.475 ;
        RECT 99.995 106.675 100.325 107.305 ;
        RECT 99.030 105.935 99.380 106.585 ;
        RECT 99.995 106.075 100.245 106.675 ;
        RECT 100.495 106.655 100.725 107.475 ;
        RECT 100.935 106.725 102.145 107.475 ;
        RECT 100.415 106.235 100.745 106.485 ;
        RECT 98.630 105.595 99.380 105.765 ;
        RECT 98.625 104.925 98.955 105.425 ;
        RECT 99.125 105.095 99.380 105.595 ;
        RECT 99.615 104.925 99.825 106.065 ;
        RECT 99.995 105.095 100.325 106.075 ;
        RECT 100.495 104.925 100.725 106.065 ;
        RECT 100.935 106.015 101.455 106.555 ;
        RECT 101.625 106.185 102.145 106.725 ;
        RECT 102.355 106.655 102.585 107.475 ;
        RECT 102.755 106.675 103.085 107.305 ;
        RECT 102.335 106.235 102.665 106.485 ;
        RECT 102.835 106.075 103.085 106.675 ;
        RECT 103.255 106.655 103.465 107.475 ;
        RECT 104.005 107.005 104.175 107.475 ;
        RECT 104.345 106.825 104.675 107.305 ;
        RECT 104.845 107.005 105.015 107.475 ;
        RECT 105.185 106.825 105.515 107.305 ;
        RECT 103.750 106.655 105.515 106.825 ;
        RECT 105.685 106.665 105.855 107.475 ;
        RECT 106.055 107.095 107.125 107.265 ;
        RECT 106.055 106.740 106.375 107.095 ;
        RECT 100.935 104.925 102.145 106.015 ;
        RECT 102.355 104.925 102.585 106.065 ;
        RECT 102.755 105.095 103.085 106.075 ;
        RECT 103.750 106.105 104.160 106.655 ;
        RECT 106.050 106.485 106.375 106.740 ;
        RECT 104.345 106.275 106.375 106.485 ;
        RECT 106.030 106.265 106.375 106.275 ;
        RECT 106.545 106.525 106.785 106.925 ;
        RECT 106.955 106.865 107.125 107.095 ;
        RECT 107.295 107.035 107.485 107.475 ;
        RECT 107.655 107.025 108.605 107.305 ;
        RECT 108.825 107.115 109.175 107.285 ;
        RECT 106.955 106.695 107.485 106.865 ;
        RECT 103.255 104.925 103.465 106.065 ;
        RECT 103.750 105.935 105.475 106.105 ;
        RECT 104.005 104.925 104.175 105.765 ;
        RECT 104.385 105.095 104.635 105.935 ;
        RECT 104.845 104.925 105.015 105.765 ;
        RECT 105.185 105.095 105.475 105.935 ;
        RECT 105.685 104.925 105.855 105.985 ;
        RECT 106.030 105.645 106.200 106.265 ;
        RECT 106.545 106.155 107.085 106.525 ;
        RECT 107.265 106.415 107.485 106.695 ;
        RECT 107.655 106.245 107.825 107.025 ;
        RECT 107.420 106.075 107.825 106.245 ;
        RECT 107.995 106.235 108.345 106.855 ;
        RECT 107.420 105.985 107.590 106.075 ;
        RECT 108.515 106.065 108.725 106.855 ;
        RECT 106.370 105.815 107.590 105.985 ;
        RECT 108.050 105.905 108.725 106.065 ;
        RECT 106.030 105.475 106.830 105.645 ;
        RECT 106.150 104.925 106.480 105.305 ;
        RECT 106.660 105.185 106.830 105.475 ;
        RECT 107.420 105.435 107.590 105.815 ;
        RECT 107.760 105.895 108.725 105.905 ;
        RECT 108.915 106.725 109.175 107.115 ;
        RECT 109.385 107.015 109.715 107.475 ;
        RECT 110.590 107.085 111.445 107.255 ;
        RECT 111.650 107.085 112.145 107.255 ;
        RECT 112.315 107.115 112.645 107.475 ;
        RECT 108.915 106.035 109.085 106.725 ;
        RECT 109.255 106.375 109.425 106.555 ;
        RECT 109.595 106.545 110.385 106.795 ;
        RECT 110.590 106.375 110.760 107.085 ;
        RECT 110.930 106.575 111.285 106.795 ;
        RECT 109.255 106.205 110.945 106.375 ;
        RECT 107.760 105.605 108.220 105.895 ;
        RECT 108.915 105.865 110.415 106.035 ;
        RECT 108.915 105.725 109.085 105.865 ;
        RECT 108.525 105.555 109.085 105.725 ;
        RECT 107.000 104.925 107.250 105.385 ;
        RECT 107.420 105.095 108.290 105.435 ;
        RECT 108.525 105.095 108.695 105.555 ;
        RECT 109.530 105.525 110.605 105.695 ;
        RECT 108.865 104.925 109.235 105.385 ;
        RECT 109.530 105.185 109.700 105.525 ;
        RECT 109.870 104.925 110.200 105.355 ;
        RECT 110.435 105.185 110.605 105.525 ;
        RECT 110.775 105.425 110.945 106.205 ;
        RECT 111.115 105.985 111.285 106.575 ;
        RECT 111.455 106.175 111.805 106.795 ;
        RECT 111.115 105.595 111.580 105.985 ;
        RECT 111.975 105.725 112.145 107.085 ;
        RECT 112.315 105.895 112.775 106.945 ;
        RECT 111.750 105.555 112.145 105.725 ;
        RECT 111.750 105.425 111.920 105.555 ;
        RECT 110.775 105.095 111.455 105.425 ;
        RECT 111.670 105.095 111.920 105.425 ;
        RECT 112.090 104.925 112.340 105.385 ;
        RECT 112.510 105.110 112.835 105.895 ;
        RECT 113.005 105.095 113.175 107.215 ;
        RECT 113.345 107.095 113.675 107.475 ;
        RECT 113.845 106.925 114.100 107.215 ;
        RECT 113.350 106.755 114.100 106.925 ;
        RECT 113.350 105.765 113.580 106.755 ;
        RECT 114.275 106.750 114.565 107.475 ;
        RECT 115.660 106.925 115.915 107.215 ;
        RECT 116.085 107.095 116.415 107.475 ;
        RECT 115.660 106.755 116.410 106.925 ;
        RECT 113.750 105.935 114.100 106.585 ;
        RECT 113.350 105.595 114.100 105.765 ;
        RECT 113.345 104.925 113.675 105.425 ;
        RECT 113.845 105.095 114.100 105.595 ;
        RECT 114.275 104.925 114.565 106.090 ;
        RECT 115.660 105.935 116.010 106.585 ;
        RECT 116.180 105.765 116.410 106.755 ;
        RECT 115.660 105.595 116.410 105.765 ;
        RECT 115.660 105.095 115.915 105.595 ;
        RECT 116.085 104.925 116.415 105.425 ;
        RECT 116.585 105.095 116.755 107.215 ;
        RECT 117.115 107.115 117.445 107.475 ;
        RECT 117.615 107.085 118.110 107.255 ;
        RECT 118.315 107.085 119.170 107.255 ;
        RECT 116.985 105.895 117.445 106.945 ;
        RECT 116.925 105.110 117.250 105.895 ;
        RECT 117.615 105.725 117.785 107.085 ;
        RECT 117.955 106.175 118.305 106.795 ;
        RECT 118.475 106.575 118.830 106.795 ;
        RECT 118.475 105.985 118.645 106.575 ;
        RECT 119.000 106.375 119.170 107.085 ;
        RECT 120.045 107.015 120.375 107.475 ;
        RECT 120.585 107.115 120.935 107.285 ;
        RECT 119.375 106.545 120.165 106.795 ;
        RECT 120.585 106.725 120.845 107.115 ;
        RECT 121.155 107.025 122.105 107.305 ;
        RECT 122.275 107.035 122.465 107.475 ;
        RECT 122.635 107.095 123.705 107.265 ;
        RECT 120.335 106.375 120.505 106.555 ;
        RECT 117.615 105.555 118.010 105.725 ;
        RECT 118.180 105.595 118.645 105.985 ;
        RECT 118.815 106.205 120.505 106.375 ;
        RECT 117.840 105.425 118.010 105.555 ;
        RECT 118.815 105.425 118.985 106.205 ;
        RECT 120.675 106.035 120.845 106.725 ;
        RECT 119.345 105.865 120.845 106.035 ;
        RECT 121.035 106.065 121.245 106.855 ;
        RECT 121.415 106.235 121.765 106.855 ;
        RECT 121.935 106.245 122.105 107.025 ;
        RECT 122.635 106.865 122.805 107.095 ;
        RECT 122.275 106.695 122.805 106.865 ;
        RECT 122.275 106.415 122.495 106.695 ;
        RECT 122.975 106.525 123.215 106.925 ;
        RECT 121.935 106.075 122.340 106.245 ;
        RECT 122.675 106.155 123.215 106.525 ;
        RECT 123.385 106.740 123.705 107.095 ;
        RECT 123.385 106.485 123.710 106.740 ;
        RECT 123.905 106.665 124.075 107.475 ;
        RECT 124.245 106.825 124.575 107.305 ;
        RECT 124.745 107.005 124.915 107.475 ;
        RECT 125.085 106.825 125.415 107.305 ;
        RECT 125.585 107.005 125.755 107.475 ;
        RECT 124.245 106.655 126.010 106.825 ;
        RECT 126.235 106.725 127.445 107.475 ;
        RECT 123.385 106.275 125.415 106.485 ;
        RECT 123.385 106.265 123.730 106.275 ;
        RECT 121.035 105.905 121.710 106.065 ;
        RECT 122.170 105.985 122.340 106.075 ;
        RECT 121.035 105.895 122.000 105.905 ;
        RECT 120.675 105.725 120.845 105.865 ;
        RECT 117.420 104.925 117.670 105.385 ;
        RECT 117.840 105.095 118.090 105.425 ;
        RECT 118.305 105.095 118.985 105.425 ;
        RECT 119.155 105.525 120.230 105.695 ;
        RECT 120.675 105.555 121.235 105.725 ;
        RECT 121.540 105.605 122.000 105.895 ;
        RECT 122.170 105.815 123.390 105.985 ;
        RECT 119.155 105.185 119.325 105.525 ;
        RECT 119.560 104.925 119.890 105.355 ;
        RECT 120.060 105.185 120.230 105.525 ;
        RECT 120.525 104.925 120.895 105.385 ;
        RECT 121.065 105.095 121.235 105.555 ;
        RECT 122.170 105.435 122.340 105.815 ;
        RECT 123.560 105.645 123.730 106.265 ;
        RECT 125.600 106.105 126.010 106.655 ;
        RECT 121.470 105.095 122.340 105.435 ;
        RECT 122.930 105.475 123.730 105.645 ;
        RECT 122.510 104.925 122.760 105.385 ;
        RECT 122.930 105.185 123.100 105.475 ;
        RECT 123.280 104.925 123.610 105.305 ;
        RECT 123.905 104.925 124.075 105.985 ;
        RECT 124.285 105.935 126.010 106.105 ;
        RECT 126.235 106.015 126.755 106.555 ;
        RECT 126.925 106.185 127.445 106.725 ;
        RECT 124.285 105.095 124.575 105.935 ;
        RECT 124.745 104.925 124.915 105.765 ;
        RECT 125.125 105.095 125.375 105.935 ;
        RECT 125.585 104.925 125.755 105.765 ;
        RECT 126.235 104.925 127.445 106.015 ;
        RECT 14.370 104.755 127.530 104.925 ;
        RECT 14.455 103.665 15.665 104.755 ;
        RECT 14.455 102.955 14.975 103.495 ;
        RECT 15.145 103.125 15.665 103.665 ;
        RECT 15.835 103.665 18.425 104.755 ;
        RECT 18.600 104.320 23.945 104.755 ;
        RECT 15.835 103.145 17.045 103.665 ;
        RECT 17.215 102.975 18.425 103.495 ;
        RECT 20.190 103.070 20.540 104.320 ;
        RECT 24.115 103.590 24.405 104.755 ;
        RECT 24.575 103.665 27.165 104.755 ;
        RECT 14.455 102.205 15.665 102.955 ;
        RECT 15.835 102.205 18.425 102.975 ;
        RECT 22.020 102.750 22.360 103.580 ;
        RECT 24.575 103.145 25.785 103.665 ;
        RECT 27.375 103.615 27.605 104.755 ;
        RECT 27.775 103.605 28.105 104.585 ;
        RECT 28.275 103.615 28.485 104.755 ;
        RECT 28.720 104.085 28.975 104.585 ;
        RECT 29.145 104.255 29.475 104.755 ;
        RECT 28.720 103.915 29.470 104.085 ;
        RECT 25.955 102.975 27.165 103.495 ;
        RECT 27.355 103.195 27.685 103.445 ;
        RECT 18.600 102.205 23.945 102.750 ;
        RECT 24.115 102.205 24.405 102.930 ;
        RECT 24.575 102.205 27.165 102.975 ;
        RECT 27.375 102.205 27.605 103.025 ;
        RECT 27.855 103.005 28.105 103.605 ;
        RECT 28.720 103.095 29.070 103.745 ;
        RECT 27.775 102.375 28.105 103.005 ;
        RECT 28.275 102.205 28.485 103.025 ;
        RECT 29.240 102.925 29.470 103.915 ;
        RECT 28.720 102.755 29.470 102.925 ;
        RECT 28.720 102.465 28.975 102.755 ;
        RECT 29.145 102.205 29.475 102.585 ;
        RECT 29.645 102.465 29.815 104.585 ;
        RECT 29.985 103.785 30.310 104.570 ;
        RECT 30.480 104.295 30.730 104.755 ;
        RECT 30.900 104.255 31.150 104.585 ;
        RECT 31.365 104.255 32.045 104.585 ;
        RECT 30.900 104.125 31.070 104.255 ;
        RECT 30.675 103.955 31.070 104.125 ;
        RECT 30.045 102.735 30.505 103.785 ;
        RECT 30.675 102.595 30.845 103.955 ;
        RECT 31.240 103.695 31.705 104.085 ;
        RECT 31.015 102.885 31.365 103.505 ;
        RECT 31.535 103.105 31.705 103.695 ;
        RECT 31.875 103.475 32.045 104.255 ;
        RECT 32.215 104.155 32.385 104.495 ;
        RECT 32.620 104.325 32.950 104.755 ;
        RECT 33.120 104.155 33.290 104.495 ;
        RECT 33.585 104.295 33.955 104.755 ;
        RECT 32.215 103.985 33.290 104.155 ;
        RECT 34.125 104.125 34.295 104.585 ;
        RECT 34.530 104.245 35.400 104.585 ;
        RECT 35.570 104.295 35.820 104.755 ;
        RECT 33.735 103.955 34.295 104.125 ;
        RECT 33.735 103.815 33.905 103.955 ;
        RECT 32.405 103.645 33.905 103.815 ;
        RECT 34.600 103.785 35.060 104.075 ;
        RECT 31.875 103.305 33.565 103.475 ;
        RECT 31.535 102.885 31.890 103.105 ;
        RECT 32.060 102.595 32.230 103.305 ;
        RECT 32.435 102.885 33.225 103.135 ;
        RECT 33.395 103.125 33.565 103.305 ;
        RECT 33.735 102.955 33.905 103.645 ;
        RECT 30.175 102.205 30.505 102.565 ;
        RECT 30.675 102.425 31.170 102.595 ;
        RECT 31.375 102.425 32.230 102.595 ;
        RECT 33.105 102.205 33.435 102.665 ;
        RECT 33.645 102.565 33.905 102.955 ;
        RECT 34.095 103.775 35.060 103.785 ;
        RECT 35.230 103.865 35.400 104.245 ;
        RECT 35.990 104.205 36.160 104.495 ;
        RECT 36.340 104.375 36.670 104.755 ;
        RECT 35.990 104.035 36.790 104.205 ;
        RECT 34.095 103.615 34.770 103.775 ;
        RECT 35.230 103.695 36.450 103.865 ;
        RECT 34.095 102.825 34.305 103.615 ;
        RECT 35.230 103.605 35.400 103.695 ;
        RECT 34.475 102.825 34.825 103.445 ;
        RECT 34.995 103.435 35.400 103.605 ;
        RECT 34.995 102.655 35.165 103.435 ;
        RECT 35.335 102.985 35.555 103.265 ;
        RECT 35.735 103.155 36.275 103.525 ;
        RECT 36.620 103.415 36.790 104.035 ;
        RECT 36.965 103.695 37.135 104.755 ;
        RECT 37.345 103.745 37.635 104.585 ;
        RECT 37.805 103.915 37.975 104.755 ;
        RECT 38.185 103.745 38.435 104.585 ;
        RECT 38.645 103.915 38.815 104.755 ;
        RECT 39.605 103.915 39.775 104.755 ;
        RECT 39.985 103.745 40.235 104.585 ;
        RECT 40.445 103.915 40.615 104.755 ;
        RECT 40.785 103.745 41.075 104.585 ;
        RECT 37.345 103.575 39.070 103.745 ;
        RECT 35.335 102.815 35.865 102.985 ;
        RECT 33.645 102.395 33.995 102.565 ;
        RECT 34.215 102.375 35.165 102.655 ;
        RECT 35.335 102.205 35.525 102.645 ;
        RECT 35.695 102.585 35.865 102.815 ;
        RECT 36.035 102.755 36.275 103.155 ;
        RECT 36.445 103.405 36.790 103.415 ;
        RECT 36.445 103.195 38.475 103.405 ;
        RECT 36.445 102.940 36.770 103.195 ;
        RECT 38.660 103.025 39.070 103.575 ;
        RECT 36.445 102.585 36.765 102.940 ;
        RECT 35.695 102.415 36.765 102.585 ;
        RECT 36.965 102.205 37.135 103.015 ;
        RECT 37.305 102.855 39.070 103.025 ;
        RECT 39.350 103.575 41.075 103.745 ;
        RECT 41.285 103.695 41.455 104.755 ;
        RECT 41.750 104.375 42.080 104.755 ;
        RECT 42.260 104.205 42.430 104.495 ;
        RECT 42.600 104.295 42.850 104.755 ;
        RECT 41.630 104.035 42.430 104.205 ;
        RECT 43.020 104.245 43.890 104.585 ;
        RECT 39.350 103.025 39.760 103.575 ;
        RECT 41.630 103.415 41.800 104.035 ;
        RECT 43.020 103.865 43.190 104.245 ;
        RECT 44.125 104.125 44.295 104.585 ;
        RECT 44.465 104.295 44.835 104.755 ;
        RECT 45.130 104.155 45.300 104.495 ;
        RECT 45.470 104.325 45.800 104.755 ;
        RECT 46.035 104.155 46.205 104.495 ;
        RECT 41.970 103.695 43.190 103.865 ;
        RECT 43.360 103.785 43.820 104.075 ;
        RECT 44.125 103.955 44.685 104.125 ;
        RECT 45.130 103.985 46.205 104.155 ;
        RECT 46.375 104.255 47.055 104.585 ;
        RECT 47.270 104.255 47.520 104.585 ;
        RECT 47.690 104.295 47.940 104.755 ;
        RECT 44.515 103.815 44.685 103.955 ;
        RECT 43.360 103.775 44.325 103.785 ;
        RECT 43.020 103.605 43.190 103.695 ;
        RECT 43.650 103.615 44.325 103.775 ;
        RECT 41.630 103.405 41.975 103.415 ;
        RECT 39.945 103.195 41.975 103.405 ;
        RECT 39.350 102.855 41.115 103.025 ;
        RECT 37.305 102.375 37.635 102.855 ;
        RECT 37.805 102.205 37.975 102.675 ;
        RECT 38.145 102.375 38.475 102.855 ;
        RECT 38.645 102.205 38.815 102.675 ;
        RECT 39.605 102.205 39.775 102.675 ;
        RECT 39.945 102.375 40.275 102.855 ;
        RECT 40.445 102.205 40.615 102.675 ;
        RECT 40.785 102.375 41.115 102.855 ;
        RECT 41.285 102.205 41.455 103.015 ;
        RECT 41.650 102.940 41.975 103.195 ;
        RECT 41.655 102.585 41.975 102.940 ;
        RECT 42.145 103.155 42.685 103.525 ;
        RECT 43.020 103.435 43.425 103.605 ;
        RECT 42.145 102.755 42.385 103.155 ;
        RECT 42.865 102.985 43.085 103.265 ;
        RECT 42.555 102.815 43.085 102.985 ;
        RECT 42.555 102.585 42.725 102.815 ;
        RECT 43.255 102.655 43.425 103.435 ;
        RECT 43.595 102.825 43.945 103.445 ;
        RECT 44.115 102.825 44.325 103.615 ;
        RECT 44.515 103.645 46.015 103.815 ;
        RECT 44.515 102.955 44.685 103.645 ;
        RECT 46.375 103.475 46.545 104.255 ;
        RECT 47.350 104.125 47.520 104.255 ;
        RECT 44.855 103.305 46.545 103.475 ;
        RECT 46.715 103.695 47.180 104.085 ;
        RECT 47.350 103.955 47.745 104.125 ;
        RECT 44.855 103.125 45.025 103.305 ;
        RECT 41.655 102.415 42.725 102.585 ;
        RECT 42.895 102.205 43.085 102.645 ;
        RECT 43.255 102.375 44.205 102.655 ;
        RECT 44.515 102.565 44.775 102.955 ;
        RECT 45.195 102.885 45.985 103.135 ;
        RECT 44.425 102.395 44.775 102.565 ;
        RECT 44.985 102.205 45.315 102.665 ;
        RECT 46.190 102.595 46.360 103.305 ;
        RECT 46.715 103.105 46.885 103.695 ;
        RECT 46.530 102.885 46.885 103.105 ;
        RECT 47.055 102.885 47.405 103.505 ;
        RECT 47.575 102.595 47.745 103.955 ;
        RECT 48.110 103.785 48.435 104.570 ;
        RECT 47.915 102.735 48.375 103.785 ;
        RECT 46.190 102.425 47.045 102.595 ;
        RECT 47.250 102.425 47.745 102.595 ;
        RECT 47.915 102.205 48.245 102.565 ;
        RECT 48.605 102.465 48.775 104.585 ;
        RECT 48.945 104.255 49.275 104.755 ;
        RECT 49.445 104.085 49.700 104.585 ;
        RECT 48.950 103.915 49.700 104.085 ;
        RECT 48.950 102.925 49.180 103.915 ;
        RECT 49.350 103.095 49.700 103.745 ;
        RECT 49.875 103.590 50.165 104.755 ;
        RECT 51.315 103.615 51.525 104.755 ;
        RECT 51.695 103.605 52.025 104.585 ;
        RECT 52.195 103.615 52.425 104.755 ;
        RECT 52.945 103.915 53.115 104.755 ;
        RECT 53.325 103.745 53.575 104.585 ;
        RECT 53.785 103.915 53.955 104.755 ;
        RECT 54.125 103.745 54.415 104.585 ;
        RECT 48.950 102.755 49.700 102.925 ;
        RECT 48.945 102.205 49.275 102.585 ;
        RECT 49.445 102.465 49.700 102.755 ;
        RECT 49.875 102.205 50.165 102.930 ;
        RECT 51.315 102.205 51.525 103.025 ;
        RECT 51.695 103.005 51.945 103.605 ;
        RECT 52.690 103.575 54.415 103.745 ;
        RECT 54.625 103.695 54.795 104.755 ;
        RECT 55.090 104.375 55.420 104.755 ;
        RECT 55.600 104.205 55.770 104.495 ;
        RECT 55.940 104.295 56.190 104.755 ;
        RECT 54.970 104.035 55.770 104.205 ;
        RECT 56.360 104.245 57.230 104.585 ;
        RECT 52.115 103.195 52.445 103.445 ;
        RECT 52.690 103.025 53.100 103.575 ;
        RECT 54.970 103.415 55.140 104.035 ;
        RECT 56.360 103.865 56.530 104.245 ;
        RECT 57.465 104.125 57.635 104.585 ;
        RECT 57.805 104.295 58.175 104.755 ;
        RECT 58.470 104.155 58.640 104.495 ;
        RECT 58.810 104.325 59.140 104.755 ;
        RECT 59.375 104.155 59.545 104.495 ;
        RECT 55.310 103.695 56.530 103.865 ;
        RECT 56.700 103.785 57.160 104.075 ;
        RECT 57.465 103.955 58.025 104.125 ;
        RECT 58.470 103.985 59.545 104.155 ;
        RECT 59.715 104.255 60.395 104.585 ;
        RECT 60.610 104.255 60.860 104.585 ;
        RECT 61.030 104.295 61.280 104.755 ;
        RECT 57.855 103.815 58.025 103.955 ;
        RECT 56.700 103.775 57.665 103.785 ;
        RECT 56.360 103.605 56.530 103.695 ;
        RECT 56.990 103.615 57.665 103.775 ;
        RECT 54.970 103.405 55.315 103.415 ;
        RECT 53.285 103.195 55.315 103.405 ;
        RECT 51.695 102.375 52.025 103.005 ;
        RECT 52.195 102.205 52.425 103.025 ;
        RECT 52.690 102.855 54.455 103.025 ;
        RECT 52.945 102.205 53.115 102.675 ;
        RECT 53.285 102.375 53.615 102.855 ;
        RECT 53.785 102.205 53.955 102.675 ;
        RECT 54.125 102.375 54.455 102.855 ;
        RECT 54.625 102.205 54.795 103.015 ;
        RECT 54.990 102.940 55.315 103.195 ;
        RECT 54.995 102.585 55.315 102.940 ;
        RECT 55.485 103.155 56.025 103.525 ;
        RECT 56.360 103.435 56.765 103.605 ;
        RECT 55.485 102.755 55.725 103.155 ;
        RECT 56.205 102.985 56.425 103.265 ;
        RECT 55.895 102.815 56.425 102.985 ;
        RECT 55.895 102.585 56.065 102.815 ;
        RECT 56.595 102.655 56.765 103.435 ;
        RECT 56.935 102.825 57.285 103.445 ;
        RECT 57.455 102.825 57.665 103.615 ;
        RECT 57.855 103.645 59.355 103.815 ;
        RECT 57.855 102.955 58.025 103.645 ;
        RECT 59.715 103.475 59.885 104.255 ;
        RECT 60.690 104.125 60.860 104.255 ;
        RECT 58.195 103.305 59.885 103.475 ;
        RECT 60.055 103.695 60.520 104.085 ;
        RECT 60.690 103.955 61.085 104.125 ;
        RECT 58.195 103.125 58.365 103.305 ;
        RECT 54.995 102.415 56.065 102.585 ;
        RECT 56.235 102.205 56.425 102.645 ;
        RECT 56.595 102.375 57.545 102.655 ;
        RECT 57.855 102.565 58.115 102.955 ;
        RECT 58.535 102.885 59.325 103.135 ;
        RECT 57.765 102.395 58.115 102.565 ;
        RECT 58.325 102.205 58.655 102.665 ;
        RECT 59.530 102.595 59.700 103.305 ;
        RECT 60.055 103.105 60.225 103.695 ;
        RECT 59.870 102.885 60.225 103.105 ;
        RECT 60.395 102.885 60.745 103.505 ;
        RECT 60.915 102.595 61.085 103.955 ;
        RECT 61.450 103.785 61.775 104.570 ;
        RECT 61.255 102.735 61.715 103.785 ;
        RECT 59.530 102.425 60.385 102.595 ;
        RECT 60.590 102.425 61.085 102.595 ;
        RECT 61.255 102.205 61.585 102.565 ;
        RECT 61.945 102.465 62.115 104.585 ;
        RECT 62.285 104.255 62.615 104.755 ;
        RECT 62.785 104.085 63.040 104.585 ;
        RECT 62.290 103.915 63.040 104.085 ;
        RECT 63.525 103.915 63.695 104.755 ;
        RECT 62.290 102.925 62.520 103.915 ;
        RECT 63.905 103.745 64.155 104.585 ;
        RECT 64.365 103.915 64.535 104.755 ;
        RECT 64.705 103.745 64.995 104.585 ;
        RECT 62.690 103.095 63.040 103.745 ;
        RECT 63.270 103.575 64.995 103.745 ;
        RECT 65.205 103.695 65.375 104.755 ;
        RECT 65.670 104.375 66.000 104.755 ;
        RECT 66.180 104.205 66.350 104.495 ;
        RECT 66.520 104.295 66.770 104.755 ;
        RECT 65.550 104.035 66.350 104.205 ;
        RECT 66.940 104.245 67.810 104.585 ;
        RECT 63.270 103.025 63.680 103.575 ;
        RECT 65.550 103.415 65.720 104.035 ;
        RECT 66.940 103.865 67.110 104.245 ;
        RECT 68.045 104.125 68.215 104.585 ;
        RECT 68.385 104.295 68.755 104.755 ;
        RECT 69.050 104.155 69.220 104.495 ;
        RECT 69.390 104.325 69.720 104.755 ;
        RECT 69.955 104.155 70.125 104.495 ;
        RECT 65.890 103.695 67.110 103.865 ;
        RECT 67.280 103.785 67.740 104.075 ;
        RECT 68.045 103.955 68.605 104.125 ;
        RECT 69.050 103.985 70.125 104.155 ;
        RECT 70.295 104.255 70.975 104.585 ;
        RECT 71.190 104.255 71.440 104.585 ;
        RECT 71.610 104.295 71.860 104.755 ;
        RECT 68.435 103.815 68.605 103.955 ;
        RECT 67.280 103.775 68.245 103.785 ;
        RECT 66.940 103.605 67.110 103.695 ;
        RECT 67.570 103.615 68.245 103.775 ;
        RECT 65.550 103.405 65.895 103.415 ;
        RECT 63.865 103.195 65.895 103.405 ;
        RECT 62.290 102.755 63.040 102.925 ;
        RECT 63.270 102.855 65.035 103.025 ;
        RECT 62.285 102.205 62.615 102.585 ;
        RECT 62.785 102.465 63.040 102.755 ;
        RECT 63.525 102.205 63.695 102.675 ;
        RECT 63.865 102.375 64.195 102.855 ;
        RECT 64.365 102.205 64.535 102.675 ;
        RECT 64.705 102.375 65.035 102.855 ;
        RECT 65.205 102.205 65.375 103.015 ;
        RECT 65.570 102.940 65.895 103.195 ;
        RECT 65.575 102.585 65.895 102.940 ;
        RECT 66.065 103.155 66.605 103.525 ;
        RECT 66.940 103.435 67.345 103.605 ;
        RECT 66.065 102.755 66.305 103.155 ;
        RECT 66.785 102.985 67.005 103.265 ;
        RECT 66.475 102.815 67.005 102.985 ;
        RECT 66.475 102.585 66.645 102.815 ;
        RECT 67.175 102.655 67.345 103.435 ;
        RECT 67.515 102.825 67.865 103.445 ;
        RECT 68.035 102.825 68.245 103.615 ;
        RECT 68.435 103.645 69.935 103.815 ;
        RECT 68.435 102.955 68.605 103.645 ;
        RECT 70.295 103.475 70.465 104.255 ;
        RECT 71.270 104.125 71.440 104.255 ;
        RECT 68.775 103.305 70.465 103.475 ;
        RECT 70.635 103.695 71.100 104.085 ;
        RECT 71.270 103.955 71.665 104.125 ;
        RECT 68.775 103.125 68.945 103.305 ;
        RECT 65.575 102.415 66.645 102.585 ;
        RECT 66.815 102.205 67.005 102.645 ;
        RECT 67.175 102.375 68.125 102.655 ;
        RECT 68.435 102.565 68.695 102.955 ;
        RECT 69.115 102.885 69.905 103.135 ;
        RECT 68.345 102.395 68.695 102.565 ;
        RECT 68.905 102.205 69.235 102.665 ;
        RECT 70.110 102.595 70.280 103.305 ;
        RECT 70.635 103.105 70.805 103.695 ;
        RECT 70.450 102.885 70.805 103.105 ;
        RECT 70.975 102.885 71.325 103.505 ;
        RECT 71.495 102.595 71.665 103.955 ;
        RECT 72.030 103.785 72.355 104.570 ;
        RECT 71.835 102.735 72.295 103.785 ;
        RECT 70.110 102.425 70.965 102.595 ;
        RECT 71.170 102.425 71.665 102.595 ;
        RECT 71.835 102.205 72.165 102.565 ;
        RECT 72.525 102.465 72.695 104.585 ;
        RECT 72.865 104.255 73.195 104.755 ;
        RECT 73.365 104.085 73.620 104.585 ;
        RECT 72.870 103.915 73.620 104.085 ;
        RECT 72.870 102.925 73.100 103.915 ;
        RECT 73.270 103.095 73.620 103.745 ;
        RECT 73.795 103.665 75.465 104.755 ;
        RECT 73.795 103.145 74.545 103.665 ;
        RECT 75.635 103.590 75.925 104.755 ;
        RECT 76.405 103.915 76.575 104.755 ;
        RECT 76.785 103.745 77.035 104.585 ;
        RECT 77.245 103.915 77.415 104.755 ;
        RECT 77.585 103.745 77.875 104.585 ;
        RECT 76.150 103.575 77.875 103.745 ;
        RECT 78.085 103.695 78.255 104.755 ;
        RECT 78.550 104.375 78.880 104.755 ;
        RECT 79.060 104.205 79.230 104.495 ;
        RECT 79.400 104.295 79.650 104.755 ;
        RECT 78.430 104.035 79.230 104.205 ;
        RECT 79.820 104.245 80.690 104.585 ;
        RECT 74.715 102.975 75.465 103.495 ;
        RECT 72.870 102.755 73.620 102.925 ;
        RECT 72.865 102.205 73.195 102.585 ;
        RECT 73.365 102.465 73.620 102.755 ;
        RECT 73.795 102.205 75.465 102.975 ;
        RECT 76.150 103.025 76.560 103.575 ;
        RECT 78.430 103.415 78.600 104.035 ;
        RECT 79.820 103.865 79.990 104.245 ;
        RECT 80.925 104.125 81.095 104.585 ;
        RECT 81.265 104.295 81.635 104.755 ;
        RECT 81.930 104.155 82.100 104.495 ;
        RECT 82.270 104.325 82.600 104.755 ;
        RECT 82.835 104.155 83.005 104.495 ;
        RECT 78.770 103.695 79.990 103.865 ;
        RECT 80.160 103.785 80.620 104.075 ;
        RECT 80.925 103.955 81.485 104.125 ;
        RECT 81.930 103.985 83.005 104.155 ;
        RECT 83.175 104.255 83.855 104.585 ;
        RECT 84.070 104.255 84.320 104.585 ;
        RECT 84.490 104.295 84.740 104.755 ;
        RECT 81.315 103.815 81.485 103.955 ;
        RECT 80.160 103.775 81.125 103.785 ;
        RECT 79.820 103.605 79.990 103.695 ;
        RECT 80.450 103.615 81.125 103.775 ;
        RECT 78.430 103.405 78.775 103.415 ;
        RECT 76.745 103.195 78.775 103.405 ;
        RECT 75.635 102.205 75.925 102.930 ;
        RECT 76.150 102.855 77.915 103.025 ;
        RECT 76.405 102.205 76.575 102.675 ;
        RECT 76.745 102.375 77.075 102.855 ;
        RECT 77.245 102.205 77.415 102.675 ;
        RECT 77.585 102.375 77.915 102.855 ;
        RECT 78.085 102.205 78.255 103.015 ;
        RECT 78.450 102.940 78.775 103.195 ;
        RECT 78.455 102.585 78.775 102.940 ;
        RECT 78.945 103.155 79.485 103.525 ;
        RECT 79.820 103.435 80.225 103.605 ;
        RECT 78.945 102.755 79.185 103.155 ;
        RECT 79.665 102.985 79.885 103.265 ;
        RECT 79.355 102.815 79.885 102.985 ;
        RECT 79.355 102.585 79.525 102.815 ;
        RECT 80.055 102.655 80.225 103.435 ;
        RECT 80.395 102.825 80.745 103.445 ;
        RECT 80.915 102.825 81.125 103.615 ;
        RECT 81.315 103.645 82.815 103.815 ;
        RECT 81.315 102.955 81.485 103.645 ;
        RECT 83.175 103.475 83.345 104.255 ;
        RECT 84.150 104.125 84.320 104.255 ;
        RECT 81.655 103.305 83.345 103.475 ;
        RECT 83.515 103.695 83.980 104.085 ;
        RECT 84.150 103.955 84.545 104.125 ;
        RECT 81.655 103.125 81.825 103.305 ;
        RECT 78.455 102.415 79.525 102.585 ;
        RECT 79.695 102.205 79.885 102.645 ;
        RECT 80.055 102.375 81.005 102.655 ;
        RECT 81.315 102.565 81.575 102.955 ;
        RECT 81.995 102.885 82.785 103.135 ;
        RECT 81.225 102.395 81.575 102.565 ;
        RECT 81.785 102.205 82.115 102.665 ;
        RECT 82.990 102.595 83.160 103.305 ;
        RECT 83.515 103.105 83.685 103.695 ;
        RECT 83.330 102.885 83.685 103.105 ;
        RECT 83.855 102.885 84.205 103.505 ;
        RECT 84.375 102.595 84.545 103.955 ;
        RECT 84.910 103.785 85.235 104.570 ;
        RECT 84.715 102.735 85.175 103.785 ;
        RECT 82.990 102.425 83.845 102.595 ;
        RECT 84.050 102.425 84.545 102.595 ;
        RECT 84.715 102.205 85.045 102.565 ;
        RECT 85.405 102.465 85.575 104.585 ;
        RECT 85.745 104.255 86.075 104.755 ;
        RECT 86.245 104.085 86.500 104.585 ;
        RECT 85.750 103.915 86.500 104.085 ;
        RECT 86.985 103.915 87.155 104.755 ;
        RECT 85.750 102.925 85.980 103.915 ;
        RECT 87.365 103.745 87.615 104.585 ;
        RECT 87.825 103.915 87.995 104.755 ;
        RECT 88.165 103.745 88.455 104.585 ;
        RECT 86.150 103.095 86.500 103.745 ;
        RECT 86.730 103.575 88.455 103.745 ;
        RECT 88.665 103.695 88.835 104.755 ;
        RECT 89.130 104.375 89.460 104.755 ;
        RECT 89.640 104.205 89.810 104.495 ;
        RECT 89.980 104.295 90.230 104.755 ;
        RECT 89.010 104.035 89.810 104.205 ;
        RECT 90.400 104.245 91.270 104.585 ;
        RECT 86.730 103.025 87.140 103.575 ;
        RECT 89.010 103.415 89.180 104.035 ;
        RECT 90.400 103.865 90.570 104.245 ;
        RECT 91.505 104.125 91.675 104.585 ;
        RECT 91.845 104.295 92.215 104.755 ;
        RECT 92.510 104.155 92.680 104.495 ;
        RECT 92.850 104.325 93.180 104.755 ;
        RECT 93.415 104.155 93.585 104.495 ;
        RECT 89.350 103.695 90.570 103.865 ;
        RECT 90.740 103.785 91.200 104.075 ;
        RECT 91.505 103.955 92.065 104.125 ;
        RECT 92.510 103.985 93.585 104.155 ;
        RECT 93.755 104.255 94.435 104.585 ;
        RECT 94.650 104.255 94.900 104.585 ;
        RECT 95.070 104.295 95.320 104.755 ;
        RECT 91.895 103.815 92.065 103.955 ;
        RECT 90.740 103.775 91.705 103.785 ;
        RECT 90.400 103.605 90.570 103.695 ;
        RECT 91.030 103.615 91.705 103.775 ;
        RECT 89.010 103.405 89.355 103.415 ;
        RECT 87.325 103.195 89.355 103.405 ;
        RECT 85.750 102.755 86.500 102.925 ;
        RECT 86.730 102.855 88.495 103.025 ;
        RECT 85.745 102.205 86.075 102.585 ;
        RECT 86.245 102.465 86.500 102.755 ;
        RECT 86.985 102.205 87.155 102.675 ;
        RECT 87.325 102.375 87.655 102.855 ;
        RECT 87.825 102.205 87.995 102.675 ;
        RECT 88.165 102.375 88.495 102.855 ;
        RECT 88.665 102.205 88.835 103.015 ;
        RECT 89.030 102.940 89.355 103.195 ;
        RECT 89.035 102.585 89.355 102.940 ;
        RECT 89.525 103.155 90.065 103.525 ;
        RECT 90.400 103.435 90.805 103.605 ;
        RECT 89.525 102.755 89.765 103.155 ;
        RECT 90.245 102.985 90.465 103.265 ;
        RECT 89.935 102.815 90.465 102.985 ;
        RECT 89.935 102.585 90.105 102.815 ;
        RECT 90.635 102.655 90.805 103.435 ;
        RECT 90.975 102.825 91.325 103.445 ;
        RECT 91.495 102.825 91.705 103.615 ;
        RECT 91.895 103.645 93.395 103.815 ;
        RECT 91.895 102.955 92.065 103.645 ;
        RECT 93.755 103.475 93.925 104.255 ;
        RECT 94.730 104.125 94.900 104.255 ;
        RECT 92.235 103.305 93.925 103.475 ;
        RECT 94.095 103.695 94.560 104.085 ;
        RECT 94.730 103.955 95.125 104.125 ;
        RECT 92.235 103.125 92.405 103.305 ;
        RECT 89.035 102.415 90.105 102.585 ;
        RECT 90.275 102.205 90.465 102.645 ;
        RECT 90.635 102.375 91.585 102.655 ;
        RECT 91.895 102.565 92.155 102.955 ;
        RECT 92.575 102.885 93.365 103.135 ;
        RECT 91.805 102.395 92.155 102.565 ;
        RECT 92.365 102.205 92.695 102.665 ;
        RECT 93.570 102.595 93.740 103.305 ;
        RECT 94.095 103.105 94.265 103.695 ;
        RECT 93.910 102.885 94.265 103.105 ;
        RECT 94.435 102.885 94.785 103.505 ;
        RECT 94.955 102.595 95.125 103.955 ;
        RECT 95.490 103.785 95.815 104.570 ;
        RECT 95.295 102.735 95.755 103.785 ;
        RECT 93.570 102.425 94.425 102.595 ;
        RECT 94.630 102.425 95.125 102.595 ;
        RECT 95.295 102.205 95.625 102.565 ;
        RECT 95.985 102.465 96.155 104.585 ;
        RECT 96.325 104.255 96.655 104.755 ;
        RECT 96.825 104.085 97.080 104.585 ;
        RECT 96.330 103.915 97.080 104.085 ;
        RECT 96.330 102.925 96.560 103.915 ;
        RECT 96.730 103.095 97.080 103.745 ;
        RECT 97.715 103.665 101.225 104.755 ;
        RECT 97.715 103.145 99.405 103.665 ;
        RECT 101.395 103.590 101.685 104.755 ;
        RECT 102.165 103.915 102.335 104.755 ;
        RECT 102.545 103.745 102.795 104.585 ;
        RECT 103.005 103.915 103.175 104.755 ;
        RECT 103.345 103.745 103.635 104.585 ;
        RECT 101.910 103.575 103.635 103.745 ;
        RECT 103.845 103.695 104.015 104.755 ;
        RECT 104.310 104.375 104.640 104.755 ;
        RECT 104.820 104.205 104.990 104.495 ;
        RECT 105.160 104.295 105.410 104.755 ;
        RECT 104.190 104.035 104.990 104.205 ;
        RECT 105.580 104.245 106.450 104.585 ;
        RECT 99.575 102.975 101.225 103.495 ;
        RECT 96.330 102.755 97.080 102.925 ;
        RECT 96.325 102.205 96.655 102.585 ;
        RECT 96.825 102.465 97.080 102.755 ;
        RECT 97.715 102.205 101.225 102.975 ;
        RECT 101.910 103.025 102.320 103.575 ;
        RECT 104.190 103.415 104.360 104.035 ;
        RECT 105.580 103.865 105.750 104.245 ;
        RECT 106.685 104.125 106.855 104.585 ;
        RECT 107.025 104.295 107.395 104.755 ;
        RECT 107.690 104.155 107.860 104.495 ;
        RECT 108.030 104.325 108.360 104.755 ;
        RECT 108.595 104.155 108.765 104.495 ;
        RECT 104.530 103.695 105.750 103.865 ;
        RECT 105.920 103.785 106.380 104.075 ;
        RECT 106.685 103.955 107.245 104.125 ;
        RECT 107.690 103.985 108.765 104.155 ;
        RECT 108.935 104.255 109.615 104.585 ;
        RECT 109.830 104.255 110.080 104.585 ;
        RECT 110.250 104.295 110.500 104.755 ;
        RECT 107.075 103.815 107.245 103.955 ;
        RECT 105.920 103.775 106.885 103.785 ;
        RECT 105.580 103.605 105.750 103.695 ;
        RECT 106.210 103.615 106.885 103.775 ;
        RECT 104.190 103.405 104.535 103.415 ;
        RECT 102.505 103.195 104.535 103.405 ;
        RECT 101.395 102.205 101.685 102.930 ;
        RECT 101.910 102.855 103.675 103.025 ;
        RECT 102.165 102.205 102.335 102.675 ;
        RECT 102.505 102.375 102.835 102.855 ;
        RECT 103.005 102.205 103.175 102.675 ;
        RECT 103.345 102.375 103.675 102.855 ;
        RECT 103.845 102.205 104.015 103.015 ;
        RECT 104.210 102.940 104.535 103.195 ;
        RECT 104.215 102.585 104.535 102.940 ;
        RECT 104.705 103.155 105.245 103.525 ;
        RECT 105.580 103.435 105.985 103.605 ;
        RECT 104.705 102.755 104.945 103.155 ;
        RECT 105.425 102.985 105.645 103.265 ;
        RECT 105.115 102.815 105.645 102.985 ;
        RECT 105.115 102.585 105.285 102.815 ;
        RECT 105.815 102.655 105.985 103.435 ;
        RECT 106.155 102.825 106.505 103.445 ;
        RECT 106.675 102.825 106.885 103.615 ;
        RECT 107.075 103.645 108.575 103.815 ;
        RECT 107.075 102.955 107.245 103.645 ;
        RECT 108.935 103.475 109.105 104.255 ;
        RECT 109.910 104.125 110.080 104.255 ;
        RECT 107.415 103.305 109.105 103.475 ;
        RECT 109.275 103.695 109.740 104.085 ;
        RECT 109.910 103.955 110.305 104.125 ;
        RECT 107.415 103.125 107.585 103.305 ;
        RECT 104.215 102.415 105.285 102.585 ;
        RECT 105.455 102.205 105.645 102.645 ;
        RECT 105.815 102.375 106.765 102.655 ;
        RECT 107.075 102.565 107.335 102.955 ;
        RECT 107.755 102.885 108.545 103.135 ;
        RECT 106.985 102.395 107.335 102.565 ;
        RECT 107.545 102.205 107.875 102.665 ;
        RECT 108.750 102.595 108.920 103.305 ;
        RECT 109.275 103.105 109.445 103.695 ;
        RECT 109.090 102.885 109.445 103.105 ;
        RECT 109.615 102.885 109.965 103.505 ;
        RECT 110.135 102.595 110.305 103.955 ;
        RECT 110.670 103.785 110.995 104.570 ;
        RECT 110.475 102.735 110.935 103.785 ;
        RECT 108.750 102.425 109.605 102.595 ;
        RECT 109.810 102.425 110.305 102.595 ;
        RECT 110.475 102.205 110.805 102.565 ;
        RECT 111.165 102.465 111.335 104.585 ;
        RECT 111.505 104.255 111.835 104.755 ;
        RECT 112.005 104.085 112.260 104.585 ;
        RECT 111.510 103.915 112.260 104.085 ;
        RECT 112.440 104.085 112.695 104.585 ;
        RECT 112.865 104.255 113.195 104.755 ;
        RECT 112.440 103.915 113.190 104.085 ;
        RECT 111.510 102.925 111.740 103.915 ;
        RECT 111.910 103.095 112.260 103.745 ;
        RECT 112.440 103.095 112.790 103.745 ;
        RECT 112.960 102.925 113.190 103.915 ;
        RECT 111.510 102.755 112.260 102.925 ;
        RECT 111.505 102.205 111.835 102.585 ;
        RECT 112.005 102.465 112.260 102.755 ;
        RECT 112.440 102.755 113.190 102.925 ;
        RECT 112.440 102.465 112.695 102.755 ;
        RECT 112.865 102.205 113.195 102.585 ;
        RECT 113.365 102.465 113.535 104.585 ;
        RECT 113.705 103.785 114.030 104.570 ;
        RECT 114.200 104.295 114.450 104.755 ;
        RECT 114.620 104.255 114.870 104.585 ;
        RECT 115.085 104.255 115.765 104.585 ;
        RECT 114.620 104.125 114.790 104.255 ;
        RECT 114.395 103.955 114.790 104.125 ;
        RECT 113.765 102.735 114.225 103.785 ;
        RECT 114.395 102.595 114.565 103.955 ;
        RECT 114.960 103.695 115.425 104.085 ;
        RECT 114.735 102.885 115.085 103.505 ;
        RECT 115.255 103.105 115.425 103.695 ;
        RECT 115.595 103.475 115.765 104.255 ;
        RECT 115.935 104.155 116.105 104.495 ;
        RECT 116.340 104.325 116.670 104.755 ;
        RECT 116.840 104.155 117.010 104.495 ;
        RECT 117.305 104.295 117.675 104.755 ;
        RECT 115.935 103.985 117.010 104.155 ;
        RECT 117.845 104.125 118.015 104.585 ;
        RECT 118.250 104.245 119.120 104.585 ;
        RECT 119.290 104.295 119.540 104.755 ;
        RECT 117.455 103.955 118.015 104.125 ;
        RECT 117.455 103.815 117.625 103.955 ;
        RECT 116.125 103.645 117.625 103.815 ;
        RECT 118.320 103.785 118.780 104.075 ;
        RECT 115.595 103.305 117.285 103.475 ;
        RECT 115.255 102.885 115.610 103.105 ;
        RECT 115.780 102.595 115.950 103.305 ;
        RECT 116.155 102.885 116.945 103.135 ;
        RECT 117.115 103.125 117.285 103.305 ;
        RECT 117.455 102.955 117.625 103.645 ;
        RECT 113.895 102.205 114.225 102.565 ;
        RECT 114.395 102.425 114.890 102.595 ;
        RECT 115.095 102.425 115.950 102.595 ;
        RECT 116.825 102.205 117.155 102.665 ;
        RECT 117.365 102.565 117.625 102.955 ;
        RECT 117.815 103.775 118.780 103.785 ;
        RECT 118.950 103.865 119.120 104.245 ;
        RECT 119.710 104.205 119.880 104.495 ;
        RECT 120.060 104.375 120.390 104.755 ;
        RECT 119.710 104.035 120.510 104.205 ;
        RECT 117.815 103.615 118.490 103.775 ;
        RECT 118.950 103.695 120.170 103.865 ;
        RECT 117.815 102.825 118.025 103.615 ;
        RECT 118.950 103.605 119.120 103.695 ;
        RECT 118.195 102.825 118.545 103.445 ;
        RECT 118.715 103.435 119.120 103.605 ;
        RECT 118.715 102.655 118.885 103.435 ;
        RECT 119.055 102.985 119.275 103.265 ;
        RECT 119.455 103.155 119.995 103.525 ;
        RECT 120.340 103.415 120.510 104.035 ;
        RECT 120.685 103.695 120.855 104.755 ;
        RECT 121.065 103.745 121.355 104.585 ;
        RECT 121.525 103.915 121.695 104.755 ;
        RECT 121.905 103.745 122.155 104.585 ;
        RECT 122.365 103.915 122.535 104.755 ;
        RECT 121.065 103.575 122.790 103.745 ;
        RECT 119.055 102.815 119.585 102.985 ;
        RECT 117.365 102.395 117.715 102.565 ;
        RECT 117.935 102.375 118.885 102.655 ;
        RECT 119.055 102.205 119.245 102.645 ;
        RECT 119.415 102.585 119.585 102.815 ;
        RECT 119.755 102.755 119.995 103.155 ;
        RECT 120.165 103.405 120.510 103.415 ;
        RECT 120.165 103.195 122.195 103.405 ;
        RECT 120.165 102.940 120.490 103.195 ;
        RECT 122.380 103.025 122.790 103.575 ;
        RECT 123.015 103.665 124.685 104.755 ;
        RECT 124.855 103.680 125.125 104.585 ;
        RECT 125.295 103.995 125.625 104.755 ;
        RECT 125.805 103.825 125.985 104.585 ;
        RECT 123.015 103.145 123.765 103.665 ;
        RECT 120.165 102.585 120.485 102.940 ;
        RECT 119.415 102.415 120.485 102.585 ;
        RECT 120.685 102.205 120.855 103.015 ;
        RECT 121.025 102.855 122.790 103.025 ;
        RECT 123.935 102.975 124.685 103.495 ;
        RECT 121.025 102.375 121.355 102.855 ;
        RECT 121.525 102.205 121.695 102.675 ;
        RECT 121.865 102.375 122.195 102.855 ;
        RECT 122.365 102.205 122.535 102.675 ;
        RECT 123.015 102.205 124.685 102.975 ;
        RECT 124.855 102.880 125.035 103.680 ;
        RECT 125.310 103.655 125.985 103.825 ;
        RECT 126.235 103.665 127.445 104.755 ;
        RECT 125.310 103.510 125.480 103.655 ;
        RECT 125.205 103.180 125.480 103.510 ;
        RECT 125.310 102.925 125.480 103.180 ;
        RECT 125.705 103.105 126.045 103.475 ;
        RECT 126.235 103.125 126.755 103.665 ;
        RECT 126.925 102.955 127.445 103.495 ;
        RECT 124.855 102.375 125.115 102.880 ;
        RECT 125.310 102.755 125.975 102.925 ;
        RECT 125.295 102.205 125.625 102.585 ;
        RECT 125.805 102.375 125.975 102.755 ;
        RECT 126.235 102.205 127.445 102.955 ;
        RECT 14.370 102.035 127.530 102.205 ;
        RECT 14.455 101.285 15.665 102.035 ;
        RECT 14.455 100.745 14.975 101.285 ;
        RECT 15.835 101.265 18.425 102.035 ;
        RECT 18.600 101.490 23.945 102.035 ;
        RECT 15.145 100.575 15.665 101.115 ;
        RECT 14.455 99.485 15.665 100.575 ;
        RECT 15.835 100.575 17.045 101.095 ;
        RECT 17.215 100.745 18.425 101.265 ;
        RECT 15.835 99.485 18.425 100.575 ;
        RECT 20.190 99.920 20.540 101.170 ;
        RECT 22.020 100.660 22.360 101.490 ;
        RECT 24.115 101.310 24.405 102.035 ;
        RECT 24.885 101.565 25.055 102.035 ;
        RECT 25.225 101.385 25.555 101.865 ;
        RECT 25.725 101.565 25.895 102.035 ;
        RECT 26.065 101.385 26.395 101.865 ;
        RECT 24.630 101.215 26.395 101.385 ;
        RECT 26.565 101.225 26.735 102.035 ;
        RECT 26.935 101.655 28.005 101.825 ;
        RECT 26.935 101.300 27.255 101.655 ;
        RECT 24.630 100.665 25.040 101.215 ;
        RECT 26.930 101.045 27.255 101.300 ;
        RECT 25.225 100.835 27.255 101.045 ;
        RECT 26.910 100.825 27.255 100.835 ;
        RECT 27.425 101.085 27.665 101.485 ;
        RECT 27.835 101.425 28.005 101.655 ;
        RECT 28.175 101.595 28.365 102.035 ;
        RECT 28.535 101.585 29.485 101.865 ;
        RECT 29.705 101.675 30.055 101.845 ;
        RECT 27.835 101.255 28.365 101.425 ;
        RECT 18.600 99.485 23.945 99.920 ;
        RECT 24.115 99.485 24.405 100.650 ;
        RECT 24.630 100.495 26.355 100.665 ;
        RECT 24.885 99.485 25.055 100.325 ;
        RECT 25.265 99.655 25.515 100.495 ;
        RECT 25.725 99.485 25.895 100.325 ;
        RECT 26.065 99.655 26.355 100.495 ;
        RECT 26.565 99.485 26.735 100.545 ;
        RECT 26.910 100.205 27.080 100.825 ;
        RECT 27.425 100.715 27.965 101.085 ;
        RECT 28.145 100.975 28.365 101.255 ;
        RECT 28.535 100.805 28.705 101.585 ;
        RECT 28.300 100.635 28.705 100.805 ;
        RECT 28.875 100.795 29.225 101.415 ;
        RECT 28.300 100.545 28.470 100.635 ;
        RECT 29.395 100.625 29.605 101.415 ;
        RECT 27.250 100.375 28.470 100.545 ;
        RECT 28.930 100.465 29.605 100.625 ;
        RECT 26.910 100.035 27.710 100.205 ;
        RECT 27.030 99.485 27.360 99.865 ;
        RECT 27.540 99.745 27.710 100.035 ;
        RECT 28.300 99.995 28.470 100.375 ;
        RECT 28.640 100.455 29.605 100.465 ;
        RECT 29.795 101.285 30.055 101.675 ;
        RECT 30.265 101.575 30.595 102.035 ;
        RECT 31.470 101.645 32.325 101.815 ;
        RECT 32.530 101.645 33.025 101.815 ;
        RECT 33.195 101.675 33.525 102.035 ;
        RECT 29.795 100.595 29.965 101.285 ;
        RECT 30.135 100.935 30.305 101.115 ;
        RECT 30.475 101.105 31.265 101.355 ;
        RECT 31.470 100.935 31.640 101.645 ;
        RECT 31.810 101.135 32.165 101.355 ;
        RECT 30.135 100.765 31.825 100.935 ;
        RECT 28.640 100.165 29.100 100.455 ;
        RECT 29.795 100.425 31.295 100.595 ;
        RECT 29.795 100.285 29.965 100.425 ;
        RECT 29.405 100.115 29.965 100.285 ;
        RECT 27.880 99.485 28.130 99.945 ;
        RECT 28.300 99.655 29.170 99.995 ;
        RECT 29.405 99.655 29.575 100.115 ;
        RECT 30.410 100.085 31.485 100.255 ;
        RECT 29.745 99.485 30.115 99.945 ;
        RECT 30.410 99.745 30.580 100.085 ;
        RECT 30.750 99.485 31.080 99.915 ;
        RECT 31.315 99.745 31.485 100.085 ;
        RECT 31.655 99.985 31.825 100.765 ;
        RECT 31.995 100.545 32.165 101.135 ;
        RECT 32.335 100.735 32.685 101.355 ;
        RECT 31.995 100.155 32.460 100.545 ;
        RECT 32.855 100.285 33.025 101.645 ;
        RECT 33.195 100.455 33.655 101.505 ;
        RECT 32.630 100.115 33.025 100.285 ;
        RECT 32.630 99.985 32.800 100.115 ;
        RECT 31.655 99.655 32.335 99.985 ;
        RECT 32.550 99.655 32.800 99.985 ;
        RECT 32.970 99.485 33.220 99.945 ;
        RECT 33.390 99.670 33.715 100.455 ;
        RECT 33.885 99.655 34.055 101.775 ;
        RECT 34.225 101.655 34.555 102.035 ;
        RECT 34.725 101.485 34.980 101.775 ;
        RECT 34.230 101.315 34.980 101.485 ;
        RECT 34.230 100.325 34.460 101.315 ;
        RECT 35.155 101.265 36.825 102.035 ;
        RECT 36.995 101.310 37.285 102.035 ;
        RECT 37.455 101.285 38.665 102.035 ;
        RECT 38.840 101.490 44.185 102.035 ;
        RECT 44.360 101.490 49.705 102.035 ;
        RECT 34.630 100.495 34.980 101.145 ;
        RECT 35.155 100.575 35.905 101.095 ;
        RECT 36.075 100.745 36.825 101.265 ;
        RECT 34.230 100.155 34.980 100.325 ;
        RECT 34.225 99.485 34.555 99.985 ;
        RECT 34.725 99.655 34.980 100.155 ;
        RECT 35.155 99.485 36.825 100.575 ;
        RECT 36.995 99.485 37.285 100.650 ;
        RECT 37.455 100.575 37.975 101.115 ;
        RECT 38.145 100.745 38.665 101.285 ;
        RECT 37.455 99.485 38.665 100.575 ;
        RECT 40.430 99.920 40.780 101.170 ;
        RECT 42.260 100.660 42.600 101.490 ;
        RECT 45.950 99.920 46.300 101.170 ;
        RECT 47.780 100.660 48.120 101.490 ;
        RECT 49.875 101.310 50.165 102.035 ;
        RECT 50.335 101.285 51.545 102.035 ;
        RECT 51.720 101.490 57.065 102.035 ;
        RECT 57.240 101.490 62.585 102.035 ;
        RECT 38.840 99.485 44.185 99.920 ;
        RECT 44.360 99.485 49.705 99.920 ;
        RECT 49.875 99.485 50.165 100.650 ;
        RECT 50.335 100.575 50.855 101.115 ;
        RECT 51.025 100.745 51.545 101.285 ;
        RECT 50.335 99.485 51.545 100.575 ;
        RECT 53.310 99.920 53.660 101.170 ;
        RECT 55.140 100.660 55.480 101.490 ;
        RECT 58.830 99.920 59.180 101.170 ;
        RECT 60.660 100.660 61.000 101.490 ;
        RECT 62.755 101.310 63.045 102.035 ;
        RECT 63.215 101.285 64.425 102.035 ;
        RECT 64.600 101.490 69.945 102.035 ;
        RECT 70.120 101.490 75.465 102.035 ;
        RECT 51.720 99.485 57.065 99.920 ;
        RECT 57.240 99.485 62.585 99.920 ;
        RECT 62.755 99.485 63.045 100.650 ;
        RECT 63.215 100.575 63.735 101.115 ;
        RECT 63.905 100.745 64.425 101.285 ;
        RECT 63.215 99.485 64.425 100.575 ;
        RECT 66.190 99.920 66.540 101.170 ;
        RECT 68.020 100.660 68.360 101.490 ;
        RECT 71.710 99.920 72.060 101.170 ;
        RECT 73.540 100.660 73.880 101.490 ;
        RECT 75.635 101.310 75.925 102.035 ;
        RECT 76.095 101.285 77.305 102.035 ;
        RECT 77.480 101.490 82.825 102.035 ;
        RECT 83.000 101.490 88.345 102.035 ;
        RECT 64.600 99.485 69.945 99.920 ;
        RECT 70.120 99.485 75.465 99.920 ;
        RECT 75.635 99.485 75.925 100.650 ;
        RECT 76.095 100.575 76.615 101.115 ;
        RECT 76.785 100.745 77.305 101.285 ;
        RECT 76.095 99.485 77.305 100.575 ;
        RECT 79.070 99.920 79.420 101.170 ;
        RECT 80.900 100.660 81.240 101.490 ;
        RECT 84.590 99.920 84.940 101.170 ;
        RECT 86.420 100.660 86.760 101.490 ;
        RECT 88.515 101.310 88.805 102.035 ;
        RECT 88.975 101.265 90.645 102.035 ;
        RECT 91.125 101.565 91.295 102.035 ;
        RECT 91.465 101.385 91.795 101.865 ;
        RECT 91.965 101.565 92.135 102.035 ;
        RECT 92.305 101.385 92.635 101.865 ;
        RECT 77.480 99.485 82.825 99.920 ;
        RECT 83.000 99.485 88.345 99.920 ;
        RECT 88.515 99.485 88.805 100.650 ;
        RECT 88.975 100.575 89.725 101.095 ;
        RECT 89.895 100.745 90.645 101.265 ;
        RECT 90.870 101.215 92.635 101.385 ;
        RECT 92.805 101.225 92.975 102.035 ;
        RECT 93.175 101.655 94.245 101.825 ;
        RECT 93.175 101.300 93.495 101.655 ;
        RECT 90.870 100.665 91.280 101.215 ;
        RECT 93.170 101.045 93.495 101.300 ;
        RECT 91.465 100.835 93.495 101.045 ;
        RECT 93.150 100.825 93.495 100.835 ;
        RECT 93.665 101.085 93.905 101.485 ;
        RECT 94.075 101.425 94.245 101.655 ;
        RECT 94.415 101.595 94.605 102.035 ;
        RECT 94.775 101.585 95.725 101.865 ;
        RECT 95.945 101.675 96.295 101.845 ;
        RECT 94.075 101.255 94.605 101.425 ;
        RECT 88.975 99.485 90.645 100.575 ;
        RECT 90.870 100.495 92.595 100.665 ;
        RECT 91.125 99.485 91.295 100.325 ;
        RECT 91.505 99.655 91.755 100.495 ;
        RECT 91.965 99.485 92.135 100.325 ;
        RECT 92.305 99.655 92.595 100.495 ;
        RECT 92.805 99.485 92.975 100.545 ;
        RECT 93.150 100.205 93.320 100.825 ;
        RECT 93.665 100.715 94.205 101.085 ;
        RECT 94.385 100.975 94.605 101.255 ;
        RECT 94.775 100.805 94.945 101.585 ;
        RECT 94.540 100.635 94.945 100.805 ;
        RECT 95.115 100.795 95.465 101.415 ;
        RECT 94.540 100.545 94.710 100.635 ;
        RECT 95.635 100.625 95.845 101.415 ;
        RECT 93.490 100.375 94.710 100.545 ;
        RECT 95.170 100.465 95.845 100.625 ;
        RECT 93.150 100.035 93.950 100.205 ;
        RECT 93.270 99.485 93.600 99.865 ;
        RECT 93.780 99.745 93.950 100.035 ;
        RECT 94.540 99.995 94.710 100.375 ;
        RECT 94.880 100.455 95.845 100.465 ;
        RECT 96.035 101.285 96.295 101.675 ;
        RECT 96.505 101.575 96.835 102.035 ;
        RECT 97.710 101.645 98.565 101.815 ;
        RECT 98.770 101.645 99.265 101.815 ;
        RECT 99.435 101.675 99.765 102.035 ;
        RECT 96.035 100.595 96.205 101.285 ;
        RECT 96.375 100.935 96.545 101.115 ;
        RECT 96.715 101.105 97.505 101.355 ;
        RECT 97.710 100.935 97.880 101.645 ;
        RECT 98.050 101.135 98.405 101.355 ;
        RECT 96.375 100.765 98.065 100.935 ;
        RECT 94.880 100.165 95.340 100.455 ;
        RECT 96.035 100.425 97.535 100.595 ;
        RECT 96.035 100.285 96.205 100.425 ;
        RECT 95.645 100.115 96.205 100.285 ;
        RECT 94.120 99.485 94.370 99.945 ;
        RECT 94.540 99.655 95.410 99.995 ;
        RECT 95.645 99.655 95.815 100.115 ;
        RECT 96.650 100.085 97.725 100.255 ;
        RECT 95.985 99.485 96.355 99.945 ;
        RECT 96.650 99.745 96.820 100.085 ;
        RECT 96.990 99.485 97.320 99.915 ;
        RECT 97.555 99.745 97.725 100.085 ;
        RECT 97.895 99.985 98.065 100.765 ;
        RECT 98.235 100.545 98.405 101.135 ;
        RECT 98.575 100.735 98.925 101.355 ;
        RECT 98.235 100.155 98.700 100.545 ;
        RECT 99.095 100.285 99.265 101.645 ;
        RECT 99.435 100.455 99.895 101.505 ;
        RECT 98.870 100.115 99.265 100.285 ;
        RECT 98.870 99.985 99.040 100.115 ;
        RECT 97.895 99.655 98.575 99.985 ;
        RECT 98.790 99.655 99.040 99.985 ;
        RECT 99.210 99.485 99.460 99.945 ;
        RECT 99.630 99.670 99.955 100.455 ;
        RECT 100.125 99.655 100.295 101.775 ;
        RECT 100.465 101.655 100.795 102.035 ;
        RECT 100.965 101.485 101.220 101.775 ;
        RECT 100.470 101.315 101.220 101.485 ;
        RECT 100.470 100.325 100.700 101.315 ;
        RECT 101.395 101.310 101.685 102.035 ;
        RECT 101.855 101.285 103.065 102.035 ;
        RECT 103.240 101.490 108.585 102.035 ;
        RECT 108.760 101.490 114.105 102.035 ;
        RECT 100.870 100.495 101.220 101.145 ;
        RECT 100.470 100.155 101.220 100.325 ;
        RECT 100.465 99.485 100.795 99.985 ;
        RECT 100.965 99.655 101.220 100.155 ;
        RECT 101.395 99.485 101.685 100.650 ;
        RECT 101.855 100.575 102.375 101.115 ;
        RECT 102.545 100.745 103.065 101.285 ;
        RECT 101.855 99.485 103.065 100.575 ;
        RECT 104.830 99.920 105.180 101.170 ;
        RECT 106.660 100.660 107.000 101.490 ;
        RECT 110.350 99.920 110.700 101.170 ;
        RECT 112.180 100.660 112.520 101.490 ;
        RECT 114.275 101.310 114.565 102.035 ;
        RECT 115.655 101.265 119.165 102.035 ;
        RECT 103.240 99.485 108.585 99.920 ;
        RECT 108.760 99.485 114.105 99.920 ;
        RECT 114.275 99.485 114.565 100.650 ;
        RECT 115.655 100.575 117.345 101.095 ;
        RECT 117.515 100.745 119.165 101.265 ;
        RECT 119.375 101.215 119.605 102.035 ;
        RECT 119.775 101.235 120.105 101.865 ;
        RECT 119.355 100.795 119.685 101.045 ;
        RECT 119.855 100.635 120.105 101.235 ;
        RECT 120.275 101.215 120.485 102.035 ;
        RECT 120.720 101.490 126.065 102.035 ;
        RECT 115.655 99.485 119.165 100.575 ;
        RECT 119.375 99.485 119.605 100.625 ;
        RECT 119.775 99.655 120.105 100.635 ;
        RECT 120.275 99.485 120.485 100.625 ;
        RECT 122.310 99.920 122.660 101.170 ;
        RECT 124.140 100.660 124.480 101.490 ;
        RECT 126.235 101.285 127.445 102.035 ;
        RECT 126.235 100.575 126.755 101.115 ;
        RECT 126.925 100.745 127.445 101.285 ;
        RECT 120.720 99.485 126.065 99.920 ;
        RECT 126.235 99.485 127.445 100.575 ;
        RECT 14.370 99.315 127.530 99.485 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 14.370 210.680 127.530 211.160 ;
        RECT 14.370 207.960 127.530 208.440 ;
        RECT 73.320 207.420 73.640 207.480 ;
        RECT 74.715 207.420 75.005 207.465 ;
        RECT 73.320 207.280 79.070 207.420 ;
        RECT 73.320 207.220 73.640 207.280 ;
        RECT 74.715 207.235 75.005 207.280 ;
        RECT 65.960 206.740 66.280 206.800 ;
        RECT 72.415 206.740 72.705 206.785 ;
        RECT 65.960 206.600 72.705 206.740 ;
        RECT 65.960 206.540 66.280 206.600 ;
        RECT 72.415 206.555 72.705 206.600 ;
        RECT 72.860 206.740 73.180 206.800 ;
        RECT 78.930 206.785 79.070 207.280 ;
        RECT 79.300 206.880 79.620 207.140 ;
        RECT 73.795 206.740 74.085 206.785 ;
        RECT 72.860 206.600 74.085 206.740 ;
        RECT 72.860 206.540 73.180 206.600 ;
        RECT 73.795 206.555 74.085 206.600 ;
        RECT 78.855 206.555 79.145 206.785 ;
        RECT 72.875 206.060 73.165 206.105 ;
        RECT 73.780 206.060 74.100 206.120 ;
        RECT 72.875 205.920 74.100 206.060 ;
        RECT 72.875 205.875 73.165 205.920 ;
        RECT 73.780 205.860 74.100 205.920 ;
        RECT 75.620 206.060 75.940 206.120 ;
        RECT 77.015 206.060 77.305 206.105 ;
        RECT 75.620 205.920 77.305 206.060 ;
        RECT 75.620 205.860 75.940 205.920 ;
        RECT 77.015 205.875 77.305 205.920 ;
        RECT 14.370 205.240 127.530 205.720 ;
        RECT 73.780 205.040 74.100 205.100 ;
        RECT 73.780 204.900 76.310 205.040 ;
        RECT 73.780 204.840 74.100 204.900 ;
        RECT 67.355 204.700 67.645 204.745 ;
        RECT 69.755 204.700 70.045 204.745 ;
        RECT 72.995 204.700 73.645 204.745 ;
        RECT 67.355 204.560 73.645 204.700 ;
        RECT 67.355 204.515 67.645 204.560 ;
        RECT 69.755 204.515 70.345 204.560 ;
        RECT 72.995 204.515 73.645 204.560 ;
        RECT 65.515 204.360 65.805 204.405 ;
        RECT 65.960 204.360 66.280 204.420 ;
        RECT 66.895 204.360 67.185 204.405 ;
        RECT 65.515 204.220 67.185 204.360 ;
        RECT 65.515 204.175 65.805 204.220 ;
        RECT 65.960 204.160 66.280 204.220 ;
        RECT 66.895 204.175 67.185 204.220 ;
        RECT 70.055 204.200 70.345 204.515 ;
        RECT 75.620 204.500 75.940 204.760 ;
        RECT 76.170 204.700 76.310 204.900 ;
        RECT 78.955 204.700 79.245 204.745 ;
        RECT 82.195 204.700 82.845 204.745 ;
        RECT 76.170 204.560 82.845 204.700 ;
        RECT 78.955 204.515 79.545 204.560 ;
        RECT 82.195 204.515 82.845 204.560 ;
        RECT 83.440 204.700 83.760 204.760 ;
        RECT 84.835 204.700 85.125 204.745 ;
        RECT 83.440 204.560 85.125 204.700 ;
        RECT 71.135 204.360 71.425 204.405 ;
        RECT 74.715 204.360 75.005 204.405 ;
        RECT 76.550 204.360 76.840 204.405 ;
        RECT 71.135 204.220 76.840 204.360 ;
        RECT 71.135 204.175 71.425 204.220 ;
        RECT 74.715 204.175 75.005 204.220 ;
        RECT 76.550 204.175 76.840 204.220 ;
        RECT 79.255 204.200 79.545 204.515 ;
        RECT 83.440 204.500 83.760 204.560 ;
        RECT 84.835 204.515 85.125 204.560 ;
        RECT 80.335 204.360 80.625 204.405 ;
        RECT 83.915 204.360 84.205 204.405 ;
        RECT 85.750 204.360 86.040 204.405 ;
        RECT 80.335 204.220 86.040 204.360 ;
        RECT 80.335 204.175 80.625 204.220 ;
        RECT 83.915 204.175 84.205 204.220 ;
        RECT 85.750 204.175 86.040 204.220 ;
        RECT 63.660 204.020 63.980 204.080 ;
        RECT 77.015 204.020 77.305 204.065 ;
        RECT 63.660 203.880 77.305 204.020 ;
        RECT 63.660 203.820 63.980 203.880 ;
        RECT 77.015 203.835 77.305 203.880 ;
        RECT 86.215 204.020 86.505 204.065 ;
        RECT 88.040 204.020 88.360 204.080 ;
        RECT 86.215 203.880 88.360 204.020 ;
        RECT 86.215 203.835 86.505 203.880 ;
        RECT 88.040 203.820 88.360 203.880 ;
        RECT 71.135 203.680 71.425 203.725 ;
        RECT 74.255 203.680 74.545 203.725 ;
        RECT 76.145 203.680 76.435 203.725 ;
        RECT 71.135 203.540 76.435 203.680 ;
        RECT 71.135 203.495 71.425 203.540 ;
        RECT 74.255 203.495 74.545 203.540 ;
        RECT 76.145 203.495 76.435 203.540 ;
        RECT 80.335 203.680 80.625 203.725 ;
        RECT 83.455 203.680 83.745 203.725 ;
        RECT 85.345 203.680 85.635 203.725 ;
        RECT 80.335 203.540 85.635 203.680 ;
        RECT 80.335 203.495 80.625 203.540 ;
        RECT 83.455 203.495 83.745 203.540 ;
        RECT 85.345 203.495 85.635 203.540 ;
        RECT 64.580 203.340 64.900 203.400 ;
        RECT 65.055 203.340 65.345 203.385 ;
        RECT 64.580 203.200 65.345 203.340 ;
        RECT 64.580 203.140 64.900 203.200 ;
        RECT 65.055 203.155 65.345 203.200 ;
        RECT 68.275 203.340 68.565 203.385 ;
        RECT 72.860 203.340 73.180 203.400 ;
        RECT 68.275 203.200 73.180 203.340 ;
        RECT 68.275 203.155 68.565 203.200 ;
        RECT 72.860 203.140 73.180 203.200 ;
        RECT 73.780 203.340 74.100 203.400 ;
        RECT 77.475 203.340 77.765 203.385 ;
        RECT 73.780 203.200 77.765 203.340 ;
        RECT 73.780 203.140 74.100 203.200 ;
        RECT 77.475 203.155 77.765 203.200 ;
        RECT 14.370 202.520 127.530 203.000 ;
        RECT 63.660 202.320 63.980 202.380 ;
        RECT 60.070 202.180 63.980 202.320 ;
        RECT 59.535 201.640 59.825 201.685 ;
        RECT 60.070 201.640 60.210 202.180 ;
        RECT 63.660 202.120 63.980 202.180 ;
        RECT 66.420 202.320 66.740 202.380 ;
        RECT 70.115 202.320 70.405 202.365 ;
        RECT 66.420 202.180 70.405 202.320 ;
        RECT 66.420 202.120 66.740 202.180 ;
        RECT 70.115 202.135 70.405 202.180 ;
        RECT 77.475 202.135 77.765 202.365 ;
        RECT 60.405 201.980 60.695 202.025 ;
        RECT 62.295 201.980 62.585 202.025 ;
        RECT 65.415 201.980 65.705 202.025 ;
        RECT 76.080 201.980 76.400 202.040 ;
        RECT 77.550 201.980 77.690 202.135 ;
        RECT 60.405 201.840 65.705 201.980 ;
        RECT 60.405 201.795 60.695 201.840 ;
        RECT 62.295 201.795 62.585 201.840 ;
        RECT 65.415 201.795 65.705 201.840 ;
        RECT 69.730 201.840 73.550 201.980 ;
        RECT 59.535 201.500 60.210 201.640 ;
        RECT 59.535 201.455 59.825 201.500 ;
        RECT 60.900 201.440 61.220 201.700 ;
        RECT 69.730 201.685 69.870 201.840 ;
        RECT 69.655 201.455 69.945 201.685 ;
        RECT 71.955 201.640 72.245 201.685 ;
        RECT 72.860 201.640 73.180 201.700 ;
        RECT 73.410 201.685 73.550 201.840 ;
        RECT 76.080 201.840 77.690 201.980 ;
        RECT 82.175 201.980 82.465 202.025 ;
        RECT 85.295 201.980 85.585 202.025 ;
        RECT 87.185 201.980 87.475 202.025 ;
        RECT 82.175 201.840 87.475 201.980 ;
        RECT 76.080 201.780 76.400 201.840 ;
        RECT 82.175 201.795 82.465 201.840 ;
        RECT 85.295 201.795 85.585 201.840 ;
        RECT 87.185 201.795 87.475 201.840 ;
        RECT 71.955 201.500 73.180 201.640 ;
        RECT 71.955 201.455 72.245 201.500 ;
        RECT 72.860 201.440 73.180 201.500 ;
        RECT 73.335 201.640 73.625 201.685 ;
        RECT 74.240 201.640 74.560 201.700 ;
        RECT 73.335 201.500 74.560 201.640 ;
        RECT 73.335 201.455 73.625 201.500 ;
        RECT 74.240 201.440 74.560 201.500 ;
        RECT 78.840 201.640 79.160 201.700 ;
        RECT 79.315 201.640 79.605 201.685 ;
        RECT 78.840 201.500 79.605 201.640 ;
        RECT 78.840 201.440 79.160 201.500 ;
        RECT 79.315 201.455 79.605 201.500 ;
        RECT 84.360 201.640 84.680 201.700 ;
        RECT 86.675 201.640 86.965 201.685 ;
        RECT 84.360 201.500 86.965 201.640 ;
        RECT 84.360 201.440 84.680 201.500 ;
        RECT 86.675 201.455 86.965 201.500 ;
        RECT 60.000 201.300 60.290 201.345 ;
        RECT 61.835 201.300 62.125 201.345 ;
        RECT 65.415 201.300 65.705 201.345 ;
        RECT 60.000 201.160 65.705 201.300 ;
        RECT 60.000 201.115 60.290 201.160 ;
        RECT 61.835 201.115 62.125 201.160 ;
        RECT 65.415 201.115 65.705 201.160 ;
        RECT 63.195 200.960 63.845 201.005 ;
        RECT 64.580 200.960 64.900 201.020 ;
        RECT 66.495 201.005 66.785 201.320 ;
        RECT 70.910 201.300 71.200 201.345 ;
        RECT 73.780 201.300 74.100 201.360 ;
        RECT 70.910 201.160 74.100 201.300 ;
        RECT 70.910 201.115 71.200 201.160 ;
        RECT 73.780 201.100 74.100 201.160 ;
        RECT 66.495 200.960 67.085 201.005 ;
        RECT 63.195 200.820 67.085 200.960 ;
        RECT 63.195 200.775 63.845 200.820 ;
        RECT 64.580 200.760 64.900 200.820 ;
        RECT 66.795 200.775 67.085 200.820 ;
        RECT 74.700 200.760 75.020 201.020 ;
        RECT 75.160 200.960 75.480 201.020 ;
        RECT 77.315 200.960 77.605 201.005 ;
        RECT 75.160 200.820 77.605 200.960 ;
        RECT 75.160 200.760 75.480 200.820 ;
        RECT 77.315 200.775 77.605 200.820 ;
        RECT 78.395 200.960 78.685 201.005 ;
        RECT 79.300 200.960 79.620 201.020 ;
        RECT 81.095 201.005 81.385 201.320 ;
        RECT 82.175 201.300 82.465 201.345 ;
        RECT 85.755 201.300 86.045 201.345 ;
        RECT 87.590 201.300 87.880 201.345 ;
        RECT 82.175 201.160 87.880 201.300 ;
        RECT 82.175 201.115 82.465 201.160 ;
        RECT 85.755 201.115 86.045 201.160 ;
        RECT 87.590 201.115 87.880 201.160 ;
        RECT 88.040 201.300 88.360 201.360 ;
        RECT 96.320 201.300 96.640 201.360 ;
        RECT 88.040 201.160 96.640 201.300 ;
        RECT 88.040 201.100 88.360 201.160 ;
        RECT 96.320 201.100 96.640 201.160 ;
        RECT 78.395 200.820 79.620 200.960 ;
        RECT 78.395 200.775 78.685 200.820 ;
        RECT 79.300 200.760 79.620 200.820 ;
        RECT 80.795 200.960 81.385 201.005 ;
        RECT 84.035 200.960 84.685 201.005 ;
        RECT 85.280 200.960 85.600 201.020 ;
        RECT 80.795 200.820 85.600 200.960 ;
        RECT 80.795 200.775 81.085 200.820 ;
        RECT 84.035 200.775 84.685 200.820 ;
        RECT 85.280 200.760 85.600 200.820 ;
        RECT 71.480 200.420 71.800 200.680 ;
        RECT 72.400 200.620 72.720 200.680 ;
        RECT 74.255 200.620 74.545 200.665 ;
        RECT 72.400 200.480 74.545 200.620 ;
        RECT 72.400 200.420 72.720 200.480 ;
        RECT 74.255 200.435 74.545 200.480 ;
        RECT 75.620 200.620 75.940 200.680 ;
        RECT 76.555 200.620 76.845 200.665 ;
        RECT 75.620 200.480 76.845 200.620 ;
        RECT 75.620 200.420 75.940 200.480 ;
        RECT 76.555 200.435 76.845 200.480 ;
        RECT 14.370 199.800 127.530 200.280 ;
        RECT 60.900 199.600 61.220 199.660 ;
        RECT 67.355 199.600 67.645 199.645 ;
        RECT 71.955 199.600 72.245 199.645 ;
        RECT 73.780 199.600 74.100 199.660 ;
        RECT 60.900 199.460 67.645 199.600 ;
        RECT 60.900 199.400 61.220 199.460 ;
        RECT 67.355 199.415 67.645 199.460 ;
        RECT 70.880 199.460 74.100 199.600 ;
        RECT 69.655 199.260 69.945 199.305 ;
        RECT 70.880 199.260 71.020 199.460 ;
        RECT 71.955 199.415 72.245 199.460 ;
        RECT 73.780 199.400 74.100 199.460 ;
        RECT 74.700 199.600 75.020 199.660 ;
        RECT 75.175 199.600 75.465 199.645 ;
        RECT 74.700 199.460 75.465 199.600 ;
        RECT 74.700 199.400 75.020 199.460 ;
        RECT 75.175 199.415 75.465 199.460 ;
        RECT 76.080 199.600 76.400 199.660 ;
        RECT 78.855 199.600 79.145 199.645 ;
        RECT 76.080 199.460 79.145 199.600 ;
        RECT 76.080 199.400 76.400 199.460 ;
        RECT 78.855 199.415 79.145 199.460 ;
        RECT 79.300 199.600 79.620 199.660 ;
        RECT 81.155 199.600 81.445 199.645 ;
        RECT 79.300 199.460 81.445 199.600 ;
        RECT 79.300 199.400 79.620 199.460 ;
        RECT 81.155 199.415 81.445 199.460 ;
        RECT 83.440 199.400 83.760 199.660 ;
        RECT 84.360 199.400 84.680 199.660 ;
        RECT 85.280 199.600 85.600 199.660 ;
        RECT 85.755 199.600 86.045 199.645 ;
        RECT 85.280 199.460 86.045 199.600 ;
        RECT 85.280 199.400 85.600 199.460 ;
        RECT 85.755 199.415 86.045 199.460 ;
        RECT 69.655 199.120 71.020 199.260 ;
        RECT 69.655 199.075 69.945 199.120 ;
        RECT 74.240 199.060 74.560 199.320 ;
        RECT 80.680 199.260 81.000 199.320 ;
        RECT 97.700 199.260 98.020 199.320 ;
        RECT 98.275 199.260 98.565 199.305 ;
        RECT 101.515 199.260 102.165 199.305 ;
        RECT 80.680 199.120 84.130 199.260 ;
        RECT 80.680 199.060 81.000 199.120 ;
        RECT 68.260 198.720 68.580 198.980 ;
        RECT 71.480 198.920 71.800 198.980 ;
        RECT 78.395 198.920 78.685 198.965 ;
        RECT 78.840 198.920 79.160 198.980 ;
        RECT 71.480 198.780 79.160 198.920 ;
        RECT 71.480 198.720 71.800 198.780 ;
        RECT 78.395 198.735 78.685 198.780 ;
        RECT 78.840 198.720 79.160 198.780 ;
        RECT 79.760 198.920 80.080 198.980 ;
        RECT 82.150 198.965 82.290 199.120 ;
        RECT 83.990 198.965 84.130 199.120 ;
        RECT 97.700 199.120 102.165 199.260 ;
        RECT 97.700 199.060 98.020 199.120 ;
        RECT 98.275 199.075 98.865 199.120 ;
        RECT 101.515 199.075 102.165 199.120 ;
        RECT 81.155 198.920 81.445 198.965 ;
        RECT 79.760 198.780 81.445 198.920 ;
        RECT 79.760 198.720 80.080 198.780 ;
        RECT 81.155 198.735 81.445 198.780 ;
        RECT 82.075 198.735 82.365 198.965 ;
        RECT 82.535 198.735 82.825 198.965 ;
        RECT 83.915 198.735 84.205 198.965 ;
        RECT 86.215 198.920 86.505 198.965 ;
        RECT 86.660 198.920 86.980 198.980 ;
        RECT 86.215 198.780 86.980 198.920 ;
        RECT 86.215 198.735 86.505 198.780 ;
        RECT 75.620 198.580 75.940 198.640 ;
        RECT 82.610 198.580 82.750 198.735 ;
        RECT 86.660 198.720 86.980 198.780 ;
        RECT 98.575 198.760 98.865 199.075 ;
        RECT 99.655 198.920 99.945 198.965 ;
        RECT 103.235 198.920 103.525 198.965 ;
        RECT 105.070 198.920 105.360 198.965 ;
        RECT 99.655 198.780 105.360 198.920 ;
        RECT 99.655 198.735 99.945 198.780 ;
        RECT 103.235 198.735 103.525 198.780 ;
        RECT 105.070 198.735 105.360 198.780 ;
        RECT 75.620 198.440 82.750 198.580 ;
        RECT 75.620 198.380 75.940 198.440 ;
        RECT 104.140 198.380 104.460 198.640 ;
        RECT 105.520 198.380 105.840 198.640 ;
        RECT 68.735 198.240 69.025 198.285 ;
        RECT 72.860 198.240 73.180 198.300 ;
        RECT 68.735 198.100 73.180 198.240 ;
        RECT 68.735 198.055 69.025 198.100 ;
        RECT 72.860 198.040 73.180 198.100 ;
        RECT 73.320 198.240 73.640 198.300 ;
        RECT 74.255 198.240 74.545 198.285 ;
        RECT 73.320 198.100 74.545 198.240 ;
        RECT 73.320 198.040 73.640 198.100 ;
        RECT 74.255 198.055 74.545 198.100 ;
        RECT 99.655 198.240 99.945 198.285 ;
        RECT 102.775 198.240 103.065 198.285 ;
        RECT 104.665 198.240 104.955 198.285 ;
        RECT 99.655 198.100 104.955 198.240 ;
        RECT 99.655 198.055 99.945 198.100 ;
        RECT 102.775 198.055 103.065 198.100 ;
        RECT 104.665 198.055 104.955 198.100 ;
        RECT 64.580 197.900 64.900 197.960 ;
        RECT 70.575 197.900 70.865 197.945 ;
        RECT 64.580 197.760 70.865 197.900 ;
        RECT 64.580 197.700 64.900 197.760 ;
        RECT 70.575 197.715 70.865 197.760 ;
        RECT 72.400 197.900 72.720 197.960 ;
        RECT 80.680 197.900 81.000 197.960 ;
        RECT 72.400 197.760 81.000 197.900 ;
        RECT 72.400 197.700 72.720 197.760 ;
        RECT 80.680 197.700 81.000 197.760 ;
        RECT 96.795 197.900 97.085 197.945 ;
        RECT 98.160 197.900 98.480 197.960 ;
        RECT 96.795 197.760 98.480 197.900 ;
        RECT 96.795 197.715 97.085 197.760 ;
        RECT 98.160 197.700 98.480 197.760 ;
        RECT 14.370 197.080 127.530 197.560 ;
        RECT 68.260 196.880 68.580 196.940 ;
        RECT 68.735 196.880 69.025 196.925 ;
        RECT 68.260 196.740 69.025 196.880 ;
        RECT 68.260 196.680 68.580 196.740 ;
        RECT 68.735 196.695 69.025 196.740 ;
        RECT 69.640 196.680 69.960 196.940 ;
        RECT 73.320 196.880 73.640 196.940 ;
        RECT 72.030 196.740 73.640 196.880 ;
        RECT 50.320 196.200 50.640 196.260 ;
        RECT 54.015 196.200 54.305 196.245 ;
        RECT 50.320 196.060 54.305 196.200 ;
        RECT 50.320 196.000 50.640 196.060 ;
        RECT 54.015 196.015 54.305 196.060 ;
        RECT 70.100 196.200 70.420 196.260 ;
        RECT 72.030 196.245 72.170 196.740 ;
        RECT 73.320 196.680 73.640 196.740 ;
        RECT 79.760 196.540 80.080 196.600 ;
        RECT 73.410 196.400 80.080 196.540 ;
        RECT 71.955 196.200 72.245 196.245 ;
        RECT 70.100 196.060 72.245 196.200 ;
        RECT 70.100 196.000 70.420 196.060 ;
        RECT 71.955 196.015 72.245 196.060 ;
        RECT 72.400 196.000 72.720 196.260 ;
        RECT 72.860 196.200 73.180 196.260 ;
        RECT 73.410 196.200 73.550 196.400 ;
        RECT 79.760 196.340 80.080 196.400 ;
        RECT 89.390 196.540 89.680 196.585 ;
        RECT 92.170 196.540 92.460 196.585 ;
        RECT 94.030 196.540 94.320 196.585 ;
        RECT 89.390 196.400 94.320 196.540 ;
        RECT 89.390 196.355 89.680 196.400 ;
        RECT 92.170 196.355 92.460 196.400 ;
        RECT 94.030 196.355 94.320 196.400 ;
        RECT 112.995 196.540 113.285 196.585 ;
        RECT 116.115 196.540 116.405 196.585 ;
        RECT 118.005 196.540 118.295 196.585 ;
        RECT 112.995 196.400 118.295 196.540 ;
        RECT 112.995 196.355 113.285 196.400 ;
        RECT 116.115 196.355 116.405 196.400 ;
        RECT 118.005 196.355 118.295 196.400 ;
        RECT 72.860 196.060 73.550 196.200 ;
        RECT 92.655 196.200 92.945 196.245 ;
        RECT 93.560 196.200 93.880 196.260 ;
        RECT 92.655 196.060 93.880 196.200 ;
        RECT 72.860 196.000 73.180 196.060 ;
        RECT 92.655 196.015 92.945 196.060 ;
        RECT 93.560 196.000 93.880 196.060 ;
        RECT 48.940 195.860 49.260 195.920 ;
        RECT 53.555 195.860 53.845 195.905 ;
        RECT 48.940 195.720 53.845 195.860 ;
        RECT 48.940 195.660 49.260 195.720 ;
        RECT 53.555 195.675 53.845 195.720 ;
        RECT 68.720 195.860 69.040 195.920 ;
        RECT 73.335 195.860 73.625 195.905 ;
        RECT 74.240 195.860 74.560 195.920 ;
        RECT 68.720 195.720 74.560 195.860 ;
        RECT 68.720 195.660 69.040 195.720 ;
        RECT 73.335 195.675 73.625 195.720 ;
        RECT 74.240 195.660 74.560 195.720 ;
        RECT 89.390 195.860 89.680 195.905 ;
        RECT 94.495 195.860 94.785 195.905 ;
        RECT 96.320 195.860 96.640 195.920 ;
        RECT 89.390 195.720 91.925 195.860 ;
        RECT 89.390 195.675 89.680 195.720 ;
        RECT 70.575 195.520 70.865 195.565 ;
        RECT 71.480 195.520 71.800 195.580 ;
        RECT 75.160 195.520 75.480 195.580 ;
        RECT 70.575 195.380 75.480 195.520 ;
        RECT 70.575 195.335 70.865 195.380 ;
        RECT 71.480 195.320 71.800 195.380 ;
        RECT 75.160 195.320 75.480 195.380 ;
        RECT 87.530 195.520 87.820 195.565 ;
        RECT 89.880 195.520 90.200 195.580 ;
        RECT 91.710 195.565 91.925 195.720 ;
        RECT 94.495 195.720 96.640 195.860 ;
        RECT 94.495 195.675 94.785 195.720 ;
        RECT 96.320 195.660 96.640 195.720 ;
        RECT 98.160 195.660 98.480 195.920 ;
        RECT 111.915 195.565 112.205 195.880 ;
        RECT 112.995 195.860 113.285 195.905 ;
        RECT 116.575 195.860 116.865 195.905 ;
        RECT 118.410 195.860 118.700 195.905 ;
        RECT 112.995 195.720 118.700 195.860 ;
        RECT 112.995 195.675 113.285 195.720 ;
        RECT 116.575 195.675 116.865 195.720 ;
        RECT 118.410 195.675 118.700 195.720 ;
        RECT 118.875 195.675 119.165 195.905 ;
        RECT 115.180 195.565 115.500 195.580 ;
        RECT 90.790 195.520 91.080 195.565 ;
        RECT 87.530 195.380 91.080 195.520 ;
        RECT 87.530 195.335 87.820 195.380 ;
        RECT 89.880 195.320 90.200 195.380 ;
        RECT 90.790 195.335 91.080 195.380 ;
        RECT 91.710 195.520 92.000 195.565 ;
        RECT 93.570 195.520 93.860 195.565 ;
        RECT 91.710 195.380 93.860 195.520 ;
        RECT 91.710 195.335 92.000 195.380 ;
        RECT 93.570 195.335 93.860 195.380 ;
        RECT 111.615 195.520 112.205 195.565 ;
        RECT 114.855 195.520 115.505 195.565 ;
        RECT 111.615 195.380 115.505 195.520 ;
        RECT 111.615 195.335 111.905 195.380 ;
        RECT 114.855 195.335 115.505 195.380 ;
        RECT 115.180 195.320 115.500 195.335 ;
        RECT 117.480 195.320 117.800 195.580 ;
        RECT 117.940 195.520 118.260 195.580 ;
        RECT 118.950 195.520 119.090 195.675 ;
        RECT 117.940 195.380 119.090 195.520 ;
        RECT 117.940 195.320 118.260 195.380 ;
        RECT 53.080 194.980 53.400 195.240 ;
        RECT 57.235 195.180 57.525 195.225 ;
        RECT 57.680 195.180 58.000 195.240 ;
        RECT 85.280 195.225 85.600 195.240 ;
        RECT 57.235 195.040 58.000 195.180 ;
        RECT 57.235 194.995 57.525 195.040 ;
        RECT 57.680 194.980 58.000 195.040 ;
        RECT 69.575 195.180 69.865 195.225 ;
        RECT 71.035 195.180 71.325 195.225 ;
        RECT 69.575 195.040 71.325 195.180 ;
        RECT 69.575 194.995 69.865 195.040 ;
        RECT 71.035 194.995 71.325 195.040 ;
        RECT 85.280 194.995 85.815 195.225 ;
        RECT 85.280 194.980 85.600 194.995 ;
        RECT 100.920 194.980 101.240 195.240 ;
        RECT 108.740 195.180 109.060 195.240 ;
        RECT 110.135 195.180 110.425 195.225 ;
        RECT 108.740 195.040 110.425 195.180 ;
        RECT 108.740 194.980 109.060 195.040 ;
        RECT 110.135 194.995 110.425 195.040 ;
        RECT 14.370 194.360 127.530 194.840 ;
        RECT 50.320 194.160 50.640 194.220 ;
        RECT 57.695 194.160 57.985 194.205 ;
        RECT 50.320 194.020 57.985 194.160 ;
        RECT 50.320 193.960 50.640 194.020 ;
        RECT 57.695 193.975 57.985 194.020 ;
        RECT 71.480 193.960 71.800 194.220 ;
        RECT 85.280 194.160 85.600 194.220 ;
        RECT 85.755 194.160 86.045 194.205 ;
        RECT 72.030 194.020 85.050 194.160 ;
        RECT 48.940 193.820 49.260 193.880 ;
        RECT 53.080 193.865 53.400 193.880 ;
        RECT 48.570 193.680 49.260 193.820 ;
        RECT 45.720 193.480 46.040 193.540 ;
        RECT 48.570 193.525 48.710 193.680 ;
        RECT 48.940 193.620 49.260 193.680 ;
        RECT 52.615 193.820 53.400 193.865 ;
        RECT 56.215 193.820 56.505 193.865 ;
        RECT 72.030 193.820 72.170 194.020 ;
        RECT 52.615 193.680 56.505 193.820 ;
        RECT 52.615 193.635 53.400 193.680 ;
        RECT 53.080 193.620 53.400 193.635 ;
        RECT 55.915 193.635 56.505 193.680 ;
        RECT 66.050 193.680 72.170 193.820 ;
        RECT 72.400 193.820 72.720 193.880 ;
        RECT 84.910 193.820 85.050 194.020 ;
        RECT 85.280 194.020 86.045 194.160 ;
        RECT 85.280 193.960 85.600 194.020 ;
        RECT 85.755 193.975 86.045 194.020 ;
        RECT 89.435 194.160 89.725 194.205 ;
        RECT 89.880 194.160 90.200 194.220 ;
        RECT 89.435 194.020 90.200 194.160 ;
        RECT 89.435 193.975 89.725 194.020 ;
        RECT 89.880 193.960 90.200 194.020 ;
        RECT 93.575 194.160 93.865 194.205 ;
        RECT 97.700 194.160 98.020 194.220 ;
        RECT 93.575 194.020 98.020 194.160 ;
        RECT 93.575 193.975 93.865 194.020 ;
        RECT 97.700 193.960 98.020 194.020 ;
        RECT 111.975 194.160 112.265 194.205 ;
        RECT 112.420 194.160 112.740 194.220 ;
        RECT 111.975 194.020 112.740 194.160 ;
        RECT 111.975 193.975 112.265 194.020 ;
        RECT 112.420 193.960 112.740 194.020 ;
        RECT 115.180 193.960 115.500 194.220 ;
        RECT 86.660 193.820 86.980 193.880 ;
        RECT 96.320 193.820 96.640 193.880 ;
        RECT 103.235 193.820 103.525 193.865 ;
        RECT 105.520 193.820 105.840 193.880 ;
        RECT 117.940 193.820 118.260 193.880 ;
        RECT 72.400 193.680 74.930 193.820 ;
        RECT 84.910 193.680 95.170 193.820 ;
        RECT 48.495 193.480 48.785 193.525 ;
        RECT 45.720 193.340 48.785 193.480 ;
        RECT 45.720 193.280 46.040 193.340 ;
        RECT 48.495 193.295 48.785 193.340 ;
        RECT 49.420 193.480 49.710 193.525 ;
        RECT 51.255 193.480 51.545 193.525 ;
        RECT 54.835 193.480 55.125 193.525 ;
        RECT 49.420 193.340 55.125 193.480 ;
        RECT 49.420 193.295 49.710 193.340 ;
        RECT 51.255 193.295 51.545 193.340 ;
        RECT 54.835 193.295 55.125 193.340 ;
        RECT 55.915 193.320 56.205 193.635 ;
        RECT 66.050 193.540 66.190 193.680 ;
        RECT 72.400 193.620 72.720 193.680 ;
        RECT 65.960 193.280 66.280 193.540 ;
        RECT 68.720 193.280 69.040 193.540 ;
        RECT 72.860 193.280 73.180 193.540 ;
        RECT 74.790 193.525 74.930 193.680 ;
        RECT 86.660 193.620 86.980 193.680 ;
        RECT 74.715 193.480 75.005 193.525 ;
        RECT 76.080 193.480 76.400 193.540 ;
        RECT 74.715 193.340 76.400 193.480 ;
        RECT 74.715 193.295 75.005 193.340 ;
        RECT 76.080 193.280 76.400 193.340 ;
        RECT 85.740 193.480 86.060 193.540 ;
        RECT 86.215 193.480 86.505 193.525 ;
        RECT 85.740 193.340 86.505 193.480 ;
        RECT 85.740 193.280 86.060 193.340 ;
        RECT 86.215 193.295 86.505 193.340 ;
        RECT 89.880 193.280 90.200 193.540 ;
        RECT 93.190 193.525 93.330 193.680 ;
        RECT 93.115 193.295 93.405 193.525 ;
        RECT 94.480 193.280 94.800 193.540 ;
        RECT 95.030 193.480 95.170 193.680 ;
        RECT 96.320 193.680 118.260 193.820 ;
        RECT 96.320 193.620 96.640 193.680 ;
        RECT 103.235 193.635 103.525 193.680 ;
        RECT 105.520 193.620 105.840 193.680 ;
        RECT 117.940 193.620 118.260 193.680 ;
        RECT 108.755 193.480 109.045 193.525 ;
        RECT 115.640 193.480 115.960 193.540 ;
        RECT 95.030 193.340 115.960 193.480 ;
        RECT 108.755 193.295 109.045 193.340 ;
        RECT 115.640 193.280 115.960 193.340 ;
        RECT 48.940 192.940 49.260 193.200 ;
        RECT 50.320 192.940 50.640 193.200 ;
        RECT 70.115 193.140 70.405 193.185 ;
        RECT 70.115 193.000 72.170 193.140 ;
        RECT 70.115 192.955 70.405 193.000 ;
        RECT 72.030 192.845 72.170 193.000 ;
        RECT 84.820 192.940 85.140 193.200 ;
        RECT 107.820 193.140 108.140 193.200 ;
        RECT 110.580 193.140 110.900 193.200 ;
        RECT 107.820 193.000 110.900 193.140 ;
        RECT 107.820 192.940 108.140 193.000 ;
        RECT 110.580 192.940 110.900 193.000 ;
        RECT 111.515 192.955 111.805 193.185 ;
        RECT 49.825 192.800 50.115 192.845 ;
        RECT 51.715 192.800 52.005 192.845 ;
        RECT 54.835 192.800 55.125 192.845 ;
        RECT 49.825 192.660 55.125 192.800 ;
        RECT 49.825 192.615 50.115 192.660 ;
        RECT 51.715 192.615 52.005 192.660 ;
        RECT 54.835 192.615 55.125 192.660 ;
        RECT 71.955 192.615 72.245 192.845 ;
        RECT 111.590 192.800 111.730 192.955 ;
        RECT 111.960 192.800 112.280 192.860 ;
        RECT 111.590 192.660 112.280 192.800 ;
        RECT 111.960 192.600 112.280 192.660 ;
        RECT 48.035 192.460 48.325 192.505 ;
        RECT 54.000 192.460 54.320 192.520 ;
        RECT 48.035 192.320 54.320 192.460 ;
        RECT 48.035 192.275 48.325 192.320 ;
        RECT 54.000 192.260 54.320 192.320 ;
        RECT 65.500 192.260 65.820 192.520 ;
        RECT 70.100 192.260 70.420 192.520 ;
        RECT 72.400 192.460 72.720 192.520 ;
        RECT 72.875 192.460 73.165 192.505 ;
        RECT 72.400 192.320 73.165 192.460 ;
        RECT 72.400 192.260 72.720 192.320 ;
        RECT 72.875 192.275 73.165 192.320 ;
        RECT 88.055 192.460 88.345 192.505 ;
        RECT 90.800 192.460 91.120 192.520 ;
        RECT 88.055 192.320 91.120 192.460 ;
        RECT 88.055 192.275 88.345 192.320 ;
        RECT 90.800 192.260 91.120 192.320 ;
        RECT 109.200 192.260 109.520 192.520 ;
        RECT 113.815 192.460 114.105 192.505 ;
        RECT 118.860 192.460 119.180 192.520 ;
        RECT 113.815 192.320 119.180 192.460 ;
        RECT 113.815 192.275 114.105 192.320 ;
        RECT 118.860 192.260 119.180 192.320 ;
        RECT 14.370 191.640 127.530 192.120 ;
        RECT 50.320 191.440 50.640 191.500 ;
        RECT 50.795 191.440 51.085 191.485 ;
        RECT 50.320 191.300 51.085 191.440 ;
        RECT 50.320 191.240 50.640 191.300 ;
        RECT 50.795 191.255 51.085 191.300 ;
        RECT 85.280 191.440 85.600 191.500 ;
        RECT 85.280 191.300 93.330 191.440 ;
        RECT 85.280 191.240 85.600 191.300 ;
        RECT 40.170 191.100 40.460 191.145 ;
        RECT 42.950 191.100 43.240 191.145 ;
        RECT 44.810 191.100 45.100 191.145 ;
        RECT 40.170 190.960 45.100 191.100 ;
        RECT 40.170 190.915 40.460 190.960 ;
        RECT 42.950 190.915 43.240 190.960 ;
        RECT 44.810 190.915 45.100 190.960 ;
        RECT 49.415 190.915 49.705 191.145 ;
        RECT 55.035 191.100 55.325 191.145 ;
        RECT 58.155 191.100 58.445 191.145 ;
        RECT 60.045 191.100 60.335 191.145 ;
        RECT 55.035 190.960 60.335 191.100 ;
        RECT 55.035 190.915 55.325 190.960 ;
        RECT 58.155 190.915 58.445 190.960 ;
        RECT 60.045 190.915 60.335 190.960 ;
        RECT 36.305 190.760 36.595 190.805 ;
        RECT 41.120 190.760 41.440 190.820 ;
        RECT 36.305 190.620 45.950 190.760 ;
        RECT 36.305 190.575 36.595 190.620 ;
        RECT 41.120 190.560 41.440 190.620 ;
        RECT 40.170 190.420 40.460 190.465 ;
        RECT 43.435 190.420 43.725 190.465 ;
        RECT 44.800 190.420 45.120 190.480 ;
        RECT 40.170 190.280 42.705 190.420 ;
        RECT 40.170 190.235 40.460 190.280 ;
        RECT 38.310 190.080 38.600 190.125 ;
        RECT 38.820 190.080 39.140 190.140 ;
        RECT 42.490 190.125 42.705 190.280 ;
        RECT 43.435 190.280 45.120 190.420 ;
        RECT 43.435 190.235 43.725 190.280 ;
        RECT 44.800 190.220 45.120 190.280 ;
        RECT 45.275 190.235 45.565 190.465 ;
        RECT 45.810 190.420 45.950 190.620 ;
        RECT 46.180 190.560 46.500 190.820 ;
        RECT 47.575 190.420 47.865 190.465 ;
        RECT 45.810 190.280 47.865 190.420 ;
        RECT 49.490 190.420 49.630 190.915 ;
        RECT 63.660 190.900 63.980 191.160 ;
        RECT 64.695 191.100 64.985 191.145 ;
        RECT 67.815 191.100 68.105 191.145 ;
        RECT 69.705 191.100 69.995 191.145 ;
        RECT 76.555 191.100 76.845 191.145 ;
        RECT 64.695 190.960 69.995 191.100 ;
        RECT 64.695 190.915 64.985 190.960 ;
        RECT 67.815 190.915 68.105 190.960 ;
        RECT 69.705 190.915 69.995 190.960 ;
        RECT 73.410 190.960 76.845 191.100 ;
        RECT 52.160 190.560 52.480 190.820 ;
        RECT 59.060 190.760 59.380 190.820 ;
        RECT 60.915 190.760 61.205 190.805 ;
        RECT 63.750 190.760 63.890 190.900 ;
        RECT 70.575 190.760 70.865 190.805 ;
        RECT 59.060 190.620 70.865 190.760 ;
        RECT 59.060 190.560 59.380 190.620 ;
        RECT 60.915 190.575 61.205 190.620 ;
        RECT 70.575 190.575 70.865 190.620 ;
        RECT 71.020 190.760 71.340 190.820 ;
        RECT 73.410 190.805 73.550 190.960 ;
        RECT 76.555 190.915 76.845 190.960 ;
        RECT 87.090 191.100 87.380 191.145 ;
        RECT 89.870 191.100 90.160 191.145 ;
        RECT 91.730 191.100 92.020 191.145 ;
        RECT 87.090 190.960 92.020 191.100 ;
        RECT 93.190 191.100 93.330 191.300 ;
        RECT 93.560 191.240 93.880 191.500 ;
        RECT 102.775 191.440 103.065 191.485 ;
        RECT 104.140 191.440 104.460 191.500 ;
        RECT 112.420 191.440 112.740 191.500 ;
        RECT 102.775 191.300 104.460 191.440 ;
        RECT 102.775 191.255 103.065 191.300 ;
        RECT 104.140 191.240 104.460 191.300 ;
        RECT 108.370 191.300 112.740 191.440 ;
        RECT 107.820 191.100 108.140 191.160 ;
        RECT 93.190 190.960 97.010 191.100 ;
        RECT 87.090 190.915 87.380 190.960 ;
        RECT 89.870 190.915 90.160 190.960 ;
        RECT 91.730 190.915 92.020 190.960 ;
        RECT 73.335 190.760 73.625 190.805 ;
        RECT 71.020 190.620 73.625 190.760 ;
        RECT 71.020 190.560 71.340 190.620 ;
        RECT 73.335 190.575 73.625 190.620 ;
        RECT 77.935 190.760 78.225 190.805 ;
        RECT 79.760 190.760 80.080 190.820 ;
        RECT 77.935 190.620 80.080 190.760 ;
        RECT 77.935 190.575 78.225 190.620 ;
        RECT 79.760 190.560 80.080 190.620 ;
        RECT 92.195 190.760 92.485 190.805 ;
        RECT 93.560 190.760 93.880 190.820 ;
        RECT 92.195 190.620 96.550 190.760 ;
        RECT 92.195 190.575 92.485 190.620 ;
        RECT 93.560 190.560 93.880 190.620 ;
        RECT 96.410 190.480 96.550 190.620 ;
        RECT 51.715 190.420 52.005 190.465 ;
        RECT 54.000 190.440 54.320 190.480 ;
        RECT 49.490 190.280 52.005 190.420 ;
        RECT 47.575 190.235 47.865 190.280 ;
        RECT 51.715 190.235 52.005 190.280 ;
        RECT 41.570 190.080 41.860 190.125 ;
        RECT 38.310 189.940 41.860 190.080 ;
        RECT 38.310 189.895 38.600 189.940 ;
        RECT 38.820 189.880 39.140 189.940 ;
        RECT 41.570 189.895 41.860 189.940 ;
        RECT 42.490 190.080 42.780 190.125 ;
        RECT 44.350 190.080 44.640 190.125 ;
        RECT 42.490 189.940 44.640 190.080 ;
        RECT 45.350 190.080 45.490 190.235 ;
        RECT 53.955 190.220 54.320 190.440 ;
        RECT 55.035 190.420 55.325 190.465 ;
        RECT 58.615 190.420 58.905 190.465 ;
        RECT 60.450 190.420 60.740 190.465 ;
        RECT 55.035 190.280 60.740 190.420 ;
        RECT 55.035 190.235 55.325 190.280 ;
        RECT 58.615 190.235 58.905 190.280 ;
        RECT 60.450 190.235 60.740 190.280 ;
        RECT 48.940 190.080 49.260 190.140 ;
        RECT 53.955 190.125 54.245 190.220 ;
        RECT 45.350 189.940 49.260 190.080 ;
        RECT 42.490 189.895 42.780 189.940 ;
        RECT 44.350 189.895 44.640 189.940 ;
        RECT 48.940 189.880 49.260 189.940 ;
        RECT 53.655 190.080 54.245 190.125 ;
        RECT 56.895 190.080 57.545 190.125 ;
        RECT 53.655 189.940 57.545 190.080 ;
        RECT 53.655 189.895 53.945 189.940 ;
        RECT 56.895 189.895 57.545 189.940 ;
        RECT 59.535 190.080 59.825 190.125 ;
        RECT 59.980 190.080 60.300 190.140 ;
        RECT 63.615 190.125 63.905 190.440 ;
        RECT 64.695 190.420 64.985 190.465 ;
        RECT 68.275 190.420 68.565 190.465 ;
        RECT 70.110 190.420 70.400 190.465 ;
        RECT 64.695 190.280 70.400 190.420 ;
        RECT 64.695 190.235 64.985 190.280 ;
        RECT 68.275 190.235 68.565 190.280 ;
        RECT 70.110 190.235 70.400 190.280 ;
        RECT 72.860 190.220 73.180 190.480 ;
        RECT 74.240 190.420 74.560 190.480 ;
        RECT 76.095 190.420 76.385 190.465 ;
        RECT 74.240 190.280 76.385 190.420 ;
        RECT 74.240 190.220 74.560 190.280 ;
        RECT 76.095 190.235 76.385 190.280 ;
        RECT 87.090 190.420 87.380 190.465 ;
        RECT 87.090 190.280 89.625 190.420 ;
        RECT 87.090 190.235 87.380 190.280 ;
        RECT 59.535 189.940 60.300 190.080 ;
        RECT 59.535 189.895 59.825 189.940 ;
        RECT 59.980 189.880 60.300 189.940 ;
        RECT 63.315 190.080 63.905 190.125 ;
        RECT 65.500 190.080 65.820 190.140 ;
        RECT 66.555 190.080 67.205 190.125 ;
        RECT 63.315 189.940 67.205 190.080 ;
        RECT 63.315 189.895 63.605 189.940 ;
        RECT 65.500 189.880 65.820 189.940 ;
        RECT 66.555 189.895 67.205 189.940 ;
        RECT 69.195 190.080 69.485 190.125 ;
        RECT 73.320 190.080 73.640 190.140 ;
        RECT 76.555 190.080 76.845 190.125 ;
        RECT 69.195 189.940 71.250 190.080 ;
        RECT 69.195 189.895 69.485 189.940 ;
        RECT 47.115 189.740 47.405 189.785 ;
        RECT 57.680 189.740 58.000 189.800 ;
        RECT 47.115 189.600 58.000 189.740 ;
        RECT 47.115 189.555 47.405 189.600 ;
        RECT 57.680 189.540 58.000 189.600 ;
        RECT 61.820 189.540 62.140 189.800 ;
        RECT 65.960 189.740 66.280 189.800 ;
        RECT 69.640 189.740 69.960 189.800 ;
        RECT 71.110 189.785 71.250 189.940 ;
        RECT 73.320 189.940 76.845 190.080 ;
        RECT 73.320 189.880 73.640 189.940 ;
        RECT 76.555 189.895 76.845 189.940 ;
        RECT 85.230 190.080 85.520 190.125 ;
        RECT 87.580 190.080 87.900 190.140 ;
        RECT 89.410 190.125 89.625 190.280 ;
        RECT 90.340 190.220 90.660 190.480 ;
        RECT 90.800 190.420 91.120 190.480 ;
        RECT 92.655 190.420 92.945 190.465 ;
        RECT 90.800 190.280 92.945 190.420 ;
        RECT 90.800 190.220 91.120 190.280 ;
        RECT 92.655 190.235 92.945 190.280 ;
        RECT 96.320 190.220 96.640 190.480 ;
        RECT 96.870 190.420 97.010 190.960 ;
        RECT 97.790 190.960 108.140 191.100 ;
        RECT 97.790 190.820 97.930 190.960 ;
        RECT 97.700 190.560 98.020 190.820 ;
        RECT 98.635 190.760 98.925 190.805 ;
        RECT 100.920 190.760 101.240 190.820 ;
        RECT 105.150 190.805 105.290 190.960 ;
        RECT 107.820 190.900 108.140 190.960 ;
        RECT 98.635 190.620 102.530 190.760 ;
        RECT 98.635 190.575 98.925 190.620 ;
        RECT 100.920 190.560 101.240 190.620 ;
        RECT 99.095 190.420 99.385 190.465 ;
        RECT 101.855 190.420 102.145 190.465 ;
        RECT 96.870 190.280 99.385 190.420 ;
        RECT 99.095 190.235 99.385 190.280 ;
        RECT 101.010 190.280 102.145 190.420 ;
        RECT 102.390 190.420 102.530 190.620 ;
        RECT 105.075 190.575 105.365 190.805 ;
        RECT 105.980 190.760 106.300 190.820 ;
        RECT 108.370 190.760 108.510 191.300 ;
        RECT 112.420 191.240 112.740 191.300 ;
        RECT 117.480 191.440 117.800 191.500 ;
        RECT 117.955 191.440 118.245 191.485 ;
        RECT 117.480 191.300 118.245 191.440 ;
        RECT 117.480 191.240 117.800 191.300 ;
        RECT 117.955 191.255 118.245 191.300 ;
        RECT 111.615 191.100 111.905 191.145 ;
        RECT 114.735 191.100 115.025 191.145 ;
        RECT 116.625 191.100 116.915 191.145 ;
        RECT 111.615 190.960 116.915 191.100 ;
        RECT 111.615 190.915 111.905 190.960 ;
        RECT 114.735 190.915 115.025 190.960 ;
        RECT 116.625 190.915 116.915 190.960 ;
        RECT 105.980 190.620 108.510 190.760 ;
        RECT 108.755 190.760 109.045 190.805 ;
        RECT 109.660 190.760 109.980 190.820 ;
        RECT 108.755 190.620 109.980 190.760 ;
        RECT 105.980 190.560 106.300 190.620 ;
        RECT 108.755 190.575 109.045 190.620 ;
        RECT 109.660 190.560 109.980 190.620 ;
        RECT 106.455 190.420 106.745 190.465 ;
        RECT 102.390 190.280 106.745 190.420 ;
        RECT 88.490 190.080 88.780 190.125 ;
        RECT 85.230 189.940 88.780 190.080 ;
        RECT 85.230 189.895 85.520 189.940 ;
        RECT 87.580 189.880 87.900 189.940 ;
        RECT 88.490 189.895 88.780 189.940 ;
        RECT 89.410 190.080 89.700 190.125 ;
        RECT 91.270 190.080 91.560 190.125 ;
        RECT 89.410 189.940 91.560 190.080 ;
        RECT 89.410 189.895 89.700 189.940 ;
        RECT 91.270 189.895 91.560 189.940 ;
        RECT 65.960 189.600 69.960 189.740 ;
        RECT 65.960 189.540 66.280 189.600 ;
        RECT 69.640 189.540 69.960 189.600 ;
        RECT 71.035 189.555 71.325 189.785 ;
        RECT 76.080 189.740 76.400 189.800 ;
        RECT 77.015 189.740 77.305 189.785 ;
        RECT 76.080 189.600 77.305 189.740 ;
        RECT 76.080 189.540 76.400 189.600 ;
        RECT 77.015 189.555 77.305 189.600 ;
        RECT 83.225 189.740 83.515 189.785 ;
        RECT 85.740 189.740 86.060 189.800 ;
        RECT 101.010 189.785 101.150 190.280 ;
        RECT 101.855 190.235 102.145 190.280 ;
        RECT 106.455 190.235 106.745 190.280 ;
        RECT 109.200 190.080 109.520 190.140 ;
        RECT 110.535 190.125 110.825 190.440 ;
        RECT 111.615 190.420 111.905 190.465 ;
        RECT 115.195 190.420 115.485 190.465 ;
        RECT 117.030 190.420 117.320 190.465 ;
        RECT 111.615 190.280 117.320 190.420 ;
        RECT 111.615 190.235 111.905 190.280 ;
        RECT 115.195 190.235 115.485 190.280 ;
        RECT 117.030 190.235 117.320 190.280 ;
        RECT 117.495 190.420 117.785 190.465 ;
        RECT 117.940 190.420 118.260 190.480 ;
        RECT 117.495 190.280 118.260 190.420 ;
        RECT 117.495 190.235 117.785 190.280 ;
        RECT 117.940 190.220 118.260 190.280 ;
        RECT 118.860 190.220 119.180 190.480 ;
        RECT 110.235 190.080 110.825 190.125 ;
        RECT 113.475 190.080 114.125 190.125 ;
        RECT 109.200 189.940 114.125 190.080 ;
        RECT 109.200 189.880 109.520 189.940 ;
        RECT 110.235 189.895 110.525 189.940 ;
        RECT 113.475 189.895 114.125 189.940 ;
        RECT 116.100 189.880 116.420 190.140 ;
        RECT 83.225 189.600 86.060 189.740 ;
        RECT 83.225 189.555 83.515 189.600 ;
        RECT 85.740 189.540 86.060 189.600 ;
        RECT 100.935 189.555 101.225 189.785 ;
        RECT 108.295 189.740 108.585 189.785 ;
        RECT 112.880 189.740 113.200 189.800 ;
        RECT 108.295 189.600 113.200 189.740 ;
        RECT 108.295 189.555 108.585 189.600 ;
        RECT 112.880 189.540 113.200 189.600 ;
        RECT 14.370 188.920 127.530 189.400 ;
        RECT 57.680 188.520 58.000 188.780 ;
        RECT 59.535 188.535 59.825 188.765 ;
        RECT 36.075 188.380 36.365 188.425 ;
        RECT 38.935 188.380 39.225 188.425 ;
        RECT 42.175 188.380 42.825 188.425 ;
        RECT 36.075 188.240 42.825 188.380 ;
        RECT 36.075 188.195 36.365 188.240 ;
        RECT 38.935 188.195 39.525 188.240 ;
        RECT 42.175 188.195 42.825 188.240 ;
        RECT 30.095 188.040 30.385 188.085 ;
        RECT 35.615 188.040 35.905 188.085 ;
        RECT 30.095 187.900 36.290 188.040 ;
        RECT 30.095 187.855 30.385 187.900 ;
        RECT 35.615 187.855 35.905 187.900 ;
        RECT 36.150 187.760 36.290 187.900 ;
        RECT 39.235 187.880 39.525 188.195 ;
        RECT 40.315 188.040 40.605 188.085 ;
        RECT 43.895 188.040 44.185 188.085 ;
        RECT 45.730 188.040 46.020 188.085 ;
        RECT 40.315 187.900 46.020 188.040 ;
        RECT 40.315 187.855 40.605 187.900 ;
        RECT 43.895 187.855 44.185 187.900 ;
        RECT 45.730 187.855 46.020 187.900 ;
        RECT 55.380 187.840 55.700 188.100 ;
        RECT 56.300 188.040 56.620 188.100 ;
        RECT 57.235 188.040 57.525 188.085 ;
        RECT 56.300 187.900 57.525 188.040 ;
        RECT 59.610 188.040 59.750 188.535 ;
        RECT 59.980 188.520 60.300 188.780 ;
        RECT 66.895 188.720 67.185 188.765 ;
        RECT 72.860 188.720 73.180 188.780 ;
        RECT 66.895 188.580 73.180 188.720 ;
        RECT 66.895 188.535 67.185 188.580 ;
        RECT 72.860 188.520 73.180 188.580 ;
        RECT 87.135 188.720 87.425 188.765 ;
        RECT 87.580 188.720 87.900 188.780 ;
        RECT 87.135 188.580 87.900 188.720 ;
        RECT 87.135 188.535 87.425 188.580 ;
        RECT 87.580 188.520 87.900 188.580 ;
        RECT 89.895 188.720 90.185 188.765 ;
        RECT 90.340 188.720 90.660 188.780 ;
        RECT 89.895 188.580 90.660 188.720 ;
        RECT 89.895 188.535 90.185 188.580 ;
        RECT 90.340 188.520 90.660 188.580 ;
        RECT 105.980 188.720 106.300 188.780 ;
        RECT 106.915 188.720 107.205 188.765 ;
        RECT 105.980 188.580 107.205 188.720 ;
        RECT 105.980 188.520 106.300 188.580 ;
        RECT 106.915 188.535 107.205 188.580 ;
        RECT 113.815 188.720 114.105 188.765 ;
        RECT 116.100 188.720 116.420 188.780 ;
        RECT 113.815 188.580 116.420 188.720 ;
        RECT 113.815 188.535 114.105 188.580 ;
        RECT 116.100 188.520 116.420 188.580 ;
        RECT 99.195 188.380 99.485 188.425 ;
        RECT 100.000 188.380 100.320 188.440 ;
        RECT 102.435 188.380 103.085 188.425 ;
        RECT 99.195 188.240 103.085 188.380 ;
        RECT 99.195 188.195 99.785 188.240 ;
        RECT 60.915 188.040 61.205 188.085 ;
        RECT 59.610 187.900 61.205 188.040 ;
        RECT 56.300 187.840 56.620 187.900 ;
        RECT 57.235 187.855 57.525 187.900 ;
        RECT 60.915 187.855 61.205 187.900 ;
        RECT 87.595 187.855 87.885 188.085 ;
        RECT 28.240 187.700 28.560 187.760 ;
        RECT 29.635 187.700 29.925 187.745 ;
        RECT 28.240 187.560 29.925 187.700 ;
        RECT 28.240 187.500 28.560 187.560 ;
        RECT 29.635 187.515 29.925 187.560 ;
        RECT 36.060 187.500 36.380 187.760 ;
        RECT 44.340 187.700 44.660 187.760 ;
        RECT 46.195 187.700 46.485 187.745 ;
        RECT 44.340 187.560 46.485 187.700 ;
        RECT 44.340 187.500 44.660 187.560 ;
        RECT 46.195 187.515 46.485 187.560 ;
        RECT 46.640 187.700 46.960 187.760 ;
        RECT 56.775 187.700 57.065 187.745 ;
        RECT 46.640 187.560 57.065 187.700 ;
        RECT 40.315 187.360 40.605 187.405 ;
        RECT 43.435 187.360 43.725 187.405 ;
        RECT 45.325 187.360 45.615 187.405 ;
        RECT 40.315 187.220 45.615 187.360 ;
        RECT 46.270 187.360 46.410 187.515 ;
        RECT 46.640 187.500 46.960 187.560 ;
        RECT 56.775 187.515 57.065 187.560 ;
        RECT 61.820 187.700 62.140 187.760 ;
        RECT 64.135 187.700 64.425 187.745 ;
        RECT 65.500 187.700 65.820 187.760 ;
        RECT 71.940 187.700 72.260 187.760 ;
        RECT 61.820 187.560 72.260 187.700 ;
        RECT 87.670 187.700 87.810 187.855 ;
        RECT 88.960 187.840 89.280 188.100 ;
        RECT 99.495 187.880 99.785 188.195 ;
        RECT 100.000 188.180 100.320 188.240 ;
        RECT 102.435 188.195 103.085 188.240 ;
        RECT 100.575 188.040 100.865 188.085 ;
        RECT 104.155 188.040 104.445 188.085 ;
        RECT 105.990 188.040 106.280 188.085 ;
        RECT 100.575 187.900 106.280 188.040 ;
        RECT 100.575 187.855 100.865 187.900 ;
        RECT 104.155 187.855 104.445 187.900 ;
        RECT 105.990 187.855 106.280 187.900 ;
        RECT 109.660 187.840 109.980 188.100 ;
        RECT 112.880 187.840 113.200 188.100 ;
        RECT 89.880 187.700 90.200 187.760 ;
        RECT 90.800 187.700 91.120 187.760 ;
        RECT 87.670 187.560 91.120 187.700 ;
        RECT 61.820 187.500 62.140 187.560 ;
        RECT 64.135 187.515 64.425 187.560 ;
        RECT 65.500 187.500 65.820 187.560 ;
        RECT 71.940 187.500 72.260 187.560 ;
        RECT 89.880 187.500 90.200 187.560 ;
        RECT 90.800 187.500 91.120 187.560 ;
        RECT 106.455 187.700 106.745 187.745 ;
        RECT 117.940 187.700 118.260 187.760 ;
        RECT 106.455 187.560 118.260 187.700 ;
        RECT 106.455 187.515 106.745 187.560 ;
        RECT 117.940 187.500 118.260 187.560 ;
        RECT 48.940 187.360 49.260 187.420 ;
        RECT 59.060 187.360 59.380 187.420 ;
        RECT 46.270 187.220 59.380 187.360 ;
        RECT 40.315 187.175 40.605 187.220 ;
        RECT 43.435 187.175 43.725 187.220 ;
        RECT 45.325 187.175 45.615 187.220 ;
        RECT 48.940 187.160 49.260 187.220 ;
        RECT 59.060 187.160 59.380 187.220 ;
        RECT 100.575 187.360 100.865 187.405 ;
        RECT 103.695 187.360 103.985 187.405 ;
        RECT 105.585 187.360 105.875 187.405 ;
        RECT 100.575 187.220 105.875 187.360 ;
        RECT 100.575 187.175 100.865 187.220 ;
        RECT 103.695 187.175 103.985 187.220 ;
        RECT 105.585 187.175 105.875 187.220 ;
        RECT 37.440 186.820 37.760 187.080 ;
        RECT 44.910 187.020 45.200 187.065 ;
        RECT 49.860 187.020 50.180 187.080 ;
        RECT 44.910 186.880 50.180 187.020 ;
        RECT 44.910 186.835 45.200 186.880 ;
        RECT 49.860 186.820 50.180 186.880 ;
        RECT 97.715 187.020 98.005 187.065 ;
        RECT 99.080 187.020 99.400 187.080 ;
        RECT 97.715 186.880 99.400 187.020 ;
        RECT 97.715 186.835 98.005 186.880 ;
        RECT 99.080 186.820 99.400 186.880 ;
        RECT 99.540 187.020 99.860 187.080 ;
        RECT 105.140 187.020 105.430 187.065 ;
        RECT 99.540 186.880 105.430 187.020 ;
        RECT 99.540 186.820 99.860 186.880 ;
        RECT 105.140 186.835 105.430 186.880 ;
        RECT 14.370 186.200 127.530 186.680 ;
        RECT 38.820 185.800 39.140 186.060 ;
        RECT 45.720 186.000 46.040 186.060 ;
        RECT 88.055 186.000 88.345 186.045 ;
        RECT 88.960 186.000 89.280 186.060 ;
        RECT 45.720 185.860 47.330 186.000 ;
        RECT 45.720 185.800 46.040 185.860 ;
        RECT 28.815 185.660 29.105 185.705 ;
        RECT 31.935 185.660 32.225 185.705 ;
        RECT 33.825 185.660 34.115 185.705 ;
        RECT 44.340 185.660 44.660 185.720 ;
        RECT 28.815 185.520 34.115 185.660 ;
        RECT 28.815 185.475 29.105 185.520 ;
        RECT 31.935 185.475 32.225 185.520 ;
        RECT 33.825 185.475 34.115 185.520 ;
        RECT 34.770 185.520 44.660 185.660 ;
        RECT 22.720 185.320 23.040 185.380 ;
        RECT 34.770 185.365 34.910 185.520 ;
        RECT 44.340 185.460 44.660 185.520 ;
        RECT 46.180 185.460 46.500 185.720 ;
        RECT 33.315 185.320 33.605 185.365 ;
        RECT 22.720 185.180 33.605 185.320 ;
        RECT 22.720 185.120 23.040 185.180 ;
        RECT 33.315 185.135 33.605 185.180 ;
        RECT 34.695 185.135 34.985 185.365 ;
        RECT 37.900 185.320 38.220 185.380 ;
        RECT 40.215 185.320 40.505 185.365 ;
        RECT 37.900 185.180 40.505 185.320 ;
        RECT 37.900 185.120 38.220 185.180 ;
        RECT 40.215 185.135 40.505 185.180 ;
        RECT 27.735 184.685 28.025 185.000 ;
        RECT 28.815 184.980 29.105 185.025 ;
        RECT 32.395 184.980 32.685 185.025 ;
        RECT 34.230 184.980 34.520 185.025 ;
        RECT 28.815 184.840 34.520 184.980 ;
        RECT 28.815 184.795 29.105 184.840 ;
        RECT 32.395 184.795 32.685 184.840 ;
        RECT 34.230 184.795 34.520 184.840 ;
        RECT 36.060 184.980 36.380 185.040 ;
        RECT 38.375 184.980 38.665 185.025 ;
        RECT 36.060 184.840 38.665 184.980 ;
        RECT 40.290 184.980 40.430 185.135 ;
        RECT 41.120 185.120 41.440 185.380 ;
        RECT 46.270 185.320 46.410 185.460 ;
        RECT 46.655 185.320 46.945 185.365 ;
        RECT 45.810 185.180 46.945 185.320 ;
        RECT 45.260 184.980 45.580 185.040 ;
        RECT 45.810 184.980 45.950 185.180 ;
        RECT 46.655 185.135 46.945 185.180 ;
        RECT 40.290 184.840 45.950 184.980 ;
        RECT 36.060 184.780 36.380 184.840 ;
        RECT 38.375 184.795 38.665 184.840 ;
        RECT 45.260 184.780 45.580 184.840 ;
        RECT 46.195 184.795 46.485 185.025 ;
        RECT 47.190 184.980 47.330 185.860 ;
        RECT 88.055 185.860 89.280 186.000 ;
        RECT 88.055 185.815 88.345 185.860 ;
        RECT 88.960 185.800 89.280 185.860 ;
        RECT 99.540 185.800 99.860 186.060 ;
        RECT 100.000 186.000 100.320 186.060 ;
        RECT 100.475 186.000 100.765 186.045 ;
        RECT 100.000 185.860 100.765 186.000 ;
        RECT 100.000 185.800 100.320 185.860 ;
        RECT 100.475 185.815 100.765 185.860 ;
        RECT 53.195 185.660 53.485 185.705 ;
        RECT 56.315 185.660 56.605 185.705 ;
        RECT 58.205 185.660 58.495 185.705 ;
        RECT 60.440 185.660 60.760 185.720 ;
        RECT 53.195 185.520 58.495 185.660 ;
        RECT 53.195 185.475 53.485 185.520 ;
        RECT 56.315 185.475 56.605 185.520 ;
        RECT 58.205 185.475 58.495 185.520 ;
        RECT 58.690 185.520 60.760 185.660 ;
        RECT 58.690 185.320 58.830 185.520 ;
        RECT 60.440 185.460 60.760 185.520 ;
        RECT 71.020 185.660 71.340 185.720 ;
        RECT 74.715 185.660 75.005 185.705 ;
        RECT 76.080 185.660 76.400 185.720 ;
        RECT 71.020 185.520 76.400 185.660 ;
        RECT 71.020 185.460 71.340 185.520 ;
        RECT 74.715 185.475 75.005 185.520 ;
        RECT 76.080 185.460 76.400 185.520 ;
        RECT 90.800 185.660 91.120 185.720 ;
        RECT 90.800 185.520 100.230 185.660 ;
        RECT 90.800 185.460 91.120 185.520 ;
        RECT 51.790 185.180 58.830 185.320 ;
        RECT 48.495 184.980 48.785 185.025 ;
        RECT 51.790 184.980 51.930 185.180 ;
        RECT 59.060 185.120 59.380 185.380 ;
        RECT 67.800 185.320 68.120 185.380 ;
        RECT 72.415 185.320 72.705 185.365 ;
        RECT 73.320 185.320 73.640 185.380 ;
        RECT 67.800 185.180 73.640 185.320 ;
        RECT 67.800 185.120 68.120 185.180 ;
        RECT 72.415 185.135 72.705 185.180 ;
        RECT 73.320 185.120 73.640 185.180 ;
        RECT 84.820 185.120 85.140 185.380 ;
        RECT 94.495 185.320 94.785 185.365 ;
        RECT 99.080 185.320 99.400 185.380 ;
        RECT 94.495 185.180 99.400 185.320 ;
        RECT 94.495 185.135 94.785 185.180 ;
        RECT 99.080 185.120 99.400 185.180 ;
        RECT 47.190 184.840 51.930 184.980 ;
        RECT 48.495 184.795 48.785 184.840 ;
        RECT 27.435 184.640 28.025 184.685 ;
        RECT 28.240 184.640 28.560 184.700 ;
        RECT 30.675 184.640 31.325 184.685 ;
        RECT 27.435 184.500 31.325 184.640 ;
        RECT 27.435 184.455 27.725 184.500 ;
        RECT 28.240 184.440 28.560 184.500 ;
        RECT 30.675 184.455 31.325 184.500 ;
        RECT 37.440 184.640 37.760 184.700 ;
        RECT 46.270 184.640 46.410 184.795 ;
        RECT 52.115 184.685 52.405 185.000 ;
        RECT 53.195 184.980 53.485 185.025 ;
        RECT 56.775 184.980 57.065 185.025 ;
        RECT 58.610 184.980 58.900 185.025 ;
        RECT 53.195 184.840 58.900 184.980 ;
        RECT 53.195 184.795 53.485 184.840 ;
        RECT 56.775 184.795 57.065 184.840 ;
        RECT 58.610 184.795 58.900 184.840 ;
        RECT 74.240 184.780 74.560 185.040 ;
        RECT 100.090 185.025 100.230 185.520 ;
        RECT 105.060 185.320 105.380 185.380 ;
        RECT 106.915 185.320 107.205 185.365 ;
        RECT 108.740 185.320 109.060 185.380 ;
        RECT 105.060 185.180 109.060 185.320 ;
        RECT 105.060 185.120 105.380 185.180 ;
        RECT 106.915 185.135 107.205 185.180 ;
        RECT 108.740 185.120 109.060 185.180 ;
        RECT 98.635 184.795 98.925 185.025 ;
        RECT 100.015 184.795 100.305 185.025 ;
        RECT 37.440 184.500 46.410 184.640 ;
        RECT 48.955 184.640 49.245 184.685 ;
        RECT 51.815 184.640 52.405 184.685 ;
        RECT 55.055 184.640 55.705 184.685 ;
        RECT 48.955 184.500 55.705 184.640 ;
        RECT 37.440 184.440 37.760 184.500 ;
        RECT 48.955 184.455 49.245 184.500 ;
        RECT 51.815 184.455 52.105 184.500 ;
        RECT 55.055 184.455 55.705 184.500 ;
        RECT 57.680 184.440 58.000 184.700 ;
        RECT 71.955 184.640 72.245 184.685 ;
        RECT 72.400 184.640 72.720 184.700 ;
        RECT 71.955 184.500 72.720 184.640 ;
        RECT 74.330 184.640 74.470 184.780 ;
        RECT 74.715 184.640 75.005 184.685 ;
        RECT 75.620 184.640 75.940 184.700 ;
        RECT 74.330 184.500 75.940 184.640 ;
        RECT 98.710 184.640 98.850 184.795 ;
        RECT 105.520 184.780 105.840 185.040 ;
        RECT 110.120 184.780 110.440 185.040 ;
        RECT 102.315 184.640 102.605 184.685 ;
        RECT 98.710 184.500 102.605 184.640 ;
        RECT 71.955 184.455 72.245 184.500 ;
        RECT 72.400 184.440 72.720 184.500 ;
        RECT 74.715 184.455 75.005 184.500 ;
        RECT 75.620 184.440 75.940 184.500 ;
        RECT 102.315 184.455 102.605 184.500 ;
        RECT 109.675 184.640 109.965 184.685 ;
        RECT 111.960 184.640 112.280 184.700 ;
        RECT 109.675 184.500 112.280 184.640 ;
        RECT 109.675 184.455 109.965 184.500 ;
        RECT 111.960 184.440 112.280 184.500 ;
        RECT 25.955 184.300 26.245 184.345 ;
        RECT 29.620 184.300 29.940 184.360 ;
        RECT 25.955 184.160 29.940 184.300 ;
        RECT 25.955 184.115 26.245 184.160 ;
        RECT 29.620 184.100 29.940 184.160 ;
        RECT 30.080 184.300 30.400 184.360 ;
        RECT 41.595 184.300 41.885 184.345 ;
        RECT 30.080 184.160 41.885 184.300 ;
        RECT 30.080 184.100 30.400 184.160 ;
        RECT 41.595 184.115 41.885 184.160 ;
        RECT 43.420 184.100 43.740 184.360 ;
        RECT 43.880 184.100 44.200 184.360 ;
        RECT 45.720 184.100 46.040 184.360 ;
        RECT 46.180 184.300 46.500 184.360 ;
        RECT 50.335 184.300 50.625 184.345 ;
        RECT 46.180 184.160 50.625 184.300 ;
        RECT 46.180 184.100 46.500 184.160 ;
        RECT 50.335 184.115 50.625 184.160 ;
        RECT 71.035 184.300 71.325 184.345 ;
        RECT 74.240 184.300 74.560 184.360 ;
        RECT 71.035 184.160 74.560 184.300 ;
        RECT 71.035 184.115 71.325 184.160 ;
        RECT 74.240 184.100 74.560 184.160 ;
        RECT 85.740 184.100 86.060 184.360 ;
        RECT 86.200 184.100 86.520 184.360 ;
        RECT 97.240 184.100 97.560 184.360 ;
        RECT 111.500 184.300 111.820 184.360 ;
        RECT 113.355 184.300 113.645 184.345 ;
        RECT 111.500 184.160 113.645 184.300 ;
        RECT 111.500 184.100 111.820 184.160 ;
        RECT 113.355 184.115 113.645 184.160 ;
        RECT 14.370 183.480 127.530 183.960 ;
        RECT 22.720 183.080 23.040 183.340 ;
        RECT 30.080 183.080 30.400 183.340 ;
        RECT 44.800 183.280 45.120 183.340 ;
        RECT 48.495 183.280 48.785 183.325 ;
        RECT 44.800 183.140 48.785 183.280 ;
        RECT 44.800 183.080 45.120 183.140 ;
        RECT 48.495 183.095 48.785 183.140 ;
        RECT 49.860 183.080 50.180 183.340 ;
        RECT 52.175 183.280 52.465 183.325 ;
        RECT 57.680 183.280 58.000 183.340 ;
        RECT 71.020 183.280 71.340 183.340 ;
        RECT 52.175 183.140 58.000 183.280 ;
        RECT 52.175 183.095 52.465 183.140 ;
        RECT 57.680 183.080 58.000 183.140 ;
        RECT 68.810 183.140 71.340 183.280 ;
        RECT 32.395 182.940 32.685 182.985 ;
        RECT 33.760 182.940 34.080 183.000 ;
        RECT 32.395 182.800 34.080 182.940 ;
        RECT 32.395 182.755 32.685 182.800 ;
        RECT 33.760 182.740 34.080 182.800 ;
        RECT 44.355 182.940 44.645 182.985 ;
        RECT 44.355 182.800 51.010 182.940 ;
        RECT 44.355 182.755 44.645 182.800 ;
        RECT 21.815 182.600 22.105 182.645 ;
        RECT 23.195 182.600 23.485 182.645 ;
        RECT 21.815 182.460 23.485 182.600 ;
        RECT 21.815 182.415 22.105 182.460 ;
        RECT 23.195 182.415 23.485 182.460 ;
        RECT 27.335 182.600 27.625 182.645 ;
        RECT 29.620 182.600 29.940 182.660 ;
        RECT 32.855 182.600 33.145 182.645 ;
        RECT 35.600 182.600 35.920 182.660 ;
        RECT 27.335 182.460 35.920 182.600 ;
        RECT 27.335 182.415 27.625 182.460 ;
        RECT 29.620 182.400 29.940 182.460 ;
        RECT 32.855 182.415 33.145 182.460 ;
        RECT 35.600 182.400 35.920 182.460 ;
        RECT 37.440 182.400 37.760 182.660 ;
        RECT 41.595 182.600 41.885 182.645 ;
        RECT 43.880 182.600 44.200 182.660 ;
        RECT 41.595 182.460 44.200 182.600 ;
        RECT 41.595 182.415 41.885 182.460 ;
        RECT 43.880 182.400 44.200 182.460 ;
        RECT 45.275 182.600 45.565 182.645 ;
        RECT 46.180 182.600 46.500 182.660 ;
        RECT 50.870 182.645 51.010 182.800 ;
        RECT 45.275 182.460 46.500 182.600 ;
        RECT 45.275 182.415 45.565 182.460 ;
        RECT 46.180 182.400 46.500 182.460 ;
        RECT 49.415 182.415 49.705 182.645 ;
        RECT 50.795 182.415 51.085 182.645 ;
        RECT 51.255 182.415 51.545 182.645 ;
        RECT 55.395 182.600 55.685 182.645 ;
        RECT 59.060 182.600 59.380 182.660 ;
        RECT 55.395 182.460 59.380 182.600 ;
        RECT 55.395 182.415 55.685 182.460 ;
        RECT 26.415 182.075 26.705 182.305 ;
        RECT 33.775 182.260 34.065 182.305 ;
        RECT 37.900 182.260 38.220 182.320 ;
        RECT 33.775 182.120 38.220 182.260 ;
        RECT 33.775 182.075 34.065 182.120 ;
        RECT 26.490 181.920 26.630 182.075 ;
        RECT 37.900 182.060 38.220 182.120 ;
        RECT 43.420 182.260 43.740 182.320 ;
        RECT 49.490 182.260 49.630 182.415 ;
        RECT 43.420 182.120 49.630 182.260 ;
        RECT 49.860 182.260 50.180 182.320 ;
        RECT 51.330 182.260 51.470 182.415 ;
        RECT 59.060 182.400 59.380 182.460 ;
        RECT 59.995 182.600 60.285 182.645 ;
        RECT 60.440 182.600 60.760 182.660 ;
        RECT 59.995 182.460 60.760 182.600 ;
        RECT 59.995 182.415 60.285 182.460 ;
        RECT 60.440 182.400 60.760 182.460 ;
        RECT 67.800 182.400 68.120 182.660 ;
        RECT 68.810 182.645 68.950 183.140 ;
        RECT 71.020 183.080 71.340 183.140 ;
        RECT 71.480 183.280 71.800 183.340 ;
        RECT 72.400 183.280 72.720 183.340 ;
        RECT 73.780 183.280 74.100 183.340 ;
        RECT 89.435 183.280 89.725 183.325 ;
        RECT 71.480 183.140 76.310 183.280 ;
        RECT 71.480 183.080 71.800 183.140 ;
        RECT 72.400 183.080 72.720 183.140 ;
        RECT 73.780 183.080 74.100 183.140 ;
        RECT 73.320 182.740 73.640 183.000 ;
        RECT 68.735 182.415 69.025 182.645 ;
        RECT 70.575 182.600 70.865 182.645 ;
        RECT 71.480 182.600 71.800 182.660 ;
        RECT 70.575 182.460 71.800 182.600 ;
        RECT 70.575 182.415 70.865 182.460 ;
        RECT 49.860 182.120 51.470 182.260 ;
        RECT 43.420 182.060 43.740 182.120 ;
        RECT 49.860 182.060 50.180 182.120 ;
        RECT 67.355 182.075 67.645 182.305 ;
        RECT 68.275 182.260 68.565 182.305 ;
        RECT 70.650 182.260 70.790 182.415 ;
        RECT 71.480 182.400 71.800 182.460 ;
        RECT 71.955 182.415 72.245 182.645 ;
        RECT 68.275 182.120 70.790 182.260 ;
        RECT 72.030 182.260 72.170 182.415 ;
        RECT 72.400 182.400 72.720 182.660 ;
        RECT 73.410 182.600 73.550 182.740 ;
        RECT 74.715 182.600 75.005 182.645 ;
        RECT 73.410 182.460 75.005 182.600 ;
        RECT 74.715 182.415 75.005 182.460 ;
        RECT 72.030 182.120 72.630 182.260 ;
        RECT 68.275 182.075 68.565 182.120 ;
        RECT 30.555 181.920 30.845 181.965 ;
        RECT 26.490 181.780 30.845 181.920 ;
        RECT 67.430 181.920 67.570 182.075 ;
        RECT 72.490 181.980 72.630 182.120 ;
        RECT 73.320 182.060 73.640 182.320 ;
        RECT 74.790 182.260 74.930 182.415 ;
        RECT 75.620 182.400 75.940 182.660 ;
        RECT 76.170 182.645 76.310 183.140 ;
        RECT 86.290 183.140 89.725 183.280 ;
        RECT 80.795 182.940 81.085 182.985 ;
        RECT 84.035 182.940 84.685 182.985 ;
        RECT 86.290 182.940 86.430 183.140 ;
        RECT 89.435 183.095 89.725 183.140 ;
        RECT 97.240 183.080 97.560 183.340 ;
        RECT 105.520 183.280 105.840 183.340 ;
        RECT 105.995 183.280 106.285 183.325 ;
        RECT 105.520 183.140 106.285 183.280 ;
        RECT 105.520 183.080 105.840 183.140 ;
        RECT 105.995 183.095 106.285 183.140 ;
        RECT 111.515 183.095 111.805 183.325 ;
        RECT 80.795 182.800 86.430 182.940 ;
        RECT 104.155 182.940 104.445 182.985 ;
        RECT 111.590 182.940 111.730 183.095 ;
        RECT 104.155 182.800 111.730 182.940 ;
        RECT 117.135 182.940 117.425 182.985 ;
        RECT 120.375 182.940 121.025 182.985 ;
        RECT 117.135 182.800 121.025 182.940 ;
        RECT 80.795 182.755 81.385 182.800 ;
        RECT 84.035 182.755 84.685 182.800 ;
        RECT 104.155 182.755 104.445 182.800 ;
        RECT 76.095 182.415 76.385 182.645 ;
        RECT 76.540 182.400 76.860 182.660 ;
        RECT 81.095 182.440 81.385 182.755 ;
        RECT 105.610 182.660 105.750 182.800 ;
        RECT 117.135 182.755 117.725 182.800 ;
        RECT 120.375 182.755 121.025 182.800 ;
        RECT 123.015 182.940 123.305 182.985 ;
        RECT 124.380 182.940 124.700 183.000 ;
        RECT 123.015 182.800 124.700 182.940 ;
        RECT 123.015 182.755 123.305 182.800 ;
        RECT 117.435 182.660 117.725 182.755 ;
        RECT 124.380 182.740 124.700 182.800 ;
        RECT 82.175 182.600 82.465 182.645 ;
        RECT 85.755 182.600 86.045 182.645 ;
        RECT 87.590 182.600 87.880 182.645 ;
        RECT 82.175 182.460 87.880 182.600 ;
        RECT 82.175 182.415 82.465 182.460 ;
        RECT 85.755 182.415 86.045 182.460 ;
        RECT 87.590 182.415 87.880 182.460 ;
        RECT 89.895 182.600 90.185 182.645 ;
        RECT 90.800 182.600 91.120 182.660 ;
        RECT 89.895 182.460 91.120 182.600 ;
        RECT 89.895 182.415 90.185 182.460 ;
        RECT 90.800 182.400 91.120 182.460 ;
        RECT 95.860 182.600 96.180 182.660 ;
        RECT 96.795 182.600 97.085 182.645 ;
        RECT 95.860 182.460 97.085 182.600 ;
        RECT 95.860 182.400 96.180 182.460 ;
        RECT 96.795 182.415 97.085 182.460 ;
        RECT 99.080 182.600 99.400 182.660 ;
        RECT 103.695 182.600 103.985 182.645 ;
        RECT 99.080 182.460 103.985 182.600 ;
        RECT 99.080 182.400 99.400 182.460 ;
        RECT 103.695 182.415 103.985 182.460 ;
        RECT 105.520 182.400 105.840 182.660 ;
        RECT 105.980 182.600 106.300 182.660 ;
        RECT 105.980 182.460 107.590 182.600 ;
        RECT 105.980 182.400 106.300 182.460 ;
        RECT 77.015 182.260 77.305 182.305 ;
        RECT 74.790 182.120 77.305 182.260 ;
        RECT 77.015 182.075 77.305 182.120 ;
        RECT 86.675 182.260 86.965 182.305 ;
        RECT 88.055 182.260 88.345 182.305 ;
        RECT 93.560 182.260 93.880 182.320 ;
        RECT 86.675 182.120 87.810 182.260 ;
        RECT 86.675 182.075 86.965 182.120 ;
        RECT 72.400 181.920 72.720 181.980 ;
        RECT 75.620 181.920 75.940 181.980 ;
        RECT 67.430 181.780 75.940 181.920 ;
        RECT 30.555 181.735 30.845 181.780 ;
        RECT 72.400 181.720 72.720 181.780 ;
        RECT 75.620 181.720 75.940 181.780 ;
        RECT 82.175 181.920 82.465 181.965 ;
        RECT 85.295 181.920 85.585 181.965 ;
        RECT 87.185 181.920 87.475 181.965 ;
        RECT 82.175 181.780 87.475 181.920 ;
        RECT 87.670 181.920 87.810 182.120 ;
        RECT 88.055 182.120 93.880 182.260 ;
        RECT 88.055 182.075 88.345 182.120 ;
        RECT 93.560 182.060 93.880 182.120 ;
        RECT 96.335 182.260 96.625 182.305 ;
        RECT 97.700 182.260 98.020 182.320 ;
        RECT 102.775 182.260 103.065 182.305 ;
        RECT 96.335 182.120 103.065 182.260 ;
        RECT 96.335 182.075 96.625 182.120 ;
        RECT 89.420 181.920 89.740 181.980 ;
        RECT 87.670 181.780 89.740 181.920 ;
        RECT 82.175 181.735 82.465 181.780 ;
        RECT 85.295 181.735 85.585 181.780 ;
        RECT 87.185 181.735 87.475 181.780 ;
        RECT 89.420 181.720 89.740 181.780 ;
        RECT 39.280 181.580 39.600 181.640 ;
        RECT 40.675 181.580 40.965 181.625 ;
        RECT 39.280 181.440 40.965 181.580 ;
        RECT 39.280 181.380 39.600 181.440 ;
        RECT 40.675 181.395 40.965 181.440 ;
        RECT 45.720 181.580 46.040 181.640 ;
        RECT 47.100 181.580 47.420 181.640 ;
        RECT 48.035 181.580 48.325 181.625 ;
        RECT 45.720 181.440 48.325 181.580 ;
        RECT 45.720 181.380 46.040 181.440 ;
        RECT 47.100 181.380 47.420 181.440 ;
        RECT 48.035 181.395 48.325 181.440 ;
        RECT 55.840 181.580 56.160 181.640 ;
        RECT 59.535 181.580 59.825 181.625 ;
        RECT 55.840 181.440 59.825 181.580 ;
        RECT 55.840 181.380 56.160 181.440 ;
        RECT 59.535 181.395 59.825 181.440 ;
        RECT 66.435 181.580 66.725 181.625 ;
        RECT 69.180 181.580 69.500 181.640 ;
        RECT 66.435 181.440 69.500 181.580 ;
        RECT 66.435 181.395 66.725 181.440 ;
        RECT 69.180 181.380 69.500 181.440 ;
        RECT 74.700 181.580 75.020 181.640 ;
        RECT 77.935 181.580 78.225 181.625 ;
        RECT 74.700 181.440 78.225 181.580 ;
        RECT 74.700 181.380 75.020 181.440 ;
        RECT 77.935 181.395 78.225 181.440 ;
        RECT 79.300 181.380 79.620 181.640 ;
        RECT 84.820 181.580 85.140 181.640 ;
        RECT 96.410 181.580 96.550 182.075 ;
        RECT 97.700 182.060 98.020 182.120 ;
        RECT 102.775 182.075 103.065 182.120 ;
        RECT 104.140 182.260 104.460 182.320 ;
        RECT 106.455 182.260 106.745 182.305 ;
        RECT 104.140 182.120 106.745 182.260 ;
        RECT 107.450 182.260 107.590 182.460 ;
        RECT 107.820 182.400 108.140 182.660 ;
        RECT 108.295 182.415 108.585 182.645 ;
        RECT 108.755 182.415 109.045 182.645 ;
        RECT 109.200 182.600 109.520 182.660 ;
        RECT 109.675 182.600 109.965 182.645 ;
        RECT 109.200 182.460 109.965 182.600 ;
        RECT 108.370 182.260 108.510 182.415 ;
        RECT 107.450 182.120 108.510 182.260 ;
        RECT 104.140 182.060 104.460 182.120 ;
        RECT 106.455 182.075 106.745 182.120 ;
        RECT 98.160 181.920 98.480 181.980 ;
        RECT 108.830 181.920 108.970 182.415 ;
        RECT 109.200 182.400 109.520 182.460 ;
        RECT 109.675 182.415 109.965 182.460 ;
        RECT 111.500 182.600 111.820 182.660 ;
        RECT 111.975 182.600 112.265 182.645 ;
        RECT 111.500 182.460 112.265 182.600 ;
        RECT 111.500 182.400 111.820 182.460 ;
        RECT 111.975 182.415 112.265 182.460 ;
        RECT 117.435 182.440 117.800 182.660 ;
        RECT 117.480 182.400 117.800 182.440 ;
        RECT 118.515 182.600 118.805 182.645 ;
        RECT 122.095 182.600 122.385 182.645 ;
        RECT 123.930 182.600 124.220 182.645 ;
        RECT 118.515 182.460 124.220 182.600 ;
        RECT 118.515 182.415 118.805 182.460 ;
        RECT 122.095 182.415 122.385 182.460 ;
        RECT 123.930 182.415 124.220 182.460 ;
        RECT 110.580 182.060 110.900 182.320 ;
        RECT 117.940 182.260 118.260 182.320 ;
        RECT 124.395 182.260 124.685 182.305 ;
        RECT 117.940 182.120 124.685 182.260 ;
        RECT 117.940 182.060 118.260 182.120 ;
        RECT 124.395 182.075 124.685 182.120 ;
        RECT 98.160 181.780 108.970 181.920 ;
        RECT 110.120 181.920 110.440 181.980 ;
        RECT 115.655 181.920 115.945 181.965 ;
        RECT 110.120 181.780 115.945 181.920 ;
        RECT 98.160 181.720 98.480 181.780 ;
        RECT 110.120 181.720 110.440 181.780 ;
        RECT 115.655 181.735 115.945 181.780 ;
        RECT 118.515 181.920 118.805 181.965 ;
        RECT 121.635 181.920 121.925 181.965 ;
        RECT 123.525 181.920 123.815 181.965 ;
        RECT 118.515 181.780 123.815 181.920 ;
        RECT 118.515 181.735 118.805 181.780 ;
        RECT 121.635 181.735 121.925 181.780 ;
        RECT 123.525 181.735 123.815 181.780 ;
        RECT 84.820 181.440 96.550 181.580 ;
        RECT 99.095 181.580 99.385 181.625 ;
        RECT 104.600 181.580 104.920 181.640 ;
        RECT 99.095 181.440 104.920 181.580 ;
        RECT 84.820 181.380 85.140 181.440 ;
        RECT 99.095 181.395 99.385 181.440 ;
        RECT 104.600 181.380 104.920 181.440 ;
        RECT 113.815 181.580 114.105 181.625 ;
        RECT 116.560 181.580 116.880 181.640 ;
        RECT 113.815 181.440 116.880 181.580 ;
        RECT 113.815 181.395 114.105 181.440 ;
        RECT 116.560 181.380 116.880 181.440 ;
        RECT 14.370 180.760 127.530 181.240 ;
        RECT 45.260 180.560 45.580 180.620 ;
        RECT 46.640 180.560 46.960 180.620 ;
        RECT 45.260 180.420 46.960 180.560 ;
        RECT 45.260 180.360 45.580 180.420 ;
        RECT 46.640 180.360 46.960 180.420 ;
        RECT 49.415 180.560 49.705 180.605 ;
        RECT 49.860 180.560 50.180 180.620 ;
        RECT 82.060 180.560 82.380 180.620 ;
        RECT 49.415 180.420 50.180 180.560 ;
        RECT 49.415 180.375 49.705 180.420 ;
        RECT 49.860 180.360 50.180 180.420 ;
        RECT 78.470 180.420 82.380 180.560 ;
        RECT 25.445 180.220 25.735 180.265 ;
        RECT 27.335 180.220 27.625 180.265 ;
        RECT 30.455 180.220 30.745 180.265 ;
        RECT 25.445 180.080 30.745 180.220 ;
        RECT 25.445 180.035 25.735 180.080 ;
        RECT 27.335 180.035 27.625 180.080 ;
        RECT 30.455 180.035 30.745 180.080 ;
        RECT 53.555 180.220 53.845 180.265 ;
        RECT 56.300 180.220 56.620 180.280 ;
        RECT 53.555 180.080 56.620 180.220 ;
        RECT 53.555 180.035 53.845 180.080 ;
        RECT 56.300 180.020 56.620 180.080 ;
        RECT 67.340 180.220 67.660 180.280 ;
        RECT 78.470 180.220 78.610 180.420 ;
        RECT 82.060 180.360 82.380 180.420 ;
        RECT 89.420 180.360 89.740 180.620 ;
        RECT 105.520 180.360 105.840 180.620 ;
        RECT 117.480 180.560 117.800 180.620 ;
        RECT 122.555 180.560 122.845 180.605 ;
        RECT 124.380 180.560 124.700 180.620 ;
        RECT 117.480 180.420 119.550 180.560 ;
        RECT 117.480 180.360 117.800 180.420 ;
        RECT 67.340 180.080 78.610 180.220 ;
        RECT 78.840 180.220 79.160 180.280 ;
        RECT 85.280 180.220 85.600 180.280 ;
        RECT 78.840 180.080 85.600 180.220 ;
        RECT 67.340 180.020 67.660 180.080 ;
        RECT 78.840 180.020 79.160 180.080 ;
        RECT 85.280 180.020 85.600 180.080 ;
        RECT 95.055 180.220 95.345 180.265 ;
        RECT 98.175 180.220 98.465 180.265 ;
        RECT 100.065 180.220 100.355 180.265 ;
        RECT 95.055 180.080 100.355 180.220 ;
        RECT 95.055 180.035 95.345 180.080 ;
        RECT 98.175 180.035 98.465 180.080 ;
        RECT 100.065 180.035 100.355 180.080 ;
        RECT 113.915 180.220 114.205 180.265 ;
        RECT 117.035 180.220 117.325 180.265 ;
        RECT 118.925 180.220 119.215 180.265 ;
        RECT 113.915 180.080 119.215 180.220 ;
        RECT 119.410 180.220 119.550 180.420 ;
        RECT 122.555 180.420 124.700 180.560 ;
        RECT 122.555 180.375 122.845 180.420 ;
        RECT 124.380 180.360 124.700 180.420 ;
        RECT 120.715 180.220 121.005 180.265 ;
        RECT 119.410 180.080 121.005 180.220 ;
        RECT 113.915 180.035 114.205 180.080 ;
        RECT 117.035 180.035 117.325 180.080 ;
        RECT 118.925 180.035 119.215 180.080 ;
        RECT 120.715 180.035 121.005 180.080 ;
        RECT 33.315 179.695 33.605 179.925 ;
        RECT 46.180 179.880 46.500 179.940 ;
        RECT 44.430 179.740 46.500 179.880 ;
        RECT 24.575 179.355 24.865 179.585 ;
        RECT 25.040 179.540 25.330 179.585 ;
        RECT 26.875 179.540 27.165 179.585 ;
        RECT 30.455 179.540 30.745 179.585 ;
        RECT 25.040 179.400 30.745 179.540 ;
        RECT 25.040 179.355 25.330 179.400 ;
        RECT 26.875 179.355 27.165 179.400 ;
        RECT 30.455 179.355 30.745 179.400 ;
        RECT 24.650 179.200 24.790 179.355 ;
        RECT 24.650 179.060 25.250 179.200 ;
        RECT 25.110 178.860 25.250 179.060 ;
        RECT 25.940 179.000 26.260 179.260 ;
        RECT 27.320 179.200 27.640 179.260 ;
        RECT 31.535 179.245 31.825 179.560 ;
        RECT 33.390 179.540 33.530 179.695 ;
        RECT 36.980 179.540 37.300 179.600 ;
        RECT 33.390 179.400 37.300 179.540 ;
        RECT 36.980 179.340 37.300 179.400 ;
        RECT 39.295 179.355 39.585 179.585 ;
        RECT 39.755 179.355 40.045 179.585 ;
        RECT 40.215 179.540 40.505 179.585 ;
        RECT 40.660 179.540 40.980 179.600 ;
        RECT 40.215 179.400 40.980 179.540 ;
        RECT 40.215 179.355 40.505 179.400 ;
        RECT 28.235 179.200 28.885 179.245 ;
        RECT 31.535 179.200 32.125 179.245 ;
        RECT 27.320 179.060 32.125 179.200 ;
        RECT 27.320 179.000 27.640 179.060 ;
        RECT 28.235 179.015 28.885 179.060 ;
        RECT 31.835 179.015 32.125 179.060 ;
        RECT 33.760 179.000 34.080 179.260 ;
        RECT 34.680 179.200 35.000 179.260 ;
        RECT 37.915 179.200 38.205 179.245 ;
        RECT 34.680 179.060 38.205 179.200 ;
        RECT 34.680 179.000 35.000 179.060 ;
        RECT 37.915 179.015 38.205 179.060 ;
        RECT 36.520 178.860 36.840 178.920 ;
        RECT 25.110 178.720 36.840 178.860 ;
        RECT 39.370 178.860 39.510 179.355 ;
        RECT 39.830 179.200 39.970 179.355 ;
        RECT 40.660 179.340 40.980 179.400 ;
        RECT 41.135 179.355 41.425 179.585 ;
        RECT 43.435 179.355 43.725 179.585 ;
        RECT 39.830 179.060 40.430 179.200 ;
        RECT 40.290 178.920 40.430 179.060 ;
        RECT 39.740 178.860 40.060 178.920 ;
        RECT 39.370 178.720 40.060 178.860 ;
        RECT 36.520 178.660 36.840 178.720 ;
        RECT 39.740 178.660 40.060 178.720 ;
        RECT 40.200 178.660 40.520 178.920 ;
        RECT 40.660 178.860 40.980 178.920 ;
        RECT 41.210 178.860 41.350 179.355 ;
        RECT 40.660 178.720 41.350 178.860 ;
        RECT 40.660 178.660 40.980 178.720 ;
        RECT 42.040 178.660 42.360 178.920 ;
        RECT 43.510 178.860 43.650 179.355 ;
        RECT 43.880 179.340 44.200 179.600 ;
        RECT 44.430 179.585 44.570 179.740 ;
        RECT 46.180 179.680 46.500 179.740 ;
        RECT 46.640 179.680 46.960 179.940 ;
        RECT 47.100 179.680 47.420 179.940 ;
        RECT 50.795 179.880 51.085 179.925 ;
        RECT 52.160 179.880 52.480 179.940 ;
        RECT 50.795 179.740 52.480 179.880 ;
        RECT 50.795 179.695 51.085 179.740 ;
        RECT 52.160 179.680 52.480 179.740 ;
        RECT 54.000 179.880 54.320 179.940 ;
        RECT 58.615 179.880 58.905 179.925 ;
        RECT 60.455 179.880 60.745 179.925 ;
        RECT 54.000 179.740 60.745 179.880 ;
        RECT 54.000 179.680 54.320 179.740 ;
        RECT 58.615 179.695 58.905 179.740 ;
        RECT 60.455 179.695 60.745 179.740 ;
        RECT 72.400 179.680 72.720 179.940 ;
        RECT 72.860 179.680 73.180 179.940 ;
        RECT 73.335 179.880 73.625 179.925 ;
        RECT 75.620 179.880 75.940 179.940 ;
        RECT 73.335 179.740 75.940 179.880 ;
        RECT 73.335 179.695 73.625 179.740 ;
        RECT 75.620 179.680 75.940 179.740 ;
        RECT 76.555 179.880 76.845 179.925 ;
        RECT 79.300 179.880 79.620 179.940 ;
        RECT 84.820 179.880 85.140 179.940 ;
        RECT 85.755 179.880 86.045 179.925 ;
        RECT 76.555 179.740 80.910 179.880 ;
        RECT 76.555 179.695 76.845 179.740 ;
        RECT 79.300 179.680 79.620 179.740 ;
        RECT 44.355 179.355 44.645 179.585 ;
        RECT 45.260 179.340 45.580 179.600 ;
        RECT 65.500 179.340 65.820 179.600 ;
        RECT 68.260 179.340 68.580 179.600 ;
        RECT 71.020 179.540 71.340 179.600 ;
        RECT 71.495 179.540 71.785 179.585 ;
        RECT 71.020 179.400 71.785 179.540 ;
        RECT 71.020 179.340 71.340 179.400 ;
        RECT 71.495 179.355 71.785 179.400 ;
        RECT 73.780 179.340 74.100 179.600 ;
        RECT 76.080 179.540 76.400 179.600 ;
        RECT 80.770 179.585 80.910 179.740 ;
        RECT 84.820 179.740 86.045 179.880 ;
        RECT 84.820 179.680 85.140 179.740 ;
        RECT 85.755 179.695 86.045 179.740 ;
        RECT 104.600 179.680 104.920 179.940 ;
        RECT 105.520 179.880 105.840 179.940 ;
        RECT 107.820 179.880 108.140 179.940 ;
        RECT 111.055 179.880 111.345 179.925 ;
        RECT 115.640 179.880 115.960 179.940 ;
        RECT 105.520 179.740 108.140 179.880 ;
        RECT 105.520 179.680 105.840 179.740 ;
        RECT 107.820 179.680 108.140 179.740 ;
        RECT 108.830 179.740 111.345 179.880 ;
        RECT 108.830 179.600 108.970 179.740 ;
        RECT 111.055 179.695 111.345 179.740 ;
        RECT 111.590 179.740 120.470 179.880 ;
        RECT 79.775 179.540 80.065 179.585 ;
        RECT 76.080 179.400 80.065 179.540 ;
        RECT 76.080 179.340 76.400 179.400 ;
        RECT 53.540 179.200 53.860 179.260 ;
        RECT 58.155 179.200 58.445 179.245 ;
        RECT 53.540 179.060 58.445 179.200 ;
        RECT 53.540 179.000 53.860 179.060 ;
        RECT 58.155 179.015 58.445 179.060 ;
        RECT 61.835 179.200 62.125 179.245 ;
        RECT 69.195 179.200 69.485 179.245 ;
        RECT 72.860 179.200 73.180 179.260 ;
        RECT 61.835 179.060 73.180 179.200 ;
        RECT 61.835 179.015 62.125 179.060 ;
        RECT 69.195 179.015 69.485 179.060 ;
        RECT 72.860 179.000 73.180 179.060 ;
        RECT 44.340 178.860 44.660 178.920 ;
        RECT 43.510 178.720 44.660 178.860 ;
        RECT 44.340 178.660 44.660 178.720 ;
        RECT 45.720 178.860 46.040 178.920 ;
        RECT 47.575 178.860 47.865 178.905 ;
        RECT 45.720 178.720 47.865 178.860 ;
        RECT 45.720 178.660 46.040 178.720 ;
        RECT 47.575 178.675 47.865 178.720 ;
        RECT 50.320 178.860 50.640 178.920 ;
        RECT 55.855 178.860 56.145 178.905 ;
        RECT 50.320 178.720 56.145 178.860 ;
        RECT 50.320 178.660 50.640 178.720 ;
        RECT 55.855 178.675 56.145 178.720 ;
        RECT 57.680 178.660 58.000 178.920 ;
        RECT 65.960 178.660 66.280 178.920 ;
        RECT 70.575 178.860 70.865 178.905 ;
        RECT 78.380 178.860 78.700 178.920 ;
        RECT 70.575 178.720 78.700 178.860 ;
        RECT 78.930 178.860 79.070 179.400 ;
        RECT 79.775 179.355 80.065 179.400 ;
        RECT 80.695 179.355 80.985 179.585 ;
        RECT 81.140 179.340 81.460 179.600 ;
        RECT 81.600 179.340 81.920 179.600 ;
        RECT 90.340 179.340 90.660 179.600 ;
        RECT 90.800 179.340 91.120 179.600 ;
        RECT 79.315 179.200 79.605 179.245 ;
        RECT 86.200 179.200 86.520 179.260 ;
        RECT 93.975 179.245 94.265 179.560 ;
        RECT 95.055 179.540 95.345 179.585 ;
        RECT 98.635 179.540 98.925 179.585 ;
        RECT 100.470 179.540 100.760 179.585 ;
        RECT 95.055 179.400 100.760 179.540 ;
        RECT 95.055 179.355 95.345 179.400 ;
        RECT 98.635 179.355 98.925 179.400 ;
        RECT 100.470 179.355 100.760 179.400 ;
        RECT 100.935 179.355 101.225 179.585 ;
        RECT 86.675 179.200 86.965 179.245 ;
        RECT 91.275 179.200 91.565 179.245 ;
        RECT 93.675 179.200 94.265 179.245 ;
        RECT 96.915 179.200 97.565 179.245 ;
        RECT 79.315 179.060 86.965 179.200 ;
        RECT 79.315 179.015 79.605 179.060 ;
        RECT 86.200 179.000 86.520 179.060 ;
        RECT 86.675 179.015 86.965 179.060 ;
        RECT 87.210 179.060 90.110 179.200 ;
        RECT 87.210 178.920 87.350 179.060 ;
        RECT 82.520 178.860 82.840 178.920 ;
        RECT 78.930 178.720 82.840 178.860 ;
        RECT 70.575 178.675 70.865 178.720 ;
        RECT 78.380 178.660 78.700 178.720 ;
        RECT 82.520 178.660 82.840 178.720 ;
        RECT 82.995 178.860 83.285 178.905 ;
        RECT 83.440 178.860 83.760 178.920 ;
        RECT 82.995 178.720 83.760 178.860 ;
        RECT 82.995 178.675 83.285 178.720 ;
        RECT 83.440 178.660 83.760 178.720 ;
        RECT 87.120 178.660 87.440 178.920 ;
        RECT 88.960 178.660 89.280 178.920 ;
        RECT 89.970 178.860 90.110 179.060 ;
        RECT 91.275 179.060 97.565 179.200 ;
        RECT 91.275 179.015 91.565 179.060 ;
        RECT 93.675 179.015 93.965 179.060 ;
        RECT 96.915 179.015 97.565 179.060 ;
        RECT 99.540 179.000 99.860 179.260 ;
        RECT 92.195 178.860 92.485 178.905 ;
        RECT 95.860 178.860 96.180 178.920 ;
        RECT 89.970 178.720 96.180 178.860 ;
        RECT 101.010 178.860 101.150 179.355 ;
        RECT 108.740 179.340 109.060 179.600 ;
        RECT 109.675 179.540 109.965 179.585 ;
        RECT 111.590 179.540 111.730 179.740 ;
        RECT 115.640 179.680 115.960 179.740 ;
        RECT 120.330 179.585 120.470 179.740 ;
        RECT 109.675 179.400 111.730 179.540 ;
        RECT 109.675 179.355 109.965 179.400 ;
        RECT 101.840 179.000 102.160 179.260 ;
        RECT 112.835 179.245 113.125 179.560 ;
        RECT 113.915 179.540 114.205 179.585 ;
        RECT 117.495 179.540 117.785 179.585 ;
        RECT 119.330 179.540 119.620 179.585 ;
        RECT 113.915 179.400 119.620 179.540 ;
        RECT 113.915 179.355 114.205 179.400 ;
        RECT 117.495 179.355 117.785 179.400 ;
        RECT 119.330 179.355 119.620 179.400 ;
        RECT 119.795 179.355 120.085 179.585 ;
        RECT 120.255 179.355 120.545 179.585 ;
        RECT 110.135 179.200 110.425 179.245 ;
        RECT 112.535 179.200 113.125 179.245 ;
        RECT 115.775 179.200 116.425 179.245 ;
        RECT 110.135 179.060 116.425 179.200 ;
        RECT 110.135 179.015 110.425 179.060 ;
        RECT 112.535 179.015 112.825 179.060 ;
        RECT 115.775 179.015 116.425 179.060 ;
        RECT 118.400 179.000 118.720 179.260 ;
        RECT 117.940 178.860 118.260 178.920 ;
        RECT 119.870 178.860 120.010 179.355 ;
        RECT 121.620 179.340 121.940 179.600 ;
        RECT 101.010 178.720 120.010 178.860 ;
        RECT 92.195 178.675 92.485 178.720 ;
        RECT 95.860 178.660 96.180 178.720 ;
        RECT 117.940 178.660 118.260 178.720 ;
        RECT 14.370 178.040 127.530 178.520 ;
        RECT 25.495 177.840 25.785 177.885 ;
        RECT 27.320 177.840 27.640 177.900 ;
        RECT 25.495 177.700 27.640 177.840 ;
        RECT 25.495 177.655 25.785 177.700 ;
        RECT 27.320 177.640 27.640 177.700 ;
        RECT 39.280 177.640 39.600 177.900 ;
        RECT 45.720 177.640 46.040 177.900 ;
        RECT 53.540 177.840 53.860 177.900 ;
        RECT 61.820 177.840 62.140 177.900 ;
        RECT 63.215 177.840 63.505 177.885 ;
        RECT 71.480 177.840 71.800 177.900 ;
        RECT 71.955 177.840 72.245 177.885 ;
        RECT 46.270 177.700 53.860 177.840 ;
        RECT 26.875 177.500 27.165 177.545 ;
        RECT 29.275 177.500 29.565 177.545 ;
        RECT 32.515 177.500 33.165 177.545 ;
        RECT 46.270 177.500 46.410 177.700 ;
        RECT 53.540 177.640 53.860 177.700 ;
        RECT 54.550 177.700 61.590 177.840 ;
        RECT 52.160 177.500 52.480 177.560 ;
        RECT 26.875 177.360 33.165 177.500 ;
        RECT 26.875 177.315 27.165 177.360 ;
        RECT 29.275 177.315 29.865 177.360 ;
        RECT 32.515 177.315 33.165 177.360 ;
        RECT 43.050 177.360 46.410 177.500 ;
        RECT 47.190 177.360 52.480 177.500 ;
        RECT 25.955 177.160 26.245 177.205 ;
        RECT 26.415 177.160 26.705 177.205 ;
        RECT 25.955 177.020 26.705 177.160 ;
        RECT 25.955 176.975 26.245 177.020 ;
        RECT 26.415 176.975 26.705 177.020 ;
        RECT 29.575 177.000 29.865 177.315 ;
        RECT 43.050 177.205 43.190 177.360 ;
        RECT 30.655 177.160 30.945 177.205 ;
        RECT 34.235 177.160 34.525 177.205 ;
        RECT 36.070 177.160 36.360 177.205 ;
        RECT 30.655 177.020 36.360 177.160 ;
        RECT 30.655 176.975 30.945 177.020 ;
        RECT 34.235 176.975 34.525 177.020 ;
        RECT 36.070 176.975 36.360 177.020 ;
        RECT 42.975 177.160 43.265 177.205 ;
        RECT 43.420 177.160 43.740 177.220 ;
        RECT 42.975 177.020 43.740 177.160 ;
        RECT 42.975 176.975 43.265 177.020 ;
        RECT 26.490 176.820 26.630 176.975 ;
        RECT 43.420 176.960 43.740 177.020 ;
        RECT 45.260 177.160 45.580 177.220 ;
        RECT 47.190 177.205 47.330 177.360 ;
        RECT 52.160 177.300 52.480 177.360 ;
        RECT 46.195 177.160 46.485 177.205 ;
        RECT 45.260 177.020 46.485 177.160 ;
        RECT 45.260 176.960 45.580 177.020 ;
        RECT 46.195 176.975 46.485 177.020 ;
        RECT 47.115 176.975 47.405 177.205 ;
        RECT 30.080 176.820 30.400 176.880 ;
        RECT 26.490 176.680 30.400 176.820 ;
        RECT 30.080 176.620 30.400 176.680 ;
        RECT 35.140 176.620 35.460 176.880 ;
        RECT 36.520 176.620 36.840 176.880 ;
        RECT 37.900 176.620 38.220 176.880 ;
        RECT 38.835 176.635 39.125 176.865 ;
        RECT 30.655 176.480 30.945 176.525 ;
        RECT 33.775 176.480 34.065 176.525 ;
        RECT 35.665 176.480 35.955 176.525 ;
        RECT 30.655 176.340 35.955 176.480 ;
        RECT 30.655 176.295 30.945 176.340 ;
        RECT 33.775 176.295 34.065 176.340 ;
        RECT 35.665 176.295 35.955 176.340 ;
        RECT 27.780 175.940 28.100 176.200 ;
        RECT 34.220 176.140 34.540 176.200 ;
        RECT 38.910 176.140 39.050 176.635 ;
        RECT 46.270 176.480 46.410 176.975 ;
        RECT 47.560 176.960 47.880 177.220 ;
        RECT 48.035 177.160 48.325 177.205 ;
        RECT 48.940 177.160 49.260 177.220 ;
        RECT 48.035 177.020 49.260 177.160 ;
        RECT 48.035 176.975 48.325 177.020 ;
        RECT 48.940 176.960 49.260 177.020 ;
        RECT 50.320 176.960 50.640 177.220 ;
        RECT 49.030 176.820 49.170 176.960 ;
        RECT 54.550 176.820 54.690 177.700 ;
        RECT 55.035 177.500 55.325 177.545 ;
        RECT 55.840 177.500 56.160 177.560 ;
        RECT 58.275 177.500 58.925 177.545 ;
        RECT 55.035 177.360 58.925 177.500 ;
        RECT 55.035 177.315 55.625 177.360 ;
        RECT 55.335 177.000 55.625 177.315 ;
        RECT 55.840 177.300 56.160 177.360 ;
        RECT 58.275 177.315 58.925 177.360 ;
        RECT 60.900 177.300 61.220 177.560 ;
        RECT 61.450 177.500 61.590 177.700 ;
        RECT 61.820 177.700 63.505 177.840 ;
        RECT 61.820 177.640 62.140 177.700 ;
        RECT 63.215 177.655 63.505 177.700 ;
        RECT 70.190 177.700 72.245 177.840 ;
        RECT 70.190 177.500 70.330 177.700 ;
        RECT 71.480 177.640 71.800 177.700 ;
        RECT 71.955 177.655 72.245 177.700 ;
        RECT 72.860 177.640 73.180 177.900 ;
        RECT 81.600 177.840 81.920 177.900 ;
        RECT 81.230 177.700 81.920 177.840 ;
        RECT 61.450 177.360 70.330 177.500 ;
        RECT 79.300 177.500 79.620 177.560 ;
        RECT 79.775 177.500 80.065 177.545 ;
        RECT 81.230 177.500 81.370 177.700 ;
        RECT 81.600 177.640 81.920 177.700 ;
        RECT 82.060 177.840 82.380 177.900 ;
        RECT 88.055 177.840 88.345 177.885 ;
        RECT 90.340 177.840 90.660 177.900 ;
        RECT 82.060 177.700 87.810 177.840 ;
        RECT 82.060 177.640 82.380 177.700 ;
        RECT 85.740 177.500 86.060 177.560 ;
        RECT 79.300 177.360 80.065 177.500 ;
        RECT 79.300 177.300 79.620 177.360 ;
        RECT 79.775 177.315 80.065 177.360 ;
        RECT 80.310 177.360 81.370 177.500 ;
        RECT 56.415 177.160 56.705 177.205 ;
        RECT 59.995 177.160 60.285 177.205 ;
        RECT 61.830 177.160 62.120 177.205 ;
        RECT 56.415 177.020 62.120 177.160 ;
        RECT 56.415 176.975 56.705 177.020 ;
        RECT 59.995 176.975 60.285 177.020 ;
        RECT 61.830 176.975 62.120 177.020 ;
        RECT 64.135 176.975 64.425 177.205 ;
        RECT 49.030 176.680 54.690 176.820 ;
        RECT 59.060 176.820 59.380 176.880 ;
        RECT 62.295 176.820 62.585 176.865 ;
        RECT 63.660 176.820 63.980 176.880 ;
        RECT 59.060 176.680 63.980 176.820 ;
        RECT 59.060 176.620 59.380 176.680 ;
        RECT 62.295 176.635 62.585 176.680 ;
        RECT 63.660 176.620 63.980 176.680 ;
        RECT 50.780 176.480 51.100 176.540 ;
        RECT 46.270 176.340 51.100 176.480 ;
        RECT 50.780 176.280 51.100 176.340 ;
        RECT 56.415 176.480 56.705 176.525 ;
        RECT 59.535 176.480 59.825 176.525 ;
        RECT 61.425 176.480 61.715 176.525 ;
        RECT 56.415 176.340 61.715 176.480 ;
        RECT 56.415 176.295 56.705 176.340 ;
        RECT 59.535 176.295 59.825 176.340 ;
        RECT 61.425 176.295 61.715 176.340 ;
        RECT 34.220 176.000 39.050 176.140 ;
        RECT 41.135 176.140 41.425 176.185 ;
        RECT 42.500 176.140 42.820 176.200 ;
        RECT 41.135 176.000 42.820 176.140 ;
        RECT 34.220 175.940 34.540 176.000 ;
        RECT 41.135 175.955 41.425 176.000 ;
        RECT 42.500 175.940 42.820 176.000 ;
        RECT 49.415 176.140 49.705 176.185 ;
        RECT 49.860 176.140 50.180 176.200 ;
        RECT 49.415 176.000 50.180 176.140 ;
        RECT 49.415 175.955 49.705 176.000 ;
        RECT 49.860 175.940 50.180 176.000 ;
        RECT 53.095 176.140 53.385 176.185 ;
        RECT 64.210 176.140 64.350 176.975 ;
        RECT 68.720 176.960 69.040 177.220 ;
        RECT 69.180 177.160 69.500 177.220 ;
        RECT 71.070 177.160 71.360 177.205 ;
        RECT 72.400 177.160 72.720 177.220 ;
        RECT 73.335 177.160 73.625 177.205 ;
        RECT 69.180 177.020 72.170 177.160 ;
        RECT 69.180 176.960 69.500 177.020 ;
        RECT 71.070 176.975 71.360 177.020 ;
        RECT 72.030 176.820 72.170 177.020 ;
        RECT 72.400 177.020 73.625 177.160 ;
        RECT 72.400 176.960 72.720 177.020 ;
        RECT 73.335 176.975 73.625 177.020 ;
        RECT 73.780 176.960 74.100 177.220 ;
        RECT 74.700 176.960 75.020 177.220 ;
        RECT 75.175 176.975 75.465 177.205 ;
        RECT 75.250 176.820 75.390 176.975 ;
        RECT 76.080 176.960 76.400 177.220 ;
        RECT 77.015 176.975 77.305 177.205 ;
        RECT 72.030 176.680 75.390 176.820 ;
        RECT 77.090 176.820 77.230 176.975 ;
        RECT 77.460 176.960 77.780 177.220 ;
        RECT 77.920 177.160 78.240 177.220 ;
        RECT 80.310 177.160 80.450 177.360 ;
        RECT 81.230 177.205 81.370 177.360 ;
        RECT 82.150 177.360 86.060 177.500 ;
        RECT 87.670 177.500 87.810 177.700 ;
        RECT 88.055 177.700 90.660 177.840 ;
        RECT 88.055 177.655 88.345 177.700 ;
        RECT 90.340 177.640 90.660 177.700 ;
        RECT 99.540 177.840 99.860 177.900 ;
        RECT 101.855 177.840 102.145 177.885 ;
        RECT 99.540 177.700 102.145 177.840 ;
        RECT 99.540 177.640 99.860 177.700 ;
        RECT 101.855 177.655 102.145 177.700 ;
        RECT 111.500 177.640 111.820 177.900 ;
        RECT 111.960 177.640 112.280 177.900 ;
        RECT 113.815 177.655 114.105 177.885 ;
        RECT 117.495 177.840 117.785 177.885 ;
        RECT 118.400 177.840 118.720 177.900 ;
        RECT 117.495 177.700 118.720 177.840 ;
        RECT 117.495 177.655 117.785 177.700 ;
        RECT 108.740 177.500 109.060 177.560 ;
        RECT 87.670 177.360 106.670 177.500 ;
        RECT 77.920 177.020 80.450 177.160 ;
        RECT 77.920 176.960 78.240 177.020 ;
        RECT 81.155 176.975 81.445 177.205 ;
        RECT 81.600 176.960 81.920 177.220 ;
        RECT 82.150 177.205 82.290 177.360 ;
        RECT 85.740 177.300 86.060 177.360 ;
        RECT 82.075 176.975 82.365 177.205 ;
        RECT 82.520 177.160 82.840 177.220 ;
        RECT 82.995 177.160 83.285 177.205 ;
        RECT 83.900 177.160 84.220 177.220 ;
        RECT 82.520 177.020 84.220 177.160 ;
        RECT 82.520 176.960 82.840 177.020 ;
        RECT 82.995 176.975 83.285 177.020 ;
        RECT 83.900 176.960 84.220 177.020 ;
        RECT 85.295 177.160 85.585 177.205 ;
        RECT 88.960 177.160 89.280 177.220 ;
        RECT 85.295 177.020 89.280 177.160 ;
        RECT 85.295 176.975 85.585 177.020 ;
        RECT 88.960 176.960 89.280 177.020 ;
        RECT 98.160 176.960 98.480 177.220 ;
        RECT 99.080 176.960 99.400 177.220 ;
        RECT 99.630 177.205 99.770 177.360 ;
        RECT 106.530 177.220 106.670 177.360 ;
        RECT 106.990 177.360 109.060 177.500 ;
        RECT 113.890 177.500 114.030 177.655 ;
        RECT 118.400 177.640 118.720 177.700 ;
        RECT 121.620 177.500 121.940 177.560 ;
        RECT 113.890 177.360 121.940 177.500 ;
        RECT 99.555 176.975 99.845 177.205 ;
        RECT 100.015 176.975 100.305 177.205 ;
        RECT 101.840 177.160 102.160 177.220 ;
        RECT 102.775 177.160 103.065 177.205 ;
        RECT 101.840 177.020 103.065 177.160 ;
        RECT 78.840 176.820 79.160 176.880 ;
        RECT 77.090 176.680 79.160 176.820 ;
        RECT 78.840 176.620 79.160 176.680 ;
        RECT 79.315 176.820 79.605 176.865 ;
        RECT 80.220 176.820 80.540 176.880 ;
        RECT 100.090 176.820 100.230 176.975 ;
        RECT 101.840 176.960 102.160 177.020 ;
        RECT 102.775 176.975 103.065 177.020 ;
        RECT 105.995 176.975 106.285 177.205 ;
        RECT 105.520 176.820 105.840 176.880 ;
        RECT 106.070 176.820 106.210 176.975 ;
        RECT 106.440 176.960 106.760 177.220 ;
        RECT 106.990 177.205 107.130 177.360 ;
        RECT 108.740 177.300 109.060 177.360 ;
        RECT 121.620 177.300 121.940 177.360 ;
        RECT 106.915 176.975 107.205 177.205 ;
        RECT 107.820 177.160 108.140 177.220 ;
        RECT 109.200 177.160 109.520 177.220 ;
        RECT 107.820 177.020 109.520 177.160 ;
        RECT 107.820 176.960 108.140 177.020 ;
        RECT 109.200 176.960 109.520 177.020 ;
        RECT 116.560 176.960 116.880 177.220 ;
        RECT 79.315 176.680 80.540 176.820 ;
        RECT 79.315 176.635 79.605 176.680 ;
        RECT 80.220 176.620 80.540 176.680 ;
        RECT 84.680 176.680 106.210 176.820 ;
        RECT 65.040 176.480 65.360 176.540 ;
        RECT 70.115 176.480 70.405 176.525 ;
        RECT 84.680 176.480 84.820 176.680 ;
        RECT 105.520 176.620 105.840 176.680 ;
        RECT 110.580 176.620 110.900 176.880 ;
        RECT 65.040 176.340 84.820 176.480 ;
        RECT 65.040 176.280 65.360 176.340 ;
        RECT 70.115 176.295 70.405 176.340 ;
        RECT 53.095 176.000 64.350 176.140 ;
        RECT 64.580 176.140 64.900 176.200 ;
        RECT 67.800 176.140 68.120 176.200 ;
        RECT 64.580 176.000 68.120 176.140 ;
        RECT 53.095 175.955 53.385 176.000 ;
        RECT 64.580 175.940 64.900 176.000 ;
        RECT 67.800 175.940 68.120 176.000 ;
        RECT 68.720 176.140 69.040 176.200 ;
        RECT 74.700 176.140 75.020 176.200 ;
        RECT 68.720 176.000 75.020 176.140 ;
        RECT 68.720 175.940 69.040 176.000 ;
        RECT 74.700 175.940 75.020 176.000 ;
        RECT 100.460 176.140 100.780 176.200 ;
        RECT 101.395 176.140 101.685 176.185 ;
        RECT 100.460 176.000 101.685 176.140 ;
        RECT 100.460 175.940 100.780 176.000 ;
        RECT 101.395 175.955 101.685 176.000 ;
        RECT 101.840 176.140 102.160 176.200 ;
        RECT 104.615 176.140 104.905 176.185 ;
        RECT 101.840 176.000 104.905 176.140 ;
        RECT 101.840 175.940 102.160 176.000 ;
        RECT 104.615 175.955 104.905 176.000 ;
        RECT 14.370 175.320 127.530 175.800 ;
        RECT 25.495 175.120 25.785 175.165 ;
        RECT 25.940 175.120 26.260 175.180 ;
        RECT 37.900 175.120 38.220 175.180 ;
        RECT 40.660 175.120 40.980 175.180 ;
        RECT 25.495 174.980 26.260 175.120 ;
        RECT 25.495 174.935 25.785 174.980 ;
        RECT 25.940 174.920 26.260 174.980 ;
        RECT 33.850 174.980 38.220 175.120 ;
        RECT 30.555 174.780 30.845 174.825 ;
        RECT 26.490 174.640 30.845 174.780 ;
        RECT 26.490 174.145 26.630 174.640 ;
        RECT 30.555 174.595 30.845 174.640 ;
        RECT 33.850 174.485 33.990 174.980 ;
        RECT 37.900 174.920 38.220 174.980 ;
        RECT 38.450 174.980 40.980 175.120 ;
        RECT 38.450 174.780 38.590 174.980 ;
        RECT 40.660 174.920 40.980 174.980 ;
        RECT 46.180 175.120 46.500 175.180 ;
        RECT 54.000 175.120 54.320 175.180 ;
        RECT 46.180 174.980 54.320 175.120 ;
        RECT 46.180 174.920 46.500 174.980 ;
        RECT 54.000 174.920 54.320 174.980 ;
        RECT 63.660 175.120 63.980 175.180 ;
        RECT 65.960 175.120 66.280 175.180 ;
        RECT 63.660 174.980 66.280 175.120 ;
        RECT 63.660 174.920 63.980 174.980 ;
        RECT 65.960 174.920 66.280 174.980 ;
        RECT 67.800 175.120 68.120 175.180 ;
        RECT 77.460 175.120 77.780 175.180 ;
        RECT 81.600 175.120 81.920 175.180 ;
        RECT 105.980 175.120 106.300 175.180 ;
        RECT 107.820 175.120 108.140 175.180 ;
        RECT 67.800 174.980 81.920 175.120 ;
        RECT 67.800 174.920 68.120 174.980 ;
        RECT 77.460 174.920 77.780 174.980 ;
        RECT 81.600 174.920 81.920 174.980 ;
        RECT 103.770 174.980 110.350 175.120 ;
        RECT 36.610 174.640 38.590 174.780 ;
        RECT 38.835 174.780 39.125 174.825 ;
        RECT 40.200 174.780 40.520 174.840 ;
        RECT 57.235 174.780 57.525 174.825 ;
        RECT 38.835 174.640 40.520 174.780 ;
        RECT 33.775 174.255 34.065 174.485 ;
        RECT 36.610 174.440 36.750 174.640 ;
        RECT 38.835 174.595 39.125 174.640 ;
        RECT 40.200 174.580 40.520 174.640 ;
        RECT 53.630 174.640 57.525 174.780 ;
        RECT 53.630 174.500 53.770 174.640 ;
        RECT 57.235 174.595 57.525 174.640 ;
        RECT 60.095 174.780 60.385 174.825 ;
        RECT 63.215 174.780 63.505 174.825 ;
        RECT 65.105 174.780 65.395 174.825 ;
        RECT 71.495 174.780 71.785 174.825 ;
        RECT 76.080 174.780 76.400 174.840 ;
        RECT 60.095 174.640 65.395 174.780 ;
        RECT 60.095 174.595 60.385 174.640 ;
        RECT 63.215 174.595 63.505 174.640 ;
        RECT 65.105 174.595 65.395 174.640 ;
        RECT 69.270 174.640 76.400 174.780 ;
        RECT 35.230 174.300 36.750 174.440 ;
        RECT 37.440 174.440 37.760 174.500 ;
        RECT 45.260 174.440 45.580 174.500 ;
        RECT 37.440 174.300 41.350 174.440 ;
        RECT 26.415 173.915 26.705 174.145 ;
        RECT 26.875 173.915 27.165 174.145 ;
        RECT 30.095 174.100 30.385 174.145 ;
        RECT 32.395 174.100 32.685 174.145 ;
        RECT 34.220 174.100 34.540 174.160 ;
        RECT 35.230 174.145 35.370 174.300 ;
        RECT 37.440 174.240 37.760 174.300 ;
        RECT 30.095 173.960 34.540 174.100 ;
        RECT 30.095 173.915 30.385 173.960 ;
        RECT 32.395 173.915 32.685 173.960 ;
        RECT 26.950 173.760 27.090 173.915 ;
        RECT 34.220 173.900 34.540 173.960 ;
        RECT 35.155 173.915 35.445 174.145 ;
        RECT 36.075 173.915 36.365 174.145 ;
        RECT 36.535 173.915 36.825 174.145 ;
        RECT 36.995 174.100 37.285 174.145 ;
        RECT 37.900 174.100 38.220 174.160 ;
        RECT 39.740 174.100 40.060 174.160 ;
        RECT 41.210 174.145 41.350 174.300 ;
        RECT 42.590 174.300 45.580 174.440 ;
        RECT 42.590 174.145 42.730 174.300 ;
        RECT 45.260 174.240 45.580 174.300 ;
        RECT 46.655 174.440 46.945 174.485 ;
        RECT 53.540 174.440 53.860 174.500 ;
        RECT 46.655 174.300 53.860 174.440 ;
        RECT 46.655 174.255 46.945 174.300 ;
        RECT 53.540 174.240 53.860 174.300 ;
        RECT 54.000 174.240 54.320 174.500 ;
        RECT 57.680 174.440 58.000 174.500 ;
        RECT 64.580 174.440 64.900 174.500 ;
        RECT 54.550 174.300 58.000 174.440 ;
        RECT 40.215 174.100 40.505 174.145 ;
        RECT 36.995 173.960 40.505 174.100 ;
        RECT 36.995 173.915 37.285 173.960 ;
        RECT 27.780 173.760 28.100 173.820 ;
        RECT 32.855 173.760 33.145 173.805 ;
        RECT 33.760 173.760 34.080 173.820 ;
        RECT 36.150 173.760 36.290 173.915 ;
        RECT 26.950 173.620 32.610 173.760 ;
        RECT 27.780 173.560 28.100 173.620 ;
        RECT 32.470 173.420 32.610 173.620 ;
        RECT 32.855 173.620 34.080 173.760 ;
        RECT 32.855 173.575 33.145 173.620 ;
        RECT 33.760 173.560 34.080 173.620 ;
        RECT 34.310 173.620 36.290 173.760 ;
        RECT 34.310 173.420 34.450 173.620 ;
        RECT 32.470 173.280 34.450 173.420 ;
        RECT 36.610 173.420 36.750 173.915 ;
        RECT 37.900 173.900 38.220 173.960 ;
        RECT 39.740 173.900 40.060 173.960 ;
        RECT 40.215 173.915 40.505 173.960 ;
        RECT 40.675 173.915 40.965 174.145 ;
        RECT 41.135 173.915 41.425 174.145 ;
        RECT 42.055 174.100 42.345 174.145 ;
        RECT 42.515 174.100 42.805 174.145 ;
        RECT 42.055 173.960 42.805 174.100 ;
        RECT 42.055 173.915 42.345 173.960 ;
        RECT 42.515 173.915 42.805 173.960 ;
        RECT 38.375 173.760 38.665 173.805 ;
        RECT 38.820 173.760 39.140 173.820 ;
        RECT 38.375 173.620 39.140 173.760 ;
        RECT 38.375 173.575 38.665 173.620 ;
        RECT 38.820 173.560 39.140 173.620 ;
        RECT 39.280 173.760 39.600 173.820 ;
        RECT 40.750 173.760 40.890 173.915 ;
        RECT 43.420 173.900 43.740 174.160 ;
        RECT 43.880 173.900 44.200 174.160 ;
        RECT 44.340 173.900 44.660 174.160 ;
        RECT 54.550 174.145 54.690 174.300 ;
        RECT 57.680 174.240 58.000 174.300 ;
        RECT 58.230 174.300 64.900 174.440 ;
        RECT 49.415 174.100 49.705 174.145 ;
        RECT 54.475 174.100 54.765 174.145 ;
        RECT 49.415 173.960 54.765 174.100 ;
        RECT 49.415 173.915 49.705 173.960 ;
        RECT 54.475 173.915 54.765 173.960 ;
        RECT 54.935 174.100 55.225 174.145 ;
        RECT 56.300 174.100 56.620 174.160 ;
        RECT 54.935 173.960 56.620 174.100 ;
        RECT 54.935 173.915 55.225 173.960 ;
        RECT 56.300 173.900 56.620 173.960 ;
        RECT 41.580 173.760 41.900 173.820 ;
        RECT 39.280 173.620 41.900 173.760 ;
        RECT 39.280 173.560 39.600 173.620 ;
        RECT 41.580 173.560 41.900 173.620 ;
        RECT 39.370 173.420 39.510 173.560 ;
        RECT 36.610 173.280 39.510 173.420 ;
        RECT 43.970 173.420 44.110 173.900 ;
        RECT 45.260 173.760 45.580 173.820 ;
        RECT 45.735 173.760 46.025 173.805 ;
        RECT 45.260 173.620 46.025 173.760 ;
        RECT 45.260 173.560 45.580 173.620 ;
        RECT 45.735 173.575 46.025 173.620 ;
        RECT 47.560 173.760 47.880 173.820 ;
        RECT 53.080 173.760 53.400 173.820 ;
        RECT 58.230 173.760 58.370 174.300 ;
        RECT 64.580 174.240 64.900 174.300 ;
        RECT 65.960 174.240 66.280 174.500 ;
        RECT 59.015 173.805 59.305 174.120 ;
        RECT 60.095 174.100 60.385 174.145 ;
        RECT 63.675 174.100 63.965 174.145 ;
        RECT 65.510 174.100 65.800 174.145 ;
        RECT 60.095 173.960 65.800 174.100 ;
        RECT 60.095 173.915 60.385 173.960 ;
        RECT 63.675 173.915 63.965 173.960 ;
        RECT 65.510 173.915 65.800 173.960 ;
        RECT 68.275 174.100 68.565 174.145 ;
        RECT 68.720 174.100 69.040 174.160 ;
        RECT 68.275 173.960 69.040 174.100 ;
        RECT 68.275 173.915 68.565 173.960 ;
        RECT 68.720 173.900 69.040 173.960 ;
        RECT 47.560 173.620 58.370 173.760 ;
        RECT 58.715 173.760 59.305 173.805 ;
        RECT 60.900 173.760 61.220 173.820 ;
        RECT 61.955 173.760 62.605 173.805 ;
        RECT 58.715 173.620 62.605 173.760 ;
        RECT 47.560 173.560 47.880 173.620 ;
        RECT 53.080 173.560 53.400 173.620 ;
        RECT 58.715 173.575 59.005 173.620 ;
        RECT 60.900 173.560 61.220 173.620 ;
        RECT 61.955 173.575 62.605 173.620 ;
        RECT 64.580 173.560 64.900 173.820 ;
        RECT 69.270 173.760 69.410 174.640 ;
        RECT 71.495 174.595 71.785 174.640 ;
        RECT 76.080 174.580 76.400 174.640 ;
        RECT 69.640 174.240 69.960 174.500 ;
        RECT 81.690 174.440 81.830 174.920 ;
        RECT 87.120 174.440 87.440 174.500 ;
        RECT 81.690 174.300 82.750 174.440 ;
        RECT 72.400 173.900 72.720 174.160 ;
        RECT 77.920 174.100 78.240 174.160 ;
        RECT 82.610 174.145 82.750 174.300 ;
        RECT 83.070 174.300 87.440 174.440 ;
        RECT 83.070 174.145 83.210 174.300 ;
        RECT 87.120 174.240 87.440 174.300 ;
        RECT 82.075 174.100 82.365 174.145 ;
        RECT 77.920 173.960 82.365 174.100 ;
        RECT 77.920 173.900 78.240 173.960 ;
        RECT 82.075 173.915 82.365 173.960 ;
        RECT 82.535 173.915 82.825 174.145 ;
        RECT 82.995 173.915 83.285 174.145 ;
        RECT 83.900 173.900 84.220 174.160 ;
        RECT 98.160 174.100 98.480 174.160 ;
        RECT 103.770 174.145 103.910 174.980 ;
        RECT 105.980 174.920 106.300 174.980 ;
        RECT 107.820 174.920 108.140 174.980 ;
        RECT 106.915 174.780 107.205 174.825 ;
        RECT 108.740 174.780 109.060 174.840 ;
        RECT 106.915 174.640 109.060 174.780 ;
        RECT 106.915 174.595 107.205 174.640 ;
        RECT 108.740 174.580 109.060 174.640 ;
        RECT 106.440 174.440 106.760 174.500 ;
        RECT 105.150 174.300 109.430 174.440 ;
        RECT 103.695 174.100 103.985 174.145 ;
        RECT 98.160 173.960 103.985 174.100 ;
        RECT 98.160 173.900 98.480 173.960 ;
        RECT 103.695 173.915 103.985 173.960 ;
        RECT 104.600 173.900 104.920 174.160 ;
        RECT 105.150 174.145 105.290 174.300 ;
        RECT 106.440 174.240 106.760 174.300 ;
        RECT 109.290 174.160 109.430 174.300 ;
        RECT 105.075 173.915 105.365 174.145 ;
        RECT 105.520 174.100 105.840 174.160 ;
        RECT 108.755 174.100 109.045 174.145 ;
        RECT 105.520 173.960 109.045 174.100 ;
        RECT 105.520 173.900 105.840 173.960 ;
        RECT 108.755 173.915 109.045 173.960 ;
        RECT 65.130 173.620 69.410 173.760 ;
        RECT 80.695 173.760 80.985 173.805 ;
        RECT 81.600 173.760 81.920 173.820 ;
        RECT 80.695 173.620 81.920 173.760 ;
        RECT 47.650 173.420 47.790 173.560 ;
        RECT 43.970 173.280 47.790 173.420 ;
        RECT 56.760 173.220 57.080 173.480 ;
        RECT 62.740 173.420 63.060 173.480 ;
        RECT 65.130 173.420 65.270 173.620 ;
        RECT 80.695 173.575 80.985 173.620 ;
        RECT 81.600 173.560 81.920 173.620 ;
        RECT 104.140 173.760 104.460 173.820 ;
        RECT 107.375 173.760 107.665 173.805 ;
        RECT 104.140 173.620 107.665 173.760 ;
        RECT 104.140 173.560 104.460 173.620 ;
        RECT 107.375 173.575 107.665 173.620 ;
        RECT 62.740 173.280 65.270 173.420 ;
        RECT 70.560 173.420 70.880 173.480 ;
        RECT 98.160 173.420 98.480 173.480 ;
        RECT 70.560 173.280 98.480 173.420 ;
        RECT 108.830 173.420 108.970 173.915 ;
        RECT 109.200 173.900 109.520 174.160 ;
        RECT 109.660 173.900 109.980 174.160 ;
        RECT 110.210 174.100 110.350 174.980 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 110.595 174.100 110.885 174.145 ;
        RECT 110.210 173.960 110.885 174.100 ;
        RECT 110.595 173.915 110.885 173.960 ;
        RECT 117.955 174.100 118.245 174.145 ;
        RECT 118.860 174.100 119.180 174.160 ;
        RECT 117.955 173.960 119.180 174.100 ;
        RECT 117.955 173.915 118.245 173.960 ;
        RECT 118.860 173.900 119.180 173.960 ;
        RECT 118.415 173.575 118.705 173.805 ;
        RECT 109.660 173.420 109.980 173.480 ;
        RECT 108.830 173.280 109.980 173.420 ;
        RECT 62.740 173.220 63.060 173.280 ;
        RECT 70.560 173.220 70.880 173.280 ;
        RECT 98.160 173.220 98.480 173.280 ;
        RECT 109.660 173.220 109.980 173.280 ;
        RECT 117.940 173.420 118.260 173.480 ;
        RECT 118.490 173.420 118.630 173.575 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 117.940 173.280 118.630 173.420 ;
        RECT 117.940 173.220 118.260 173.280 ;
        RECT 14.370 172.600 127.530 173.080 ;
        RECT 35.140 172.400 35.460 172.460 ;
        RECT 41.595 172.400 41.885 172.445 ;
        RECT 35.140 172.260 41.885 172.400 ;
        RECT 35.140 172.200 35.460 172.260 ;
        RECT 41.595 172.215 41.885 172.260 ;
        RECT 44.340 172.400 44.660 172.460 ;
        RECT 48.940 172.400 49.260 172.460 ;
        RECT 44.340 172.260 49.260 172.400 ;
        RECT 44.340 172.200 44.660 172.260 ;
        RECT 36.980 172.060 37.300 172.120 ;
        RECT 36.980 171.920 39.970 172.060 ;
        RECT 36.980 171.860 37.300 171.920 ;
        RECT 37.900 171.720 38.220 171.780 ;
        RECT 38.835 171.720 39.125 171.765 ;
        RECT 37.900 171.580 39.125 171.720 ;
        RECT 37.900 171.520 38.220 171.580 ;
        RECT 38.835 171.535 39.125 171.580 ;
        RECT 39.280 171.520 39.600 171.780 ;
        RECT 39.830 171.765 39.970 171.920 ;
        RECT 39.755 171.535 40.045 171.765 ;
        RECT 40.660 171.520 40.980 171.780 ;
        RECT 42.500 171.520 42.820 171.780 ;
        RECT 45.350 171.765 45.490 172.260 ;
        RECT 48.940 172.200 49.260 172.260 ;
        RECT 49.400 172.400 49.720 172.460 ;
        RECT 50.780 172.400 51.100 172.460 ;
        RECT 54.460 172.400 54.780 172.460 ;
        RECT 49.400 172.260 50.090 172.400 ;
        RECT 49.400 172.200 49.720 172.260 ;
        RECT 45.810 171.920 49.630 172.060 ;
        RECT 45.810 171.765 45.950 171.920 ;
        RECT 49.490 171.780 49.630 171.920 ;
        RECT 45.275 171.535 45.565 171.765 ;
        RECT 45.735 171.535 46.025 171.765 ;
        RECT 46.195 171.535 46.485 171.765 ;
        RECT 35.600 171.380 35.920 171.440 ;
        RECT 46.270 171.380 46.410 171.535 ;
        RECT 47.100 171.520 47.420 171.780 ;
        RECT 48.940 171.520 49.260 171.780 ;
        RECT 49.400 171.520 49.720 171.780 ;
        RECT 49.950 171.765 50.090 172.260 ;
        RECT 50.780 172.260 54.780 172.400 ;
        RECT 50.780 172.200 51.100 172.260 ;
        RECT 54.460 172.200 54.780 172.260 ;
        RECT 60.455 172.400 60.745 172.445 ;
        RECT 60.900 172.400 61.220 172.460 ;
        RECT 60.455 172.260 61.220 172.400 ;
        RECT 60.455 172.215 60.745 172.260 ;
        RECT 60.900 172.200 61.220 172.260 ;
        RECT 62.295 172.400 62.585 172.445 ;
        RECT 64.580 172.400 64.900 172.460 ;
        RECT 90.800 172.400 91.120 172.460 ;
        RECT 118.860 172.400 119.180 172.460 ;
        RECT 62.295 172.260 64.900 172.400 ;
        RECT 62.295 172.215 62.585 172.260 ;
        RECT 64.580 172.200 64.900 172.260 ;
        RECT 89.510 172.260 99.770 172.400 ;
        RECT 56.760 172.060 57.080 172.120 ;
        RECT 83.455 172.060 83.745 172.105 ;
        RECT 89.510 172.060 89.650 172.260 ;
        RECT 90.800 172.200 91.120 172.260 ;
        RECT 56.760 171.920 61.590 172.060 ;
        RECT 56.760 171.860 57.080 171.920 ;
        RECT 49.875 171.535 50.165 171.765 ;
        RECT 50.780 171.520 51.100 171.780 ;
        RECT 52.635 171.535 52.925 171.765 ;
        RECT 35.600 171.240 46.410 171.380 ;
        RECT 49.030 171.380 49.170 171.520 ;
        RECT 52.710 171.380 52.850 171.535 ;
        RECT 53.080 171.520 53.400 171.780 ;
        RECT 53.540 171.520 53.860 171.780 ;
        RECT 54.460 171.520 54.780 171.780 ;
        RECT 60.440 171.720 60.760 171.780 ;
        RECT 61.450 171.765 61.590 171.920 ;
        RECT 83.455 171.920 89.650 172.060 ;
        RECT 83.455 171.875 83.745 171.920 ;
        RECT 60.915 171.720 61.205 171.765 ;
        RECT 60.440 171.580 61.205 171.720 ;
        RECT 60.440 171.520 60.760 171.580 ;
        RECT 60.915 171.535 61.205 171.580 ;
        RECT 61.375 171.535 61.665 171.765 ;
        RECT 68.720 171.720 69.040 171.780 ;
        RECT 89.510 171.765 89.650 171.920 ;
        RECT 89.895 172.060 90.185 172.105 ;
        RECT 92.295 172.060 92.585 172.105 ;
        RECT 95.535 172.060 96.185 172.105 ;
        RECT 89.895 171.920 96.185 172.060 ;
        RECT 89.895 171.875 90.185 171.920 ;
        RECT 92.295 171.875 92.885 171.920 ;
        RECT 95.535 171.875 96.185 171.920 ;
        RECT 82.075 171.720 82.365 171.765 ;
        RECT 68.720 171.580 82.365 171.720 ;
        RECT 68.720 171.520 69.040 171.580 ;
        RECT 82.075 171.535 82.365 171.580 ;
        RECT 89.435 171.535 89.725 171.765 ;
        RECT 92.595 171.560 92.885 171.875 ;
        RECT 93.675 171.720 93.965 171.765 ;
        RECT 97.255 171.720 97.545 171.765 ;
        RECT 99.090 171.720 99.380 171.765 ;
        RECT 93.675 171.580 99.380 171.720 ;
        RECT 99.630 171.720 99.770 172.260 ;
        RECT 112.970 172.260 119.180 172.400 ;
        RECT 105.980 172.060 106.300 172.120 ;
        RECT 110.120 172.060 110.440 172.120 ;
        RECT 105.980 171.920 108.050 172.060 ;
        RECT 105.980 171.860 106.300 171.920 ;
        RECT 107.910 171.765 108.050 171.920 ;
        RECT 108.830 171.920 110.440 172.060 ;
        RECT 108.830 171.765 108.970 171.920 ;
        RECT 110.120 171.860 110.440 171.920 ;
        RECT 107.375 171.720 107.665 171.765 ;
        RECT 99.630 171.580 107.665 171.720 ;
        RECT 93.675 171.535 93.965 171.580 ;
        RECT 97.255 171.535 97.545 171.580 ;
        RECT 99.090 171.535 99.380 171.580 ;
        RECT 107.375 171.535 107.665 171.580 ;
        RECT 107.835 171.535 108.125 171.765 ;
        RECT 108.755 171.535 109.045 171.765 ;
        RECT 49.030 171.240 52.850 171.380 ;
        RECT 35.600 171.180 35.920 171.240 ;
        RECT 49.400 171.040 49.720 171.100 ;
        RECT 53.170 171.040 53.310 171.520 ;
        RECT 85.295 171.380 85.585 171.425 ;
        RECT 85.295 171.240 91.030 171.380 ;
        RECT 85.295 171.195 85.585 171.240 ;
        RECT 49.400 170.900 53.310 171.040 ;
        RECT 49.400 170.840 49.720 170.900 ;
        RECT 35.140 170.700 35.460 170.760 ;
        RECT 37.455 170.700 37.745 170.745 ;
        RECT 35.140 170.560 37.745 170.700 ;
        RECT 35.140 170.500 35.460 170.560 ;
        RECT 37.455 170.515 37.745 170.560 ;
        RECT 41.120 170.700 41.440 170.760 ;
        RECT 43.895 170.700 44.185 170.745 ;
        RECT 41.120 170.560 44.185 170.700 ;
        RECT 41.120 170.500 41.440 170.560 ;
        RECT 43.895 170.515 44.185 170.560 ;
        RECT 45.720 170.700 46.040 170.760 ;
        RECT 47.575 170.700 47.865 170.745 ;
        RECT 45.720 170.560 47.865 170.700 ;
        RECT 45.720 170.500 46.040 170.560 ;
        RECT 47.575 170.515 47.865 170.560 ;
        RECT 51.255 170.700 51.545 170.745 ;
        RECT 52.160 170.700 52.480 170.760 ;
        RECT 51.255 170.560 52.480 170.700 ;
        RECT 51.255 170.515 51.545 170.560 ;
        RECT 52.160 170.500 52.480 170.560 ;
        RECT 88.055 170.700 88.345 170.745 ;
        RECT 89.420 170.700 89.740 170.760 ;
        RECT 90.890 170.745 91.030 171.240 ;
        RECT 98.160 171.180 98.480 171.440 ;
        RECT 99.555 171.380 99.845 171.425 ;
        RECT 105.520 171.380 105.840 171.440 ;
        RECT 99.555 171.240 105.840 171.380 ;
        RECT 107.450 171.380 107.590 171.535 ;
        RECT 109.200 171.520 109.520 171.780 ;
        RECT 109.660 171.520 109.980 171.780 ;
        RECT 112.970 171.765 113.110 172.260 ;
        RECT 118.860 172.200 119.180 172.260 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 117.135 172.060 117.425 172.105 ;
        RECT 117.940 172.060 118.260 172.120 ;
        RECT 120.375 172.060 121.025 172.105 ;
        RECT 117.135 171.920 121.025 172.060 ;
        RECT 117.135 171.875 117.725 171.920 ;
        RECT 112.895 171.535 113.185 171.765 ;
        RECT 117.435 171.560 117.725 171.875 ;
        RECT 117.940 171.860 118.260 171.920 ;
        RECT 120.375 171.875 121.025 171.920 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 118.515 171.720 118.805 171.765 ;
        RECT 122.095 171.720 122.385 171.765 ;
        RECT 123.930 171.720 124.220 171.765 ;
        RECT 118.515 171.580 124.220 171.720 ;
        RECT 118.515 171.535 118.805 171.580 ;
        RECT 122.095 171.535 122.385 171.580 ;
        RECT 123.930 171.535 124.220 171.580 ;
        RECT 112.970 171.380 113.110 171.535 ;
        RECT 107.450 171.240 113.110 171.380 ;
        RECT 121.160 171.380 121.480 171.440 ;
        RECT 123.015 171.380 123.305 171.425 ;
        RECT 121.160 171.240 123.305 171.380 ;
        RECT 99.555 171.195 99.845 171.240 ;
        RECT 105.520 171.180 105.840 171.240 ;
        RECT 121.160 171.180 121.480 171.240 ;
        RECT 123.015 171.195 123.305 171.240 ;
        RECT 124.380 171.180 124.700 171.440 ;
        RECT 93.675 171.040 93.965 171.085 ;
        RECT 96.795 171.040 97.085 171.085 ;
        RECT 98.685 171.040 98.975 171.085 ;
        RECT 114.260 171.040 114.580 171.100 ;
        RECT 93.675 170.900 98.975 171.040 ;
        RECT 93.675 170.855 93.965 170.900 ;
        RECT 96.795 170.855 97.085 170.900 ;
        RECT 98.685 170.855 98.975 170.900 ;
        RECT 99.630 170.900 114.580 171.040 ;
        RECT 88.055 170.560 89.740 170.700 ;
        RECT 88.055 170.515 88.345 170.560 ;
        RECT 89.420 170.500 89.740 170.560 ;
        RECT 90.815 170.700 91.105 170.745 ;
        RECT 99.630 170.700 99.770 170.900 ;
        RECT 114.260 170.840 114.580 170.900 ;
        RECT 118.515 171.040 118.805 171.085 ;
        RECT 121.635 171.040 121.925 171.085 ;
        RECT 123.525 171.040 123.815 171.085 ;
        RECT 118.515 170.900 123.815 171.040 ;
        RECT 118.515 170.855 118.805 170.900 ;
        RECT 121.635 170.855 121.925 170.900 ;
        RECT 123.525 170.855 123.815 170.900 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 90.815 170.560 99.770 170.700 ;
        RECT 90.815 170.515 91.105 170.560 ;
        RECT 106.900 170.500 107.220 170.760 ;
        RECT 111.040 170.500 111.360 170.760 ;
        RECT 113.340 170.500 113.660 170.760 ;
        RECT 115.655 170.700 115.945 170.745 ;
        RECT 117.020 170.700 117.340 170.760 ;
        RECT 115.655 170.560 117.340 170.700 ;
        RECT 115.655 170.515 115.945 170.560 ;
        RECT 117.020 170.500 117.340 170.560 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 14.370 169.880 127.530 170.360 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 47.100 169.680 47.420 169.740 ;
        RECT 67.340 169.680 67.660 169.740 ;
        RECT 68.735 169.680 69.025 169.725 ;
        RECT 47.100 169.540 69.025 169.680 ;
        RECT 47.100 169.480 47.420 169.540 ;
        RECT 67.340 169.480 67.660 169.540 ;
        RECT 68.735 169.495 69.025 169.540 ;
        RECT 70.560 169.480 70.880 169.740 ;
        RECT 96.795 169.680 97.085 169.725 ;
        RECT 98.160 169.680 98.480 169.740 ;
        RECT 96.795 169.540 98.480 169.680 ;
        RECT 96.795 169.495 97.085 169.540 ;
        RECT 98.160 169.480 98.480 169.540 ;
        RECT 121.160 169.480 121.480 169.740 ;
        RECT 40.660 169.340 40.980 169.400 ;
        RECT 70.650 169.340 70.790 169.480 ;
        RECT 40.660 169.200 70.790 169.340 ;
        RECT 84.330 169.340 84.620 169.385 ;
        RECT 87.110 169.340 87.400 169.385 ;
        RECT 88.970 169.340 89.260 169.385 ;
        RECT 84.330 169.200 89.260 169.340 ;
        RECT 40.660 169.140 40.980 169.200 ;
        RECT 84.330 169.155 84.620 169.200 ;
        RECT 87.110 169.155 87.400 169.200 ;
        RECT 88.970 169.155 89.260 169.200 ;
        RECT 89.420 169.340 89.740 169.400 ;
        RECT 89.420 169.200 92.870 169.340 ;
        RECT 89.420 169.140 89.740 169.200 ;
        RECT 77.015 169.000 77.305 169.045 ;
        RECT 79.760 169.000 80.080 169.060 ;
        RECT 77.015 168.860 80.080 169.000 ;
        RECT 77.015 168.815 77.305 168.860 ;
        RECT 79.760 168.800 80.080 168.860 ;
        RECT 81.690 168.860 91.490 169.000 ;
        RECT 26.875 168.660 27.165 168.705 ;
        RECT 30.080 168.660 30.400 168.720 ;
        RECT 33.315 168.660 33.605 168.705 ;
        RECT 35.600 168.660 35.920 168.720 ;
        RECT 26.875 168.520 35.920 168.660 ;
        RECT 26.875 168.475 27.165 168.520 ;
        RECT 30.080 168.460 30.400 168.520 ;
        RECT 33.315 168.475 33.605 168.520 ;
        RECT 35.600 168.460 35.920 168.520 ;
        RECT 43.880 168.460 44.200 168.720 ;
        RECT 69.655 168.660 69.945 168.705 ;
        RECT 70.100 168.660 70.420 168.720 ;
        RECT 71.495 168.660 71.785 168.705 ;
        RECT 69.655 168.520 71.785 168.660 ;
        RECT 69.655 168.475 69.945 168.520 ;
        RECT 70.100 168.460 70.420 168.520 ;
        RECT 71.495 168.475 71.785 168.520 ;
        RECT 80.465 168.320 80.755 168.365 ;
        RECT 81.690 168.320 81.830 168.860 ;
        RECT 84.330 168.660 84.620 168.705 ;
        RECT 84.330 168.520 86.865 168.660 ;
        RECT 84.330 168.475 84.620 168.520 ;
        RECT 77.550 168.180 81.830 168.320 ;
        RECT 82.470 168.320 82.760 168.365 ;
        RECT 83.900 168.320 84.220 168.380 ;
        RECT 86.650 168.365 86.865 168.520 ;
        RECT 87.580 168.460 87.900 168.720 ;
        RECT 89.435 168.660 89.725 168.705 ;
        RECT 90.800 168.660 91.120 168.720 ;
        RECT 89.435 168.520 91.120 168.660 ;
        RECT 91.350 168.660 91.490 168.860 ;
        RECT 91.720 168.800 92.040 169.060 ;
        RECT 92.730 169.045 92.870 169.200 ;
        RECT 94.955 169.155 95.245 169.385 ;
        RECT 105.635 169.340 105.925 169.385 ;
        RECT 108.755 169.340 109.045 169.385 ;
        RECT 110.645 169.340 110.935 169.385 ;
        RECT 105.635 169.200 110.935 169.340 ;
        RECT 105.635 169.155 105.925 169.200 ;
        RECT 108.755 169.155 109.045 169.200 ;
        RECT 110.645 169.155 110.935 169.200 ;
        RECT 92.655 168.815 92.945 169.045 ;
        RECT 93.115 168.660 93.405 168.705 ;
        RECT 91.350 168.520 93.405 168.660 ;
        RECT 95.030 168.660 95.170 169.155 ;
        RECT 109.660 169.000 109.980 169.060 ;
        RECT 110.135 169.000 110.425 169.045 ;
        RECT 109.660 168.860 110.425 169.000 ;
        RECT 109.660 168.800 109.980 168.860 ;
        RECT 110.135 168.815 110.425 168.860 ;
        RECT 112.420 169.000 112.740 169.060 ;
        RECT 115.195 169.000 115.485 169.045 ;
        RECT 112.420 168.860 115.485 169.000 ;
        RECT 112.420 168.800 112.740 168.860 ;
        RECT 115.195 168.815 115.485 168.860 ;
        RECT 117.020 169.000 117.340 169.060 ;
        RECT 119.335 169.000 119.625 169.045 ;
        RECT 117.020 168.860 119.625 169.000 ;
        RECT 117.020 168.800 117.340 168.860 ;
        RECT 119.335 168.815 119.625 168.860 ;
        RECT 95.875 168.660 96.165 168.705 ;
        RECT 95.030 168.520 96.165 168.660 ;
        RECT 89.435 168.475 89.725 168.520 ;
        RECT 90.800 168.460 91.120 168.520 ;
        RECT 93.115 168.475 93.405 168.520 ;
        RECT 95.875 168.475 96.165 168.520 ;
        RECT 104.555 168.365 104.845 168.680 ;
        RECT 105.635 168.660 105.925 168.705 ;
        RECT 109.215 168.660 109.505 168.705 ;
        RECT 111.050 168.660 111.340 168.705 ;
        RECT 105.635 168.520 111.340 168.660 ;
        RECT 105.635 168.475 105.925 168.520 ;
        RECT 109.215 168.475 109.505 168.520 ;
        RECT 111.050 168.475 111.340 168.520 ;
        RECT 111.500 168.460 111.820 168.720 ;
        RECT 114.260 168.460 114.580 168.720 ;
        RECT 114.735 168.660 115.025 168.705 ;
        RECT 116.575 168.660 116.865 168.705 ;
        RECT 114.735 168.520 116.865 168.660 ;
        RECT 114.735 168.475 115.025 168.520 ;
        RECT 116.575 168.475 116.865 168.520 ;
        RECT 120.255 168.475 120.545 168.705 ;
        RECT 122.555 168.660 122.845 168.705 ;
        RECT 127.600 168.660 127.920 168.720 ;
        RECT 122.555 168.520 127.920 168.660 ;
        RECT 122.555 168.475 122.845 168.520 ;
        RECT 85.730 168.320 86.020 168.365 ;
        RECT 82.470 168.180 86.020 168.320 ;
        RECT 27.335 167.980 27.625 168.025 ;
        RECT 29.620 167.980 29.940 168.040 ;
        RECT 27.335 167.840 29.940 167.980 ;
        RECT 27.335 167.795 27.625 167.840 ;
        RECT 29.620 167.780 29.940 167.840 ;
        RECT 32.855 167.980 33.145 168.025 ;
        RECT 33.760 167.980 34.080 168.040 ;
        RECT 32.855 167.840 34.080 167.980 ;
        RECT 32.855 167.795 33.145 167.840 ;
        RECT 33.760 167.780 34.080 167.840 ;
        RECT 36.520 167.780 36.840 168.040 ;
        RECT 76.080 167.980 76.400 168.040 ;
        RECT 77.550 168.025 77.690 168.180 ;
        RECT 80.465 168.135 80.755 168.180 ;
        RECT 82.470 168.135 82.760 168.180 ;
        RECT 83.900 168.120 84.220 168.180 ;
        RECT 85.730 168.135 86.020 168.180 ;
        RECT 86.650 168.320 86.940 168.365 ;
        RECT 88.510 168.320 88.800 168.365 ;
        RECT 86.650 168.180 88.800 168.320 ;
        RECT 86.650 168.135 86.940 168.180 ;
        RECT 88.510 168.135 88.800 168.180 ;
        RECT 104.255 168.320 104.845 168.365 ;
        RECT 106.900 168.320 107.220 168.380 ;
        RECT 107.495 168.320 108.145 168.365 ;
        RECT 104.255 168.180 108.145 168.320 ;
        RECT 104.255 168.135 104.545 168.180 ;
        RECT 106.900 168.120 107.220 168.180 ;
        RECT 107.495 168.135 108.145 168.180 ;
        RECT 110.120 168.320 110.440 168.380 ;
        RECT 120.330 168.320 120.470 168.475 ;
        RECT 127.600 168.460 127.920 168.520 ;
        RECT 110.120 168.180 120.470 168.320 ;
        RECT 110.120 168.120 110.440 168.180 ;
        RECT 77.475 167.980 77.765 168.025 ;
        RECT 76.080 167.840 77.765 167.980 ;
        RECT 76.080 167.780 76.400 167.840 ;
        RECT 77.475 167.795 77.765 167.840 ;
        RECT 77.935 167.980 78.225 168.025 ;
        RECT 78.840 167.980 79.160 168.040 ;
        RECT 77.935 167.840 79.160 167.980 ;
        RECT 77.935 167.795 78.225 167.840 ;
        RECT 78.840 167.780 79.160 167.840 ;
        RECT 79.775 167.980 80.065 168.025 ;
        RECT 82.980 167.980 83.300 168.040 ;
        RECT 79.775 167.840 83.300 167.980 ;
        RECT 79.775 167.795 80.065 167.840 ;
        RECT 82.980 167.780 83.300 167.840 ;
        RECT 102.300 167.980 102.620 168.040 ;
        RECT 102.775 167.980 103.065 168.025 ;
        RECT 102.300 167.840 103.065 167.980 ;
        RECT 102.300 167.780 102.620 167.840 ;
        RECT 102.775 167.795 103.065 167.840 ;
        RECT 110.580 167.980 110.900 168.040 ;
        RECT 112.435 167.980 112.725 168.025 ;
        RECT 110.580 167.840 112.725 167.980 ;
        RECT 110.580 167.780 110.900 167.840 ;
        RECT 112.435 167.795 112.725 167.840 ;
        RECT 112.880 167.980 113.200 168.040 ;
        RECT 122.095 167.980 122.385 168.025 ;
        RECT 112.880 167.840 122.385 167.980 ;
        RECT 112.880 167.780 113.200 167.840 ;
        RECT 122.095 167.795 122.385 167.840 ;
        RECT 14.370 167.160 127.530 167.640 ;
        RECT 70.100 166.960 70.420 167.020 ;
        RECT 48.110 166.820 52.850 166.960 ;
        RECT 24.560 166.420 24.880 166.680 ;
        RECT 26.855 166.620 27.505 166.665 ;
        RECT 29.620 166.620 29.940 166.680 ;
        RECT 30.455 166.620 30.745 166.665 ;
        RECT 26.855 166.480 30.745 166.620 ;
        RECT 26.855 166.435 27.505 166.480 ;
        RECT 29.620 166.420 29.940 166.480 ;
        RECT 30.155 166.435 30.745 166.480 ;
        RECT 35.600 166.620 35.920 166.680 ;
        RECT 48.110 166.620 48.250 166.820 ;
        RECT 35.600 166.480 48.250 166.620 ;
        RECT 48.595 166.620 48.885 166.665 ;
        RECT 50.780 166.620 51.100 166.680 ;
        RECT 51.835 166.620 52.485 166.665 ;
        RECT 48.595 166.480 52.485 166.620 ;
        RECT 52.710 166.620 52.850 166.820 ;
        RECT 70.100 166.820 73.550 166.960 ;
        RECT 70.100 166.760 70.420 166.820 ;
        RECT 53.080 166.620 53.400 166.680 ;
        RECT 72.875 166.620 73.165 166.665 ;
        RECT 52.710 166.480 59.290 166.620 ;
        RECT 23.660 166.280 23.950 166.325 ;
        RECT 25.495 166.280 25.785 166.325 ;
        RECT 29.075 166.280 29.365 166.325 ;
        RECT 23.660 166.140 29.365 166.280 ;
        RECT 23.660 166.095 23.950 166.140 ;
        RECT 25.495 166.095 25.785 166.140 ;
        RECT 29.075 166.095 29.365 166.140 ;
        RECT 30.155 166.120 30.445 166.435 ;
        RECT 35.600 166.420 35.920 166.480 ;
        RECT 33.315 166.280 33.605 166.325 ;
        RECT 34.220 166.280 34.540 166.340 ;
        RECT 33.315 166.140 34.540 166.280 ;
        RECT 33.315 166.095 33.605 166.140 ;
        RECT 34.220 166.080 34.540 166.140 ;
        RECT 36.075 166.280 36.365 166.325 ;
        RECT 36.520 166.280 36.840 166.340 ;
        RECT 37.530 166.325 37.670 166.480 ;
        RECT 48.595 166.435 49.185 166.480 ;
        RECT 36.075 166.140 36.840 166.280 ;
        RECT 36.075 166.095 36.365 166.140 ;
        RECT 36.520 166.080 36.840 166.140 ;
        RECT 37.455 166.095 37.745 166.325 ;
        RECT 45.350 166.140 48.710 166.280 ;
        RECT 23.195 165.940 23.485 165.985 ;
        RECT 26.860 165.940 27.180 166.000 ;
        RECT 23.195 165.800 27.180 165.940 ;
        RECT 23.195 165.755 23.485 165.800 ;
        RECT 26.860 165.740 27.180 165.800 ;
        RECT 31.935 165.940 32.225 165.985 ;
        RECT 39.295 165.940 39.585 165.985 ;
        RECT 42.960 165.940 43.280 166.000 ;
        RECT 31.935 165.800 43.280 165.940 ;
        RECT 31.935 165.755 32.225 165.800 ;
        RECT 39.295 165.755 39.585 165.800 ;
        RECT 42.960 165.740 43.280 165.800 ;
        RECT 24.065 165.600 24.355 165.645 ;
        RECT 25.955 165.600 26.245 165.645 ;
        RECT 29.075 165.600 29.365 165.645 ;
        RECT 24.065 165.460 29.365 165.600 ;
        RECT 24.065 165.415 24.355 165.460 ;
        RECT 25.955 165.415 26.245 165.460 ;
        RECT 29.075 165.415 29.365 165.460 ;
        RECT 29.620 165.600 29.940 165.660 ;
        RECT 42.055 165.600 42.345 165.645 ;
        RECT 45.350 165.600 45.490 166.140 ;
        RECT 45.735 165.940 46.025 165.985 ;
        RECT 48.570 165.940 48.710 166.140 ;
        RECT 48.895 166.120 49.185 166.435 ;
        RECT 50.780 166.420 51.100 166.480 ;
        RECT 51.835 166.435 52.485 166.480 ;
        RECT 53.080 166.420 53.400 166.480 ;
        RECT 59.150 166.325 59.290 166.480 ;
        RECT 68.350 166.480 73.165 166.620 ;
        RECT 68.350 166.340 68.490 166.480 ;
        RECT 72.875 166.435 73.165 166.480 ;
        RECT 49.975 166.280 50.265 166.325 ;
        RECT 53.555 166.280 53.845 166.325 ;
        RECT 55.390 166.280 55.680 166.325 ;
        RECT 49.975 166.140 55.680 166.280 ;
        RECT 49.975 166.095 50.265 166.140 ;
        RECT 53.555 166.095 53.845 166.140 ;
        RECT 55.390 166.095 55.680 166.140 ;
        RECT 59.075 166.280 59.365 166.325 ;
        RECT 60.915 166.280 61.205 166.325 ;
        RECT 59.075 166.140 61.205 166.280 ;
        RECT 59.075 166.095 59.365 166.140 ;
        RECT 60.915 166.095 61.205 166.140 ;
        RECT 61.360 166.280 61.680 166.340 ;
        RECT 62.295 166.280 62.585 166.325 ;
        RECT 66.895 166.280 67.185 166.325 ;
        RECT 61.360 166.140 67.185 166.280 ;
        RECT 61.360 166.080 61.680 166.140 ;
        RECT 62.295 166.095 62.585 166.140 ;
        RECT 66.895 166.095 67.185 166.140 ;
        RECT 68.260 166.080 68.580 166.340 ;
        RECT 70.560 166.080 70.880 166.340 ;
        RECT 72.415 166.280 72.705 166.325 ;
        RECT 73.410 166.280 73.550 166.820 ;
        RECT 110.120 166.760 110.440 167.020 ;
        RECT 77.410 166.620 77.700 166.665 ;
        RECT 80.670 166.620 80.960 166.665 ;
        RECT 77.410 166.480 80.960 166.620 ;
        RECT 77.410 166.435 77.700 166.480 ;
        RECT 72.415 166.140 73.550 166.280 ;
        RECT 72.415 166.095 72.705 166.140 ;
        RECT 54.000 165.940 54.320 166.000 ;
        RECT 45.735 165.800 47.330 165.940 ;
        RECT 48.570 165.800 54.320 165.940 ;
        RECT 45.735 165.755 46.025 165.800 ;
        RECT 29.620 165.460 45.490 165.600 ;
        RECT 29.620 165.400 29.940 165.460 ;
        RECT 42.055 165.415 42.345 165.460 ;
        RECT 28.240 165.260 28.560 165.320 ;
        RECT 32.395 165.260 32.685 165.305 ;
        RECT 28.240 165.120 32.685 165.260 ;
        RECT 28.240 165.060 28.560 165.120 ;
        RECT 32.395 165.075 32.685 165.120 ;
        RECT 37.900 165.060 38.220 165.320 ;
        RECT 42.500 165.060 42.820 165.320 ;
        RECT 47.190 165.305 47.330 165.800 ;
        RECT 54.000 165.740 54.320 165.800 ;
        RECT 54.460 165.740 54.780 166.000 ;
        RECT 55.855 165.940 56.145 165.985 ;
        RECT 57.220 165.940 57.540 166.000 ;
        RECT 63.660 165.940 63.980 166.000 ;
        RECT 55.855 165.800 63.980 165.940 ;
        RECT 55.855 165.755 56.145 165.800 ;
        RECT 57.220 165.740 57.540 165.800 ;
        RECT 63.660 165.740 63.980 165.800 ;
        RECT 66.420 165.940 66.740 166.000 ;
        RECT 71.035 165.940 71.325 165.985 ;
        RECT 66.420 165.800 71.325 165.940 ;
        RECT 66.420 165.740 66.740 165.800 ;
        RECT 71.035 165.755 71.325 165.800 ;
        RECT 71.955 165.940 72.245 165.985 ;
        RECT 73.780 165.940 74.100 166.000 ;
        RECT 74.700 165.940 75.020 166.000 ;
        RECT 71.955 165.800 75.020 165.940 ;
        RECT 78.930 165.940 79.070 166.480 ;
        RECT 80.670 166.435 80.960 166.480 ;
        RECT 81.590 166.620 81.880 166.665 ;
        RECT 83.450 166.620 83.740 166.665 ;
        RECT 81.590 166.480 83.740 166.620 ;
        RECT 81.590 166.435 81.880 166.480 ;
        RECT 83.450 166.435 83.740 166.480 ;
        RECT 83.900 166.620 84.220 166.680 ;
        RECT 86.675 166.620 86.965 166.665 ;
        RECT 83.900 166.480 86.965 166.620 ;
        RECT 79.270 166.280 79.560 166.325 ;
        RECT 81.590 166.280 81.805 166.435 ;
        RECT 83.900 166.420 84.220 166.480 ;
        RECT 86.675 166.435 86.965 166.480 ;
        RECT 99.490 166.620 99.780 166.665 ;
        RECT 100.000 166.620 100.320 166.680 ;
        RECT 102.750 166.620 103.040 166.665 ;
        RECT 99.490 166.480 103.040 166.620 ;
        RECT 99.490 166.435 99.780 166.480 ;
        RECT 100.000 166.420 100.320 166.480 ;
        RECT 102.750 166.435 103.040 166.480 ;
        RECT 103.670 166.620 103.960 166.665 ;
        RECT 105.530 166.620 105.820 166.665 ;
        RECT 103.670 166.480 105.820 166.620 ;
        RECT 103.670 166.435 103.960 166.480 ;
        RECT 105.530 166.435 105.820 166.480 ;
        RECT 117.135 166.620 117.425 166.665 ;
        RECT 119.320 166.620 119.640 166.680 ;
        RECT 120.375 166.620 121.025 166.665 ;
        RECT 117.135 166.480 121.025 166.620 ;
        RECT 117.135 166.435 117.725 166.480 ;
        RECT 85.295 166.280 85.585 166.325 ;
        RECT 79.270 166.140 81.805 166.280 ;
        RECT 82.150 166.140 85.585 166.280 ;
        RECT 79.270 166.095 79.560 166.140 ;
        RECT 82.150 165.940 82.290 166.140 ;
        RECT 85.295 166.095 85.585 166.140 ;
        RECT 85.755 166.280 86.045 166.325 ;
        RECT 87.135 166.280 87.425 166.325 ;
        RECT 88.500 166.280 88.820 166.340 ;
        RECT 85.755 166.140 88.820 166.280 ;
        RECT 85.755 166.095 86.045 166.140 ;
        RECT 87.135 166.095 87.425 166.140 ;
        RECT 88.500 166.080 88.820 166.140 ;
        RECT 94.955 166.095 95.245 166.325 ;
        RECT 101.350 166.280 101.640 166.325 ;
        RECT 103.670 166.280 103.885 166.435 ;
        RECT 101.350 166.140 103.885 166.280 ;
        RECT 107.375 166.280 107.665 166.325 ;
        RECT 110.580 166.280 110.900 166.340 ;
        RECT 107.375 166.140 110.900 166.280 ;
        RECT 101.350 166.095 101.640 166.140 ;
        RECT 107.375 166.095 107.665 166.140 ;
        RECT 78.930 165.800 82.290 165.940 ;
        RECT 71.955 165.755 72.245 165.800 ;
        RECT 73.780 165.740 74.100 165.800 ;
        RECT 74.700 165.740 75.020 165.800 ;
        RECT 82.520 165.740 82.840 166.000 ;
        RECT 84.375 165.940 84.665 165.985 ;
        RECT 90.800 165.940 91.120 166.000 ;
        RECT 84.375 165.800 91.120 165.940 ;
        RECT 84.375 165.755 84.665 165.800 ;
        RECT 90.800 165.740 91.120 165.800 ;
        RECT 91.720 165.940 92.040 166.000 ;
        RECT 93.560 165.940 93.880 166.000 ;
        RECT 91.720 165.800 93.880 165.940 ;
        RECT 91.720 165.740 92.040 165.800 ;
        RECT 93.560 165.740 93.880 165.800 ;
        RECT 94.480 165.740 94.800 166.000 ;
        RECT 95.030 165.940 95.170 166.095 ;
        RECT 110.580 166.080 110.900 166.140 ;
        RECT 111.055 166.280 111.345 166.325 ;
        RECT 111.960 166.280 112.280 166.340 ;
        RECT 111.055 166.140 112.280 166.280 ;
        RECT 111.055 166.095 111.345 166.140 ;
        RECT 111.960 166.080 112.280 166.140 ;
        RECT 117.435 166.120 117.725 166.435 ;
        RECT 119.320 166.420 119.640 166.480 ;
        RECT 120.375 166.435 121.025 166.480 ;
        RECT 118.515 166.280 118.805 166.325 ;
        RECT 122.095 166.280 122.385 166.325 ;
        RECT 123.930 166.280 124.220 166.325 ;
        RECT 118.515 166.140 124.220 166.280 ;
        RECT 118.515 166.095 118.805 166.140 ;
        RECT 122.095 166.095 122.385 166.140 ;
        RECT 123.930 166.095 124.220 166.140 ;
        RECT 124.380 166.080 124.700 166.340 ;
        RECT 97.485 165.940 97.775 165.985 ;
        RECT 98.160 165.940 98.480 166.000 ;
        RECT 95.030 165.800 98.480 165.940 ;
        RECT 97.485 165.755 97.775 165.800 ;
        RECT 98.160 165.740 98.480 165.800 ;
        RECT 104.600 165.740 104.920 166.000 ;
        RECT 105.520 165.940 105.840 166.000 ;
        RECT 106.455 165.940 106.745 165.985 ;
        RECT 111.500 165.940 111.820 166.000 ;
        RECT 124.470 165.940 124.610 166.080 ;
        RECT 105.520 165.800 124.610 165.940 ;
        RECT 105.520 165.740 105.840 165.800 ;
        RECT 106.455 165.755 106.745 165.800 ;
        RECT 111.500 165.740 111.820 165.800 ;
        RECT 49.975 165.600 50.265 165.645 ;
        RECT 53.095 165.600 53.385 165.645 ;
        RECT 54.985 165.600 55.275 165.645 ;
        RECT 49.975 165.460 55.275 165.600 ;
        RECT 49.975 165.415 50.265 165.460 ;
        RECT 53.095 165.415 53.385 165.460 ;
        RECT 54.985 165.415 55.275 165.460 ;
        RECT 69.655 165.600 69.945 165.645 ;
        RECT 78.380 165.600 78.700 165.660 ;
        RECT 69.655 165.460 78.700 165.600 ;
        RECT 69.655 165.415 69.945 165.460 ;
        RECT 78.380 165.400 78.700 165.460 ;
        RECT 79.270 165.600 79.560 165.645 ;
        RECT 82.050 165.600 82.340 165.645 ;
        RECT 83.910 165.600 84.200 165.645 ;
        RECT 79.270 165.460 84.200 165.600 ;
        RECT 79.270 165.415 79.560 165.460 ;
        RECT 82.050 165.415 82.340 165.460 ;
        RECT 83.910 165.415 84.200 165.460 ;
        RECT 101.350 165.600 101.640 165.645 ;
        RECT 104.130 165.600 104.420 165.645 ;
        RECT 105.990 165.600 106.280 165.645 ;
        RECT 101.350 165.460 106.280 165.600 ;
        RECT 101.350 165.415 101.640 165.460 ;
        RECT 104.130 165.415 104.420 165.460 ;
        RECT 105.990 165.415 106.280 165.460 ;
        RECT 108.740 165.600 109.060 165.660 ;
        RECT 110.580 165.600 110.900 165.660 ;
        RECT 108.740 165.460 110.900 165.600 ;
        RECT 108.740 165.400 109.060 165.460 ;
        RECT 110.580 165.400 110.900 165.460 ;
        RECT 111.960 165.600 112.280 165.660 ;
        RECT 115.655 165.600 115.945 165.645 ;
        RECT 111.960 165.460 115.945 165.600 ;
        RECT 111.960 165.400 112.280 165.460 ;
        RECT 115.655 165.415 115.945 165.460 ;
        RECT 118.515 165.600 118.805 165.645 ;
        RECT 121.635 165.600 121.925 165.645 ;
        RECT 123.525 165.600 123.815 165.645 ;
        RECT 118.515 165.460 123.815 165.600 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 118.515 165.415 118.805 165.460 ;
        RECT 121.635 165.415 121.925 165.460 ;
        RECT 123.525 165.415 123.815 165.460 ;
        RECT 47.115 165.260 47.405 165.305 ;
        RECT 49.400 165.260 49.720 165.320 ;
        RECT 47.115 165.120 49.720 165.260 ;
        RECT 47.115 165.075 47.405 165.120 ;
        RECT 49.400 165.060 49.720 165.120 ;
        RECT 58.600 165.060 58.920 165.320 ;
        RECT 66.435 165.260 66.725 165.305 ;
        RECT 68.720 165.260 69.040 165.320 ;
        RECT 66.435 165.120 69.040 165.260 ;
        RECT 66.435 165.075 66.725 165.120 ;
        RECT 68.720 165.060 69.040 165.120 ;
        RECT 72.860 165.260 73.180 165.320 ;
        RECT 75.405 165.260 75.695 165.305 ;
        RECT 72.860 165.120 75.695 165.260 ;
        RECT 78.470 165.260 78.610 165.400 ;
        RECT 79.760 165.260 80.080 165.320 ;
        RECT 91.720 165.260 92.040 165.320 ;
        RECT 78.470 165.120 92.040 165.260 ;
        RECT 72.860 165.060 73.180 165.120 ;
        RECT 75.405 165.075 75.695 165.120 ;
        RECT 79.760 165.060 80.080 165.120 ;
        RECT 91.720 165.060 92.040 165.120 ;
        RECT 96.320 165.260 96.640 165.320 ;
        RECT 96.795 165.260 97.085 165.305 ;
        RECT 96.320 165.120 97.085 165.260 ;
        RECT 96.320 165.060 96.640 165.120 ;
        RECT 96.795 165.075 97.085 165.120 ;
        RECT 113.800 165.060 114.120 165.320 ;
        RECT 121.160 165.260 121.480 165.320 ;
        RECT 123.080 165.260 123.370 165.305 ;
        RECT 121.160 165.120 123.370 165.260 ;
        RECT 121.160 165.060 121.480 165.120 ;
        RECT 123.080 165.075 123.370 165.120 ;
        RECT 14.370 164.440 127.530 164.920 ;
        RECT 24.560 164.240 24.880 164.300 ;
        RECT 25.495 164.240 25.785 164.285 ;
        RECT 24.560 164.100 25.785 164.240 ;
        RECT 24.560 164.040 24.880 164.100 ;
        RECT 25.495 164.055 25.785 164.100 ;
        RECT 50.780 164.040 51.100 164.300 ;
        RECT 54.460 164.040 54.780 164.300 ;
        RECT 61.360 164.240 61.680 164.300 ;
        RECT 82.520 164.240 82.840 164.300 ;
        RECT 82.995 164.240 83.285 164.285 ;
        RECT 61.360 164.100 71.020 164.240 ;
        RECT 61.360 164.040 61.680 164.100 ;
        RECT 27.745 163.900 28.035 163.945 ;
        RECT 29.635 163.900 29.925 163.945 ;
        RECT 32.755 163.900 33.045 163.945 ;
        RECT 27.745 163.760 33.045 163.900 ;
        RECT 27.745 163.715 28.035 163.760 ;
        RECT 29.635 163.715 29.925 163.760 ;
        RECT 32.755 163.715 33.045 163.760 ;
        RECT 38.935 163.900 39.225 163.945 ;
        RECT 42.055 163.900 42.345 163.945 ;
        RECT 43.945 163.900 44.235 163.945 ;
        RECT 57.220 163.900 57.540 163.960 ;
        RECT 38.935 163.760 44.235 163.900 ;
        RECT 38.935 163.715 39.225 163.760 ;
        RECT 42.055 163.715 42.345 163.760 ;
        RECT 43.945 163.715 44.235 163.760 ;
        RECT 44.890 163.760 57.540 163.900 ;
        RECT 28.240 163.360 28.560 163.620 ;
        RECT 28.700 163.560 29.020 163.620 ;
        RECT 36.520 163.560 36.840 163.620 ;
        RECT 44.890 163.605 45.030 163.760 ;
        RECT 57.220 163.700 57.540 163.760 ;
        RECT 57.795 163.900 58.085 163.945 ;
        RECT 60.915 163.900 61.205 163.945 ;
        RECT 62.805 163.900 63.095 163.945 ;
        RECT 57.795 163.760 63.095 163.900 ;
        RECT 57.795 163.715 58.085 163.760 ;
        RECT 60.915 163.715 61.205 163.760 ;
        RECT 62.805 163.715 63.095 163.760 ;
        RECT 44.815 163.560 45.105 163.605 ;
        RECT 28.700 163.420 45.105 163.560 ;
        RECT 28.700 163.360 29.020 163.420 ;
        RECT 36.520 163.360 36.840 163.420 ;
        RECT 44.815 163.375 45.105 163.420 ;
        RECT 49.415 163.560 49.705 163.605 ;
        RECT 60.440 163.560 60.760 163.620 ;
        RECT 49.415 163.420 53.770 163.560 ;
        RECT 49.415 163.375 49.705 163.420 ;
        RECT 26.400 163.020 26.720 163.280 ;
        RECT 26.860 163.020 27.180 163.280 ;
        RECT 27.340 163.220 27.630 163.265 ;
        RECT 29.175 163.220 29.465 163.265 ;
        RECT 32.755 163.220 33.045 163.265 ;
        RECT 27.340 163.080 33.045 163.220 ;
        RECT 27.340 163.035 27.630 163.080 ;
        RECT 29.175 163.035 29.465 163.080 ;
        RECT 32.755 163.035 33.045 163.080 ;
        RECT 33.760 163.240 34.080 163.280 ;
        RECT 37.900 163.240 38.220 163.280 ;
        RECT 33.760 163.020 34.125 163.240 ;
        RECT 26.950 162.880 27.090 163.020 ;
        RECT 28.700 162.880 29.020 162.940 ;
        RECT 33.835 162.925 34.125 163.020 ;
        RECT 37.855 163.020 38.220 163.240 ;
        RECT 38.935 163.220 39.225 163.265 ;
        RECT 42.515 163.220 42.805 163.265 ;
        RECT 44.350 163.220 44.640 163.265 ;
        RECT 38.935 163.080 44.640 163.220 ;
        RECT 38.935 163.035 39.225 163.080 ;
        RECT 42.515 163.035 42.805 163.080 ;
        RECT 44.350 163.035 44.640 163.080 ;
        RECT 46.655 163.220 46.945 163.265 ;
        RECT 48.940 163.220 49.260 163.280 ;
        RECT 46.655 163.080 49.260 163.220 ;
        RECT 46.655 163.035 46.945 163.080 ;
        RECT 48.940 163.020 49.260 163.080 ;
        RECT 51.255 163.220 51.545 163.265 ;
        RECT 53.080 163.220 53.400 163.280 ;
        RECT 53.630 163.265 53.770 163.420 ;
        RECT 60.440 163.420 65.270 163.560 ;
        RECT 60.440 163.360 60.760 163.420 ;
        RECT 51.255 163.080 53.400 163.220 ;
        RECT 51.255 163.035 51.545 163.080 ;
        RECT 53.080 163.020 53.400 163.080 ;
        RECT 53.555 163.035 53.845 163.265 ;
        RECT 37.855 162.925 38.145 163.020 ;
        RECT 26.950 162.740 29.020 162.880 ;
        RECT 28.700 162.680 29.020 162.740 ;
        RECT 30.535 162.880 31.185 162.925 ;
        RECT 33.835 162.880 34.425 162.925 ;
        RECT 30.535 162.740 34.425 162.880 ;
        RECT 30.535 162.695 31.185 162.740 ;
        RECT 34.135 162.695 34.425 162.740 ;
        RECT 37.555 162.880 38.145 162.925 ;
        RECT 40.795 162.880 41.445 162.925 ;
        RECT 37.555 162.740 41.445 162.880 ;
        RECT 37.555 162.695 37.845 162.740 ;
        RECT 40.795 162.695 41.445 162.740 ;
        RECT 43.435 162.880 43.725 162.925 ;
        RECT 46.180 162.880 46.500 162.940 ;
        RECT 56.715 162.925 57.005 163.240 ;
        RECT 57.795 163.220 58.085 163.265 ;
        RECT 61.375 163.220 61.665 163.265 ;
        RECT 63.210 163.220 63.500 163.265 ;
        RECT 57.795 163.080 63.500 163.220 ;
        RECT 57.795 163.035 58.085 163.080 ;
        RECT 61.375 163.035 61.665 163.080 ;
        RECT 63.210 163.035 63.500 163.080 ;
        RECT 63.660 163.020 63.980 163.280 ;
        RECT 43.435 162.740 46.500 162.880 ;
        RECT 43.435 162.695 43.725 162.740 ;
        RECT 46.180 162.680 46.500 162.740 ;
        RECT 56.415 162.880 57.005 162.925 ;
        RECT 58.600 162.880 58.920 162.940 ;
        RECT 59.655 162.880 60.305 162.925 ;
        RECT 56.415 162.740 60.305 162.880 ;
        RECT 56.415 162.695 56.705 162.740 ;
        RECT 58.600 162.680 58.920 162.740 ;
        RECT 59.655 162.695 60.305 162.740 ;
        RECT 62.280 162.680 62.600 162.940 ;
        RECT 65.130 162.925 65.270 163.420 ;
        RECT 65.590 163.220 65.730 164.100 ;
        RECT 70.880 163.900 71.020 164.100 ;
        RECT 82.520 164.100 83.285 164.240 ;
        RECT 82.520 164.040 82.840 164.100 ;
        RECT 82.995 164.055 83.285 164.100 ;
        RECT 86.215 164.240 86.505 164.285 ;
        RECT 87.580 164.240 87.900 164.300 ;
        RECT 112.880 164.240 113.200 164.300 ;
        RECT 86.215 164.100 87.900 164.240 ;
        RECT 86.215 164.055 86.505 164.100 ;
        RECT 87.580 164.040 87.900 164.100 ;
        RECT 105.610 164.100 113.200 164.240 ;
        RECT 105.610 163.900 105.750 164.100 ;
        RECT 112.880 164.040 113.200 164.100 ;
        RECT 70.880 163.760 105.750 163.900 ;
        RECT 106.455 163.900 106.745 163.945 ;
        RECT 108.740 163.900 109.060 163.960 ;
        RECT 106.455 163.760 109.060 163.900 ;
        RECT 106.455 163.715 106.745 163.760 ;
        RECT 108.740 163.700 109.060 163.760 ;
        RECT 116.215 163.900 116.505 163.945 ;
        RECT 119.335 163.900 119.625 163.945 ;
        RECT 121.225 163.900 121.515 163.945 ;
        RECT 116.215 163.760 121.515 163.900 ;
        RECT 116.215 163.715 116.505 163.760 ;
        RECT 119.335 163.715 119.625 163.760 ;
        RECT 121.225 163.715 121.515 163.760 ;
        RECT 78.380 163.360 78.700 163.620 ;
        RECT 93.560 163.560 93.880 163.620 ;
        RECT 102.315 163.560 102.605 163.605 ;
        RECT 109.215 163.560 109.505 163.605 ;
        RECT 93.560 163.420 109.505 163.560 ;
        RECT 93.560 163.360 93.880 163.420 ;
        RECT 102.315 163.375 102.605 163.420 ;
        RECT 109.215 163.375 109.505 163.420 ;
        RECT 110.120 163.560 110.440 163.620 ;
        RECT 113.355 163.560 113.645 163.605 ;
        RECT 110.120 163.420 113.645 163.560 ;
        RECT 66.435 163.220 66.725 163.265 ;
        RECT 65.590 163.080 66.725 163.220 ;
        RECT 66.435 163.035 66.725 163.080 ;
        RECT 68.260 163.220 68.580 163.280 ;
        RECT 68.735 163.220 69.025 163.265 ;
        RECT 68.260 163.080 69.025 163.220 ;
        RECT 68.260 163.020 68.580 163.080 ;
        RECT 68.735 163.035 69.025 163.080 ;
        RECT 72.860 163.220 73.180 163.280 ;
        RECT 79.315 163.220 79.605 163.265 ;
        RECT 82.075 163.220 82.365 163.265 ;
        RECT 72.860 163.080 79.605 163.220 ;
        RECT 72.860 163.020 73.180 163.080 ;
        RECT 78.930 162.940 79.070 163.080 ;
        RECT 79.315 163.035 79.605 163.080 ;
        RECT 81.690 163.080 82.365 163.220 ;
        RECT 65.055 162.880 65.345 162.925 ;
        RECT 75.160 162.880 75.480 162.940 ;
        RECT 65.055 162.740 75.480 162.880 ;
        RECT 65.055 162.695 65.345 162.740 ;
        RECT 75.160 162.680 75.480 162.740 ;
        RECT 78.840 162.680 79.160 162.940 ;
        RECT 35.600 162.340 35.920 162.600 ;
        RECT 36.060 162.340 36.380 162.600 ;
        RECT 52.620 162.540 52.940 162.600 ;
        RECT 54.935 162.540 55.225 162.585 ;
        RECT 52.620 162.400 55.225 162.540 ;
        RECT 52.620 162.340 52.940 162.400 ;
        RECT 54.935 162.355 55.225 162.400 ;
        RECT 66.880 162.540 67.200 162.600 ;
        RECT 67.355 162.540 67.645 162.585 ;
        RECT 66.880 162.400 67.645 162.540 ;
        RECT 66.880 162.340 67.200 162.400 ;
        RECT 67.355 162.355 67.645 162.400 ;
        RECT 79.775 162.540 80.065 162.585 ;
        RECT 80.680 162.540 81.000 162.600 ;
        RECT 81.690 162.585 81.830 163.080 ;
        RECT 82.075 163.035 82.365 163.080 ;
        RECT 82.980 163.220 83.300 163.280 ;
        RECT 85.295 163.220 85.585 163.265 ;
        RECT 82.980 163.080 85.585 163.220 ;
        RECT 82.980 163.020 83.300 163.080 ;
        RECT 85.295 163.035 85.585 163.080 ;
        RECT 100.920 163.020 101.240 163.280 ;
        RECT 109.290 163.220 109.430 163.375 ;
        RECT 110.120 163.360 110.440 163.420 ;
        RECT 113.355 163.375 113.645 163.420 ;
        RECT 122.095 163.560 122.385 163.605 ;
        RECT 124.380 163.560 124.700 163.620 ;
        RECT 122.095 163.420 124.700 163.560 ;
        RECT 122.095 163.375 122.385 163.420 ;
        RECT 124.380 163.360 124.700 163.420 ;
        RECT 112.420 163.220 112.740 163.280 ;
        RECT 109.290 163.080 112.740 163.220 ;
        RECT 112.420 163.020 112.740 163.080 ;
        RECT 112.880 163.020 113.200 163.280 ;
        RECT 98.160 162.880 98.480 162.940 ;
        RECT 103.235 162.880 103.525 162.925 ;
        RECT 98.160 162.740 103.525 162.880 ;
        RECT 98.160 162.680 98.480 162.740 ;
        RECT 103.235 162.695 103.525 162.740 ;
        RECT 103.695 162.880 103.985 162.925 ;
        RECT 105.980 162.880 106.300 162.940 ;
        RECT 108.755 162.880 109.045 162.925 ;
        RECT 103.695 162.740 109.045 162.880 ;
        RECT 103.695 162.695 103.985 162.740 ;
        RECT 105.980 162.680 106.300 162.740 ;
        RECT 108.755 162.695 109.045 162.740 ;
        RECT 111.500 162.680 111.820 162.940 ;
        RECT 113.340 162.880 113.660 162.940 ;
        RECT 115.135 162.925 115.425 163.240 ;
        RECT 116.215 163.220 116.505 163.265 ;
        RECT 119.795 163.220 120.085 163.265 ;
        RECT 121.630 163.220 121.920 163.265 ;
        RECT 116.215 163.080 121.920 163.220 ;
        RECT 116.215 163.035 116.505 163.080 ;
        RECT 119.795 163.035 120.085 163.080 ;
        RECT 121.630 163.035 121.920 163.080 ;
        RECT 123.460 163.020 123.780 163.280 ;
        RECT 114.835 162.880 115.425 162.925 ;
        RECT 118.075 162.880 118.725 162.925 ;
        RECT 113.340 162.740 118.725 162.880 ;
        RECT 113.340 162.680 113.660 162.740 ;
        RECT 114.835 162.695 115.125 162.740 ;
        RECT 118.075 162.695 118.725 162.740 ;
        RECT 120.715 162.695 121.005 162.925 ;
        RECT 79.775 162.400 81.000 162.540 ;
        RECT 79.775 162.355 80.065 162.400 ;
        RECT 80.680 162.340 81.000 162.400 ;
        RECT 81.615 162.355 81.905 162.585 ;
        RECT 90.800 162.540 91.120 162.600 ;
        RECT 94.495 162.540 94.785 162.585 ;
        RECT 97.240 162.540 97.560 162.600 ;
        RECT 90.800 162.400 97.560 162.540 ;
        RECT 90.800 162.340 91.120 162.400 ;
        RECT 94.495 162.355 94.785 162.400 ;
        RECT 97.240 162.340 97.560 162.400 ;
        RECT 105.060 162.540 105.380 162.600 ;
        RECT 105.535 162.540 105.825 162.585 ;
        RECT 105.060 162.400 105.825 162.540 ;
        RECT 105.060 162.340 105.380 162.400 ;
        RECT 105.535 162.355 105.825 162.400 ;
        RECT 108.295 162.540 108.585 162.585 ;
        RECT 109.660 162.540 109.980 162.600 ;
        RECT 108.295 162.400 109.980 162.540 ;
        RECT 120.790 162.540 120.930 162.695 ;
        RECT 122.555 162.540 122.845 162.585 ;
        RECT 120.790 162.400 122.845 162.540 ;
        RECT 108.295 162.355 108.585 162.400 ;
        RECT 109.660 162.340 109.980 162.400 ;
        RECT 122.555 162.355 122.845 162.400 ;
        RECT 14.370 161.720 127.530 162.200 ;
        RECT 26.400 161.520 26.720 161.580 ;
        RECT 27.335 161.520 27.625 161.565 ;
        RECT 26.400 161.380 27.625 161.520 ;
        RECT 26.400 161.320 26.720 161.380 ;
        RECT 27.335 161.335 27.625 161.380 ;
        RECT 29.620 161.320 29.940 161.580 ;
        RECT 32.855 161.520 33.145 161.565 ;
        RECT 34.220 161.520 34.540 161.580 ;
        RECT 32.855 161.380 34.540 161.520 ;
        RECT 32.855 161.335 33.145 161.380 ;
        RECT 34.220 161.320 34.540 161.380 ;
        RECT 42.500 161.520 42.820 161.580 ;
        RECT 45.275 161.520 45.565 161.565 ;
        RECT 42.500 161.380 45.565 161.520 ;
        RECT 42.500 161.320 42.820 161.380 ;
        RECT 45.275 161.335 45.565 161.380 ;
        RECT 46.180 161.520 46.500 161.580 ;
        RECT 47.575 161.520 47.865 161.565 ;
        RECT 46.180 161.380 47.865 161.520 ;
        RECT 46.180 161.320 46.500 161.380 ;
        RECT 47.575 161.335 47.865 161.380 ;
        RECT 48.940 161.320 49.260 161.580 ;
        RECT 49.400 161.320 49.720 161.580 ;
        RECT 54.000 161.520 54.320 161.580 ;
        RECT 54.935 161.520 55.225 161.565 ;
        RECT 54.000 161.380 55.225 161.520 ;
        RECT 54.000 161.320 54.320 161.380 ;
        RECT 54.935 161.335 55.225 161.380 ;
        RECT 56.775 161.335 57.065 161.565 ;
        RECT 60.455 161.520 60.745 161.565 ;
        RECT 62.280 161.520 62.600 161.580 ;
        RECT 60.455 161.380 62.600 161.520 ;
        RECT 60.455 161.335 60.745 161.380 ;
        RECT 18.580 161.180 18.900 161.240 ;
        RECT 19.910 161.180 20.200 161.225 ;
        RECT 23.170 161.180 23.460 161.225 ;
        RECT 18.580 161.040 23.460 161.180 ;
        RECT 18.580 160.980 18.900 161.040 ;
        RECT 19.910 160.995 20.200 161.040 ;
        RECT 23.170 160.995 23.460 161.040 ;
        RECT 24.090 161.180 24.380 161.225 ;
        RECT 25.950 161.180 26.240 161.225 ;
        RECT 24.090 161.040 26.240 161.180 ;
        RECT 24.090 160.995 24.380 161.040 ;
        RECT 25.950 160.995 26.240 161.040 ;
        RECT 29.175 160.995 29.465 161.225 ;
        RECT 31.000 161.180 31.320 161.240 ;
        RECT 34.695 161.180 34.985 161.225 ;
        RECT 31.000 161.040 34.985 161.180 ;
        RECT 21.770 160.840 22.060 160.885 ;
        RECT 24.090 160.840 24.305 160.995 ;
        RECT 21.770 160.700 24.305 160.840 ;
        RECT 26.860 160.840 27.180 160.900 ;
        RECT 28.700 160.840 29.020 160.900 ;
        RECT 26.860 160.700 29.020 160.840 ;
        RECT 21.770 160.655 22.060 160.700 ;
        RECT 26.860 160.640 27.180 160.700 ;
        RECT 28.700 160.640 29.020 160.700 ;
        RECT 25.035 160.500 25.325 160.545 ;
        RECT 25.480 160.500 25.800 160.560 ;
        RECT 25.035 160.360 25.800 160.500 ;
        RECT 25.035 160.315 25.325 160.360 ;
        RECT 25.480 160.300 25.800 160.360 ;
        RECT 21.770 160.160 22.060 160.205 ;
        RECT 24.550 160.160 24.840 160.205 ;
        RECT 26.410 160.160 26.700 160.205 ;
        RECT 21.770 160.020 26.700 160.160 ;
        RECT 21.770 159.975 22.060 160.020 ;
        RECT 24.550 159.975 24.840 160.020 ;
        RECT 26.410 159.975 26.700 160.020 ;
        RECT 29.250 160.160 29.390 160.995 ;
        RECT 31.000 160.980 31.320 161.040 ;
        RECT 34.695 160.995 34.985 161.040 ;
        RECT 35.155 160.995 35.445 161.225 ;
        RECT 36.060 161.180 36.380 161.240 ;
        RECT 45.735 161.180 46.025 161.225 ;
        RECT 49.490 161.180 49.630 161.320 ;
        RECT 36.060 161.040 46.025 161.180 ;
        RECT 33.760 160.840 34.080 160.900 ;
        RECT 35.230 160.840 35.370 160.995 ;
        RECT 36.060 160.980 36.380 161.040 ;
        RECT 45.735 160.995 46.025 161.040 ;
        RECT 49.030 161.040 49.630 161.180 ;
        RECT 42.975 160.840 43.265 160.885 ;
        RECT 48.495 160.840 48.785 160.885 ;
        RECT 33.760 160.700 35.370 160.840 ;
        RECT 39.830 160.700 40.890 160.840 ;
        RECT 33.760 160.640 34.080 160.700 ;
        RECT 30.540 160.500 30.860 160.560 ;
        RECT 36.075 160.500 36.365 160.545 ;
        RECT 39.830 160.500 39.970 160.700 ;
        RECT 30.540 160.360 39.970 160.500 ;
        RECT 30.540 160.300 30.860 160.360 ;
        RECT 36.075 160.315 36.365 160.360 ;
        RECT 40.215 160.315 40.505 160.545 ;
        RECT 40.750 160.500 40.890 160.700 ;
        RECT 42.975 160.700 48.785 160.840 ;
        RECT 42.975 160.655 43.265 160.700 ;
        RECT 48.495 160.655 48.785 160.700 ;
        RECT 49.030 160.560 49.170 161.040 ;
        RECT 49.400 160.840 49.720 160.900 ;
        RECT 50.795 160.840 51.085 160.885 ;
        RECT 54.475 160.840 54.765 160.885 ;
        RECT 49.400 160.700 54.765 160.840 ;
        RECT 56.850 160.840 56.990 161.335 ;
        RECT 62.280 161.320 62.600 161.380 ;
        RECT 82.520 161.520 82.840 161.580 ;
        RECT 89.665 161.520 89.955 161.565 ;
        RECT 94.480 161.520 94.800 161.580 ;
        RECT 82.520 161.380 84.130 161.520 ;
        RECT 82.520 161.320 82.840 161.380 ;
        RECT 83.990 161.225 84.130 161.380 ;
        RECT 87.670 161.380 94.800 161.520 ;
        RECT 83.915 161.180 84.205 161.225 ;
        RECT 87.670 161.180 87.810 161.380 ;
        RECT 89.665 161.335 89.955 161.380 ;
        RECT 94.480 161.320 94.800 161.380 ;
        RECT 105.535 161.520 105.825 161.565 ;
        RECT 105.980 161.520 106.300 161.580 ;
        RECT 105.535 161.380 106.300 161.520 ;
        RECT 105.535 161.335 105.825 161.380 ;
        RECT 105.980 161.320 106.300 161.380 ;
        RECT 109.660 161.520 109.980 161.580 ;
        RECT 111.515 161.520 111.805 161.565 ;
        RECT 109.660 161.380 111.805 161.520 ;
        RECT 109.660 161.320 109.980 161.380 ;
        RECT 111.515 161.335 111.805 161.380 ;
        RECT 113.815 161.335 114.105 161.565 ;
        RECT 116.100 161.520 116.420 161.580 ;
        RECT 116.575 161.520 116.865 161.565 ;
        RECT 117.020 161.520 117.340 161.580 ;
        RECT 116.100 161.380 117.340 161.520 ;
        RECT 67.890 161.040 70.330 161.180 ;
        RECT 59.535 160.840 59.825 160.885 ;
        RECT 56.850 160.700 59.825 160.840 ;
        RECT 49.400 160.640 49.720 160.700 ;
        RECT 50.795 160.655 51.085 160.700 ;
        RECT 54.475 160.655 54.765 160.700 ;
        RECT 59.535 160.655 59.825 160.700 ;
        RECT 65.975 160.840 66.265 160.885 ;
        RECT 66.420 160.840 66.740 160.900 ;
        RECT 67.890 160.885 68.030 161.040 ;
        RECT 70.190 160.885 70.330 161.040 ;
        RECT 83.915 161.040 87.810 161.180 ;
        RECT 91.670 161.180 91.960 161.225 ;
        RECT 94.020 161.180 94.340 161.240 ;
        RECT 94.930 161.180 95.220 161.225 ;
        RECT 91.670 161.040 95.220 161.180 ;
        RECT 83.915 160.995 84.205 161.040 ;
        RECT 91.670 160.995 91.960 161.040 ;
        RECT 94.020 160.980 94.340 161.040 ;
        RECT 94.930 160.995 95.220 161.040 ;
        RECT 95.850 161.180 96.140 161.225 ;
        RECT 97.710 161.180 98.000 161.225 ;
        RECT 95.850 161.040 98.000 161.180 ;
        RECT 113.890 161.180 114.030 161.335 ;
        RECT 116.100 161.320 116.420 161.380 ;
        RECT 116.575 161.335 116.865 161.380 ;
        RECT 117.020 161.320 117.340 161.380 ;
        RECT 119.320 161.320 119.640 161.580 ;
        RECT 121.160 161.520 121.480 161.580 ;
        RECT 121.635 161.520 121.925 161.565 ;
        RECT 121.160 161.380 121.925 161.520 ;
        RECT 121.160 161.320 121.480 161.380 ;
        RECT 121.635 161.335 121.925 161.380 ;
        RECT 123.460 161.180 123.780 161.240 ;
        RECT 113.890 161.040 123.780 161.180 ;
        RECT 95.850 160.995 96.140 161.040 ;
        RECT 97.710 160.995 98.000 161.040 ;
        RECT 65.975 160.700 67.570 160.840 ;
        RECT 65.975 160.655 66.265 160.700 ;
        RECT 66.420 160.640 66.740 160.700 ;
        RECT 46.655 160.500 46.945 160.545 ;
        RECT 40.750 160.360 46.945 160.500 ;
        RECT 46.655 160.315 46.945 160.360 ;
        RECT 48.940 160.500 49.260 160.560 ;
        RECT 51.255 160.500 51.545 160.545 ;
        RECT 48.940 160.360 51.545 160.500 ;
        RECT 37.440 160.160 37.760 160.220 ;
        RECT 29.250 160.020 37.760 160.160 ;
        RECT 40.290 160.160 40.430 160.315 ;
        RECT 43.435 160.160 43.725 160.205 ;
        RECT 40.290 160.020 43.725 160.160 ;
        RECT 46.730 160.160 46.870 160.315 ;
        RECT 48.940 160.300 49.260 160.360 ;
        RECT 51.255 160.315 51.545 160.360 ;
        RECT 52.175 160.500 52.465 160.545 ;
        RECT 54.015 160.500 54.305 160.545 ;
        RECT 66.880 160.500 67.200 160.560 ;
        RECT 52.175 160.360 67.200 160.500 ;
        RECT 67.430 160.500 67.570 160.700 ;
        RECT 67.815 160.655 68.105 160.885 ;
        RECT 68.275 160.655 68.565 160.885 ;
        RECT 70.115 160.840 70.405 160.885 ;
        RECT 71.020 160.840 71.340 160.900 ;
        RECT 70.115 160.700 71.340 160.840 ;
        RECT 70.115 160.655 70.405 160.700 ;
        RECT 68.350 160.500 68.490 160.655 ;
        RECT 71.020 160.640 71.340 160.700 ;
        RECT 81.615 160.840 81.905 160.885 ;
        RECT 86.215 160.840 86.505 160.885 ;
        RECT 81.615 160.700 85.510 160.840 ;
        RECT 81.615 160.655 81.905 160.700 ;
        RECT 67.430 160.360 68.490 160.500 ;
        RECT 79.760 160.500 80.080 160.560 ;
        RECT 82.535 160.500 82.825 160.545 ;
        RECT 79.760 160.360 82.825 160.500 ;
        RECT 52.175 160.315 52.465 160.360 ;
        RECT 54.015 160.315 54.305 160.360 ;
        RECT 52.250 160.160 52.390 160.315 ;
        RECT 66.880 160.300 67.200 160.360 ;
        RECT 79.760 160.300 80.080 160.360 ;
        RECT 82.535 160.315 82.825 160.360 ;
        RECT 83.455 160.315 83.745 160.545 ;
        RECT 46.730 160.020 52.390 160.160 ;
        RECT 53.080 160.160 53.400 160.220 ;
        RECT 65.055 160.160 65.345 160.205 ;
        RECT 70.560 160.160 70.880 160.220 ;
        RECT 53.080 160.020 70.880 160.160 ;
        RECT 17.905 159.820 18.195 159.865 ;
        RECT 21.340 159.820 21.660 159.880 ;
        RECT 29.250 159.820 29.390 160.020 ;
        RECT 37.440 159.960 37.760 160.020 ;
        RECT 43.435 159.975 43.725 160.020 ;
        RECT 53.080 159.960 53.400 160.020 ;
        RECT 65.055 159.975 65.345 160.020 ;
        RECT 70.560 159.960 70.880 160.020 ;
        RECT 80.680 160.160 81.000 160.220 ;
        RECT 83.530 160.160 83.670 160.315 ;
        RECT 80.680 160.020 83.670 160.160 ;
        RECT 80.680 159.960 81.000 160.020 ;
        RECT 17.905 159.680 29.390 159.820 ;
        RECT 33.760 159.820 34.080 159.880 ;
        RECT 34.680 159.820 35.000 159.880 ;
        RECT 33.760 159.680 35.000 159.820 ;
        RECT 17.905 159.635 18.195 159.680 ;
        RECT 21.340 159.620 21.660 159.680 ;
        RECT 33.760 159.620 34.080 159.680 ;
        RECT 34.680 159.620 35.000 159.680 ;
        RECT 66.880 159.620 67.200 159.880 ;
        RECT 69.195 159.820 69.485 159.865 ;
        RECT 69.640 159.820 69.960 159.880 ;
        RECT 69.195 159.680 69.960 159.820 ;
        RECT 69.195 159.635 69.485 159.680 ;
        RECT 69.640 159.620 69.960 159.680 ;
        RECT 71.035 159.820 71.325 159.865 ;
        RECT 73.780 159.820 74.100 159.880 ;
        RECT 71.035 159.680 74.100 159.820 ;
        RECT 71.035 159.635 71.325 159.680 ;
        RECT 73.780 159.620 74.100 159.680 ;
        RECT 81.155 159.820 81.445 159.865 ;
        RECT 82.980 159.820 83.300 159.880 ;
        RECT 81.155 159.680 83.300 159.820 ;
        RECT 85.370 159.820 85.510 160.700 ;
        RECT 85.830 160.700 86.505 160.840 ;
        RECT 85.830 160.205 85.970 160.700 ;
        RECT 86.215 160.655 86.505 160.700 ;
        RECT 93.530 160.840 93.820 160.885 ;
        RECT 95.850 160.840 96.065 160.995 ;
        RECT 123.460 160.980 123.780 161.040 ;
        RECT 93.530 160.700 96.065 160.840 ;
        RECT 97.240 160.840 97.560 160.900 ;
        RECT 98.635 160.840 98.925 160.885 ;
        RECT 101.855 160.840 102.145 160.885 ;
        RECT 97.240 160.700 102.145 160.840 ;
        RECT 93.530 160.655 93.820 160.700 ;
        RECT 97.240 160.640 97.560 160.700 ;
        RECT 98.635 160.655 98.925 160.700 ;
        RECT 101.855 160.655 102.145 160.700 ;
        RECT 96.780 160.300 97.100 160.560 ;
        RECT 101.930 160.500 102.070 160.655 ;
        RECT 102.300 160.640 102.620 160.900 ;
        RECT 106.915 160.840 107.205 160.885 ;
        RECT 110.120 160.840 110.440 160.900 ;
        RECT 106.915 160.700 110.440 160.840 ;
        RECT 106.915 160.655 107.205 160.700 ;
        RECT 110.120 160.640 110.440 160.700 ;
        RECT 111.975 160.840 112.265 160.885 ;
        RECT 113.800 160.840 114.120 160.900 ;
        RECT 116.115 160.840 116.405 160.885 ;
        RECT 111.975 160.700 116.405 160.840 ;
        RECT 111.975 160.655 112.265 160.700 ;
        RECT 113.800 160.640 114.120 160.700 ;
        RECT 116.115 160.655 116.405 160.700 ;
        RECT 118.860 160.640 119.180 160.900 ;
        RECT 120.700 160.640 121.020 160.900 ;
        RECT 105.520 160.500 105.840 160.560 ;
        RECT 101.930 160.360 105.840 160.500 ;
        RECT 105.520 160.300 105.840 160.360 ;
        RECT 85.755 159.975 86.045 160.205 ;
        RECT 88.500 160.160 88.820 160.220 ;
        RECT 86.290 160.020 88.820 160.160 ;
        RECT 86.290 159.820 86.430 160.020 ;
        RECT 88.500 159.960 88.820 160.020 ;
        RECT 93.530 160.160 93.820 160.205 ;
        RECT 96.310 160.160 96.600 160.205 ;
        RECT 98.170 160.160 98.460 160.205 ;
        RECT 93.530 160.020 98.460 160.160 ;
        RECT 93.530 159.975 93.820 160.020 ;
        RECT 96.310 159.975 96.600 160.020 ;
        RECT 98.170 159.975 98.460 160.020 ;
        RECT 85.370 159.680 86.430 159.820 ;
        RECT 87.135 159.820 87.425 159.865 ;
        RECT 88.040 159.820 88.360 159.880 ;
        RECT 87.135 159.680 88.360 159.820 ;
        RECT 110.210 159.820 110.350 160.640 ;
        RECT 111.055 160.500 111.345 160.545 ;
        RECT 112.420 160.500 112.740 160.560 ;
        RECT 115.195 160.500 115.485 160.545 ;
        RECT 111.055 160.360 115.485 160.500 ;
        RECT 111.055 160.315 111.345 160.360 ;
        RECT 112.420 160.300 112.740 160.360 ;
        RECT 115.195 160.315 115.485 160.360 ;
        RECT 110.580 159.820 110.900 159.880 ;
        RECT 110.210 159.680 110.900 159.820 ;
        RECT 81.155 159.635 81.445 159.680 ;
        RECT 82.980 159.620 83.300 159.680 ;
        RECT 87.135 159.635 87.425 159.680 ;
        RECT 88.040 159.620 88.360 159.680 ;
        RECT 110.580 159.620 110.900 159.680 ;
        RECT 116.560 159.820 116.880 159.880 ;
        RECT 118.415 159.820 118.705 159.865 ;
        RECT 116.560 159.680 118.705 159.820 ;
        RECT 116.560 159.620 116.880 159.680 ;
        RECT 118.415 159.635 118.705 159.680 ;
        RECT 14.370 159.000 127.530 159.480 ;
        RECT 17.675 158.800 17.965 158.845 ;
        RECT 18.580 158.800 18.900 158.860 ;
        RECT 17.675 158.660 18.900 158.800 ;
        RECT 17.675 158.615 17.965 158.660 ;
        RECT 18.580 158.600 18.900 158.660 ;
        RECT 25.480 158.600 25.800 158.860 ;
        RECT 31.000 158.600 31.320 158.860 ;
        RECT 49.400 158.600 49.720 158.860 ;
        RECT 50.320 158.800 50.640 158.860 ;
        RECT 52.620 158.800 52.940 158.860 ;
        RECT 50.320 158.660 52.940 158.800 ;
        RECT 50.320 158.600 50.640 158.660 ;
        RECT 52.620 158.600 52.940 158.660 ;
        RECT 71.035 158.800 71.325 158.845 ;
        RECT 71.480 158.800 71.800 158.860 ;
        RECT 71.035 158.660 71.800 158.800 ;
        RECT 71.035 158.615 71.325 158.660 ;
        RECT 71.480 158.600 71.800 158.660 ;
        RECT 79.760 158.600 80.080 158.860 ;
        RECT 80.680 158.845 81.000 158.860 ;
        RECT 80.680 158.615 81.215 158.845 ;
        RECT 93.115 158.800 93.405 158.845 ;
        RECT 94.020 158.800 94.340 158.860 ;
        RECT 93.115 158.660 94.340 158.800 ;
        RECT 93.115 158.615 93.405 158.660 ;
        RECT 80.680 158.600 81.000 158.615 ;
        RECT 94.020 158.600 94.340 158.660 ;
        RECT 96.780 158.800 97.100 158.860 ;
        RECT 97.255 158.800 97.545 158.845 ;
        RECT 96.780 158.660 97.545 158.800 ;
        RECT 96.780 158.600 97.100 158.660 ;
        RECT 97.255 158.615 97.545 158.660 ;
        RECT 100.000 158.600 100.320 158.860 ;
        RECT 104.155 158.800 104.445 158.845 ;
        RECT 104.600 158.800 104.920 158.860 ;
        RECT 111.960 158.800 112.280 158.860 ;
        RECT 104.155 158.660 104.920 158.800 ;
        RECT 104.155 158.615 104.445 158.660 ;
        RECT 104.600 158.600 104.920 158.660 ;
        RECT 110.210 158.660 112.280 158.800 ;
        RECT 30.540 158.460 30.860 158.520 ;
        RECT 20.970 158.320 30.860 158.460 ;
        RECT 20.970 158.180 21.110 158.320 ;
        RECT 30.540 158.260 30.860 158.320 ;
        RECT 42.360 158.320 53.770 158.460 ;
        RECT 20.880 157.920 21.200 158.180 ;
        RECT 21.340 157.920 21.660 158.180 ;
        RECT 29.620 158.120 29.940 158.180 ;
        RECT 42.360 158.120 42.500 158.320 ;
        RECT 22.580 157.980 29.940 158.120 ;
        RECT 18.135 157.780 18.425 157.825 ;
        RECT 18.595 157.780 18.885 157.825 ;
        RECT 22.580 157.780 22.720 157.980 ;
        RECT 29.620 157.920 29.940 157.980 ;
        RECT 38.910 157.980 42.500 158.120 ;
        RECT 24.575 157.780 24.865 157.825 ;
        RECT 18.135 157.640 22.720 157.780 ;
        RECT 23.730 157.640 24.865 157.780 ;
        RECT 18.135 157.595 18.425 157.640 ;
        RECT 18.595 157.595 18.885 157.640 ;
        RECT 19.040 156.900 19.360 157.160 ;
        RECT 21.800 156.900 22.120 157.160 ;
        RECT 23.730 157.145 23.870 157.640 ;
        RECT 24.575 157.595 24.865 157.640 ;
        RECT 28.255 157.595 28.545 157.825 ;
        RECT 31.920 157.780 32.240 157.840 ;
        RECT 35.600 157.780 35.920 157.840 ;
        RECT 38.910 157.825 39.050 157.980 ;
        RECT 31.920 157.640 35.920 157.780 ;
        RECT 28.330 157.440 28.470 157.595 ;
        RECT 31.920 157.580 32.240 157.640 ;
        RECT 35.600 157.580 35.920 157.640 ;
        RECT 38.835 157.595 39.125 157.825 ;
        RECT 39.755 157.595 40.045 157.825 ;
        RECT 40.215 157.595 40.505 157.825 ;
        RECT 40.675 157.780 40.965 157.825 ;
        RECT 41.580 157.780 41.900 157.840 ;
        RECT 40.675 157.640 41.900 157.780 ;
        RECT 42.360 157.825 42.500 157.980 ;
        RECT 46.655 158.120 46.945 158.165 ;
        RECT 50.320 158.120 50.640 158.180 ;
        RECT 53.630 158.120 53.770 158.320 ;
        RECT 69.195 158.275 69.485 158.505 ;
        RECT 70.560 158.460 70.880 158.520 ;
        RECT 84.790 158.460 85.080 158.505 ;
        RECT 87.570 158.460 87.860 158.505 ;
        RECT 89.430 158.460 89.720 158.505 ;
        RECT 70.560 158.320 78.150 158.460 ;
        RECT 69.270 158.120 69.410 158.275 ;
        RECT 70.560 158.260 70.880 158.320 ;
        RECT 46.655 157.980 50.640 158.120 ;
        RECT 46.655 157.935 46.945 157.980 ;
        RECT 50.320 157.920 50.640 157.980 ;
        RECT 51.790 157.980 53.310 158.120 ;
        RECT 42.360 157.640 42.745 157.825 ;
        RECT 40.675 157.595 40.965 157.640 ;
        RECT 36.060 157.440 36.380 157.500 ;
        RECT 39.830 157.440 39.970 157.595 ;
        RECT 28.330 157.300 39.970 157.440 ;
        RECT 40.290 157.440 40.430 157.595 ;
        RECT 41.580 157.580 41.900 157.640 ;
        RECT 42.455 157.595 42.745 157.640 ;
        RECT 42.960 157.780 43.280 157.840 ;
        RECT 43.435 157.780 43.725 157.825 ;
        RECT 42.960 157.640 43.725 157.780 ;
        RECT 42.960 157.580 43.280 157.640 ;
        RECT 43.435 157.595 43.725 157.640 ;
        RECT 43.895 157.595 44.185 157.825 ;
        RECT 44.355 157.780 44.645 157.825 ;
        RECT 44.800 157.780 45.120 157.840 ;
        RECT 51.790 157.825 51.930 157.980 ;
        RECT 51.715 157.780 52.005 157.825 ;
        RECT 44.355 157.640 52.005 157.780 ;
        RECT 44.355 157.595 44.645 157.640 ;
        RECT 43.970 157.440 44.110 157.595 ;
        RECT 44.800 157.580 45.120 157.640 ;
        RECT 51.715 157.595 52.005 157.640 ;
        RECT 52.175 157.595 52.465 157.825 ;
        RECT 52.250 157.440 52.390 157.595 ;
        RECT 52.620 157.580 52.940 157.840 ;
        RECT 40.290 157.300 52.390 157.440 ;
        RECT 53.170 157.440 53.310 157.980 ;
        RECT 53.630 157.980 72.170 158.120 ;
        RECT 53.630 157.840 53.770 157.980 ;
        RECT 53.540 157.580 53.860 157.840 ;
        RECT 56.760 157.780 57.080 157.840 ;
        RECT 60.915 157.780 61.205 157.825 ;
        RECT 62.295 157.780 62.585 157.825 ;
        RECT 56.760 157.640 62.585 157.780 ;
        RECT 56.760 157.580 57.080 157.640 ;
        RECT 60.915 157.595 61.205 157.640 ;
        RECT 62.295 157.595 62.585 157.640 ;
        RECT 62.740 157.780 63.060 157.840 ;
        RECT 63.675 157.780 63.965 157.825 ;
        RECT 62.740 157.640 63.965 157.780 ;
        RECT 62.740 157.580 63.060 157.640 ;
        RECT 63.675 157.595 63.965 157.640 ;
        RECT 68.275 157.780 68.565 157.825 ;
        RECT 69.180 157.780 69.500 157.840 ;
        RECT 70.100 157.780 70.420 157.840 ;
        RECT 72.030 157.825 72.170 157.980 ;
        RECT 68.275 157.640 70.420 157.780 ;
        RECT 68.275 157.595 68.565 157.640 ;
        RECT 69.180 157.580 69.500 157.640 ;
        RECT 70.100 157.580 70.420 157.640 ;
        RECT 71.955 157.595 72.245 157.825 ;
        RECT 72.030 157.440 72.170 157.595 ;
        RECT 72.860 157.580 73.180 157.840 ;
        RECT 73.410 157.825 73.550 158.320 ;
        RECT 76.080 158.120 76.400 158.180 ;
        RECT 76.080 157.980 77.690 158.120 ;
        RECT 76.080 157.920 76.400 157.980 ;
        RECT 73.335 157.595 73.625 157.825 ;
        RECT 73.780 157.580 74.100 157.840 ;
        RECT 77.550 157.825 77.690 157.980 ;
        RECT 78.010 157.825 78.150 158.320 ;
        RECT 84.790 158.320 89.720 158.460 ;
        RECT 84.790 158.275 85.080 158.320 ;
        RECT 87.570 158.275 87.860 158.320 ;
        RECT 89.430 158.275 89.720 158.320 ;
        RECT 106.455 158.460 106.745 158.505 ;
        RECT 109.200 158.460 109.520 158.520 ;
        RECT 106.455 158.320 109.520 158.460 ;
        RECT 106.455 158.275 106.745 158.320 ;
        RECT 109.200 158.260 109.520 158.320 ;
        RECT 88.040 157.920 88.360 158.180 ;
        RECT 88.500 158.120 88.820 158.180 ;
        RECT 88.500 157.980 92.870 158.120 ;
        RECT 88.500 157.920 88.820 157.980 ;
        RECT 76.555 157.780 76.845 157.825 ;
        RECT 76.170 157.640 76.845 157.780 ;
        RECT 76.170 157.500 76.310 157.640 ;
        RECT 76.555 157.595 76.845 157.640 ;
        RECT 77.475 157.595 77.765 157.825 ;
        RECT 77.935 157.595 78.225 157.825 ;
        RECT 78.395 157.780 78.685 157.825 ;
        RECT 78.840 157.780 79.160 157.840 ;
        RECT 81.600 157.780 81.920 157.840 ;
        RECT 78.395 157.640 81.920 157.780 ;
        RECT 78.395 157.595 78.685 157.640 ;
        RECT 76.080 157.440 76.400 157.500 ;
        RECT 53.170 157.300 61.130 157.440 ;
        RECT 72.030 157.300 76.400 157.440 ;
        RECT 78.010 157.440 78.150 157.595 ;
        RECT 78.840 157.580 79.160 157.640 ;
        RECT 81.600 157.580 81.920 157.640 ;
        RECT 84.790 157.780 85.080 157.825 ;
        RECT 89.895 157.780 90.185 157.825 ;
        RECT 90.800 157.780 91.120 157.840 ;
        RECT 92.730 157.825 92.870 157.980 ;
        RECT 84.790 157.640 87.325 157.780 ;
        RECT 84.790 157.595 85.080 157.640 ;
        RECT 82.060 157.440 82.380 157.500 ;
        RECT 82.980 157.485 83.300 157.500 ;
        RECT 87.110 157.485 87.325 157.640 ;
        RECT 89.895 157.640 91.120 157.780 ;
        RECT 89.895 157.595 90.185 157.640 ;
        RECT 90.800 157.580 91.120 157.640 ;
        RECT 92.655 157.595 92.945 157.825 ;
        RECT 78.010 157.300 82.380 157.440 ;
        RECT 36.060 157.240 36.380 157.300 ;
        RECT 43.050 157.160 43.190 157.300 ;
        RECT 23.655 156.915 23.945 157.145 ;
        RECT 34.680 156.900 35.000 157.160 ;
        RECT 42.040 156.900 42.360 157.160 ;
        RECT 42.960 156.900 43.280 157.160 ;
        RECT 45.720 156.900 46.040 157.160 ;
        RECT 49.860 157.100 50.180 157.160 ;
        RECT 50.335 157.100 50.625 157.145 ;
        RECT 49.860 156.960 50.625 157.100 ;
        RECT 52.250 157.100 52.390 157.300 ;
        RECT 53.080 157.100 53.400 157.160 ;
        RECT 52.250 156.960 53.400 157.100 ;
        RECT 49.860 156.900 50.180 156.960 ;
        RECT 50.335 156.915 50.625 156.960 ;
        RECT 53.080 156.900 53.400 156.960 ;
        RECT 58.600 157.100 58.920 157.160 ;
        RECT 60.455 157.100 60.745 157.145 ;
        RECT 58.600 156.960 60.745 157.100 ;
        RECT 60.990 157.100 61.130 157.300 ;
        RECT 76.080 157.240 76.400 157.300 ;
        RECT 82.060 157.240 82.380 157.300 ;
        RECT 82.930 157.440 83.300 157.485 ;
        RECT 86.190 157.440 86.480 157.485 ;
        RECT 82.930 157.300 86.480 157.440 ;
        RECT 82.930 157.255 83.300 157.300 ;
        RECT 86.190 157.255 86.480 157.300 ;
        RECT 87.110 157.440 87.400 157.485 ;
        RECT 88.970 157.440 89.260 157.485 ;
        RECT 87.110 157.300 89.260 157.440 ;
        RECT 92.730 157.440 92.870 157.595 ;
        RECT 96.320 157.580 96.640 157.840 ;
        RECT 99.555 157.595 99.845 157.825 ;
        RECT 94.940 157.440 95.260 157.500 ;
        RECT 99.630 157.440 99.770 157.595 ;
        RECT 105.060 157.580 105.380 157.840 ;
        RECT 105.535 157.780 105.825 157.825 ;
        RECT 108.740 157.780 109.060 157.840 ;
        RECT 105.535 157.640 109.060 157.780 ;
        RECT 105.535 157.595 105.825 157.640 ;
        RECT 108.740 157.580 109.060 157.640 ;
        RECT 109.200 157.580 109.520 157.840 ;
        RECT 109.660 157.580 109.980 157.840 ;
        RECT 110.210 157.825 110.350 158.660 ;
        RECT 111.960 158.600 112.280 158.660 ;
        RECT 119.335 158.800 119.625 158.845 ;
        RECT 120.700 158.800 121.020 158.860 ;
        RECT 119.335 158.660 121.020 158.800 ;
        RECT 119.335 158.615 119.625 158.660 ;
        RECT 120.700 158.600 121.020 158.660 ;
        RECT 116.560 157.920 116.880 158.180 ;
        RECT 110.135 157.595 110.425 157.825 ;
        RECT 111.055 157.780 111.345 157.825 ;
        RECT 111.500 157.780 111.820 157.840 ;
        RECT 111.055 157.640 111.820 157.780 ;
        RECT 111.055 157.595 111.345 157.640 ;
        RECT 111.500 157.580 111.820 157.640 ;
        RECT 111.960 157.440 112.280 157.500 ;
        RECT 92.730 157.300 112.280 157.440 ;
        RECT 87.110 157.255 87.400 157.300 ;
        RECT 88.970 157.255 89.260 157.300 ;
        RECT 82.980 157.240 83.300 157.255 ;
        RECT 94.940 157.240 95.260 157.300 ;
        RECT 111.960 157.240 112.280 157.300 ;
        RECT 73.780 157.100 74.100 157.160 ;
        RECT 60.990 156.960 74.100 157.100 ;
        RECT 58.600 156.900 58.920 156.960 ;
        RECT 60.455 156.915 60.745 156.960 ;
        RECT 73.780 156.900 74.100 156.960 ;
        RECT 75.175 157.100 75.465 157.145 ;
        RECT 75.620 157.100 75.940 157.160 ;
        RECT 75.175 156.960 75.940 157.100 ;
        RECT 75.175 156.915 75.465 156.960 ;
        RECT 75.620 156.900 75.940 156.960 ;
        RECT 107.835 157.100 108.125 157.145 ;
        RECT 108.740 157.100 109.060 157.160 ;
        RECT 107.835 156.960 109.060 157.100 ;
        RECT 107.835 156.915 108.125 156.960 ;
        RECT 108.740 156.900 109.060 156.960 ;
        RECT 14.370 156.280 127.530 156.760 ;
        RECT 16.985 156.080 17.275 156.125 ;
        RECT 21.800 156.080 22.120 156.140 ;
        RECT 33.300 156.080 33.620 156.140 ;
        RECT 34.235 156.080 34.525 156.125 ;
        RECT 16.985 155.940 32.610 156.080 ;
        RECT 16.985 155.895 17.275 155.940 ;
        RECT 21.800 155.880 22.120 155.940 ;
        RECT 19.040 155.785 19.360 155.800 ;
        RECT 18.990 155.740 19.360 155.785 ;
        RECT 22.250 155.740 22.540 155.785 ;
        RECT 18.990 155.600 22.540 155.740 ;
        RECT 18.990 155.555 19.360 155.600 ;
        RECT 22.250 155.555 22.540 155.600 ;
        RECT 23.170 155.740 23.460 155.785 ;
        RECT 25.030 155.740 25.320 155.785 ;
        RECT 23.170 155.600 25.320 155.740 ;
        RECT 32.470 155.740 32.610 155.940 ;
        RECT 33.300 155.940 34.525 156.080 ;
        RECT 33.300 155.880 33.620 155.940 ;
        RECT 34.235 155.895 34.525 155.940 ;
        RECT 34.680 155.880 35.000 156.140 ;
        RECT 41.580 156.080 41.900 156.140 ;
        RECT 44.800 156.080 45.120 156.140 ;
        RECT 40.290 155.940 45.120 156.080 ;
        RECT 32.470 155.600 34.450 155.740 ;
        RECT 23.170 155.555 23.460 155.600 ;
        RECT 25.030 155.555 25.320 155.600 ;
        RECT 19.040 155.540 19.360 155.555 ;
        RECT 20.850 155.400 21.140 155.445 ;
        RECT 23.170 155.400 23.385 155.555 ;
        RECT 20.850 155.260 23.385 155.400 ;
        RECT 25.955 155.400 26.245 155.445 ;
        RECT 26.860 155.400 27.180 155.460 ;
        RECT 25.955 155.260 27.180 155.400 ;
        RECT 20.850 155.215 21.140 155.260 ;
        RECT 25.955 155.215 26.245 155.260 ;
        RECT 26.860 155.200 27.180 155.260 ;
        RECT 27.320 155.200 27.640 155.460 ;
        RECT 31.000 155.400 31.320 155.460 ;
        RECT 33.300 155.400 33.620 155.460 ;
        RECT 31.000 155.260 33.620 155.400 ;
        RECT 31.000 155.200 31.320 155.260 ;
        RECT 33.300 155.200 33.620 155.260 ;
        RECT 24.115 155.060 24.405 155.105 ;
        RECT 30.540 155.060 30.860 155.120 ;
        RECT 33.760 155.060 34.080 155.120 ;
        RECT 24.115 154.920 26.630 155.060 ;
        RECT 24.115 154.875 24.405 154.920 ;
        RECT 26.490 154.765 26.630 154.920 ;
        RECT 30.540 154.920 34.080 155.060 ;
        RECT 34.310 155.060 34.450 155.600 ;
        RECT 40.290 155.400 40.430 155.940 ;
        RECT 41.580 155.880 41.900 155.940 ;
        RECT 44.800 155.880 45.120 155.940 ;
        RECT 48.940 156.080 49.260 156.140 ;
        RECT 50.320 156.080 50.640 156.140 ;
        RECT 66.880 156.080 67.200 156.140 ;
        RECT 102.300 156.080 102.620 156.140 ;
        RECT 108.280 156.080 108.600 156.140 ;
        RECT 111.500 156.080 111.820 156.140 ;
        RECT 48.940 155.940 49.630 156.080 ;
        RECT 48.940 155.880 49.260 155.940 ;
        RECT 40.660 155.740 40.980 155.800 ;
        RECT 44.890 155.740 45.030 155.880 ;
        RECT 40.660 155.600 43.190 155.740 ;
        RECT 40.660 155.540 40.980 155.600 ;
        RECT 41.135 155.400 41.425 155.445 ;
        RECT 40.290 155.260 41.425 155.400 ;
        RECT 41.135 155.215 41.425 155.260 ;
        RECT 41.580 155.200 41.900 155.460 ;
        RECT 43.050 155.445 43.190 155.600 ;
        RECT 44.890 155.600 48.710 155.740 ;
        RECT 44.890 155.445 45.030 155.600 ;
        RECT 42.055 155.215 42.345 155.445 ;
        RECT 42.975 155.215 43.265 155.445 ;
        RECT 44.815 155.215 45.105 155.445 ;
        RECT 45.260 155.215 45.550 155.445 ;
        RECT 45.760 155.215 46.050 155.445 ;
        RECT 42.130 155.060 42.270 155.215 ;
        RECT 34.310 154.920 42.270 155.060 ;
        RECT 43.420 155.060 43.740 155.120 ;
        RECT 45.350 155.060 45.490 155.215 ;
        RECT 43.420 154.920 45.490 155.060 ;
        RECT 30.540 154.860 30.860 154.920 ;
        RECT 33.760 154.860 34.080 154.920 ;
        RECT 43.420 154.860 43.740 154.920 ;
        RECT 20.850 154.720 21.140 154.765 ;
        RECT 23.630 154.720 23.920 154.765 ;
        RECT 25.490 154.720 25.780 154.765 ;
        RECT 20.850 154.580 25.780 154.720 ;
        RECT 20.850 154.535 21.140 154.580 ;
        RECT 23.630 154.535 23.920 154.580 ;
        RECT 25.490 154.535 25.780 154.580 ;
        RECT 26.415 154.535 26.705 154.765 ;
        RECT 31.920 154.720 32.240 154.780 ;
        RECT 45.810 154.720 45.950 155.215 ;
        RECT 46.640 155.200 46.960 155.460 ;
        RECT 48.570 155.445 48.710 155.600 ;
        RECT 49.490 155.445 49.630 155.940 ;
        RECT 50.320 155.940 84.820 156.080 ;
        RECT 50.320 155.880 50.640 155.940 ;
        RECT 66.880 155.880 67.200 155.940 ;
        RECT 53.080 155.740 53.400 155.800 ;
        RECT 58.600 155.785 58.920 155.800 ;
        RECT 49.950 155.600 53.400 155.740 ;
        RECT 48.495 155.215 48.785 155.445 ;
        RECT 48.955 155.215 49.245 155.445 ;
        RECT 49.415 155.215 49.705 155.445 ;
        RECT 49.030 155.060 49.170 155.215 ;
        RECT 49.950 155.060 50.090 155.600 ;
        RECT 53.080 155.540 53.400 155.600 ;
        RECT 55.330 155.740 55.620 155.785 ;
        RECT 58.590 155.740 58.920 155.785 ;
        RECT 55.330 155.600 58.920 155.740 ;
        RECT 55.330 155.555 55.620 155.600 ;
        RECT 58.590 155.555 58.920 155.600 ;
        RECT 58.600 155.540 58.920 155.555 ;
        RECT 59.510 155.740 59.800 155.785 ;
        RECT 61.370 155.740 61.660 155.785 ;
        RECT 59.510 155.600 61.660 155.740 ;
        RECT 59.510 155.555 59.800 155.600 ;
        RECT 61.370 155.555 61.660 155.600 ;
        RECT 73.780 155.740 74.100 155.800 ;
        RECT 80.680 155.740 81.000 155.800 ;
        RECT 73.780 155.600 78.150 155.740 ;
        RECT 50.335 155.400 50.625 155.445 ;
        RECT 53.540 155.400 53.860 155.460 ;
        RECT 50.335 155.260 53.860 155.400 ;
        RECT 50.335 155.215 50.625 155.260 ;
        RECT 49.030 154.920 50.090 155.060 ;
        RECT 31.920 154.580 45.950 154.720 ;
        RECT 46.640 154.720 46.960 154.780 ;
        RECT 50.410 154.720 50.550 155.215 ;
        RECT 53.540 155.200 53.860 155.260 ;
        RECT 57.190 155.400 57.480 155.445 ;
        RECT 59.510 155.400 59.725 155.555 ;
        RECT 73.780 155.540 74.100 155.600 ;
        RECT 78.010 155.460 78.150 155.600 ;
        RECT 79.390 155.600 81.000 155.740 ;
        RECT 84.680 155.740 84.820 155.940 ;
        RECT 102.300 155.940 111.820 156.080 ;
        RECT 102.300 155.880 102.620 155.940 ;
        RECT 102.760 155.740 103.080 155.800 ;
        RECT 84.680 155.600 97.930 155.740 ;
        RECT 57.190 155.260 59.725 155.400 ;
        RECT 62.295 155.400 62.585 155.445 ;
        RECT 63.660 155.400 63.980 155.460 ;
        RECT 62.295 155.260 63.980 155.400 ;
        RECT 57.190 155.215 57.480 155.260 ;
        RECT 62.295 155.215 62.585 155.260 ;
        RECT 63.660 155.200 63.980 155.260 ;
        RECT 74.240 155.200 74.560 155.460 ;
        RECT 77.920 155.200 78.240 155.460 ;
        RECT 78.380 155.200 78.700 155.460 ;
        RECT 78.855 155.400 79.145 155.445 ;
        RECT 79.390 155.400 79.530 155.600 ;
        RECT 80.680 155.540 81.000 155.600 ;
        RECT 78.855 155.260 79.530 155.400 ;
        RECT 78.855 155.215 79.145 155.260 ;
        RECT 79.775 155.215 80.065 155.445 ;
        RECT 60.455 155.060 60.745 155.105 ;
        RECT 60.900 155.060 61.220 155.120 ;
        RECT 60.455 154.920 61.220 155.060 ;
        RECT 60.455 154.875 60.745 154.920 ;
        RECT 60.900 154.860 61.220 154.920 ;
        RECT 65.500 154.860 65.820 155.120 ;
        RECT 76.080 155.060 76.400 155.120 ;
        RECT 79.850 155.060 79.990 155.215 ;
        RECT 81.600 155.200 81.920 155.460 ;
        RECT 82.060 155.200 82.380 155.460 ;
        RECT 82.520 155.200 82.840 155.460 ;
        RECT 83.455 155.215 83.745 155.445 ;
        RECT 84.360 155.400 84.680 155.460 ;
        RECT 97.255 155.400 97.545 155.445 ;
        RECT 84.360 155.260 97.545 155.400 ;
        RECT 83.530 155.060 83.670 155.215 ;
        RECT 84.360 155.200 84.680 155.260 ;
        RECT 97.255 155.215 97.545 155.260 ;
        RECT 76.080 154.920 83.670 155.060 ;
        RECT 76.080 154.860 76.400 154.920 ;
        RECT 46.640 154.580 50.550 154.720 ;
        RECT 57.190 154.720 57.480 154.765 ;
        RECT 59.970 154.720 60.260 154.765 ;
        RECT 61.830 154.720 62.120 154.765 ;
        RECT 57.190 154.580 62.120 154.720 ;
        RECT 31.920 154.520 32.240 154.580 ;
        RECT 46.640 154.520 46.960 154.580 ;
        RECT 57.190 154.535 57.480 154.580 ;
        RECT 59.970 154.535 60.260 154.580 ;
        RECT 61.830 154.535 62.120 154.580 ;
        RECT 78.380 154.720 78.700 154.780 ;
        RECT 82.060 154.720 82.380 154.780 ;
        RECT 78.380 154.580 82.380 154.720 ;
        RECT 97.330 154.720 97.470 155.215 ;
        RECT 97.790 155.060 97.930 155.600 ;
        RECT 102.760 155.600 106.210 155.740 ;
        RECT 102.760 155.540 103.080 155.600 ;
        RECT 98.160 155.200 98.480 155.460 ;
        RECT 98.620 155.200 98.940 155.460 ;
        RECT 99.095 155.400 99.385 155.445 ;
        RECT 104.615 155.400 104.905 155.445 ;
        RECT 99.095 155.260 104.905 155.400 ;
        RECT 99.095 155.215 99.385 155.260 ;
        RECT 104.615 155.215 104.905 155.260 ;
        RECT 99.170 155.060 99.310 155.215 ;
        RECT 97.790 154.920 99.310 155.060 ;
        RECT 102.300 154.720 102.620 154.780 ;
        RECT 97.330 154.580 102.620 154.720 ;
        RECT 78.380 154.520 78.700 154.580 ;
        RECT 82.060 154.520 82.380 154.580 ;
        RECT 102.300 154.520 102.620 154.580 ;
        RECT 35.600 154.380 35.920 154.440 ;
        RECT 36.535 154.380 36.825 154.425 ;
        RECT 35.600 154.240 36.825 154.380 ;
        RECT 35.600 154.180 35.920 154.240 ;
        RECT 36.535 154.195 36.825 154.240 ;
        RECT 39.740 154.180 40.060 154.440 ;
        RECT 43.420 154.180 43.740 154.440 ;
        RECT 44.800 154.380 45.120 154.440 ;
        RECT 46.730 154.380 46.870 154.520 ;
        RECT 44.800 154.240 46.870 154.380 ;
        RECT 47.115 154.380 47.405 154.425 ;
        RECT 48.940 154.380 49.260 154.440 ;
        RECT 53.540 154.425 53.860 154.440 ;
        RECT 47.115 154.240 49.260 154.380 ;
        RECT 44.800 154.180 45.120 154.240 ;
        RECT 47.115 154.195 47.405 154.240 ;
        RECT 48.940 154.180 49.260 154.240 ;
        RECT 53.325 154.195 53.860 154.425 ;
        RECT 53.540 154.180 53.860 154.195 ;
        RECT 54.000 154.380 54.320 154.440 ;
        RECT 69.640 154.380 69.960 154.440 ;
        RECT 54.000 154.240 69.960 154.380 ;
        RECT 54.000 154.180 54.320 154.240 ;
        RECT 69.640 154.180 69.960 154.240 ;
        RECT 76.080 154.380 76.400 154.440 ;
        RECT 76.555 154.380 76.845 154.425 ;
        RECT 76.080 154.240 76.845 154.380 ;
        RECT 76.080 154.180 76.400 154.240 ;
        RECT 76.555 154.195 76.845 154.240 ;
        RECT 80.220 154.180 80.540 154.440 ;
        RECT 99.540 154.380 99.860 154.440 ;
        RECT 100.475 154.380 100.765 154.425 ;
        RECT 99.540 154.240 100.765 154.380 ;
        RECT 99.540 154.180 99.860 154.240 ;
        RECT 100.475 154.195 100.765 154.240 ;
        RECT 103.235 154.380 103.525 154.425 ;
        RECT 103.680 154.380 104.000 154.440 ;
        RECT 103.235 154.240 104.000 154.380 ;
        RECT 104.690 154.380 104.830 155.215 ;
        RECT 105.060 155.200 105.380 155.460 ;
        RECT 105.535 155.400 105.825 155.445 ;
        RECT 106.070 155.400 106.210 155.600 ;
        RECT 106.530 155.445 106.670 155.940 ;
        RECT 108.280 155.880 108.600 155.940 ;
        RECT 111.500 155.880 111.820 155.940 ;
        RECT 110.580 155.740 110.900 155.800 ;
        RECT 107.910 155.600 110.900 155.740 ;
        RECT 107.910 155.445 108.050 155.600 ;
        RECT 110.580 155.540 110.900 155.600 ;
        RECT 105.535 155.260 106.210 155.400 ;
        RECT 106.455 155.400 106.745 155.445 ;
        RECT 106.915 155.400 107.205 155.445 ;
        RECT 106.455 155.260 107.205 155.400 ;
        RECT 105.535 155.215 105.825 155.260 ;
        RECT 106.455 155.215 106.745 155.260 ;
        RECT 106.915 155.215 107.205 155.260 ;
        RECT 107.835 155.215 108.125 155.445 ;
        RECT 108.295 155.215 108.585 155.445 ;
        RECT 108.755 155.400 109.045 155.445 ;
        RECT 109.200 155.400 109.520 155.460 ;
        RECT 108.755 155.260 109.520 155.400 ;
        RECT 108.755 155.215 109.045 155.260 ;
        RECT 105.150 155.060 105.290 155.200 ;
        RECT 108.370 155.060 108.510 155.215 ;
        RECT 105.150 154.920 108.510 155.060 ;
        RECT 108.830 154.720 108.970 155.215 ;
        RECT 109.200 155.200 109.520 155.260 ;
        RECT 112.880 155.400 113.200 155.460 ;
        RECT 116.115 155.400 116.405 155.445 ;
        RECT 112.880 155.260 116.405 155.400 ;
        RECT 112.880 155.200 113.200 155.260 ;
        RECT 116.115 155.215 116.405 155.260 ;
        RECT 117.480 154.860 117.800 155.120 ;
        RECT 108.370 154.580 108.970 154.720 ;
        RECT 106.440 154.380 106.760 154.440 ;
        RECT 108.370 154.380 108.510 154.580 ;
        RECT 104.690 154.240 108.510 154.380 ;
        RECT 110.135 154.380 110.425 154.425 ;
        RECT 110.580 154.380 110.900 154.440 ;
        RECT 110.135 154.240 110.900 154.380 ;
        RECT 103.235 154.195 103.525 154.240 ;
        RECT 103.680 154.180 104.000 154.240 ;
        RECT 106.440 154.180 106.760 154.240 ;
        RECT 110.135 154.195 110.425 154.240 ;
        RECT 110.580 154.180 110.900 154.240 ;
        RECT 14.370 153.560 127.530 154.040 ;
        RECT 23.655 153.360 23.945 153.405 ;
        RECT 27.320 153.360 27.640 153.420 ;
        RECT 23.655 153.220 27.640 153.360 ;
        RECT 23.655 153.175 23.945 153.220 ;
        RECT 27.320 153.160 27.640 153.220 ;
        RECT 70.100 153.360 70.420 153.420 ;
        RECT 71.955 153.360 72.245 153.405 ;
        RECT 70.100 153.220 72.245 153.360 ;
        RECT 70.100 153.160 70.420 153.220 ;
        RECT 71.955 153.175 72.245 153.220 ;
        RECT 73.320 153.160 73.640 153.420 ;
        RECT 98.620 153.360 98.940 153.420 ;
        RECT 84.680 153.220 98.940 153.360 ;
        RECT 33.730 153.020 34.020 153.065 ;
        RECT 36.510 153.020 36.800 153.065 ;
        RECT 38.370 153.020 38.660 153.065 ;
        RECT 54.000 153.020 54.320 153.080 ;
        RECT 33.730 152.880 38.660 153.020 ;
        RECT 33.730 152.835 34.020 152.880 ;
        RECT 36.510 152.835 36.800 152.880 ;
        RECT 38.370 152.835 38.660 152.880 ;
        RECT 42.130 152.880 54.320 153.020 ;
        RECT 20.880 152.480 21.200 152.740 ;
        RECT 21.355 152.680 21.645 152.725 ;
        RECT 21.800 152.680 22.120 152.740 ;
        RECT 21.355 152.540 22.120 152.680 ;
        RECT 21.355 152.495 21.645 152.540 ;
        RECT 21.800 152.480 22.120 152.540 ;
        RECT 36.980 152.480 37.300 152.740 ;
        RECT 37.440 152.680 37.760 152.740 ;
        RECT 37.440 152.540 41.810 152.680 ;
        RECT 37.440 152.480 37.760 152.540 ;
        RECT 33.730 152.340 34.020 152.385 ;
        RECT 36.520 152.340 36.840 152.400 ;
        RECT 41.670 152.385 41.810 152.540 ;
        RECT 38.835 152.340 39.125 152.385 ;
        RECT 33.730 152.200 36.265 152.340 ;
        RECT 33.730 152.155 34.020 152.200 ;
        RECT 31.870 152.000 32.160 152.045 ;
        RECT 33.300 152.000 33.620 152.060 ;
        RECT 36.050 152.045 36.265 152.200 ;
        RECT 36.520 152.200 39.125 152.340 ;
        RECT 36.520 152.140 36.840 152.200 ;
        RECT 38.835 152.155 39.125 152.200 ;
        RECT 40.675 152.155 40.965 152.385 ;
        RECT 41.135 152.155 41.425 152.385 ;
        RECT 41.595 152.155 41.885 152.385 ;
        RECT 35.130 152.000 35.420 152.045 ;
        RECT 31.870 151.860 35.420 152.000 ;
        RECT 31.870 151.815 32.160 151.860 ;
        RECT 33.300 151.800 33.620 151.860 ;
        RECT 35.130 151.815 35.420 151.860 ;
        RECT 36.050 152.000 36.340 152.045 ;
        RECT 37.910 152.000 38.200 152.045 ;
        RECT 36.050 151.860 38.200 152.000 ;
        RECT 36.050 151.815 36.340 151.860 ;
        RECT 37.910 151.815 38.200 151.860 ;
        RECT 21.815 151.660 22.105 151.705 ;
        RECT 22.260 151.660 22.580 151.720 ;
        RECT 21.815 151.520 22.580 151.660 ;
        RECT 21.815 151.475 22.105 151.520 ;
        RECT 22.260 151.460 22.580 151.520 ;
        RECT 29.865 151.660 30.155 151.705 ;
        RECT 31.000 151.660 31.320 151.720 ;
        RECT 29.865 151.520 31.320 151.660 ;
        RECT 29.865 151.475 30.155 151.520 ;
        RECT 31.000 151.460 31.320 151.520 ;
        RECT 34.680 151.660 35.000 151.720 ;
        RECT 39.295 151.660 39.585 151.705 ;
        RECT 34.680 151.520 39.585 151.660 ;
        RECT 40.750 151.660 40.890 152.155 ;
        RECT 41.210 152.000 41.350 152.155 ;
        RECT 42.130 152.000 42.270 152.880 ;
        RECT 54.000 152.820 54.320 152.880 ;
        RECT 62.250 153.020 62.540 153.065 ;
        RECT 65.030 153.020 65.320 153.065 ;
        RECT 66.890 153.020 67.180 153.065 ;
        RECT 62.250 152.880 67.180 153.020 ;
        RECT 62.250 152.835 62.540 152.880 ;
        RECT 65.030 152.835 65.320 152.880 ;
        RECT 66.890 152.835 67.180 152.880 ;
        RECT 69.640 153.020 69.960 153.080 ;
        RECT 84.680 153.020 84.820 153.220 ;
        RECT 98.620 153.160 98.940 153.220 ;
        RECT 102.760 153.360 103.080 153.420 ;
        RECT 103.235 153.360 103.525 153.405 ;
        RECT 109.660 153.360 109.980 153.420 ;
        RECT 102.760 153.220 103.525 153.360 ;
        RECT 102.760 153.160 103.080 153.220 ;
        RECT 103.235 153.175 103.525 153.220 ;
        RECT 106.990 153.220 109.980 153.360 ;
        RECT 69.640 152.880 84.820 153.020 ;
        RECT 90.310 153.020 90.600 153.065 ;
        RECT 93.090 153.020 93.380 153.065 ;
        RECT 94.950 153.020 95.240 153.065 ;
        RECT 90.310 152.880 95.240 153.020 ;
        RECT 98.710 153.020 98.850 153.160 ;
        RECT 105.060 153.020 105.380 153.080 ;
        RECT 98.710 152.880 105.380 153.020 ;
        RECT 69.640 152.820 69.960 152.880 ;
        RECT 90.310 152.835 90.600 152.880 ;
        RECT 93.090 152.835 93.380 152.880 ;
        RECT 94.950 152.835 95.240 152.880 ;
        RECT 105.060 152.820 105.380 152.880 ;
        RECT 64.120 152.680 64.440 152.740 ;
        RECT 69.180 152.680 69.500 152.740 ;
        RECT 73.780 152.680 74.100 152.740 ;
        RECT 74.255 152.680 74.545 152.725 ;
        RECT 64.120 152.540 68.950 152.680 ;
        RECT 64.120 152.480 64.440 152.540 ;
        RECT 42.515 152.340 42.805 152.385 ;
        RECT 44.340 152.340 44.660 152.400 ;
        RECT 42.515 152.200 44.660 152.340 ;
        RECT 42.515 152.155 42.805 152.200 ;
        RECT 44.340 152.140 44.660 152.200 ;
        RECT 50.780 152.340 51.100 152.400 ;
        RECT 56.760 152.340 57.080 152.400 ;
        RECT 50.780 152.200 57.080 152.340 ;
        RECT 50.780 152.140 51.100 152.200 ;
        RECT 56.760 152.140 57.080 152.200 ;
        RECT 62.250 152.340 62.540 152.385 ;
        RECT 62.250 152.200 64.785 152.340 ;
        RECT 62.250 152.155 62.540 152.200 ;
        RECT 42.960 152.000 43.280 152.060 ;
        RECT 64.570 152.045 64.785 152.200 ;
        RECT 65.500 152.140 65.820 152.400 ;
        RECT 67.355 152.340 67.645 152.385 ;
        RECT 68.260 152.340 68.580 152.400 ;
        RECT 67.355 152.200 68.580 152.340 ;
        RECT 68.810 152.340 68.950 152.540 ;
        RECT 69.180 152.540 73.550 152.680 ;
        RECT 69.180 152.480 69.500 152.540 ;
        RECT 70.560 152.340 70.880 152.400 ;
        RECT 68.810 152.200 70.880 152.340 ;
        RECT 67.355 152.155 67.645 152.200 ;
        RECT 68.260 152.140 68.580 152.200 ;
        RECT 70.560 152.140 70.880 152.200 ;
        RECT 71.035 152.155 71.325 152.385 ;
        RECT 71.480 152.340 71.800 152.400 ;
        RECT 72.875 152.340 73.165 152.385 ;
        RECT 71.480 152.200 73.165 152.340 ;
        RECT 73.410 152.340 73.550 152.540 ;
        RECT 73.780 152.540 74.545 152.680 ;
        RECT 73.780 152.480 74.100 152.540 ;
        RECT 74.255 152.495 74.545 152.540 ;
        RECT 91.720 152.680 92.040 152.740 ;
        RECT 91.720 152.540 93.330 152.680 ;
        RECT 91.720 152.480 92.040 152.540 ;
        RECT 74.715 152.340 75.005 152.385 ;
        RECT 73.410 152.200 75.005 152.340 ;
        RECT 41.210 151.860 43.280 152.000 ;
        RECT 42.960 151.800 43.280 151.860 ;
        RECT 57.235 152.000 57.525 152.045 ;
        RECT 60.390 152.000 60.680 152.045 ;
        RECT 63.650 152.000 63.940 152.045 ;
        RECT 57.235 151.860 63.940 152.000 ;
        RECT 57.235 151.815 57.525 151.860 ;
        RECT 60.390 151.815 60.680 151.860 ;
        RECT 63.650 151.815 63.940 151.860 ;
        RECT 64.570 152.000 64.860 152.045 ;
        RECT 66.430 152.000 66.720 152.045 ;
        RECT 64.570 151.860 66.720 152.000 ;
        RECT 71.110 152.000 71.250 152.155 ;
        RECT 71.480 152.140 71.800 152.200 ;
        RECT 72.875 152.155 73.165 152.200 ;
        RECT 74.715 152.155 75.005 152.200 ;
        RECT 90.310 152.340 90.600 152.385 ;
        RECT 93.190 152.340 93.330 152.540 ;
        RECT 93.560 152.480 93.880 152.740 ;
        RECT 104.140 152.480 104.460 152.740 ;
        RECT 105.150 152.680 105.290 152.820 ;
        RECT 106.990 152.680 107.130 153.220 ;
        RECT 109.660 153.160 109.980 153.220 ;
        RECT 107.820 153.020 108.140 153.080 ;
        RECT 114.260 153.020 114.580 153.080 ;
        RECT 107.820 152.880 114.580 153.020 ;
        RECT 107.820 152.820 108.140 152.880 ;
        RECT 114.260 152.820 114.580 152.880 ;
        RECT 105.150 152.540 107.130 152.680 ;
        RECT 95.415 152.340 95.705 152.385 ;
        RECT 90.310 152.200 92.845 152.340 ;
        RECT 93.190 152.200 95.705 152.340 ;
        RECT 90.310 152.155 90.600 152.200 ;
        RECT 71.940 152.000 72.260 152.060 ;
        RECT 73.320 152.000 73.640 152.060 ;
        RECT 87.580 152.000 87.900 152.060 ;
        RECT 92.630 152.045 92.845 152.200 ;
        RECT 95.415 152.155 95.705 152.200 ;
        RECT 103.235 152.340 103.525 152.385 ;
        RECT 103.235 152.200 106.210 152.340 ;
        RECT 103.235 152.155 103.525 152.200 ;
        RECT 71.110 151.860 73.640 152.000 ;
        RECT 64.570 151.815 64.860 151.860 ;
        RECT 66.430 151.815 66.720 151.860 ;
        RECT 71.940 151.800 72.260 151.860 ;
        RECT 73.320 151.800 73.640 151.860 ;
        RECT 74.330 151.860 87.900 152.000 ;
        RECT 41.580 151.660 41.900 151.720 ;
        RECT 50.320 151.660 50.640 151.720 ;
        RECT 58.600 151.705 58.920 151.720 ;
        RECT 40.750 151.520 50.640 151.660 ;
        RECT 34.680 151.460 35.000 151.520 ;
        RECT 39.295 151.475 39.585 151.520 ;
        RECT 41.580 151.460 41.900 151.520 ;
        RECT 50.320 151.460 50.640 151.520 ;
        RECT 58.385 151.475 58.920 151.705 ;
        RECT 58.600 151.460 58.920 151.475 ;
        RECT 70.100 151.660 70.420 151.720 ;
        RECT 74.330 151.660 74.470 151.860 ;
        RECT 87.580 151.800 87.900 151.860 ;
        RECT 88.450 152.000 88.740 152.045 ;
        RECT 91.710 152.000 92.000 152.045 ;
        RECT 92.630 152.000 92.920 152.045 ;
        RECT 94.490 152.000 94.780 152.045 ;
        RECT 88.450 151.860 92.410 152.000 ;
        RECT 88.450 151.815 88.740 151.860 ;
        RECT 91.710 151.815 92.000 151.860 ;
        RECT 70.100 151.520 74.470 151.660 ;
        RECT 70.100 151.460 70.420 151.520 ;
        RECT 74.700 151.460 75.020 151.720 ;
        RECT 86.200 151.705 86.520 151.720 ;
        RECT 86.200 151.475 86.735 151.705 ;
        RECT 92.270 151.660 92.410 151.860 ;
        RECT 92.630 151.860 94.780 152.000 ;
        RECT 92.630 151.815 92.920 151.860 ;
        RECT 94.490 151.815 94.780 151.860 ;
        RECT 104.600 151.800 104.920 152.060 ;
        RECT 106.070 152.000 106.210 152.200 ;
        RECT 106.440 152.140 106.760 152.400 ;
        RECT 106.990 152.385 107.130 152.540 ;
        RECT 109.660 152.680 109.980 152.740 ;
        RECT 116.100 152.680 116.420 152.740 ;
        RECT 109.660 152.540 110.810 152.680 ;
        RECT 109.660 152.480 109.980 152.540 ;
        RECT 106.915 152.155 107.205 152.385 ;
        RECT 107.360 152.140 107.680 152.400 ;
        RECT 108.280 152.140 108.600 152.400 ;
        RECT 109.200 152.340 109.520 152.400 ;
        RECT 110.670 152.385 110.810 152.540 ;
        RECT 111.130 152.540 116.420 152.680 ;
        RECT 111.130 152.385 111.270 152.540 ;
        RECT 116.100 152.480 116.420 152.540 ;
        RECT 110.135 152.340 110.425 152.385 ;
        RECT 109.200 152.200 110.425 152.340 ;
        RECT 109.200 152.140 109.520 152.200 ;
        RECT 110.135 152.155 110.425 152.200 ;
        RECT 110.595 152.155 110.885 152.385 ;
        RECT 111.055 152.155 111.345 152.385 ;
        RECT 111.975 152.340 112.265 152.385 ;
        RECT 119.320 152.340 119.640 152.400 ;
        RECT 111.590 152.200 112.265 152.340 ;
        RECT 108.755 152.000 109.045 152.045 ;
        RECT 106.070 151.860 109.045 152.000 ;
        RECT 108.755 151.815 109.045 151.860 ;
        RECT 93.560 151.660 93.880 151.720 ;
        RECT 92.270 151.520 93.880 151.660 ;
        RECT 86.200 151.460 86.520 151.475 ;
        RECT 93.560 151.460 93.880 151.520 ;
        RECT 101.380 151.660 101.700 151.720 ;
        RECT 102.315 151.660 102.605 151.705 ;
        RECT 101.380 151.520 102.605 151.660 ;
        RECT 101.380 151.460 101.700 151.520 ;
        RECT 102.315 151.475 102.605 151.520 ;
        RECT 105.060 151.460 105.380 151.720 ;
        RECT 108.280 151.660 108.600 151.720 ;
        RECT 111.590 151.660 111.730 152.200 ;
        RECT 111.975 152.155 112.265 152.200 ;
        RECT 112.510 152.200 119.640 152.340 ;
        RECT 108.280 151.520 111.730 151.660 ;
        RECT 111.960 151.660 112.280 151.720 ;
        RECT 112.510 151.660 112.650 152.200 ;
        RECT 119.320 152.140 119.640 152.200 ;
        RECT 120.255 152.155 120.545 152.385 ;
        RECT 115.640 152.000 115.960 152.060 ;
        RECT 120.330 152.000 120.470 152.155 ;
        RECT 115.640 151.860 120.470 152.000 ;
        RECT 115.640 151.800 115.960 151.860 ;
        RECT 111.960 151.520 112.650 151.660 ;
        RECT 117.940 151.660 118.260 151.720 ;
        RECT 118.875 151.660 119.165 151.705 ;
        RECT 117.940 151.520 119.165 151.660 ;
        RECT 108.280 151.460 108.600 151.520 ;
        RECT 111.960 151.460 112.280 151.520 ;
        RECT 117.940 151.460 118.260 151.520 ;
        RECT 118.875 151.475 119.165 151.520 ;
        RECT 121.175 151.660 121.465 151.705 ;
        RECT 123.000 151.660 123.320 151.720 ;
        RECT 121.175 151.520 123.320 151.660 ;
        RECT 121.175 151.475 121.465 151.520 ;
        RECT 123.000 151.460 123.320 151.520 ;
        RECT 14.370 150.840 127.530 151.320 ;
        RECT 33.300 150.440 33.620 150.700 ;
        RECT 36.535 150.640 36.825 150.685 ;
        RECT 36.980 150.640 37.300 150.700 ;
        RECT 36.535 150.500 37.300 150.640 ;
        RECT 36.535 150.455 36.825 150.500 ;
        RECT 36.980 150.440 37.300 150.500 ;
        RECT 60.455 150.455 60.745 150.685 ;
        RECT 60.900 150.640 61.220 150.700 ;
        RECT 61.375 150.640 61.665 150.685 ;
        RECT 60.900 150.500 61.665 150.640 ;
        RECT 18.530 150.300 18.820 150.345 ;
        RECT 19.960 150.300 20.280 150.360 ;
        RECT 21.790 150.300 22.080 150.345 ;
        RECT 18.530 150.160 22.080 150.300 ;
        RECT 18.530 150.115 18.820 150.160 ;
        RECT 19.960 150.100 20.280 150.160 ;
        RECT 21.790 150.115 22.080 150.160 ;
        RECT 22.710 150.300 23.000 150.345 ;
        RECT 24.570 150.300 24.860 150.345 ;
        RECT 22.710 150.160 24.860 150.300 ;
        RECT 22.710 150.115 23.000 150.160 ;
        RECT 24.570 150.115 24.860 150.160 ;
        RECT 31.000 150.300 31.320 150.360 ;
        RECT 58.155 150.300 58.445 150.345 ;
        RECT 31.000 150.160 43.650 150.300 ;
        RECT 20.390 149.960 20.680 150.005 ;
        RECT 22.710 149.960 22.925 150.115 ;
        RECT 31.000 150.100 31.320 150.160 ;
        RECT 20.390 149.820 22.925 149.960 ;
        RECT 29.620 149.960 29.940 150.020 ;
        RECT 32.855 149.960 33.145 150.005 ;
        RECT 29.620 149.820 33.145 149.960 ;
        RECT 20.390 149.775 20.680 149.820 ;
        RECT 29.620 149.760 29.940 149.820 ;
        RECT 32.855 149.775 33.145 149.820 ;
        RECT 35.600 149.760 35.920 150.020 ;
        RECT 41.580 149.960 41.900 150.020 ;
        RECT 42.515 149.960 42.805 150.005 ;
        RECT 41.580 149.820 42.805 149.960 ;
        RECT 41.580 149.760 41.900 149.820 ;
        RECT 42.515 149.775 42.805 149.820 ;
        RECT 42.960 149.760 43.280 150.020 ;
        RECT 43.510 150.005 43.650 150.160 ;
        RECT 53.630 150.160 58.445 150.300 ;
        RECT 53.630 150.020 53.770 150.160 ;
        RECT 58.155 150.115 58.445 150.160 ;
        RECT 43.435 149.775 43.725 150.005 ;
        RECT 44.355 149.960 44.645 150.005 ;
        RECT 44.800 149.960 45.120 150.020 ;
        RECT 44.355 149.820 45.120 149.960 ;
        RECT 44.355 149.775 44.645 149.820 ;
        RECT 44.800 149.760 45.120 149.820 ;
        RECT 48.495 149.775 48.785 150.005 ;
        RECT 16.525 149.620 16.815 149.665 ;
        RECT 22.260 149.620 22.580 149.680 ;
        RECT 16.525 149.480 22.580 149.620 ;
        RECT 16.525 149.435 16.815 149.480 ;
        RECT 22.260 149.420 22.580 149.480 ;
        RECT 23.655 149.620 23.945 149.665 ;
        RECT 24.560 149.620 24.880 149.680 ;
        RECT 23.655 149.480 24.880 149.620 ;
        RECT 23.655 149.435 23.945 149.480 ;
        RECT 24.560 149.420 24.880 149.480 ;
        RECT 25.495 149.620 25.785 149.665 ;
        RECT 36.060 149.620 36.380 149.680 ;
        RECT 25.495 149.480 36.380 149.620 ;
        RECT 48.570 149.620 48.710 149.775 ;
        RECT 49.400 149.760 49.720 150.020 ;
        RECT 49.860 149.760 50.180 150.020 ;
        RECT 52.635 149.775 52.925 150.005 ;
        RECT 50.320 149.620 50.640 149.680 ;
        RECT 48.570 149.480 50.640 149.620 ;
        RECT 52.710 149.620 52.850 149.775 ;
        RECT 53.080 149.760 53.400 150.020 ;
        RECT 53.540 149.760 53.860 150.020 ;
        RECT 54.475 149.960 54.765 150.005 ;
        RECT 56.300 149.960 56.620 150.020 ;
        RECT 54.475 149.820 56.620 149.960 ;
        RECT 54.475 149.775 54.765 149.820 ;
        RECT 56.300 149.760 56.620 149.820 ;
        RECT 58.600 149.760 58.920 150.020 ;
        RECT 60.530 149.960 60.670 150.455 ;
        RECT 60.900 150.440 61.220 150.500 ;
        RECT 61.375 150.455 61.665 150.500 ;
        RECT 64.595 150.640 64.885 150.685 ;
        RECT 65.500 150.640 65.820 150.700 ;
        RECT 64.595 150.500 65.820 150.640 ;
        RECT 64.595 150.455 64.885 150.500 ;
        RECT 65.500 150.440 65.820 150.500 ;
        RECT 68.275 150.640 68.565 150.685 ;
        RECT 85.755 150.640 86.045 150.685 ;
        RECT 86.200 150.640 86.520 150.700 ;
        RECT 88.055 150.640 88.345 150.685 ;
        RECT 92.655 150.640 92.945 150.685 ;
        RECT 93.100 150.640 93.420 150.700 ;
        RECT 68.275 150.500 71.250 150.640 ;
        RECT 68.275 150.455 68.565 150.500 ;
        RECT 62.295 149.960 62.585 150.005 ;
        RECT 60.530 149.820 62.585 149.960 ;
        RECT 62.295 149.775 62.585 149.820 ;
        RECT 63.660 149.760 63.980 150.020 ;
        RECT 67.355 149.960 67.645 150.005 ;
        RECT 69.180 149.960 69.500 150.020 ;
        RECT 67.355 149.820 69.500 149.960 ;
        RECT 67.355 149.775 67.645 149.820 ;
        RECT 69.180 149.760 69.500 149.820 ;
        RECT 70.560 149.760 70.880 150.020 ;
        RECT 54.000 149.620 54.320 149.680 ;
        RECT 52.710 149.480 54.320 149.620 ;
        RECT 25.495 149.435 25.785 149.480 ;
        RECT 36.060 149.420 36.380 149.480 ;
        RECT 50.320 149.420 50.640 149.480 ;
        RECT 54.000 149.420 54.320 149.480 ;
        RECT 57.695 149.620 57.985 149.665 ;
        RECT 65.500 149.620 65.820 149.680 ;
        RECT 57.695 149.480 64.810 149.620 ;
        RECT 57.695 149.435 57.985 149.480 ;
        RECT 64.670 149.340 64.810 149.480 ;
        RECT 65.500 149.480 70.790 149.620 ;
        RECT 65.500 149.420 65.820 149.480 ;
        RECT 20.390 149.280 20.680 149.325 ;
        RECT 23.170 149.280 23.460 149.325 ;
        RECT 25.030 149.280 25.320 149.325 ;
        RECT 20.390 149.140 25.320 149.280 ;
        RECT 20.390 149.095 20.680 149.140 ;
        RECT 23.170 149.095 23.460 149.140 ;
        RECT 25.030 149.095 25.320 149.140 ;
        RECT 50.795 149.280 51.085 149.325 ;
        RECT 59.980 149.280 60.300 149.340 ;
        RECT 50.795 149.140 60.300 149.280 ;
        RECT 50.795 149.095 51.085 149.140 ;
        RECT 59.980 149.080 60.300 149.140 ;
        RECT 64.580 149.280 64.900 149.340 ;
        RECT 70.650 149.280 70.790 149.480 ;
        RECT 71.110 149.280 71.250 150.500 ;
        RECT 85.755 150.500 86.890 150.640 ;
        RECT 85.755 150.455 86.045 150.500 ;
        RECT 86.200 150.440 86.520 150.500 ;
        RECT 72.875 150.300 73.165 150.345 ;
        RECT 74.700 150.300 75.020 150.360 ;
        RECT 75.175 150.300 75.465 150.345 ;
        RECT 72.875 150.160 75.465 150.300 ;
        RECT 72.875 150.115 73.165 150.160 ;
        RECT 74.700 150.100 75.020 150.160 ;
        RECT 75.175 150.115 75.465 150.160 ;
        RECT 77.015 150.300 77.305 150.345 ;
        RECT 77.015 150.160 85.050 150.300 ;
        RECT 77.015 150.115 77.305 150.160 ;
        RECT 75.620 149.960 75.940 150.020 ;
        RECT 78.395 149.960 78.685 150.005 ;
        RECT 75.620 149.820 78.685 149.960 ;
        RECT 75.620 149.760 75.940 149.820 ;
        RECT 78.395 149.775 78.685 149.820 ;
        RECT 79.760 149.760 80.080 150.020 ;
        RECT 84.910 149.680 85.050 150.160 ;
        RECT 85.740 149.960 86.060 150.020 ;
        RECT 86.215 149.960 86.505 150.005 ;
        RECT 85.740 149.820 86.505 149.960 ;
        RECT 85.740 149.760 86.060 149.820 ;
        RECT 86.215 149.775 86.505 149.820 ;
        RECT 79.300 149.420 79.620 149.680 ;
        RECT 84.820 149.420 85.140 149.680 ;
        RECT 77.920 149.280 78.240 149.340 ;
        RECT 64.580 149.140 70.330 149.280 ;
        RECT 70.650 149.140 78.240 149.280 ;
        RECT 86.750 149.280 86.890 150.500 ;
        RECT 88.055 150.500 91.950 150.640 ;
        RECT 88.055 150.455 88.345 150.500 ;
        RECT 91.810 150.125 91.950 150.500 ;
        RECT 92.655 150.500 93.420 150.640 ;
        RECT 92.655 150.455 92.945 150.500 ;
        RECT 93.100 150.440 93.420 150.500 ;
        RECT 93.560 150.440 93.880 150.700 ;
        RECT 104.600 150.640 104.920 150.700 ;
        RECT 106.915 150.640 107.205 150.685 ;
        RECT 94.110 150.500 104.370 150.640 ;
        RECT 90.355 149.775 90.645 150.005 ;
        RECT 91.735 149.895 92.025 150.125 ;
        RECT 94.110 150.005 94.250 150.500 ;
        RECT 95.400 150.300 95.720 150.360 ;
        RECT 97.815 150.300 98.105 150.345 ;
        RECT 101.055 150.300 101.705 150.345 ;
        RECT 95.400 150.160 101.705 150.300 ;
        RECT 95.400 150.100 95.720 150.160 ;
        RECT 97.815 150.115 98.405 150.160 ;
        RECT 101.055 150.115 101.705 150.160 ;
        RECT 103.220 150.300 103.540 150.360 ;
        RECT 103.695 150.300 103.985 150.345 ;
        RECT 103.220 150.160 103.985 150.300 ;
        RECT 104.230 150.300 104.370 150.500 ;
        RECT 104.600 150.500 107.205 150.640 ;
        RECT 104.600 150.440 104.920 150.500 ;
        RECT 106.915 150.455 107.205 150.500 ;
        RECT 116.560 150.300 116.880 150.360 ;
        RECT 104.230 150.160 116.880 150.300 ;
        RECT 94.035 149.960 94.325 150.005 ;
        RECT 92.270 149.820 94.325 149.960 ;
        RECT 90.430 149.620 90.570 149.775 ;
        RECT 92.270 149.620 92.410 149.820 ;
        RECT 94.035 149.775 94.325 149.820 ;
        RECT 98.115 149.800 98.405 150.115 ;
        RECT 103.220 150.100 103.540 150.160 ;
        RECT 103.695 150.115 103.985 150.160 ;
        RECT 116.560 150.100 116.880 150.160 ;
        RECT 117.135 150.300 117.425 150.345 ;
        RECT 117.940 150.300 118.260 150.360 ;
        RECT 120.375 150.300 121.025 150.345 ;
        RECT 117.135 150.160 121.025 150.300 ;
        RECT 117.135 150.115 117.725 150.160 ;
        RECT 99.195 149.960 99.485 150.005 ;
        RECT 102.775 149.960 103.065 150.005 ;
        RECT 104.610 149.960 104.900 150.005 ;
        RECT 99.195 149.820 104.900 149.960 ;
        RECT 99.195 149.775 99.485 149.820 ;
        RECT 102.775 149.775 103.065 149.820 ;
        RECT 104.610 149.775 104.900 149.820 ;
        RECT 107.820 149.960 108.140 150.020 ;
        RECT 108.295 149.960 108.585 150.005 ;
        RECT 107.820 149.820 108.585 149.960 ;
        RECT 107.820 149.760 108.140 149.820 ;
        RECT 108.295 149.775 108.585 149.820 ;
        RECT 108.755 149.775 109.045 150.005 ;
        RECT 109.215 149.775 109.505 150.005 ;
        RECT 109.660 149.960 109.980 150.020 ;
        RECT 110.135 149.960 110.425 150.005 ;
        RECT 109.660 149.820 110.425 149.960 ;
        RECT 105.075 149.620 105.365 149.665 ;
        RECT 90.430 149.480 92.410 149.620 ;
        RECT 94.110 149.480 105.365 149.620 ;
        RECT 94.110 149.340 94.250 149.480 ;
        RECT 105.075 149.435 105.365 149.480 ;
        RECT 107.360 149.620 107.680 149.680 ;
        RECT 108.830 149.620 108.970 149.775 ;
        RECT 107.360 149.480 108.970 149.620 ;
        RECT 109.290 149.620 109.430 149.775 ;
        RECT 109.660 149.760 109.980 149.820 ;
        RECT 110.135 149.775 110.425 149.820 ;
        RECT 117.435 149.800 117.725 150.115 ;
        RECT 117.940 150.100 118.260 150.160 ;
        RECT 120.375 150.115 121.025 150.160 ;
        RECT 123.000 150.100 123.320 150.360 ;
        RECT 118.515 149.960 118.805 150.005 ;
        RECT 122.095 149.960 122.385 150.005 ;
        RECT 123.930 149.960 124.220 150.005 ;
        RECT 118.515 149.820 124.220 149.960 ;
        RECT 118.515 149.775 118.805 149.820 ;
        RECT 122.095 149.775 122.385 149.820 ;
        RECT 123.930 149.775 124.220 149.820 ;
        RECT 111.055 149.620 111.345 149.665 ;
        RECT 115.655 149.620 115.945 149.665 ;
        RECT 109.290 149.480 115.945 149.620 ;
        RECT 107.360 149.420 107.680 149.480 ;
        RECT 93.560 149.280 93.880 149.340 ;
        RECT 86.750 149.140 93.880 149.280 ;
        RECT 64.580 149.080 64.900 149.140 ;
        RECT 40.660 148.940 40.980 149.000 ;
        RECT 41.135 148.940 41.425 148.985 ;
        RECT 40.660 148.800 41.425 148.940 ;
        RECT 40.660 148.740 40.980 148.800 ;
        RECT 41.135 148.755 41.425 148.800 ;
        RECT 43.880 148.940 44.200 149.000 ;
        RECT 48.495 148.940 48.785 148.985 ;
        RECT 43.880 148.800 48.785 148.940 ;
        RECT 43.880 148.740 44.200 148.800 ;
        RECT 48.495 148.755 48.785 148.800 ;
        RECT 51.240 148.740 51.560 149.000 ;
        RECT 65.040 148.940 65.360 149.000 ;
        RECT 69.655 148.940 69.945 148.985 ;
        RECT 65.040 148.800 69.945 148.940 ;
        RECT 70.190 148.940 70.330 149.140 ;
        RECT 77.920 149.080 78.240 149.140 ;
        RECT 93.560 149.080 93.880 149.140 ;
        RECT 94.020 149.080 94.340 149.340 ;
        RECT 99.195 149.280 99.485 149.325 ;
        RECT 102.315 149.280 102.605 149.325 ;
        RECT 104.205 149.280 104.495 149.325 ;
        RECT 99.195 149.140 104.495 149.280 ;
        RECT 108.830 149.280 108.970 149.480 ;
        RECT 111.055 149.435 111.345 149.480 ;
        RECT 115.655 149.435 115.945 149.480 ;
        RECT 124.395 149.620 124.685 149.665 ;
        RECT 125.760 149.620 126.080 149.680 ;
        RECT 124.395 149.480 126.080 149.620 ;
        RECT 124.395 149.435 124.685 149.480 ;
        RECT 125.760 149.420 126.080 149.480 ;
        RECT 111.500 149.280 111.820 149.340 ;
        RECT 108.830 149.140 111.820 149.280 ;
        RECT 99.195 149.095 99.485 149.140 ;
        RECT 102.315 149.095 102.605 149.140 ;
        RECT 104.205 149.095 104.495 149.140 ;
        RECT 111.500 149.080 111.820 149.140 ;
        RECT 118.515 149.280 118.805 149.325 ;
        RECT 121.635 149.280 121.925 149.325 ;
        RECT 123.525 149.280 123.815 149.325 ;
        RECT 118.515 149.140 123.815 149.280 ;
        RECT 118.515 149.095 118.805 149.140 ;
        RECT 121.635 149.095 121.925 149.140 ;
        RECT 123.525 149.095 123.815 149.140 ;
        RECT 71.495 148.940 71.785 148.985 ;
        RECT 70.190 148.800 71.785 148.940 ;
        RECT 65.040 148.740 65.360 148.800 ;
        RECT 69.655 148.755 69.945 148.800 ;
        RECT 71.495 148.755 71.785 148.800 ;
        RECT 75.620 148.940 75.940 149.000 ;
        RECT 77.475 148.940 77.765 148.985 ;
        RECT 75.620 148.800 77.765 148.940 ;
        RECT 75.620 148.740 75.940 148.800 ;
        RECT 77.475 148.755 77.765 148.800 ;
        RECT 79.775 148.940 80.065 148.985 ;
        RECT 81.600 148.940 81.920 149.000 ;
        RECT 79.775 148.800 81.920 148.940 ;
        RECT 79.775 148.755 80.065 148.800 ;
        RECT 81.600 148.740 81.920 148.800 ;
        RECT 89.895 148.940 90.185 148.985 ;
        RECT 90.340 148.940 90.660 149.000 ;
        RECT 89.895 148.800 90.660 148.940 ;
        RECT 89.895 148.755 90.185 148.800 ;
        RECT 90.340 148.740 90.660 148.800 ;
        RECT 96.320 148.740 96.640 149.000 ;
        RECT 113.800 148.740 114.120 149.000 ;
        RECT 14.370 148.120 127.530 148.600 ;
        RECT 24.560 147.720 24.880 147.980 ;
        RECT 35.600 147.920 35.920 147.980 ;
        RECT 48.495 147.920 48.785 147.965 ;
        RECT 48.940 147.920 49.260 147.980 ;
        RECT 35.600 147.780 42.730 147.920 ;
        RECT 35.600 147.720 35.920 147.780 ;
        RECT 23.655 147.395 23.945 147.625 ;
        RECT 28.240 147.580 28.560 147.640 ;
        RECT 28.240 147.440 34.450 147.580 ;
        RECT 20.880 147.040 21.200 147.300 ;
        RECT 23.730 146.900 23.870 147.395 ;
        RECT 28.240 147.380 28.560 147.440 ;
        RECT 32.395 147.240 32.685 147.285 ;
        RECT 33.760 147.240 34.080 147.300 ;
        RECT 26.030 147.100 31.690 147.240 ;
        RECT 25.495 146.900 25.785 146.945 ;
        RECT 23.730 146.760 25.785 146.900 ;
        RECT 25.495 146.715 25.785 146.760 ;
        RECT 21.815 146.560 22.105 146.605 ;
        RECT 22.720 146.560 23.040 146.620 ;
        RECT 26.030 146.560 26.170 147.100 ;
        RECT 27.795 146.900 28.085 146.945 ;
        RECT 27.795 146.760 29.850 146.900 ;
        RECT 27.795 146.715 28.085 146.760 ;
        RECT 21.815 146.420 26.170 146.560 ;
        RECT 21.815 146.375 22.105 146.420 ;
        RECT 22.720 146.360 23.040 146.420 ;
        RECT 21.355 146.220 21.645 146.265 ;
        RECT 22.260 146.220 22.580 146.280 ;
        RECT 28.240 146.220 28.560 146.280 ;
        RECT 21.355 146.080 28.560 146.220 ;
        RECT 21.355 146.035 21.645 146.080 ;
        RECT 22.260 146.020 22.580 146.080 ;
        RECT 28.240 146.020 28.560 146.080 ;
        RECT 28.700 146.020 29.020 146.280 ;
        RECT 29.175 146.220 29.465 146.265 ;
        RECT 29.710 146.220 29.850 146.760 ;
        RECT 31.000 146.700 31.320 146.960 ;
        RECT 31.550 146.605 31.690 147.100 ;
        RECT 32.395 147.100 34.080 147.240 ;
        RECT 34.310 147.240 34.450 147.440 ;
        RECT 36.610 147.440 41.810 147.580 ;
        RECT 36.610 147.240 36.750 147.440 ;
        RECT 34.310 147.100 36.750 147.240 ;
        RECT 37.070 147.100 41.350 147.240 ;
        RECT 32.395 147.055 32.685 147.100 ;
        RECT 33.760 147.040 34.080 147.100 ;
        RECT 35.600 146.700 35.920 146.960 ;
        RECT 37.070 146.945 37.210 147.100 ;
        RECT 41.210 146.945 41.350 147.100 ;
        RECT 41.670 146.945 41.810 147.440 ;
        RECT 42.590 146.945 42.730 147.780 ;
        RECT 48.495 147.780 49.260 147.920 ;
        RECT 48.495 147.735 48.785 147.780 ;
        RECT 48.940 147.720 49.260 147.780 ;
        RECT 50.320 147.920 50.640 147.980 ;
        RECT 53.095 147.920 53.385 147.965 ;
        RECT 50.320 147.780 53.385 147.920 ;
        RECT 50.320 147.720 50.640 147.780 ;
        RECT 53.095 147.735 53.385 147.780 ;
        RECT 54.460 147.920 54.780 147.980 ;
        RECT 73.320 147.920 73.640 147.980 ;
        RECT 54.460 147.780 73.640 147.920 ;
        RECT 54.460 147.720 54.780 147.780 ;
        RECT 73.320 147.720 73.640 147.780 ;
        RECT 79.760 147.720 80.080 147.980 ;
        RECT 84.820 147.920 85.140 147.980 ;
        RECT 84.820 147.780 95.170 147.920 ;
        RECT 84.820 147.720 85.140 147.780 ;
        RECT 49.415 147.580 49.705 147.625 ;
        RECT 56.760 147.580 57.080 147.640 ;
        RECT 77.920 147.580 78.240 147.640 ;
        RECT 82.980 147.580 83.300 147.640 ;
        RECT 49.415 147.440 57.080 147.580 ;
        RECT 49.415 147.395 49.705 147.440 ;
        RECT 56.760 147.380 57.080 147.440 ;
        RECT 57.310 147.440 66.190 147.580 ;
        RECT 48.035 147.240 48.325 147.285 ;
        RECT 52.160 147.240 52.480 147.300 ;
        RECT 48.035 147.100 52.480 147.240 ;
        RECT 48.035 147.055 48.325 147.100 ;
        RECT 52.160 147.040 52.480 147.100 ;
        RECT 53.080 147.240 53.400 147.300 ;
        RECT 57.310 147.240 57.450 147.440 ;
        RECT 53.080 147.100 57.450 147.240 ;
        RECT 60.455 147.240 60.745 147.285 ;
        RECT 64.580 147.240 64.900 147.300 ;
        RECT 60.455 147.100 64.900 147.240 ;
        RECT 53.080 147.040 53.400 147.100 ;
        RECT 36.535 146.715 36.825 146.945 ;
        RECT 36.995 146.715 37.285 146.945 ;
        RECT 37.455 146.900 37.745 146.945 ;
        RECT 40.675 146.900 40.965 146.945 ;
        RECT 37.455 146.760 40.965 146.900 ;
        RECT 37.455 146.715 37.745 146.760 ;
        RECT 40.675 146.715 40.965 146.760 ;
        RECT 41.135 146.715 41.425 146.945 ;
        RECT 41.595 146.715 41.885 146.945 ;
        RECT 42.515 146.900 42.805 146.945 ;
        RECT 44.340 146.900 44.660 146.960 ;
        RECT 42.515 146.760 44.660 146.900 ;
        RECT 42.515 146.715 42.805 146.760 ;
        RECT 31.475 146.560 31.765 146.605 ;
        RECT 36.610 146.560 36.750 146.715 ;
        RECT 39.295 146.560 39.585 146.605 ;
        RECT 31.475 146.420 36.750 146.560 ;
        RECT 37.530 146.420 39.585 146.560 ;
        RECT 31.475 146.375 31.765 146.420 ;
        RECT 29.175 146.080 29.850 146.220 ;
        RECT 36.520 146.220 36.840 146.280 ;
        RECT 37.530 146.220 37.670 146.420 ;
        RECT 39.295 146.375 39.585 146.420 ;
        RECT 36.520 146.080 37.670 146.220 ;
        RECT 38.360 146.220 38.680 146.280 ;
        RECT 38.835 146.220 39.125 146.265 ;
        RECT 38.360 146.080 39.125 146.220 ;
        RECT 40.750 146.220 40.890 146.715 ;
        RECT 41.210 146.560 41.350 146.715 ;
        RECT 44.340 146.700 44.660 146.760 ;
        RECT 48.480 146.700 48.800 146.960 ;
        RECT 51.700 146.700 52.020 146.960 ;
        RECT 54.460 146.700 54.780 146.960 ;
        RECT 55.010 146.945 55.150 147.100 ;
        RECT 60.455 147.055 60.745 147.100 ;
        RECT 64.580 147.040 64.900 147.100 ;
        RECT 54.935 146.715 55.225 146.945 ;
        RECT 55.395 146.715 55.685 146.945 ;
        RECT 56.300 146.900 56.620 146.960 ;
        RECT 65.500 146.900 65.820 146.960 ;
        RECT 56.300 146.760 65.820 146.900 ;
        RECT 66.050 146.900 66.190 147.440 ;
        RECT 76.170 147.440 83.300 147.580 ;
        RECT 70.560 147.240 70.880 147.300 ;
        RECT 70.560 147.100 72.630 147.240 ;
        RECT 70.560 147.040 70.880 147.100 ;
        RECT 66.050 146.760 71.020 146.900 ;
        RECT 42.960 146.560 43.280 146.620 ;
        RECT 41.210 146.420 43.280 146.560 ;
        RECT 42.960 146.360 43.280 146.420 ;
        RECT 47.115 146.560 47.405 146.605 ;
        RECT 51.240 146.560 51.560 146.620 ;
        RECT 47.115 146.420 51.560 146.560 ;
        RECT 55.470 146.560 55.610 146.715 ;
        RECT 56.300 146.700 56.620 146.760 ;
        RECT 65.500 146.700 65.820 146.760 ;
        RECT 58.600 146.560 58.920 146.620 ;
        RECT 60.915 146.560 61.205 146.605 ;
        RECT 55.470 146.420 61.205 146.560 ;
        RECT 70.880 146.560 71.020 146.760 ;
        RECT 71.940 146.700 72.260 146.960 ;
        RECT 72.490 146.945 72.630 147.100 ;
        RECT 76.170 146.945 76.310 147.440 ;
        RECT 77.920 147.380 78.240 147.440 ;
        RECT 82.980 147.380 83.300 147.440 ;
        RECT 88.930 147.580 89.220 147.625 ;
        RECT 91.710 147.580 92.000 147.625 ;
        RECT 93.570 147.580 93.860 147.625 ;
        RECT 88.930 147.440 93.860 147.580 ;
        RECT 95.030 147.580 95.170 147.780 ;
        RECT 95.400 147.720 95.720 147.980 ;
        RECT 96.320 147.920 96.640 147.980 ;
        RECT 102.775 147.920 103.065 147.965 ;
        RECT 103.220 147.920 103.540 147.980 ;
        RECT 96.320 147.780 100.690 147.920 ;
        RECT 96.320 147.720 96.640 147.780 ;
        RECT 95.030 147.440 97.010 147.580 ;
        RECT 88.930 147.395 89.220 147.440 ;
        RECT 91.710 147.395 92.000 147.440 ;
        RECT 93.570 147.395 93.860 147.440 ;
        RECT 86.200 147.240 86.520 147.300 ;
        RECT 77.090 147.100 86.520 147.240 ;
        RECT 77.090 146.945 77.230 147.100 ;
        RECT 86.200 147.040 86.520 147.100 ;
        RECT 90.800 147.240 91.120 147.300 ;
        RECT 96.870 147.285 97.010 147.440 ;
        RECT 100.015 147.395 100.305 147.625 ;
        RECT 100.550 147.580 100.690 147.780 ;
        RECT 102.775 147.780 103.540 147.920 ;
        RECT 102.775 147.735 103.065 147.780 ;
        RECT 103.220 147.720 103.540 147.780 ;
        RECT 103.695 147.920 103.985 147.965 ;
        RECT 104.140 147.920 104.460 147.980 ;
        RECT 103.695 147.780 104.460 147.920 ;
        RECT 103.695 147.735 103.985 147.780 ;
        RECT 104.140 147.720 104.460 147.780 ;
        RECT 105.980 147.720 106.300 147.980 ;
        RECT 115.640 147.720 115.960 147.980 ;
        RECT 120.210 147.580 120.500 147.625 ;
        RECT 122.990 147.580 123.280 147.625 ;
        RECT 124.850 147.580 125.140 147.625 ;
        RECT 100.550 147.440 108.970 147.580 ;
        RECT 92.195 147.240 92.485 147.285 ;
        RECT 90.800 147.100 92.485 147.240 ;
        RECT 90.800 147.040 91.120 147.100 ;
        RECT 92.195 147.055 92.485 147.100 ;
        RECT 96.795 147.055 97.085 147.285 ;
        RECT 72.415 146.715 72.705 146.945 ;
        RECT 76.095 146.715 76.385 146.945 ;
        RECT 77.015 146.715 77.305 146.945 ;
        RECT 77.475 146.715 77.765 146.945 ;
        RECT 77.920 146.900 78.240 146.960 ;
        RECT 79.760 146.900 80.080 146.960 ;
        RECT 81.155 146.900 81.445 146.945 ;
        RECT 77.920 146.760 81.445 146.900 ;
        RECT 77.550 146.560 77.690 146.715 ;
        RECT 77.920 146.700 78.240 146.760 ;
        RECT 79.760 146.700 80.080 146.760 ;
        RECT 81.155 146.715 81.445 146.760 ;
        RECT 81.615 146.715 81.905 146.945 ;
        RECT 81.690 146.560 81.830 146.715 ;
        RECT 82.060 146.700 82.380 146.960 ;
        RECT 82.980 146.700 83.300 146.960 ;
        RECT 88.930 146.900 89.220 146.945 ;
        RECT 88.930 146.760 91.465 146.900 ;
        RECT 88.930 146.715 89.220 146.760 ;
        RECT 82.520 146.560 82.840 146.620 ;
        RECT 90.340 146.605 90.660 146.620 ;
        RECT 70.880 146.420 82.840 146.560 ;
        RECT 47.115 146.375 47.405 146.420 ;
        RECT 51.240 146.360 51.560 146.420 ;
        RECT 58.600 146.360 58.920 146.420 ;
        RECT 60.915 146.375 61.205 146.420 ;
        RECT 41.580 146.220 41.900 146.280 ;
        RECT 40.750 146.080 41.900 146.220 ;
        RECT 29.175 146.035 29.465 146.080 ;
        RECT 36.520 146.020 36.840 146.080 ;
        RECT 38.360 146.020 38.680 146.080 ;
        RECT 38.835 146.035 39.125 146.080 ;
        RECT 41.580 146.020 41.900 146.080 ;
        RECT 49.400 146.220 49.720 146.280 ;
        RECT 50.795 146.220 51.085 146.265 ;
        RECT 49.400 146.080 51.085 146.220 ;
        RECT 49.400 146.020 49.720 146.080 ;
        RECT 50.795 146.035 51.085 146.080 ;
        RECT 59.060 146.220 59.380 146.280 ;
        RECT 61.375 146.220 61.665 146.265 ;
        RECT 59.060 146.080 61.665 146.220 ;
        RECT 59.060 146.020 59.380 146.080 ;
        RECT 61.375 146.035 61.665 146.080 ;
        RECT 63.215 146.220 63.505 146.265 ;
        RECT 63.660 146.220 63.980 146.280 ;
        RECT 71.110 146.265 71.250 146.420 ;
        RECT 82.520 146.360 82.840 146.420 ;
        RECT 87.070 146.560 87.360 146.605 ;
        RECT 90.330 146.560 90.660 146.605 ;
        RECT 87.070 146.420 90.660 146.560 ;
        RECT 87.070 146.375 87.360 146.420 ;
        RECT 90.330 146.375 90.660 146.420 ;
        RECT 91.250 146.605 91.465 146.760 ;
        RECT 94.020 146.700 94.340 146.960 ;
        RECT 94.940 146.700 95.260 146.960 ;
        RECT 98.175 146.715 98.465 146.945 ;
        RECT 100.090 146.900 100.230 147.395 ;
        RECT 102.760 147.240 103.080 147.300 ;
        RECT 105.535 147.240 105.825 147.285 ;
        RECT 102.760 147.100 105.825 147.240 ;
        RECT 102.760 147.040 103.080 147.100 ;
        RECT 105.535 147.055 105.825 147.100 ;
        RECT 107.360 147.240 107.680 147.300 ;
        RECT 107.360 147.100 108.510 147.240 ;
        RECT 107.360 147.040 107.680 147.100 ;
        RECT 101.855 146.900 102.145 146.945 ;
        RECT 100.090 146.760 102.145 146.900 ;
        RECT 101.855 146.715 102.145 146.760 ;
        RECT 104.615 146.900 104.905 146.945 ;
        RECT 105.060 146.900 105.380 146.960 ;
        RECT 104.615 146.760 105.380 146.900 ;
        RECT 104.615 146.715 104.905 146.760 ;
        RECT 91.250 146.560 91.540 146.605 ;
        RECT 93.110 146.560 93.400 146.605 ;
        RECT 91.250 146.420 93.400 146.560 ;
        RECT 91.250 146.375 91.540 146.420 ;
        RECT 93.110 146.375 93.400 146.420 ;
        RECT 93.560 146.560 93.880 146.620 ;
        RECT 98.250 146.560 98.390 146.715 ;
        RECT 105.060 146.700 105.380 146.760 ;
        RECT 107.820 146.700 108.140 146.960 ;
        RECT 108.370 146.945 108.510 147.100 ;
        RECT 108.830 146.945 108.970 147.440 ;
        RECT 120.210 147.440 125.140 147.580 ;
        RECT 120.210 147.395 120.500 147.440 ;
        RECT 122.990 147.395 123.280 147.440 ;
        RECT 124.850 147.395 125.140 147.440 ;
        RECT 112.880 147.040 113.200 147.300 ;
        RECT 108.295 146.715 108.585 146.945 ;
        RECT 108.755 146.715 109.045 146.945 ;
        RECT 109.660 146.900 109.980 146.960 ;
        RECT 111.960 146.900 112.280 146.960 ;
        RECT 109.660 146.760 112.280 146.900 ;
        RECT 109.660 146.700 109.980 146.760 ;
        RECT 111.960 146.700 112.280 146.760 ;
        RECT 113.815 146.715 114.105 146.945 ;
        RECT 120.210 146.900 120.500 146.945 ;
        RECT 120.210 146.760 122.745 146.900 ;
        RECT 120.210 146.715 120.500 146.760 ;
        RECT 93.560 146.420 98.390 146.560 ;
        RECT 105.995 146.560 106.285 146.605 ;
        RECT 106.455 146.560 106.745 146.605 ;
        RECT 113.890 146.560 114.030 146.715 ;
        RECT 105.995 146.420 106.745 146.560 ;
        RECT 90.340 146.360 90.660 146.375 ;
        RECT 93.560 146.360 93.880 146.420 ;
        RECT 105.995 146.375 106.285 146.420 ;
        RECT 106.455 146.375 106.745 146.420 ;
        RECT 106.990 146.420 114.030 146.560 ;
        RECT 116.345 146.560 116.635 146.605 ;
        RECT 117.480 146.560 117.800 146.620 ;
        RECT 116.345 146.420 117.800 146.560 ;
        RECT 63.215 146.080 63.980 146.220 ;
        RECT 63.215 146.035 63.505 146.080 ;
        RECT 63.660 146.020 63.980 146.080 ;
        RECT 71.035 146.035 71.325 146.265 ;
        RECT 73.320 146.220 73.640 146.280 ;
        RECT 77.920 146.220 78.240 146.280 ;
        RECT 73.320 146.080 78.240 146.220 ;
        RECT 73.320 146.020 73.640 146.080 ;
        RECT 77.920 146.020 78.240 146.080 ;
        RECT 79.300 146.020 79.620 146.280 ;
        RECT 82.060 146.220 82.380 146.280 ;
        RECT 85.065 146.220 85.355 146.265 ;
        RECT 85.740 146.220 86.060 146.280 ;
        RECT 82.060 146.080 86.060 146.220 ;
        RECT 82.060 146.020 82.380 146.080 ;
        RECT 85.065 146.035 85.355 146.080 ;
        RECT 85.740 146.020 86.060 146.080 ;
        RECT 96.780 146.220 97.100 146.280 ;
        RECT 97.715 146.220 98.005 146.265 ;
        RECT 106.990 146.220 107.130 146.420 ;
        RECT 116.345 146.375 116.635 146.420 ;
        RECT 117.480 146.360 117.800 146.420 ;
        RECT 118.350 146.560 118.640 146.605 ;
        RECT 119.780 146.560 120.100 146.620 ;
        RECT 122.530 146.605 122.745 146.760 ;
        RECT 123.460 146.700 123.780 146.960 ;
        RECT 125.315 146.900 125.605 146.945 ;
        RECT 125.760 146.900 126.080 146.960 ;
        RECT 125.315 146.760 126.080 146.900 ;
        RECT 125.315 146.715 125.605 146.760 ;
        RECT 125.760 146.700 126.080 146.760 ;
        RECT 121.610 146.560 121.900 146.605 ;
        RECT 118.350 146.420 121.900 146.560 ;
        RECT 118.350 146.375 118.640 146.420 ;
        RECT 119.780 146.360 120.100 146.420 ;
        RECT 121.610 146.375 121.900 146.420 ;
        RECT 122.530 146.560 122.820 146.605 ;
        RECT 124.390 146.560 124.680 146.605 ;
        RECT 122.530 146.420 124.680 146.560 ;
        RECT 122.530 146.375 122.820 146.420 ;
        RECT 124.390 146.375 124.680 146.420 ;
        RECT 96.780 146.080 107.130 146.220 ;
        RECT 107.820 146.220 108.140 146.280 ;
        RECT 109.200 146.220 109.520 146.280 ;
        RECT 107.820 146.080 109.520 146.220 ;
        RECT 96.780 146.020 97.100 146.080 ;
        RECT 97.715 146.035 98.005 146.080 ;
        RECT 107.820 146.020 108.140 146.080 ;
        RECT 109.200 146.020 109.520 146.080 ;
        RECT 113.355 146.220 113.645 146.265 ;
        RECT 113.800 146.220 114.120 146.280 ;
        RECT 117.020 146.220 117.340 146.280 ;
        RECT 113.355 146.080 117.340 146.220 ;
        RECT 113.355 146.035 113.645 146.080 ;
        RECT 113.800 146.020 114.120 146.080 ;
        RECT 117.020 146.020 117.340 146.080 ;
        RECT 14.370 145.400 127.530 145.880 ;
        RECT 19.960 145.000 20.280 145.260 ;
        RECT 22.720 145.245 23.040 145.260 ;
        RECT 22.505 145.015 23.040 145.245 ;
        RECT 50.780 145.200 51.100 145.260 ;
        RECT 22.720 145.000 23.040 145.015 ;
        RECT 40.750 145.060 51.100 145.200 ;
        RECT 21.355 144.860 21.645 144.905 ;
        RECT 24.510 144.860 24.800 144.905 ;
        RECT 27.770 144.860 28.060 144.905 ;
        RECT 21.355 144.720 28.060 144.860 ;
        RECT 21.355 144.675 21.645 144.720 ;
        RECT 24.510 144.675 24.800 144.720 ;
        RECT 27.770 144.675 28.060 144.720 ;
        RECT 28.690 144.860 28.980 144.905 ;
        RECT 30.550 144.860 30.840 144.905 ;
        RECT 28.690 144.720 30.840 144.860 ;
        RECT 28.690 144.675 28.980 144.720 ;
        RECT 30.550 144.675 30.840 144.720 ;
        RECT 19.515 144.520 19.805 144.565 ;
        RECT 20.895 144.520 21.185 144.565 ;
        RECT 19.515 144.380 21.185 144.520 ;
        RECT 19.515 144.335 19.805 144.380 ;
        RECT 20.895 144.335 21.185 144.380 ;
        RECT 26.370 144.520 26.660 144.565 ;
        RECT 28.690 144.520 28.905 144.675 ;
        RECT 26.370 144.380 28.905 144.520 ;
        RECT 30.080 144.520 30.400 144.580 ;
        RECT 40.750 144.565 40.890 145.060 ;
        RECT 50.780 145.000 51.100 145.060 ;
        RECT 51.700 145.000 52.020 145.260 ;
        RECT 53.540 145.000 53.860 145.260 ;
        RECT 80.680 145.200 81.000 145.260 ;
        RECT 80.310 145.060 81.000 145.200 ;
        RECT 41.135 144.860 41.425 144.905 ;
        RECT 44.290 144.860 44.580 144.905 ;
        RECT 47.550 144.860 47.840 144.905 ;
        RECT 41.135 144.720 47.840 144.860 ;
        RECT 41.135 144.675 41.425 144.720 ;
        RECT 44.290 144.675 44.580 144.720 ;
        RECT 47.550 144.675 47.840 144.720 ;
        RECT 48.470 144.860 48.760 144.905 ;
        RECT 50.330 144.860 50.620 144.905 ;
        RECT 48.470 144.720 50.620 144.860 ;
        RECT 50.870 144.860 51.010 145.000 ;
        RECT 54.920 144.860 55.240 144.920 ;
        RECT 59.060 144.860 59.380 144.920 ;
        RECT 65.055 144.860 65.345 144.905 ;
        RECT 50.870 144.720 58.370 144.860 ;
        RECT 48.470 144.675 48.760 144.720 ;
        RECT 50.330 144.675 50.620 144.720 ;
        RECT 40.675 144.520 40.965 144.565 ;
        RECT 30.080 144.380 40.965 144.520 ;
        RECT 26.370 144.335 26.660 144.380 ;
        RECT 20.970 143.500 21.110 144.335 ;
        RECT 30.080 144.320 30.400 144.380 ;
        RECT 40.675 144.335 40.965 144.380 ;
        RECT 46.150 144.520 46.440 144.565 ;
        RECT 48.470 144.520 48.685 144.675 ;
        RECT 54.920 144.660 55.240 144.720 ;
        RECT 46.150 144.380 48.685 144.520 ;
        RECT 46.150 144.335 46.440 144.380 ;
        RECT 49.400 144.320 49.720 144.580 ;
        RECT 58.230 144.565 58.370 144.720 ;
        RECT 59.060 144.720 65.345 144.860 ;
        RECT 59.060 144.660 59.380 144.720 ;
        RECT 65.055 144.675 65.345 144.720 ;
        RECT 79.300 144.660 79.620 144.920 ;
        RECT 54.015 144.520 54.305 144.565 ;
        RECT 49.950 144.380 54.305 144.520 ;
        RECT 28.700 144.180 29.020 144.240 ;
        RECT 29.635 144.180 29.925 144.225 ;
        RECT 28.700 144.040 29.925 144.180 ;
        RECT 28.700 143.980 29.020 144.040 ;
        RECT 29.635 143.995 29.925 144.040 ;
        RECT 31.475 144.180 31.765 144.225 ;
        RECT 36.060 144.180 36.380 144.240 ;
        RECT 31.475 144.040 36.380 144.180 ;
        RECT 31.475 143.995 31.765 144.040 ;
        RECT 36.060 143.980 36.380 144.040 ;
        RECT 42.285 144.180 42.575 144.225 ;
        RECT 49.950 144.180 50.090 144.380 ;
        RECT 54.015 144.335 54.305 144.380 ;
        RECT 58.155 144.335 58.445 144.565 ;
        RECT 65.500 144.320 65.820 144.580 ;
        RECT 80.310 144.565 80.450 145.060 ;
        RECT 80.680 145.000 81.000 145.060 ;
        RECT 85.740 145.000 86.060 145.260 ;
        RECT 90.800 145.000 91.120 145.260 ;
        RECT 96.780 145.000 97.100 145.260 ;
        RECT 117.020 145.000 117.340 145.260 ;
        RECT 119.780 145.000 120.100 145.260 ;
        RECT 122.095 145.200 122.385 145.245 ;
        RECT 123.460 145.200 123.780 145.260 ;
        RECT 122.095 145.060 123.780 145.200 ;
        RECT 122.095 145.015 122.385 145.060 ;
        RECT 123.460 145.000 123.780 145.060 ;
        RECT 106.915 144.860 107.205 144.905 ;
        RECT 109.675 144.860 109.965 144.905 ;
        RECT 106.915 144.720 109.965 144.860 ;
        RECT 106.915 144.675 107.205 144.720 ;
        RECT 109.675 144.675 109.965 144.720 ;
        RECT 112.050 144.720 116.790 144.860 ;
        RECT 80.235 144.335 80.525 144.565 ;
        RECT 80.695 144.520 80.985 144.565 ;
        RECT 81.140 144.520 81.460 144.580 ;
        RECT 80.695 144.380 81.460 144.520 ;
        RECT 80.695 144.335 80.985 144.380 ;
        RECT 81.140 144.320 81.460 144.380 ;
        RECT 84.360 144.520 84.680 144.580 ;
        RECT 86.215 144.520 86.505 144.565 ;
        RECT 89.895 144.520 90.185 144.565 ;
        RECT 84.360 144.380 86.505 144.520 ;
        RECT 84.360 144.320 84.680 144.380 ;
        RECT 86.215 144.335 86.505 144.380 ;
        RECT 88.130 144.380 90.185 144.520 ;
        RECT 50.320 144.180 50.640 144.240 ;
        RECT 42.285 144.040 50.640 144.180 ;
        RECT 42.285 143.995 42.575 144.040 ;
        RECT 50.320 143.980 50.640 144.040 ;
        RECT 51.255 143.995 51.545 144.225 ;
        RECT 54.460 144.180 54.780 144.240 ;
        RECT 54.935 144.180 55.225 144.225 ;
        RECT 64.580 144.180 64.900 144.240 ;
        RECT 69.180 144.180 69.500 144.240 ;
        RECT 54.460 144.040 69.500 144.180 ;
        RECT 26.370 143.840 26.660 143.885 ;
        RECT 29.150 143.840 29.440 143.885 ;
        RECT 31.010 143.840 31.300 143.885 ;
        RECT 26.370 143.700 31.300 143.840 ;
        RECT 26.370 143.655 26.660 143.700 ;
        RECT 29.150 143.655 29.440 143.700 ;
        RECT 31.010 143.655 31.300 143.700 ;
        RECT 46.150 143.840 46.440 143.885 ;
        RECT 48.930 143.840 49.220 143.885 ;
        RECT 50.790 143.840 51.080 143.885 ;
        RECT 46.150 143.700 51.080 143.840 ;
        RECT 51.330 143.840 51.470 143.995 ;
        RECT 54.460 143.980 54.780 144.040 ;
        RECT 54.935 143.995 55.225 144.040 ;
        RECT 64.580 143.980 64.900 144.040 ;
        RECT 69.180 143.980 69.500 144.040 ;
        RECT 84.820 143.980 85.140 144.240 ;
        RECT 63.660 143.840 63.980 143.900 ;
        RECT 51.330 143.700 63.980 143.840 ;
        RECT 46.150 143.655 46.440 143.700 ;
        RECT 48.930 143.655 49.220 143.700 ;
        RECT 50.790 143.655 51.080 143.700 ;
        RECT 63.660 143.640 63.980 143.700 ;
        RECT 68.720 143.840 69.040 143.900 ;
        RECT 70.560 143.840 70.880 143.900 ;
        RECT 68.720 143.700 70.880 143.840 ;
        RECT 68.720 143.640 69.040 143.700 ;
        RECT 70.560 143.640 70.880 143.700 ;
        RECT 75.160 143.840 75.480 143.900 ;
        RECT 88.130 143.885 88.270 144.380 ;
        RECT 89.895 144.335 90.185 144.380 ;
        RECT 94.035 144.520 94.325 144.565 ;
        RECT 96.320 144.520 96.640 144.580 ;
        RECT 94.035 144.380 96.640 144.520 ;
        RECT 94.035 144.335 94.325 144.380 ;
        RECT 96.320 144.320 96.640 144.380 ;
        RECT 108.295 144.520 108.585 144.565 ;
        RECT 108.740 144.520 109.060 144.580 ;
        RECT 108.295 144.380 109.060 144.520 ;
        RECT 108.295 144.335 108.585 144.380 ;
        RECT 108.740 144.320 109.060 144.380 ;
        RECT 109.200 144.520 109.520 144.580 ;
        RECT 111.055 144.520 111.345 144.565 ;
        RECT 109.200 144.380 111.345 144.520 ;
        RECT 109.200 144.320 109.520 144.380 ;
        RECT 111.055 144.335 111.345 144.380 ;
        RECT 107.835 144.180 108.125 144.225 ;
        RECT 110.120 144.180 110.440 144.240 ;
        RECT 107.835 144.040 110.440 144.180 ;
        RECT 107.835 143.995 108.125 144.040 ;
        RECT 110.120 143.980 110.440 144.040 ;
        RECT 81.615 143.840 81.905 143.885 ;
        RECT 75.160 143.700 81.905 143.840 ;
        RECT 75.160 143.640 75.480 143.700 ;
        RECT 81.615 143.655 81.905 143.700 ;
        RECT 88.055 143.655 88.345 143.885 ;
        RECT 108.740 143.840 109.060 143.900 ;
        RECT 109.215 143.840 109.505 143.885 ;
        RECT 111.130 143.840 111.270 144.335 ;
        RECT 111.500 144.320 111.820 144.580 ;
        RECT 112.050 144.565 112.190 144.720 ;
        RECT 111.975 144.335 112.265 144.565 ;
        RECT 112.420 144.520 112.740 144.580 ;
        RECT 112.895 144.520 113.185 144.565 ;
        RECT 112.420 144.380 113.185 144.520 ;
        RECT 112.420 144.320 112.740 144.380 ;
        RECT 112.895 144.335 113.185 144.380 ;
        RECT 113.340 144.180 113.660 144.240 ;
        RECT 116.650 144.225 116.790 144.720 ;
        RECT 119.320 144.320 119.640 144.580 ;
        RECT 121.175 144.335 121.465 144.565 ;
        RECT 115.655 144.180 115.945 144.225 ;
        RECT 113.340 144.040 115.945 144.180 ;
        RECT 113.340 143.980 113.660 144.040 ;
        RECT 115.655 143.995 115.945 144.040 ;
        RECT 116.575 144.180 116.865 144.225 ;
        RECT 117.480 144.180 117.800 144.240 ;
        RECT 121.250 144.180 121.390 144.335 ;
        RECT 116.575 144.040 117.800 144.180 ;
        RECT 116.575 143.995 116.865 144.040 ;
        RECT 117.480 143.980 117.800 144.040 ;
        RECT 118.950 144.040 121.390 144.180 ;
        RECT 118.950 143.885 119.090 144.040 ;
        RECT 108.740 143.700 109.505 143.840 ;
        RECT 108.740 143.640 109.060 143.700 ;
        RECT 109.215 143.655 109.505 143.700 ;
        RECT 110.210 143.700 111.270 143.840 ;
        RECT 110.210 143.560 110.350 143.700 ;
        RECT 118.875 143.655 119.165 143.885 ;
        RECT 29.620 143.500 29.940 143.560 ;
        RECT 20.970 143.360 29.940 143.500 ;
        RECT 29.620 143.300 29.940 143.360 ;
        RECT 58.600 143.300 58.920 143.560 ;
        RECT 67.355 143.500 67.645 143.545 ;
        RECT 69.640 143.500 69.960 143.560 ;
        RECT 67.355 143.360 69.960 143.500 ;
        RECT 67.355 143.315 67.645 143.360 ;
        RECT 69.640 143.300 69.960 143.360 ;
        RECT 80.680 143.300 81.000 143.560 ;
        RECT 108.295 143.500 108.585 143.545 ;
        RECT 109.660 143.500 109.980 143.560 ;
        RECT 108.295 143.360 109.980 143.500 ;
        RECT 108.295 143.315 108.585 143.360 ;
        RECT 109.660 143.300 109.980 143.360 ;
        RECT 110.120 143.300 110.440 143.560 ;
        RECT 14.370 142.680 127.530 143.160 ;
        RECT 35.600 142.280 35.920 142.540 ;
        RECT 48.035 142.295 48.325 142.525 ;
        RECT 44.800 142.140 45.120 142.200 ;
        RECT 48.110 142.140 48.250 142.295 ;
        RECT 59.060 142.280 59.380 142.540 ;
        RECT 108.740 142.480 109.060 142.540 ;
        RECT 111.500 142.480 111.820 142.540 ;
        RECT 108.740 142.340 111.820 142.480 ;
        RECT 108.740 142.280 109.060 142.340 ;
        RECT 111.500 142.280 111.820 142.340 ;
        RECT 44.800 142.000 48.250 142.140 ;
        RECT 62.395 142.140 62.685 142.185 ;
        RECT 65.515 142.140 65.805 142.185 ;
        RECT 67.405 142.140 67.695 142.185 ;
        RECT 68.720 142.140 69.040 142.200 ;
        RECT 62.395 142.000 67.695 142.140 ;
        RECT 44.800 141.940 45.120 142.000 ;
        RECT 62.395 141.955 62.685 142.000 ;
        RECT 65.515 141.955 65.805 142.000 ;
        RECT 67.405 141.955 67.695 142.000 ;
        RECT 67.890 142.000 69.040 142.140 ;
        RECT 34.220 141.800 34.540 141.860 ;
        RECT 35.615 141.800 35.905 141.845 ;
        RECT 34.220 141.660 35.905 141.800 ;
        RECT 34.220 141.600 34.540 141.660 ;
        RECT 35.615 141.615 35.905 141.660 ;
        RECT 46.180 141.800 46.500 141.860 ;
        RECT 48.495 141.800 48.785 141.845 ;
        RECT 46.180 141.660 48.785 141.800 ;
        RECT 46.180 141.600 46.500 141.660 ;
        RECT 48.495 141.615 48.785 141.660 ;
        RECT 53.080 141.800 53.400 141.860 ;
        RECT 56.315 141.800 56.605 141.845 ;
        RECT 59.535 141.800 59.825 141.845 ;
        RECT 67.890 141.800 68.030 142.000 ;
        RECT 68.720 141.940 69.040 142.000 ;
        RECT 53.080 141.660 54.230 141.800 ;
        RECT 53.080 141.600 53.400 141.660 ;
        RECT 34.680 141.460 35.000 141.520 ;
        RECT 35.155 141.460 35.445 141.505 ;
        RECT 34.680 141.320 35.445 141.460 ;
        RECT 34.680 141.260 35.000 141.320 ;
        RECT 35.155 141.275 35.445 141.320 ;
        RECT 45.720 141.460 46.040 141.520 ;
        RECT 48.035 141.460 48.325 141.505 ;
        RECT 45.720 141.320 48.325 141.460 ;
        RECT 45.720 141.260 46.040 141.320 ;
        RECT 48.035 141.275 48.325 141.320 ;
        RECT 53.540 141.260 53.860 141.520 ;
        RECT 54.090 141.505 54.230 141.660 ;
        RECT 54.550 141.660 59.825 141.800 ;
        RECT 54.550 141.505 54.690 141.660 ;
        RECT 56.315 141.615 56.605 141.660 ;
        RECT 59.535 141.615 59.825 141.660 ;
        RECT 60.070 141.660 68.030 141.800 ;
        RECT 54.015 141.275 54.305 141.505 ;
        RECT 54.475 141.275 54.765 141.505 ;
        RECT 55.395 141.460 55.685 141.505 ;
        RECT 55.840 141.460 56.160 141.520 ;
        RECT 60.070 141.460 60.210 141.660 ;
        RECT 68.260 141.600 68.580 141.860 ;
        RECT 112.880 141.800 113.200 141.860 ;
        RECT 116.115 141.800 116.405 141.845 ;
        RECT 112.880 141.660 116.405 141.800 ;
        RECT 112.880 141.600 113.200 141.660 ;
        RECT 116.115 141.615 116.405 141.660 ;
        RECT 55.395 141.320 56.160 141.460 ;
        RECT 55.395 141.275 55.685 141.320 ;
        RECT 55.840 141.260 56.160 141.320 ;
        RECT 57.770 141.320 60.210 141.460 ;
        RECT 36.535 141.120 36.825 141.165 ;
        RECT 39.280 141.120 39.600 141.180 ;
        RECT 36.535 140.980 39.600 141.120 ;
        RECT 36.535 140.935 36.825 140.980 ;
        RECT 39.280 140.920 39.600 140.980 ;
        RECT 49.415 141.120 49.705 141.165 ;
        RECT 52.175 141.120 52.465 141.165 ;
        RECT 49.415 140.980 52.465 141.120 ;
        RECT 49.415 140.935 49.705 140.980 ;
        RECT 52.175 140.935 52.465 140.980 ;
        RECT 29.160 140.780 29.480 140.840 ;
        RECT 34.235 140.780 34.525 140.825 ;
        RECT 29.160 140.640 34.525 140.780 ;
        RECT 29.160 140.580 29.480 140.640 ;
        RECT 34.235 140.595 34.525 140.640 ;
        RECT 47.115 140.780 47.405 140.825 ;
        RECT 57.770 140.780 57.910 141.320 ;
        RECT 58.600 141.120 58.920 141.180 ;
        RECT 61.315 141.165 61.605 141.480 ;
        RECT 62.395 141.460 62.685 141.505 ;
        RECT 65.975 141.460 66.265 141.505 ;
        RECT 67.810 141.460 68.100 141.505 ;
        RECT 62.395 141.320 68.100 141.460 ;
        RECT 62.395 141.275 62.685 141.320 ;
        RECT 65.975 141.275 66.265 141.320 ;
        RECT 67.810 141.275 68.100 141.320 ;
        RECT 69.640 141.260 69.960 141.520 ;
        RECT 70.560 141.460 70.880 141.520 ;
        RECT 72.415 141.460 72.705 141.505 ;
        RECT 70.560 141.320 72.705 141.460 ;
        RECT 70.560 141.260 70.880 141.320 ;
        RECT 72.415 141.275 72.705 141.320 ;
        RECT 117.480 141.260 117.800 141.520 ;
        RECT 119.320 141.460 119.640 141.520 ;
        RECT 119.795 141.460 120.085 141.505 ;
        RECT 119.320 141.320 120.085 141.460 ;
        RECT 119.320 141.260 119.640 141.320 ;
        RECT 119.795 141.275 120.085 141.320 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 61.015 141.120 61.605 141.165 ;
        RECT 64.255 141.120 64.905 141.165 ;
        RECT 58.600 140.980 64.905 141.120 ;
        RECT 58.600 140.920 58.920 140.980 ;
        RECT 61.015 140.935 61.305 140.980 ;
        RECT 64.255 140.935 64.905 140.980 ;
        RECT 66.895 141.120 67.185 141.165 ;
        RECT 66.895 140.980 68.950 141.120 ;
        RECT 66.895 140.935 67.185 140.980 ;
        RECT 47.115 140.640 57.910 140.780 ;
        RECT 63.660 140.780 63.980 140.840 ;
        RECT 68.260 140.780 68.580 140.840 ;
        RECT 68.810 140.825 68.950 140.980 ;
        RECT 63.660 140.640 68.580 140.780 ;
        RECT 47.115 140.595 47.405 140.640 ;
        RECT 63.660 140.580 63.980 140.640 ;
        RECT 68.260 140.580 68.580 140.640 ;
        RECT 68.735 140.595 69.025 140.825 ;
        RECT 71.940 140.580 72.260 140.840 ;
        RECT 117.020 140.580 117.340 140.840 ;
        RECT 119.320 140.580 119.640 140.840 ;
        RECT 120.240 140.580 120.560 140.840 ;
        RECT 14.370 139.960 127.530 140.440 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 35.600 139.560 35.920 139.820 ;
        RECT 38.375 139.575 38.665 139.805 ;
        RECT 39.280 139.760 39.600 139.820 ;
        RECT 59.075 139.760 59.365 139.805 ;
        RECT 60.900 139.760 61.220 139.820 ;
        RECT 63.675 139.760 63.965 139.805 ;
        RECT 39.280 139.620 59.365 139.760 ;
        RECT 18.070 139.420 18.360 139.465 ;
        RECT 19.040 139.420 19.360 139.480 ;
        RECT 21.330 139.420 21.620 139.465 ;
        RECT 18.070 139.280 21.620 139.420 ;
        RECT 18.070 139.235 18.360 139.280 ;
        RECT 19.040 139.220 19.360 139.280 ;
        RECT 21.330 139.235 21.620 139.280 ;
        RECT 22.250 139.420 22.540 139.465 ;
        RECT 24.110 139.420 24.400 139.465 ;
        RECT 38.450 139.420 38.590 139.575 ;
        RECT 39.280 139.560 39.600 139.620 ;
        RECT 59.075 139.575 59.365 139.620 ;
        RECT 59.610 139.620 63.965 139.760 ;
        RECT 22.250 139.280 24.400 139.420 ;
        RECT 22.250 139.235 22.540 139.280 ;
        RECT 24.110 139.235 24.400 139.280 ;
        RECT 36.380 139.280 38.590 139.420 ;
        RECT 40.675 139.420 40.965 139.465 ;
        RECT 41.120 139.420 41.440 139.480 ;
        RECT 59.610 139.420 59.750 139.620 ;
        RECT 60.900 139.560 61.220 139.620 ;
        RECT 63.675 139.575 63.965 139.620 ;
        RECT 65.500 139.760 65.820 139.820 ;
        RECT 67.585 139.760 67.875 139.805 ;
        RECT 65.500 139.620 67.875 139.760 ;
        RECT 65.500 139.560 65.820 139.620 ;
        RECT 67.585 139.575 67.875 139.620 ;
        RECT 81.140 139.560 81.460 139.820 ;
        RECT 84.360 139.760 84.680 139.820 ;
        RECT 85.755 139.760 86.045 139.805 ;
        RECT 84.360 139.620 86.045 139.760 ;
        RECT 84.360 139.560 84.680 139.620 ;
        RECT 85.755 139.575 86.045 139.620 ;
        RECT 88.055 139.575 88.345 139.805 ;
        RECT 65.590 139.420 65.730 139.560 ;
        RECT 40.675 139.280 41.440 139.420 ;
        RECT 19.930 139.080 20.220 139.125 ;
        RECT 22.250 139.080 22.465 139.235 ;
        RECT 19.930 138.940 22.465 139.080 ;
        RECT 34.680 139.080 35.000 139.140 ;
        RECT 35.600 139.080 35.920 139.140 ;
        RECT 36.380 139.080 36.520 139.280 ;
        RECT 40.675 139.235 40.965 139.280 ;
        RECT 41.120 139.220 41.440 139.280 ;
        RECT 55.010 139.280 59.750 139.420 ;
        RECT 61.450 139.280 65.730 139.420 ;
        RECT 69.590 139.420 69.880 139.465 ;
        RECT 71.940 139.420 72.260 139.480 ;
        RECT 72.850 139.420 73.140 139.465 ;
        RECT 69.590 139.280 73.140 139.420 ;
        RECT 34.680 138.940 35.195 139.080 ;
        RECT 35.600 138.940 36.520 139.080 ;
        RECT 39.295 139.080 39.585 139.125 ;
        RECT 55.010 139.080 55.150 139.280 ;
        RECT 39.295 138.940 55.150 139.080 ;
        RECT 19.930 138.895 20.220 138.940 ;
        RECT 34.680 138.880 35.000 138.940 ;
        RECT 35.600 138.880 35.920 138.940 ;
        RECT 39.295 138.895 39.585 138.940 ;
        RECT 55.395 138.895 55.685 139.125 ;
        RECT 23.180 138.540 23.500 138.800 ;
        RECT 25.035 138.740 25.325 138.785 ;
        RECT 29.620 138.740 29.940 138.800 ;
        RECT 25.035 138.600 29.940 138.740 ;
        RECT 25.035 138.555 25.325 138.600 ;
        RECT 29.620 138.540 29.940 138.600 ;
        RECT 30.080 138.740 30.400 138.800 ;
        RECT 33.775 138.740 34.065 138.785 ;
        RECT 30.080 138.600 34.065 138.740 ;
        RECT 30.080 138.540 30.400 138.600 ;
        RECT 33.775 138.555 34.065 138.600 ;
        RECT 39.740 138.540 40.060 138.800 ;
        RECT 54.920 138.740 55.240 138.800 ;
        RECT 55.470 138.740 55.610 138.895 ;
        RECT 55.840 138.880 56.160 139.140 ;
        RECT 60.440 138.880 60.760 139.140 ;
        RECT 61.450 139.125 61.590 139.280 ;
        RECT 69.590 139.235 69.880 139.280 ;
        RECT 71.940 139.220 72.260 139.280 ;
        RECT 72.850 139.235 73.140 139.280 ;
        RECT 73.770 139.420 74.060 139.465 ;
        RECT 75.630 139.420 75.920 139.465 ;
        RECT 73.770 139.280 75.920 139.420 ;
        RECT 73.770 139.235 74.060 139.280 ;
        RECT 75.630 139.235 75.920 139.280 ;
        RECT 79.760 139.420 80.080 139.480 ;
        RECT 81.230 139.420 81.370 139.560 ;
        RECT 84.450 139.420 84.590 139.560 ;
        RECT 79.760 139.280 81.370 139.420 ;
        RECT 81.690 139.280 84.590 139.420 ;
        RECT 60.915 138.895 61.205 139.125 ;
        RECT 61.375 138.895 61.665 139.125 ;
        RECT 62.295 138.895 62.585 139.125 ;
        RECT 54.920 138.600 55.610 138.740 ;
        RECT 54.920 138.540 55.240 138.600 ;
        RECT 19.930 138.400 20.220 138.445 ;
        RECT 22.710 138.400 23.000 138.445 ;
        RECT 24.570 138.400 24.860 138.445 ;
        RECT 19.930 138.260 24.860 138.400 ;
        RECT 19.930 138.215 20.220 138.260 ;
        RECT 22.710 138.215 23.000 138.260 ;
        RECT 24.570 138.215 24.860 138.260 ;
        RECT 16.065 138.060 16.355 138.105 ;
        RECT 22.260 138.060 22.580 138.120 ;
        RECT 16.065 137.920 22.580 138.060 ;
        RECT 16.065 137.875 16.355 137.920 ;
        RECT 22.260 137.860 22.580 137.920 ;
        RECT 34.220 138.060 34.540 138.120 ;
        RECT 39.295 138.060 39.585 138.105 ;
        RECT 34.220 137.920 39.585 138.060 ;
        RECT 34.220 137.860 34.540 137.920 ;
        RECT 39.295 137.875 39.585 137.920 ;
        RECT 47.560 138.060 47.880 138.120 ;
        RECT 49.860 138.060 50.180 138.120 ;
        RECT 53.540 138.060 53.860 138.120 ;
        RECT 47.560 137.920 53.860 138.060 ;
        RECT 60.990 138.060 61.130 138.895 ;
        RECT 62.370 138.400 62.510 138.895 ;
        RECT 65.040 138.880 65.360 139.140 ;
        RECT 65.515 138.895 65.805 139.125 ;
        RECT 65.590 138.740 65.730 138.895 ;
        RECT 65.960 138.880 66.280 139.140 ;
        RECT 66.895 139.080 67.185 139.125 ;
        RECT 67.800 139.080 68.120 139.140 ;
        RECT 66.895 138.940 68.120 139.080 ;
        RECT 66.895 138.895 67.185 138.940 ;
        RECT 67.800 138.880 68.120 138.940 ;
        RECT 71.450 139.080 71.740 139.125 ;
        RECT 73.770 139.080 73.985 139.235 ;
        RECT 79.760 139.220 80.080 139.280 ;
        RECT 80.770 139.125 80.910 139.280 ;
        RECT 81.690 139.125 81.830 139.280 ;
        RECT 71.450 138.940 73.985 139.080 ;
        RECT 71.450 138.895 71.740 138.940 ;
        RECT 80.695 138.895 80.985 139.125 ;
        RECT 81.155 138.895 81.445 139.125 ;
        RECT 81.615 138.895 81.905 139.125 ;
        RECT 82.535 138.895 82.825 139.125 ;
        RECT 70.100 138.740 70.420 138.800 ;
        RECT 65.590 138.600 70.420 138.740 ;
        RECT 64.120 138.400 64.440 138.460 ;
        RECT 67.340 138.400 67.660 138.460 ;
        RECT 62.370 138.260 67.660 138.400 ;
        RECT 64.120 138.200 64.440 138.260 ;
        RECT 67.340 138.200 67.660 138.260 ;
        RECT 66.420 138.060 66.740 138.120 ;
        RECT 67.890 138.060 68.030 138.600 ;
        RECT 70.100 138.540 70.420 138.600 ;
        RECT 74.700 138.540 75.020 138.800 ;
        RECT 76.555 138.555 76.845 138.785 ;
        RECT 81.230 138.740 81.370 138.895 ;
        RECT 82.060 138.740 82.380 138.800 ;
        RECT 81.230 138.600 82.380 138.740 ;
        RECT 82.610 138.740 82.750 138.895 ;
        RECT 86.200 138.880 86.520 139.140 ;
        RECT 88.130 139.080 88.270 139.575 ;
        RECT 99.950 139.420 100.240 139.465 ;
        RECT 102.300 139.420 102.620 139.480 ;
        RECT 103.210 139.420 103.500 139.465 ;
        RECT 99.950 139.280 103.500 139.420 ;
        RECT 99.950 139.235 100.240 139.280 ;
        RECT 102.300 139.220 102.620 139.280 ;
        RECT 103.210 139.235 103.500 139.280 ;
        RECT 104.130 139.420 104.420 139.465 ;
        RECT 105.990 139.420 106.280 139.465 ;
        RECT 104.130 139.280 106.280 139.420 ;
        RECT 104.130 139.235 104.420 139.280 ;
        RECT 105.990 139.235 106.280 139.280 ;
        RECT 110.120 139.420 110.440 139.480 ;
        RECT 111.960 139.420 112.280 139.480 ;
        RECT 117.020 139.465 117.340 139.480 ;
        RECT 112.895 139.420 113.185 139.465 ;
        RECT 116.805 139.420 117.340 139.465 ;
        RECT 110.120 139.280 111.730 139.420 ;
        RECT 88.975 139.080 89.265 139.125 ;
        RECT 88.130 138.940 89.265 139.080 ;
        RECT 88.975 138.895 89.265 138.940 ;
        RECT 101.810 139.080 102.100 139.125 ;
        RECT 104.130 139.080 104.345 139.235 ;
        RECT 110.120 139.220 110.440 139.280 ;
        RECT 101.810 138.940 104.345 139.080 ;
        RECT 109.200 139.080 109.520 139.140 ;
        RECT 109.675 139.080 109.965 139.125 ;
        RECT 109.200 138.940 109.965 139.080 ;
        RECT 110.595 139.070 110.885 139.140 ;
        RECT 111.590 139.125 111.730 139.280 ;
        RECT 111.960 139.280 113.185 139.420 ;
        RECT 111.960 139.220 112.280 139.280 ;
        RECT 112.895 139.235 113.185 139.280 ;
        RECT 113.890 139.280 117.340 139.420 ;
        RECT 101.810 138.895 102.100 138.940 ;
        RECT 109.200 138.880 109.520 138.940 ;
        RECT 109.675 138.895 109.965 138.940 ;
        RECT 110.210 138.930 110.885 139.070 ;
        RECT 82.980 138.740 83.300 138.800 ;
        RECT 82.610 138.600 83.300 138.740 ;
        RECT 71.450 138.400 71.740 138.445 ;
        RECT 74.230 138.400 74.520 138.445 ;
        RECT 76.090 138.400 76.380 138.445 ;
        RECT 71.450 138.260 76.380 138.400 ;
        RECT 76.630 138.400 76.770 138.555 ;
        RECT 82.060 138.540 82.380 138.600 ;
        RECT 82.980 138.540 83.300 138.600 ;
        RECT 84.820 138.540 85.140 138.800 ;
        RECT 97.945 138.740 98.235 138.785 ;
        RECT 98.620 138.740 98.940 138.800 ;
        RECT 97.945 138.600 98.940 138.740 ;
        RECT 97.945 138.555 98.235 138.600 ;
        RECT 98.620 138.540 98.940 138.600 ;
        RECT 105.060 138.540 105.380 138.800 ;
        RECT 106.915 138.555 107.205 138.785 ;
        RECT 94.020 138.400 94.340 138.460 ;
        RECT 76.630 138.260 94.340 138.400 ;
        RECT 71.450 138.215 71.740 138.260 ;
        RECT 74.230 138.215 74.520 138.260 ;
        RECT 76.090 138.215 76.380 138.260 ;
        RECT 94.020 138.200 94.340 138.260 ;
        RECT 101.810 138.400 102.100 138.445 ;
        RECT 104.590 138.400 104.880 138.445 ;
        RECT 106.450 138.400 106.740 138.445 ;
        RECT 101.810 138.260 106.740 138.400 ;
        RECT 101.810 138.215 102.100 138.260 ;
        RECT 104.590 138.215 104.880 138.260 ;
        RECT 106.450 138.215 106.740 138.260 ;
        RECT 60.990 137.920 68.030 138.060 ;
        RECT 47.560 137.860 47.880 137.920 ;
        RECT 49.860 137.860 50.180 137.920 ;
        RECT 53.540 137.860 53.860 137.920 ;
        RECT 66.420 137.860 66.740 137.920 ;
        RECT 79.300 137.860 79.620 138.120 ;
        RECT 89.895 138.060 90.185 138.105 ;
        RECT 90.800 138.060 91.120 138.120 ;
        RECT 89.895 137.920 91.120 138.060 ;
        RECT 89.895 137.875 90.185 137.920 ;
        RECT 90.800 137.860 91.120 137.920 ;
        RECT 98.160 138.060 98.480 138.120 ;
        RECT 106.990 138.060 107.130 138.555 ;
        RECT 110.210 138.400 110.350 138.930 ;
        RECT 110.595 138.910 110.885 138.930 ;
        RECT 111.055 138.895 111.345 139.125 ;
        RECT 111.515 138.895 111.805 139.125 ;
        RECT 111.130 138.740 111.270 138.895 ;
        RECT 112.420 138.880 112.740 139.140 ;
        RECT 112.510 138.740 112.650 138.880 ;
        RECT 111.130 138.600 112.650 138.740 ;
        RECT 112.420 138.400 112.740 138.460 ;
        RECT 113.890 138.400 114.030 139.280 ;
        RECT 116.805 139.235 117.340 139.280 ;
        RECT 118.810 139.420 119.100 139.465 ;
        RECT 120.240 139.420 120.560 139.480 ;
        RECT 122.070 139.420 122.360 139.465 ;
        RECT 118.810 139.280 122.360 139.420 ;
        RECT 118.810 139.235 119.100 139.280 ;
        RECT 117.020 139.220 117.340 139.235 ;
        RECT 120.240 139.220 120.560 139.280 ;
        RECT 122.070 139.235 122.360 139.280 ;
        RECT 122.990 139.420 123.280 139.465 ;
        RECT 124.850 139.420 125.140 139.465 ;
        RECT 122.990 139.280 125.140 139.420 ;
        RECT 122.990 139.235 123.280 139.280 ;
        RECT 124.850 139.235 125.140 139.280 ;
        RECT 115.195 138.895 115.485 139.125 ;
        RECT 110.210 138.260 114.030 138.400 ;
        RECT 115.270 138.400 115.410 138.895 ;
        RECT 115.640 138.880 115.960 139.140 ;
        RECT 120.670 139.080 120.960 139.125 ;
        RECT 122.990 139.080 123.205 139.235 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 120.670 138.940 123.205 139.080 ;
        RECT 120.670 138.895 120.960 138.940 ;
        RECT 123.920 138.880 124.240 139.140 ;
        RECT 125.760 138.540 126.080 138.800 ;
        RECT 119.780 138.400 120.100 138.460 ;
        RECT 115.270 138.260 120.100 138.400 ;
        RECT 112.420 138.200 112.740 138.260 ;
        RECT 119.780 138.200 120.100 138.260 ;
        RECT 120.670 138.400 120.960 138.445 ;
        RECT 123.450 138.400 123.740 138.445 ;
        RECT 125.310 138.400 125.600 138.445 ;
        RECT 120.670 138.260 125.600 138.400 ;
        RECT 120.670 138.215 120.960 138.260 ;
        RECT 123.450 138.215 123.740 138.260 ;
        RECT 125.310 138.215 125.600 138.260 ;
        RECT 121.160 138.060 121.480 138.120 ;
        RECT 124.380 138.060 124.700 138.120 ;
        RECT 125.850 138.060 125.990 138.540 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 98.160 137.920 125.990 138.060 ;
        RECT 98.160 137.860 98.480 137.920 ;
        RECT 121.160 137.860 121.480 137.920 ;
        RECT 124.380 137.860 124.700 137.920 ;
        RECT 14.370 137.240 127.530 137.720 ;
        RECT 34.220 136.840 34.540 137.100 ;
        RECT 35.615 136.855 35.905 137.085 ;
        RECT 37.900 137.040 38.220 137.100 ;
        RECT 38.375 137.040 38.665 137.085 ;
        RECT 37.900 136.900 38.665 137.040 ;
        RECT 33.760 136.700 34.080 136.760 ;
        RECT 35.690 136.700 35.830 136.855 ;
        RECT 37.900 136.840 38.220 136.900 ;
        RECT 38.375 136.855 38.665 136.900 ;
        RECT 44.340 136.840 44.660 137.100 ;
        RECT 48.020 137.040 48.340 137.100 ;
        RECT 50.780 137.040 51.100 137.100 ;
        RECT 53.080 137.040 53.400 137.100 ;
        RECT 48.020 136.900 53.400 137.040 ;
        RECT 48.020 136.840 48.340 136.900 ;
        RECT 50.780 136.840 51.100 136.900 ;
        RECT 53.080 136.840 53.400 136.900 ;
        RECT 60.440 137.040 60.760 137.100 ;
        RECT 60.440 136.900 62.510 137.040 ;
        RECT 60.440 136.840 60.760 136.900 ;
        RECT 60.915 136.700 61.205 136.745 ;
        RECT 33.760 136.560 35.830 136.700 ;
        RECT 39.830 136.560 61.205 136.700 ;
        RECT 33.760 136.500 34.080 136.560 ;
        RECT 21.340 136.360 21.660 136.420 ;
        RECT 22.735 136.360 23.025 136.405 ;
        RECT 21.340 136.220 23.025 136.360 ;
        RECT 21.340 136.160 21.660 136.220 ;
        RECT 22.735 136.175 23.025 136.220 ;
        RECT 31.000 136.160 31.320 136.420 ;
        RECT 35.140 136.360 35.460 136.420 ;
        RECT 36.075 136.360 36.365 136.405 ;
        RECT 35.140 136.220 36.365 136.360 ;
        RECT 35.140 136.160 35.460 136.220 ;
        RECT 36.075 136.175 36.365 136.220 ;
        RECT 38.820 136.160 39.140 136.420 ;
        RECT 21.815 136.020 22.105 136.065 ;
        RECT 22.260 136.020 22.580 136.080 ;
        RECT 21.815 135.880 22.580 136.020 ;
        RECT 21.815 135.835 22.105 135.880 ;
        RECT 22.260 135.820 22.580 135.880 ;
        RECT 32.395 135.835 32.685 136.065 ;
        RECT 33.300 136.020 33.620 136.080 ;
        RECT 34.680 136.020 35.000 136.080 ;
        RECT 33.300 135.880 35.000 136.020 ;
        RECT 30.080 135.680 30.400 135.740 ;
        RECT 22.350 135.540 30.400 135.680 ;
        RECT 18.580 135.340 18.900 135.400 ;
        RECT 19.975 135.340 20.265 135.385 ;
        RECT 18.580 135.200 20.265 135.340 ;
        RECT 18.580 135.140 18.900 135.200 ;
        RECT 19.975 135.155 20.265 135.200 ;
        RECT 21.800 135.340 22.120 135.400 ;
        RECT 22.350 135.385 22.490 135.540 ;
        RECT 30.080 135.480 30.400 135.540 ;
        RECT 32.470 135.400 32.610 135.835 ;
        RECT 33.300 135.820 33.620 135.880 ;
        RECT 34.680 135.820 35.000 135.880 ;
        RECT 35.615 136.020 35.905 136.065 ;
        RECT 36.520 136.020 36.840 136.080 ;
        RECT 35.615 135.880 36.840 136.020 ;
        RECT 35.615 135.835 35.905 135.880 ;
        RECT 36.520 135.820 36.840 135.880 ;
        RECT 38.360 135.820 38.680 136.080 ;
        RECT 39.830 136.065 39.970 136.560 ;
        RECT 60.915 136.515 61.205 136.560 ;
        RECT 62.370 136.700 62.510 136.900 ;
        RECT 65.040 136.840 65.360 137.100 ;
        RECT 71.035 137.040 71.325 137.085 ;
        RECT 74.700 137.040 75.020 137.100 ;
        RECT 71.035 136.900 75.020 137.040 ;
        RECT 71.035 136.855 71.325 136.900 ;
        RECT 74.700 136.840 75.020 136.900 ;
        RECT 79.315 137.040 79.605 137.085 ;
        RECT 79.760 137.040 80.080 137.100 ;
        RECT 83.685 137.040 83.975 137.085 ;
        RECT 84.360 137.040 84.680 137.100 ;
        RECT 79.315 136.900 80.080 137.040 ;
        RECT 79.315 136.855 79.605 136.900 ;
        RECT 79.760 136.840 80.080 136.900 ;
        RECT 81.230 136.900 82.750 137.040 ;
        RECT 65.130 136.700 65.270 136.840 ;
        RECT 74.240 136.700 74.560 136.760 ;
        RECT 62.370 136.560 74.560 136.700 ;
        RECT 45.260 136.160 45.580 136.420 ;
        RECT 50.320 136.360 50.640 136.420 ;
        RECT 48.570 136.220 50.640 136.360 ;
        RECT 39.755 135.835 40.045 136.065 ;
        RECT 42.040 136.020 42.360 136.080 ;
        RECT 44.355 136.020 44.645 136.065 ;
        RECT 42.040 135.880 44.645 136.020 ;
        RECT 42.040 135.820 42.360 135.880 ;
        RECT 44.355 135.835 44.645 135.880 ;
        RECT 45.350 135.880 47.330 136.020 ;
        RECT 36.995 135.680 37.285 135.725 ;
        RECT 45.350 135.680 45.490 135.880 ;
        RECT 36.995 135.540 45.490 135.680 ;
        RECT 45.735 135.680 46.025 135.725 ;
        RECT 46.195 135.680 46.485 135.725 ;
        RECT 45.735 135.540 46.485 135.680 ;
        RECT 47.190 135.680 47.330 135.880 ;
        RECT 47.560 135.820 47.880 136.080 ;
        RECT 48.020 135.820 48.340 136.080 ;
        RECT 48.570 136.065 48.710 136.220 ;
        RECT 50.320 136.160 50.640 136.220 ;
        RECT 54.015 136.360 54.305 136.405 ;
        RECT 54.460 136.360 54.780 136.420 ;
        RECT 54.015 136.220 54.780 136.360 ;
        RECT 54.015 136.175 54.305 136.220 ;
        RECT 54.460 136.160 54.780 136.220 ;
        RECT 48.495 135.835 48.785 136.065 ;
        RECT 49.415 135.835 49.705 136.065 ;
        RECT 50.410 136.020 50.550 136.160 ;
        RECT 62.370 136.065 62.510 136.560 ;
        RECT 74.240 136.500 74.560 136.560 ;
        RECT 77.015 136.700 77.305 136.745 ;
        RECT 81.230 136.700 81.370 136.900 ;
        RECT 82.060 136.700 82.380 136.760 ;
        RECT 77.015 136.560 81.370 136.700 ;
        RECT 81.690 136.560 82.380 136.700 ;
        RECT 82.610 136.700 82.750 136.900 ;
        RECT 83.685 136.900 84.680 137.040 ;
        RECT 83.685 136.855 83.975 136.900 ;
        RECT 84.360 136.840 84.680 136.900 ;
        RECT 84.820 137.040 85.140 137.100 ;
        RECT 105.060 137.040 105.380 137.100 ;
        RECT 106.915 137.040 107.205 137.085 ;
        RECT 84.820 136.900 95.630 137.040 ;
        RECT 84.820 136.840 85.140 136.900 ;
        RECT 86.660 136.700 86.980 136.760 ;
        RECT 82.610 136.560 86.980 136.700 ;
        RECT 77.015 136.515 77.305 136.560 ;
        RECT 65.055 136.360 65.345 136.405 ;
        RECT 65.500 136.360 65.820 136.420 ;
        RECT 73.780 136.360 74.100 136.420 ;
        RECT 62.830 136.220 63.890 136.360 ;
        RECT 62.830 136.065 62.970 136.220 ;
        RECT 54.935 136.020 55.225 136.065 ;
        RECT 57.695 136.020 57.985 136.065 ;
        RECT 50.410 135.880 55.225 136.020 ;
        RECT 54.935 135.835 55.225 135.880 ;
        RECT 56.850 135.880 57.985 136.020 ;
        RECT 48.940 135.680 49.260 135.740 ;
        RECT 47.190 135.540 49.260 135.680 ;
        RECT 49.490 135.680 49.630 135.835 ;
        RECT 50.320 135.680 50.640 135.740 ;
        RECT 52.160 135.680 52.480 135.740 ;
        RECT 55.380 135.680 55.700 135.740 ;
        RECT 49.490 135.540 55.700 135.680 ;
        RECT 36.995 135.495 37.285 135.540 ;
        RECT 45.735 135.495 46.025 135.540 ;
        RECT 46.195 135.495 46.485 135.540 ;
        RECT 48.940 135.480 49.260 135.540 ;
        RECT 50.320 135.480 50.640 135.540 ;
        RECT 52.160 135.480 52.480 135.540 ;
        RECT 55.380 135.480 55.700 135.540 ;
        RECT 22.275 135.340 22.565 135.385 ;
        RECT 21.800 135.200 22.565 135.340 ;
        RECT 21.800 135.140 22.120 135.200 ;
        RECT 22.275 135.155 22.565 135.200 ;
        RECT 28.240 135.140 28.560 135.400 ;
        RECT 30.540 135.340 30.860 135.400 ;
        RECT 32.380 135.340 32.700 135.400 ;
        RECT 30.540 135.200 32.700 135.340 ;
        RECT 30.540 135.140 30.860 135.200 ;
        RECT 32.380 135.140 32.700 135.200 ;
        RECT 34.220 135.340 34.540 135.400 ;
        RECT 34.695 135.340 34.985 135.385 ;
        RECT 34.220 135.200 34.985 135.340 ;
        RECT 34.220 135.140 34.540 135.200 ;
        RECT 34.695 135.155 34.985 135.200 ;
        RECT 37.455 135.340 37.745 135.385 ;
        RECT 38.360 135.340 38.680 135.400 ;
        RECT 37.455 135.200 38.680 135.340 ;
        RECT 37.455 135.155 37.745 135.200 ;
        RECT 38.360 135.140 38.680 135.200 ;
        RECT 43.435 135.340 43.725 135.385 ;
        RECT 51.700 135.340 52.020 135.400 ;
        RECT 43.435 135.200 52.020 135.340 ;
        RECT 43.435 135.155 43.725 135.200 ;
        RECT 51.700 135.140 52.020 135.200 ;
        RECT 54.475 135.340 54.765 135.385 ;
        RECT 56.300 135.340 56.620 135.400 ;
        RECT 56.850 135.385 56.990 135.880 ;
        RECT 57.695 135.835 57.985 135.880 ;
        RECT 62.295 135.835 62.585 136.065 ;
        RECT 62.755 135.835 63.045 136.065 ;
        RECT 63.215 135.835 63.505 136.065 ;
        RECT 60.440 135.680 60.760 135.740 ;
        RECT 63.290 135.680 63.430 135.835 ;
        RECT 60.440 135.540 63.430 135.680 ;
        RECT 63.750 135.680 63.890 136.220 ;
        RECT 65.055 136.220 65.820 136.360 ;
        RECT 65.055 136.175 65.345 136.220 ;
        RECT 65.500 136.160 65.820 136.220 ;
        RECT 69.730 136.220 74.100 136.360 ;
        RECT 64.120 135.820 64.440 136.080 ;
        RECT 67.815 136.020 68.105 136.065 ;
        RECT 68.275 136.020 68.565 136.065 ;
        RECT 67.815 135.880 68.565 136.020 ;
        RECT 67.815 135.835 68.105 135.880 ;
        RECT 68.275 135.835 68.565 135.880 ;
        RECT 69.180 135.820 69.500 136.080 ;
        RECT 69.730 136.065 69.870 136.220 ;
        RECT 73.780 136.160 74.100 136.220 ;
        RECT 69.655 135.835 69.945 136.065 ;
        RECT 70.115 135.835 70.405 136.065 ;
        RECT 76.080 136.020 76.400 136.080 ;
        RECT 77.935 136.020 78.225 136.065 ;
        RECT 76.080 135.880 78.225 136.020 ;
        RECT 65.040 135.680 65.360 135.740 ;
        RECT 66.420 135.680 66.740 135.740 ;
        RECT 70.190 135.680 70.330 135.835 ;
        RECT 76.080 135.820 76.400 135.880 ;
        RECT 77.935 135.835 78.225 135.880 ;
        RECT 78.395 135.835 78.685 136.065 ;
        RECT 63.750 135.540 66.740 135.680 ;
        RECT 60.440 135.480 60.760 135.540 ;
        RECT 65.040 135.480 65.360 135.540 ;
        RECT 66.420 135.480 66.740 135.540 ;
        RECT 69.730 135.540 70.330 135.680 ;
        RECT 78.470 135.680 78.610 135.835 ;
        RECT 79.300 135.820 79.620 136.080 ;
        RECT 81.140 135.820 81.460 136.080 ;
        RECT 81.690 136.065 81.830 136.560 ;
        RECT 82.060 136.500 82.380 136.560 ;
        RECT 86.660 136.500 86.980 136.560 ;
        RECT 87.550 136.700 87.840 136.745 ;
        RECT 90.330 136.700 90.620 136.745 ;
        RECT 92.190 136.700 92.480 136.745 ;
        RECT 87.550 136.560 92.480 136.700 ;
        RECT 95.490 136.700 95.630 136.900 ;
        RECT 105.060 136.900 107.205 137.040 ;
        RECT 105.060 136.840 105.380 136.900 ;
        RECT 106.915 136.855 107.205 136.900 ;
        RECT 119.320 137.040 119.640 137.100 ;
        RECT 119.320 136.900 123.230 137.040 ;
        RECT 119.320 136.840 119.640 136.900 ;
        RECT 112.880 136.700 113.200 136.760 ;
        RECT 95.490 136.560 96.090 136.700 ;
        RECT 87.550 136.515 87.840 136.560 ;
        RECT 90.330 136.515 90.620 136.560 ;
        RECT 92.190 136.515 92.480 136.560 ;
        RECT 86.200 136.360 86.520 136.420 ;
        RECT 82.150 136.220 86.520 136.360 ;
        RECT 82.150 136.065 82.290 136.220 ;
        RECT 86.200 136.160 86.520 136.220 ;
        RECT 90.800 136.160 91.120 136.420 ;
        RECT 91.260 136.360 91.580 136.420 ;
        RECT 95.950 136.405 96.090 136.560 ;
        RECT 103.310 136.560 113.200 136.700 ;
        RECT 103.310 136.405 103.450 136.560 ;
        RECT 109.750 136.405 109.890 136.560 ;
        RECT 112.880 136.500 113.200 136.560 ;
        RECT 117.450 136.700 117.740 136.745 ;
        RECT 120.230 136.700 120.520 136.745 ;
        RECT 122.090 136.700 122.380 136.745 ;
        RECT 117.450 136.560 122.380 136.700 ;
        RECT 117.450 136.515 117.740 136.560 ;
        RECT 120.230 136.515 120.520 136.560 ;
        RECT 122.090 136.515 122.380 136.560 ;
        RECT 95.415 136.360 95.705 136.405 ;
        RECT 91.260 136.220 95.705 136.360 ;
        RECT 91.260 136.160 91.580 136.220 ;
        RECT 95.415 136.175 95.705 136.220 ;
        RECT 95.875 136.360 96.165 136.405 ;
        RECT 103.235 136.360 103.525 136.405 ;
        RECT 95.875 136.220 103.525 136.360 ;
        RECT 95.875 136.175 96.165 136.220 ;
        RECT 103.235 136.175 103.525 136.220 ;
        RECT 104.690 136.220 108.970 136.360 ;
        RECT 81.615 135.835 81.905 136.065 ;
        RECT 82.075 135.835 82.365 136.065 ;
        RECT 82.980 135.820 83.300 136.080 ;
        RECT 87.550 136.020 87.840 136.065 ;
        RECT 87.550 135.880 90.085 136.020 ;
        RECT 87.550 135.835 87.840 135.880 ;
        RECT 83.900 135.680 84.220 135.740 ;
        RECT 78.470 135.540 84.220 135.680 ;
        RECT 54.475 135.200 56.620 135.340 ;
        RECT 54.475 135.155 54.765 135.200 ;
        RECT 56.300 135.140 56.620 135.200 ;
        RECT 56.775 135.155 57.065 135.385 ;
        RECT 58.615 135.340 58.905 135.385 ;
        RECT 59.520 135.340 59.840 135.400 ;
        RECT 58.615 135.200 59.840 135.340 ;
        RECT 58.615 135.155 58.905 135.200 ;
        RECT 59.520 135.140 59.840 135.200 ;
        RECT 60.900 135.340 61.220 135.400 ;
        RECT 69.730 135.340 69.870 135.540 ;
        RECT 83.900 135.480 84.220 135.540 ;
        RECT 85.690 135.680 85.980 135.725 ;
        RECT 88.040 135.680 88.360 135.740 ;
        RECT 89.870 135.725 90.085 135.880 ;
        RECT 92.655 135.835 92.945 136.065 ;
        RECT 93.100 136.020 93.420 136.080 ;
        RECT 97.700 136.020 98.020 136.080 ;
        RECT 93.100 135.880 98.020 136.020 ;
        RECT 88.950 135.680 89.240 135.725 ;
        RECT 85.690 135.540 89.240 135.680 ;
        RECT 85.690 135.495 85.980 135.540 ;
        RECT 88.040 135.480 88.360 135.540 ;
        RECT 88.950 135.495 89.240 135.540 ;
        RECT 89.870 135.680 90.160 135.725 ;
        RECT 91.730 135.680 92.020 135.725 ;
        RECT 89.870 135.540 92.020 135.680 ;
        RECT 92.730 135.680 92.870 135.835 ;
        RECT 93.100 135.820 93.420 135.880 ;
        RECT 97.700 135.820 98.020 135.880 ;
        RECT 98.620 135.820 98.940 136.080 ;
        RECT 99.080 135.820 99.400 136.080 ;
        RECT 99.555 136.020 99.845 136.065 ;
        RECT 100.000 136.020 100.320 136.080 ;
        RECT 104.690 136.065 104.830 136.220 ;
        RECT 104.155 136.020 104.445 136.065 ;
        RECT 99.555 135.880 100.320 136.020 ;
        RECT 99.555 135.835 99.845 135.880 ;
        RECT 100.000 135.820 100.320 135.880 ;
        RECT 100.550 135.880 104.445 136.020 ;
        RECT 94.020 135.680 94.340 135.740 ;
        RECT 98.160 135.680 98.480 135.740 ;
        RECT 92.730 135.540 98.480 135.680 ;
        RECT 89.870 135.495 90.160 135.540 ;
        RECT 91.730 135.495 92.020 135.540 ;
        RECT 94.020 135.480 94.340 135.540 ;
        RECT 98.160 135.480 98.480 135.540 ;
        RECT 98.710 135.680 98.850 135.820 ;
        RECT 100.550 135.680 100.690 135.880 ;
        RECT 104.155 135.835 104.445 135.880 ;
        RECT 104.615 135.835 104.905 136.065 ;
        RECT 107.835 136.020 108.125 136.065 ;
        RECT 106.530 135.880 108.125 136.020 ;
        RECT 98.710 135.540 100.690 135.680 ;
        RECT 60.900 135.200 69.870 135.340 ;
        RECT 78.840 135.340 79.160 135.400 ;
        RECT 79.775 135.340 80.065 135.385 ;
        RECT 78.840 135.200 80.065 135.340 ;
        RECT 60.900 135.140 61.220 135.200 ;
        RECT 78.840 135.140 79.160 135.200 ;
        RECT 79.775 135.155 80.065 135.200 ;
        RECT 84.820 135.340 85.140 135.400 ;
        RECT 92.640 135.340 92.960 135.400 ;
        RECT 84.820 135.200 92.960 135.340 ;
        RECT 84.820 135.140 85.140 135.200 ;
        RECT 92.640 135.140 92.960 135.200 ;
        RECT 93.115 135.340 93.405 135.385 ;
        RECT 93.560 135.340 93.880 135.400 ;
        RECT 93.115 135.200 93.880 135.340 ;
        RECT 93.115 135.155 93.405 135.200 ;
        RECT 93.560 135.140 93.880 135.200 ;
        RECT 94.955 135.340 95.245 135.385 ;
        RECT 98.710 135.340 98.850 135.540 ;
        RECT 94.955 135.200 98.850 135.340 ;
        RECT 94.955 135.155 95.245 135.200 ;
        RECT 100.920 135.140 101.240 135.400 ;
        RECT 106.530 135.385 106.670 135.880 ;
        RECT 107.835 135.835 108.125 135.880 ;
        RECT 108.830 135.740 108.970 136.220 ;
        RECT 109.675 136.175 109.965 136.405 ;
        RECT 121.160 136.360 121.480 136.420 ;
        RECT 122.555 136.360 122.845 136.405 ;
        RECT 121.160 136.220 122.845 136.360 ;
        RECT 121.160 136.160 121.480 136.220 ;
        RECT 122.555 136.175 122.845 136.220 ;
        RECT 111.055 136.020 111.345 136.065 ;
        RECT 112.420 136.020 112.740 136.080 ;
        RECT 111.055 135.880 112.740 136.020 ;
        RECT 111.055 135.835 111.345 135.880 ;
        RECT 112.420 135.820 112.740 135.880 ;
        RECT 117.450 136.020 117.740 136.065 ;
        RECT 117.450 135.880 119.985 136.020 ;
        RECT 117.450 135.835 117.740 135.880 ;
        RECT 108.740 135.680 109.060 135.740 ;
        RECT 115.640 135.725 115.960 135.740 ;
        RECT 119.770 135.725 119.985 135.880 ;
        RECT 120.700 135.820 121.020 136.080 ;
        RECT 123.090 136.065 123.230 136.900 ;
        RECT 123.920 136.840 124.240 137.100 ;
        RECT 123.015 135.835 123.305 136.065 ;
        RECT 110.595 135.680 110.885 135.725 ;
        RECT 113.585 135.680 113.875 135.725 ;
        RECT 108.740 135.540 113.875 135.680 ;
        RECT 108.740 135.480 109.060 135.540 ;
        RECT 110.595 135.495 110.885 135.540 ;
        RECT 113.585 135.495 113.875 135.540 ;
        RECT 115.590 135.680 115.960 135.725 ;
        RECT 118.850 135.680 119.140 135.725 ;
        RECT 115.590 135.540 119.140 135.680 ;
        RECT 115.590 135.495 115.960 135.540 ;
        RECT 118.850 135.495 119.140 135.540 ;
        RECT 119.770 135.680 120.060 135.725 ;
        RECT 121.630 135.680 121.920 135.725 ;
        RECT 119.770 135.540 121.920 135.680 ;
        RECT 119.770 135.495 120.060 135.540 ;
        RECT 121.630 135.495 121.920 135.540 ;
        RECT 115.640 135.480 115.960 135.495 ;
        RECT 106.455 135.155 106.745 135.385 ;
        RECT 112.880 135.140 113.200 135.400 ;
        RECT 14.370 134.520 127.530 135.000 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 19.040 134.120 19.360 134.380 ;
        RECT 20.665 134.320 20.955 134.365 ;
        RECT 21.800 134.320 22.120 134.380 ;
        RECT 20.665 134.180 22.120 134.320 ;
        RECT 20.665 134.135 20.955 134.180 ;
        RECT 21.800 134.120 22.120 134.180 ;
        RECT 32.395 134.320 32.685 134.365 ;
        RECT 33.760 134.320 34.080 134.380 ;
        RECT 32.395 134.180 34.080 134.320 ;
        RECT 32.395 134.135 32.685 134.180 ;
        RECT 33.760 134.120 34.080 134.180 ;
        RECT 50.320 134.120 50.640 134.380 ;
        RECT 52.405 134.320 52.695 134.365 ;
        RECT 56.300 134.320 56.620 134.380 ;
        RECT 50.870 134.180 56.620 134.320 ;
        RECT 16.755 133.980 17.045 134.025 ;
        RECT 19.130 133.980 19.270 134.120 ;
        RECT 16.755 133.840 19.270 133.980 ;
        RECT 19.515 133.980 19.805 134.025 ;
        RECT 22.670 133.980 22.960 134.025 ;
        RECT 25.930 133.980 26.220 134.025 ;
        RECT 19.515 133.840 26.220 133.980 ;
        RECT 16.755 133.795 17.045 133.840 ;
        RECT 19.515 133.795 19.805 133.840 ;
        RECT 22.670 133.795 22.960 133.840 ;
        RECT 25.930 133.795 26.220 133.840 ;
        RECT 26.850 133.980 27.140 134.025 ;
        RECT 28.710 133.980 29.000 134.025 ;
        RECT 36.060 133.980 36.380 134.040 ;
        RECT 26.850 133.840 29.000 133.980 ;
        RECT 26.850 133.795 27.140 133.840 ;
        RECT 28.710 133.795 29.000 133.840 ;
        RECT 29.710 133.840 36.380 133.980 ;
        RECT 17.215 133.455 17.505 133.685 ;
        RECT 17.675 133.640 17.965 133.685 ;
        RECT 18.580 133.640 18.900 133.700 ;
        RECT 17.675 133.500 18.900 133.640 ;
        RECT 17.675 133.455 17.965 133.500 ;
        RECT 17.290 133.300 17.430 133.455 ;
        RECT 18.580 133.440 18.900 133.500 ;
        RECT 19.055 133.640 19.345 133.685 ;
        RECT 24.530 133.640 24.820 133.685 ;
        RECT 26.850 133.640 27.065 133.795 ;
        RECT 29.710 133.700 29.850 133.840 ;
        RECT 36.060 133.780 36.380 133.840 ;
        RECT 42.055 133.980 42.345 134.025 ;
        RECT 48.495 133.980 48.785 134.025 ;
        RECT 50.410 133.980 50.550 134.120 ;
        RECT 42.055 133.840 48.785 133.980 ;
        RECT 42.055 133.795 42.345 133.840 ;
        RECT 48.495 133.795 48.785 133.840 ;
        RECT 49.490 133.840 50.550 133.980 ;
        RECT 19.055 133.500 19.730 133.640 ;
        RECT 19.055 133.455 19.345 133.500 ;
        RECT 19.590 133.360 19.730 133.500 ;
        RECT 24.530 133.500 27.065 133.640 ;
        RECT 27.410 133.500 29.390 133.640 ;
        RECT 24.530 133.455 24.820 133.500 ;
        RECT 19.500 133.300 19.820 133.360 ;
        RECT 17.290 133.160 19.820 133.300 ;
        RECT 19.500 133.100 19.820 133.160 ;
        RECT 21.800 133.300 22.120 133.360 ;
        RECT 27.410 133.300 27.550 133.500 ;
        RECT 21.800 133.160 27.550 133.300 ;
        RECT 27.795 133.300 28.085 133.345 ;
        RECT 28.700 133.300 29.020 133.360 ;
        RECT 27.795 133.160 29.020 133.300 ;
        RECT 29.250 133.300 29.390 133.500 ;
        RECT 29.620 133.440 29.940 133.700 ;
        RECT 31.000 133.640 31.320 133.700 ;
        RECT 30.170 133.500 31.320 133.640 ;
        RECT 30.170 133.300 30.310 133.500 ;
        RECT 31.000 133.440 31.320 133.500 ;
        RECT 31.475 133.640 31.765 133.685 ;
        RECT 31.920 133.640 32.240 133.700 ;
        RECT 31.475 133.500 32.240 133.640 ;
        RECT 31.475 133.455 31.765 133.500 ;
        RECT 31.920 133.440 32.240 133.500 ;
        RECT 32.380 133.640 32.700 133.700 ;
        RECT 34.695 133.640 34.985 133.685 ;
        RECT 32.380 133.500 34.985 133.640 ;
        RECT 32.380 133.440 32.700 133.500 ;
        RECT 34.695 133.455 34.985 133.500 ;
        RECT 39.295 133.455 39.585 133.685 ;
        RECT 29.250 133.160 30.310 133.300 ;
        RECT 21.800 133.100 22.120 133.160 ;
        RECT 27.795 133.115 28.085 133.160 ;
        RECT 28.700 133.100 29.020 133.160 ;
        RECT 30.555 133.115 30.845 133.345 ;
        RECT 31.090 133.300 31.230 133.440 ;
        RECT 33.315 133.300 33.605 133.345 ;
        RECT 31.090 133.160 33.605 133.300 ;
        RECT 33.315 133.115 33.605 133.160 ;
        RECT 34.235 133.115 34.525 133.345 ;
        RECT 39.370 133.300 39.510 133.455 ;
        RECT 40.200 133.440 40.520 133.700 ;
        RECT 40.660 133.440 40.980 133.700 ;
        RECT 42.500 133.640 42.820 133.700 ;
        RECT 42.975 133.640 43.265 133.685 ;
        RECT 42.500 133.500 43.265 133.640 ;
        RECT 42.500 133.440 42.820 133.500 ;
        RECT 42.975 133.455 43.265 133.500 ;
        RECT 43.420 133.440 43.740 133.700 ;
        RECT 46.180 133.440 46.500 133.700 ;
        RECT 46.655 133.455 46.945 133.685 ;
        RECT 47.115 133.455 47.405 133.685 ;
        RECT 48.035 133.640 48.325 133.685 ;
        RECT 49.490 133.640 49.630 133.840 ;
        RECT 48.035 133.500 49.630 133.640 ;
        RECT 48.035 133.455 48.325 133.500 ;
        RECT 44.815 133.300 45.105 133.345 ;
        RECT 39.370 133.160 45.105 133.300 ;
        RECT 44.815 133.115 45.105 133.160 ;
        RECT 18.595 132.960 18.885 133.005 ;
        RECT 23.180 132.960 23.500 133.020 ;
        RECT 18.595 132.820 23.500 132.960 ;
        RECT 18.595 132.775 18.885 132.820 ;
        RECT 23.180 132.760 23.500 132.820 ;
        RECT 24.530 132.960 24.820 133.005 ;
        RECT 27.310 132.960 27.600 133.005 ;
        RECT 29.170 132.960 29.460 133.005 ;
        RECT 24.530 132.820 29.460 132.960 ;
        RECT 30.630 132.960 30.770 133.115 ;
        RECT 34.310 132.960 34.450 133.115 ;
        RECT 34.680 132.960 35.000 133.020 ;
        RECT 30.630 132.820 35.000 132.960 ;
        RECT 24.530 132.775 24.820 132.820 ;
        RECT 27.310 132.775 27.600 132.820 ;
        RECT 29.170 132.775 29.460 132.820 ;
        RECT 34.680 132.760 35.000 132.820 ;
        RECT 31.000 132.620 31.320 132.680 ;
        RECT 35.600 132.620 35.920 132.680 ;
        RECT 31.000 132.480 35.920 132.620 ;
        RECT 31.000 132.420 31.320 132.480 ;
        RECT 35.600 132.420 35.920 132.480 ;
        RECT 36.535 132.620 36.825 132.665 ;
        RECT 39.280 132.620 39.600 132.680 ;
        RECT 36.535 132.480 39.600 132.620 ;
        RECT 36.535 132.435 36.825 132.480 ;
        RECT 39.280 132.420 39.600 132.480 ;
        RECT 40.200 132.420 40.520 132.680 ;
        RECT 41.120 132.620 41.440 132.680 ;
        RECT 41.595 132.620 41.885 132.665 ;
        RECT 41.120 132.480 41.885 132.620 ;
        RECT 41.120 132.420 41.440 132.480 ;
        RECT 41.595 132.435 41.885 132.480 ;
        RECT 42.960 132.420 43.280 132.680 ;
        RECT 43.880 132.620 44.200 132.680 ;
        RECT 44.355 132.620 44.645 132.665 ;
        RECT 43.880 132.480 44.645 132.620 ;
        RECT 46.730 132.620 46.870 133.455 ;
        RECT 47.190 132.960 47.330 133.455 ;
        RECT 49.860 133.440 50.180 133.700 ;
        RECT 50.320 133.440 50.640 133.700 ;
        RECT 50.870 133.685 51.010 134.180 ;
        RECT 52.405 134.135 52.695 134.180 ;
        RECT 56.300 134.120 56.620 134.180 ;
        RECT 74.240 134.320 74.560 134.380 ;
        RECT 87.595 134.320 87.885 134.365 ;
        RECT 88.040 134.320 88.360 134.380 ;
        RECT 100.000 134.320 100.320 134.380 ;
        RECT 101.855 134.320 102.145 134.365 ;
        RECT 102.300 134.320 102.620 134.380 ;
        RECT 74.240 134.180 87.350 134.320 ;
        RECT 74.240 134.120 74.560 134.180 ;
        RECT 54.410 133.980 54.700 134.025 ;
        RECT 55.840 133.980 56.160 134.040 ;
        RECT 57.670 133.980 57.960 134.025 ;
        RECT 54.410 133.840 57.960 133.980 ;
        RECT 54.410 133.795 54.700 133.840 ;
        RECT 55.840 133.780 56.160 133.840 ;
        RECT 57.670 133.795 57.960 133.840 ;
        RECT 58.590 133.980 58.880 134.025 ;
        RECT 60.450 133.980 60.740 134.025 ;
        RECT 58.590 133.840 60.740 133.980 ;
        RECT 58.590 133.795 58.880 133.840 ;
        RECT 60.450 133.795 60.740 133.840 ;
        RECT 64.120 133.980 64.440 134.040 ;
        RECT 64.120 133.840 66.650 133.980 ;
        RECT 50.795 133.455 51.085 133.685 ;
        RECT 51.715 133.640 52.005 133.685 ;
        RECT 52.160 133.640 52.480 133.700 ;
        RECT 51.715 133.500 52.480 133.640 ;
        RECT 51.715 133.455 52.005 133.500 ;
        RECT 52.160 133.440 52.480 133.500 ;
        RECT 56.270 133.640 56.560 133.685 ;
        RECT 58.590 133.640 58.805 133.795 ;
        RECT 64.120 133.780 64.440 133.840 ;
        RECT 56.270 133.500 58.805 133.640 ;
        RECT 56.270 133.455 56.560 133.500 ;
        RECT 59.520 133.440 59.840 133.700 ;
        RECT 61.375 133.640 61.665 133.685 ;
        RECT 63.660 133.640 63.980 133.700 ;
        RECT 61.375 133.500 63.980 133.640 ;
        RECT 61.375 133.455 61.665 133.500 ;
        RECT 63.660 133.440 63.980 133.500 ;
        RECT 64.580 133.440 64.900 133.700 ;
        RECT 65.040 133.440 65.360 133.700 ;
        RECT 65.500 133.440 65.820 133.700 ;
        RECT 66.510 133.685 66.650 133.840 ;
        RECT 78.840 133.780 79.160 134.040 ;
        RECT 84.820 133.980 85.140 134.040 ;
        RECT 79.850 133.840 85.140 133.980 ;
        RECT 87.210 133.980 87.350 134.180 ;
        RECT 87.595 134.180 88.360 134.320 ;
        RECT 87.595 134.135 87.885 134.180 ;
        RECT 88.040 134.120 88.360 134.180 ;
        RECT 89.970 134.180 101.610 134.320 ;
        RECT 89.970 133.980 90.110 134.180 ;
        RECT 100.000 134.120 100.320 134.180 ;
        RECT 87.210 133.840 90.110 133.980 ;
        RECT 90.340 133.980 90.660 134.040 ;
        RECT 91.210 133.980 91.500 134.025 ;
        RECT 94.470 133.980 94.760 134.025 ;
        RECT 90.340 133.840 94.760 133.980 ;
        RECT 66.435 133.640 66.725 133.685 ;
        RECT 79.850 133.640 79.990 133.840 ;
        RECT 84.820 133.780 85.140 133.840 ;
        RECT 90.340 133.780 90.660 133.840 ;
        RECT 91.210 133.795 91.500 133.840 ;
        RECT 94.470 133.795 94.760 133.840 ;
        RECT 95.390 133.980 95.680 134.025 ;
        RECT 97.250 133.980 97.540 134.025 ;
        RECT 95.390 133.840 97.540 133.980 ;
        RECT 95.390 133.795 95.680 133.840 ;
        RECT 97.250 133.795 97.540 133.840 ;
        RECT 66.435 133.500 79.990 133.640 ;
        RECT 66.435 133.455 66.725 133.500 ;
        RECT 80.220 133.440 80.540 133.700 ;
        RECT 88.040 133.440 88.360 133.700 ;
        RECT 93.070 133.640 93.360 133.685 ;
        RECT 95.390 133.640 95.605 133.795 ;
        RECT 100.920 133.780 101.240 134.040 ;
        RECT 101.470 133.980 101.610 134.180 ;
        RECT 101.855 134.180 102.620 134.320 ;
        RECT 101.855 134.135 102.145 134.180 ;
        RECT 102.300 134.120 102.620 134.180 ;
        RECT 119.795 134.320 120.085 134.365 ;
        RECT 120.700 134.320 121.020 134.380 ;
        RECT 119.795 134.180 121.020 134.320 ;
        RECT 119.795 134.135 120.085 134.180 ;
        RECT 120.700 134.120 121.020 134.180 ;
        RECT 105.535 133.980 105.825 134.025 ;
        RECT 105.995 133.980 106.285 134.025 ;
        RECT 110.120 133.980 110.440 134.040 ;
        RECT 101.470 133.840 104.730 133.980 ;
        RECT 93.070 133.500 95.605 133.640 ;
        RECT 93.070 133.455 93.360 133.500 ;
        RECT 97.700 133.440 98.020 133.700 ;
        RECT 98.160 133.440 98.480 133.700 ;
        RECT 99.540 133.440 99.860 133.700 ;
        RECT 102.300 133.440 102.620 133.700 ;
        RECT 103.680 133.640 104.000 133.700 ;
        RECT 104.155 133.640 104.445 133.685 ;
        RECT 103.680 133.500 104.445 133.640 ;
        RECT 104.590 133.640 104.730 133.840 ;
        RECT 105.535 133.840 106.285 133.980 ;
        RECT 105.535 133.795 105.825 133.840 ;
        RECT 105.995 133.795 106.285 133.840 ;
        RECT 107.450 133.840 110.440 133.980 ;
        RECT 107.450 133.685 107.590 133.840 ;
        RECT 110.120 133.780 110.440 133.840 ;
        RECT 111.960 133.780 112.280 134.040 ;
        RECT 107.375 133.640 107.665 133.685 ;
        RECT 104.590 133.500 107.665 133.640 ;
        RECT 103.680 133.440 104.000 133.500 ;
        RECT 104.155 133.455 104.445 133.500 ;
        RECT 107.375 133.455 107.665 133.500 ;
        RECT 107.820 133.440 108.140 133.700 ;
        RECT 108.295 133.640 108.585 133.685 ;
        RECT 108.740 133.640 109.060 133.700 ;
        RECT 108.295 133.500 109.060 133.640 ;
        RECT 108.295 133.455 108.585 133.500 ;
        RECT 108.740 133.440 109.060 133.500 ;
        RECT 109.200 133.440 109.520 133.700 ;
        RECT 110.580 133.440 110.900 133.700 ;
        RECT 111.040 133.440 111.360 133.700 ;
        RECT 112.880 133.640 113.200 133.700 ;
        RECT 118.875 133.640 119.165 133.685 ;
        RECT 112.880 133.500 119.165 133.640 ;
        RECT 112.880 133.440 113.200 133.500 ;
        RECT 118.875 133.455 119.165 133.500 ;
        RECT 48.940 133.300 49.260 133.360 ;
        RECT 63.215 133.300 63.505 133.345 ;
        RECT 48.940 133.160 63.505 133.300 ;
        RECT 48.940 133.100 49.260 133.160 ;
        RECT 63.215 133.115 63.505 133.160 ;
        RECT 79.775 133.300 80.065 133.345 ;
        RECT 83.440 133.300 83.760 133.360 ;
        RECT 79.775 133.160 83.760 133.300 ;
        RECT 79.775 133.115 80.065 133.160 ;
        RECT 83.440 133.100 83.760 133.160 ;
        RECT 86.200 133.300 86.520 133.360 ;
        RECT 89.205 133.300 89.495 133.345 ;
        RECT 91.260 133.300 91.580 133.360 ;
        RECT 86.200 133.160 91.580 133.300 ;
        RECT 86.200 133.100 86.520 133.160 ;
        RECT 89.205 133.115 89.495 133.160 ;
        RECT 91.260 133.100 91.580 133.160 ;
        RECT 94.940 133.300 95.260 133.360 ;
        RECT 96.335 133.300 96.625 133.345 ;
        RECT 94.940 133.160 96.625 133.300 ;
        RECT 97.790 133.300 97.930 133.440 ;
        RECT 97.790 133.160 100.230 133.300 ;
        RECT 94.940 133.100 95.260 133.160 ;
        RECT 96.335 133.115 96.625 133.160 ;
        RECT 55.380 132.960 55.700 133.020 ;
        RECT 47.190 132.820 55.700 132.960 ;
        RECT 55.380 132.760 55.700 132.820 ;
        RECT 56.270 132.960 56.560 133.005 ;
        RECT 59.050 132.960 59.340 133.005 ;
        RECT 60.910 132.960 61.200 133.005 ;
        RECT 56.270 132.820 61.200 132.960 ;
        RECT 56.270 132.775 56.560 132.820 ;
        RECT 59.050 132.775 59.340 132.820 ;
        RECT 60.910 132.775 61.200 132.820 ;
        RECT 81.155 132.960 81.445 133.005 ;
        RECT 93.070 132.960 93.360 133.005 ;
        RECT 95.850 132.960 96.140 133.005 ;
        RECT 97.710 132.960 98.000 133.005 ;
        RECT 81.155 132.820 87.810 132.960 ;
        RECT 81.155 132.775 81.445 132.820 ;
        RECT 50.320 132.620 50.640 132.680 ;
        RECT 46.730 132.480 50.640 132.620 ;
        RECT 43.880 132.420 44.200 132.480 ;
        RECT 44.355 132.435 44.645 132.480 ;
        RECT 50.320 132.420 50.640 132.480 ;
        RECT 80.235 132.620 80.525 132.665 ;
        RECT 82.980 132.620 83.300 132.680 ;
        RECT 80.235 132.480 83.300 132.620 ;
        RECT 87.670 132.620 87.810 132.820 ;
        RECT 93.070 132.820 98.000 132.960 ;
        RECT 100.090 132.960 100.230 133.160 ;
        RECT 100.460 133.100 100.780 133.360 ;
        RECT 101.840 133.300 102.160 133.360 ;
        RECT 104.615 133.300 104.905 133.345 ;
        RECT 101.840 133.160 104.905 133.300 ;
        RECT 101.840 133.100 102.160 133.160 ;
        RECT 104.615 133.115 104.905 133.160 ;
        RECT 109.290 132.960 109.430 133.440 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 100.090 132.820 109.430 132.960 ;
        RECT 93.070 132.775 93.360 132.820 ;
        RECT 95.850 132.775 96.140 132.820 ;
        RECT 97.710 132.775 98.000 132.820 ;
        RECT 94.480 132.620 94.800 132.680 ;
        RECT 87.670 132.480 94.800 132.620 ;
        RECT 80.235 132.435 80.525 132.480 ;
        RECT 82.980 132.420 83.300 132.480 ;
        RECT 94.480 132.420 94.800 132.480 ;
        RECT 98.635 132.620 98.925 132.665 ;
        RECT 99.540 132.620 99.860 132.680 ;
        RECT 98.635 132.480 99.860 132.620 ;
        RECT 98.635 132.435 98.925 132.480 ;
        RECT 99.540 132.420 99.860 132.480 ;
        RECT 100.920 132.420 101.240 132.680 ;
        RECT 103.220 132.420 103.540 132.680 ;
        RECT 104.600 132.420 104.920 132.680 ;
        RECT 109.675 132.620 109.965 132.665 ;
        RECT 110.120 132.620 110.440 132.680 ;
        RECT 109.675 132.480 110.440 132.620 ;
        RECT 109.675 132.435 109.965 132.480 ;
        RECT 110.120 132.420 110.440 132.480 ;
        RECT 111.040 132.420 111.360 132.680 ;
        RECT 14.370 131.800 127.530 132.280 ;
        RECT 28.700 131.400 29.020 131.660 ;
        RECT 30.540 131.645 30.860 131.660 ;
        RECT 30.325 131.415 30.860 131.645 ;
        RECT 30.540 131.400 30.860 131.415 ;
        RECT 33.760 131.600 34.080 131.660 ;
        RECT 78.395 131.600 78.685 131.645 ;
        RECT 79.760 131.600 80.080 131.660 ;
        RECT 33.760 131.460 39.970 131.600 ;
        RECT 33.760 131.400 34.080 131.460 ;
        RECT 39.830 131.320 39.970 131.460 ;
        RECT 78.395 131.460 80.080 131.600 ;
        RECT 78.395 131.415 78.685 131.460 ;
        RECT 79.760 131.400 80.080 131.460 ;
        RECT 89.435 131.600 89.725 131.645 ;
        RECT 90.340 131.600 90.660 131.660 ;
        RECT 89.435 131.460 90.660 131.600 ;
        RECT 89.435 131.415 89.725 131.460 ;
        RECT 90.340 131.400 90.660 131.460 ;
        RECT 109.660 131.400 109.980 131.660 ;
        RECT 34.190 131.260 34.480 131.305 ;
        RECT 36.970 131.260 37.260 131.305 ;
        RECT 38.830 131.260 39.120 131.305 ;
        RECT 34.190 131.120 39.120 131.260 ;
        RECT 34.190 131.075 34.480 131.120 ;
        RECT 36.970 131.075 37.260 131.120 ;
        RECT 38.830 131.075 39.120 131.120 ;
        RECT 39.740 131.260 40.060 131.320 ;
        RECT 69.655 131.260 69.945 131.305 ;
        RECT 100.000 131.260 100.320 131.320 ;
        RECT 39.740 131.120 100.320 131.260 ;
        RECT 39.740 131.060 40.060 131.120 ;
        RECT 69.655 131.075 69.945 131.120 ;
        RECT 100.000 131.060 100.320 131.120 ;
        RECT 102.300 131.260 102.620 131.320 ;
        RECT 117.940 131.260 118.260 131.320 ;
        RECT 102.300 131.120 118.260 131.260 ;
        RECT 102.300 131.060 102.620 131.120 ;
        RECT 117.940 131.060 118.260 131.120 ;
        RECT 20.895 130.920 21.185 130.965 ;
        RECT 21.800 130.920 22.120 130.980 ;
        RECT 20.895 130.780 22.120 130.920 ;
        RECT 20.895 130.735 21.185 130.780 ;
        RECT 21.800 130.720 22.120 130.780 ;
        RECT 36.060 130.920 36.380 130.980 ;
        RECT 36.060 130.780 37.210 130.920 ;
        RECT 36.060 130.720 36.380 130.780 ;
        RECT 28.240 130.580 28.560 130.640 ;
        RECT 29.635 130.580 29.925 130.625 ;
        RECT 28.240 130.440 29.925 130.580 ;
        RECT 28.240 130.380 28.560 130.440 ;
        RECT 29.635 130.395 29.925 130.440 ;
        RECT 34.190 130.580 34.480 130.625 ;
        RECT 37.070 130.580 37.210 130.780 ;
        RECT 37.440 130.720 37.760 130.980 ;
        RECT 64.580 130.920 64.900 130.980 ;
        RECT 66.435 130.920 66.725 130.965 ;
        RECT 69.180 130.920 69.500 130.980 ;
        RECT 64.580 130.780 69.500 130.920 ;
        RECT 64.580 130.720 64.900 130.780 ;
        RECT 66.435 130.735 66.725 130.780 ;
        RECT 69.180 130.720 69.500 130.780 ;
        RECT 73.335 130.920 73.625 130.965 ;
        RECT 73.780 130.920 74.100 130.980 ;
        RECT 73.335 130.780 74.100 130.920 ;
        RECT 73.335 130.735 73.625 130.780 ;
        RECT 73.780 130.720 74.100 130.780 ;
        RECT 39.295 130.580 39.585 130.625 ;
        RECT 70.575 130.580 70.865 130.625 ;
        RECT 72.400 130.580 72.720 130.640 ;
        RECT 74.255 130.580 74.545 130.625 ;
        RECT 79.315 130.580 79.605 130.625 ;
        RECT 34.190 130.440 36.725 130.580 ;
        RECT 37.070 130.440 42.270 130.580 ;
        RECT 34.190 130.395 34.480 130.440 ;
        RECT 21.815 130.240 22.105 130.285 ;
        RECT 23.180 130.240 23.500 130.300 ;
        RECT 21.815 130.100 23.500 130.240 ;
        RECT 21.815 130.055 22.105 130.100 ;
        RECT 23.180 130.040 23.500 130.100 ;
        RECT 32.330 130.240 32.620 130.285 ;
        RECT 33.760 130.240 34.080 130.300 ;
        RECT 36.510 130.285 36.725 130.440 ;
        RECT 39.295 130.395 39.585 130.440 ;
        RECT 35.590 130.240 35.880 130.285 ;
        RECT 32.330 130.100 35.880 130.240 ;
        RECT 32.330 130.055 32.620 130.100 ;
        RECT 33.760 130.040 34.080 130.100 ;
        RECT 35.590 130.055 35.880 130.100 ;
        RECT 36.510 130.240 36.800 130.285 ;
        RECT 38.370 130.240 38.660 130.285 ;
        RECT 36.510 130.100 38.660 130.240 ;
        RECT 36.510 130.055 36.800 130.100 ;
        RECT 38.370 130.055 38.660 130.100 ;
        RECT 21.355 129.900 21.645 129.945 ;
        RECT 22.260 129.900 22.580 129.960 ;
        RECT 21.355 129.760 22.580 129.900 ;
        RECT 21.355 129.715 21.645 129.760 ;
        RECT 22.260 129.700 22.580 129.760 ;
        RECT 22.720 129.900 23.040 129.960 ;
        RECT 42.130 129.945 42.270 130.440 ;
        RECT 70.575 130.440 74.545 130.580 ;
        RECT 70.575 130.395 70.865 130.440 ;
        RECT 72.400 130.380 72.720 130.440 ;
        RECT 74.255 130.395 74.545 130.440 ;
        RECT 74.790 130.440 79.605 130.580 ;
        RECT 48.495 130.240 48.785 130.285 ;
        RECT 48.940 130.240 49.260 130.300 ;
        RECT 48.495 130.100 49.260 130.240 ;
        RECT 48.495 130.055 48.785 130.100 ;
        RECT 48.940 130.040 49.260 130.100 ;
        RECT 64.120 130.240 64.440 130.300 ;
        RECT 65.500 130.240 65.820 130.300 ;
        RECT 67.355 130.240 67.645 130.285 ;
        RECT 64.120 130.100 67.645 130.240 ;
        RECT 64.120 130.040 64.440 130.100 ;
        RECT 65.500 130.040 65.820 130.100 ;
        RECT 67.355 130.055 67.645 130.100 ;
        RECT 67.800 130.240 68.120 130.300 ;
        RECT 74.790 130.240 74.930 130.440 ;
        RECT 79.315 130.395 79.605 130.440 ;
        RECT 79.760 130.380 80.080 130.640 ;
        RECT 88.040 130.580 88.360 130.640 ;
        RECT 88.975 130.580 89.265 130.625 ;
        RECT 90.800 130.580 91.120 130.640 ;
        RECT 88.040 130.440 91.120 130.580 ;
        RECT 88.040 130.380 88.360 130.440 ;
        RECT 88.975 130.395 89.265 130.440 ;
        RECT 90.800 130.380 91.120 130.440 ;
        RECT 98.160 130.580 98.480 130.640 ;
        RECT 100.015 130.580 100.305 130.625 ;
        RECT 98.160 130.440 100.305 130.580 ;
        RECT 98.160 130.380 98.480 130.440 ;
        RECT 100.015 130.395 100.305 130.440 ;
        RECT 110.580 130.380 110.900 130.640 ;
        RECT 111.515 130.580 111.805 130.625 ;
        RECT 111.960 130.580 112.280 130.640 ;
        RECT 111.515 130.440 112.280 130.580 ;
        RECT 111.515 130.395 111.805 130.440 ;
        RECT 111.960 130.380 112.280 130.440 ;
        RECT 67.800 130.100 74.930 130.240 ;
        RECT 67.800 130.040 68.120 130.100 ;
        RECT 74.790 129.960 74.930 130.100 ;
        RECT 23.655 129.900 23.945 129.945 ;
        RECT 22.720 129.760 23.945 129.900 ;
        RECT 22.720 129.700 23.040 129.760 ;
        RECT 23.655 129.715 23.945 129.760 ;
        RECT 42.055 129.900 42.345 129.945 ;
        RECT 42.500 129.900 42.820 129.960 ;
        RECT 42.055 129.760 42.820 129.900 ;
        RECT 42.055 129.715 42.345 129.760 ;
        RECT 42.500 129.700 42.820 129.760 ;
        RECT 65.960 129.900 66.280 129.960 ;
        RECT 66.895 129.900 67.185 129.945 ;
        RECT 65.960 129.760 67.185 129.900 ;
        RECT 65.960 129.700 66.280 129.760 ;
        RECT 66.895 129.715 67.185 129.760 ;
        RECT 69.195 129.900 69.485 129.945 ;
        RECT 70.100 129.900 70.420 129.960 ;
        RECT 69.195 129.760 70.420 129.900 ;
        RECT 69.195 129.715 69.485 129.760 ;
        RECT 70.100 129.700 70.420 129.760 ;
        RECT 71.480 129.700 71.800 129.960 ;
        RECT 74.700 129.700 75.020 129.960 ;
        RECT 14.370 129.080 127.530 129.560 ;
        RECT 17.445 128.880 17.735 128.925 ;
        RECT 23.180 128.880 23.500 128.940 ;
        RECT 17.445 128.740 27.550 128.880 ;
        RECT 17.445 128.695 17.735 128.740 ;
        RECT 23.180 128.680 23.500 128.740 ;
        RECT 19.450 128.540 19.740 128.585 ;
        RECT 20.880 128.540 21.200 128.600 ;
        RECT 22.710 128.540 23.000 128.585 ;
        RECT 19.450 128.400 23.000 128.540 ;
        RECT 19.450 128.355 19.740 128.400 ;
        RECT 20.880 128.340 21.200 128.400 ;
        RECT 22.710 128.355 23.000 128.400 ;
        RECT 23.630 128.540 23.920 128.585 ;
        RECT 25.490 128.540 25.780 128.585 ;
        RECT 23.630 128.400 25.780 128.540 ;
        RECT 27.410 128.540 27.550 128.740 ;
        RECT 33.760 128.680 34.080 128.940 ;
        RECT 37.440 128.880 37.760 128.940 ;
        RECT 38.375 128.880 38.665 128.925 ;
        RECT 37.440 128.740 38.665 128.880 ;
        RECT 37.440 128.680 37.760 128.740 ;
        RECT 38.375 128.695 38.665 128.740 ;
        RECT 41.595 128.880 41.885 128.925 ;
        RECT 43.420 128.880 43.740 128.940 ;
        RECT 41.595 128.740 43.740 128.880 ;
        RECT 41.595 128.695 41.885 128.740 ;
        RECT 43.420 128.680 43.740 128.740 ;
        RECT 43.895 128.880 44.185 128.925 ;
        RECT 44.800 128.880 45.120 128.940 ;
        RECT 43.895 128.740 45.120 128.880 ;
        RECT 43.895 128.695 44.185 128.740 ;
        RECT 44.800 128.680 45.120 128.740 ;
        RECT 48.955 128.880 49.245 128.925 ;
        RECT 49.400 128.880 49.720 128.940 ;
        RECT 48.955 128.740 49.720 128.880 ;
        RECT 48.955 128.695 49.245 128.740 ;
        RECT 49.400 128.680 49.720 128.740 ;
        RECT 55.380 128.880 55.700 128.940 ;
        RECT 55.855 128.880 56.145 128.925 ;
        RECT 55.380 128.740 56.145 128.880 ;
        RECT 55.380 128.680 55.700 128.740 ;
        RECT 55.855 128.695 56.145 128.740 ;
        RECT 56.300 128.680 56.620 128.940 ;
        RECT 64.825 128.880 65.115 128.925 ;
        RECT 65.960 128.880 66.280 128.940 ;
        RECT 64.825 128.740 66.280 128.880 ;
        RECT 64.825 128.695 65.115 128.740 ;
        RECT 65.960 128.680 66.280 128.740 ;
        RECT 77.550 128.740 81.370 128.880 ;
        RECT 42.500 128.540 42.820 128.600 ;
        RECT 46.655 128.540 46.945 128.585 ;
        RECT 63.660 128.540 63.980 128.600 ;
        RECT 27.410 128.400 39.970 128.540 ;
        RECT 23.630 128.355 23.920 128.400 ;
        RECT 25.490 128.355 25.780 128.400 ;
        RECT 21.310 128.200 21.600 128.245 ;
        RECT 23.630 128.200 23.845 128.355 ;
        RECT 21.310 128.060 23.845 128.200 ;
        RECT 26.415 128.200 26.705 128.245 ;
        RECT 29.620 128.200 29.940 128.260 ;
        RECT 26.415 128.060 29.940 128.200 ;
        RECT 21.310 128.015 21.600 128.060 ;
        RECT 26.415 128.015 26.705 128.060 ;
        RECT 29.620 128.000 29.940 128.060 ;
        RECT 30.080 128.200 30.400 128.260 ;
        RECT 33.315 128.200 33.605 128.245 ;
        RECT 30.080 128.060 33.605 128.200 ;
        RECT 30.080 128.000 30.400 128.060 ;
        RECT 33.315 128.015 33.605 128.060 ;
        RECT 39.280 128.000 39.600 128.260 ;
        RECT 39.830 128.245 39.970 128.400 ;
        RECT 42.500 128.400 63.980 128.540 ;
        RECT 42.500 128.340 42.820 128.400 ;
        RECT 46.655 128.355 46.945 128.400 ;
        RECT 63.660 128.340 63.980 128.400 ;
        RECT 66.830 128.540 67.120 128.585 ;
        RECT 68.260 128.540 68.580 128.600 ;
        RECT 70.090 128.540 70.380 128.585 ;
        RECT 66.830 128.400 70.380 128.540 ;
        RECT 66.830 128.355 67.120 128.400 ;
        RECT 68.260 128.340 68.580 128.400 ;
        RECT 70.090 128.355 70.380 128.400 ;
        RECT 71.010 128.540 71.300 128.585 ;
        RECT 72.870 128.540 73.160 128.585 ;
        RECT 71.010 128.400 73.160 128.540 ;
        RECT 71.010 128.355 71.300 128.400 ;
        RECT 72.870 128.355 73.160 128.400 ;
        RECT 39.755 128.015 40.045 128.245 ;
        RECT 40.675 128.200 40.965 128.245 ;
        RECT 42.975 128.200 43.265 128.245 ;
        RECT 45.720 128.200 46.040 128.260 ;
        RECT 48.035 128.200 48.325 128.245 ;
        RECT 67.800 128.200 68.120 128.260 ;
        RECT 40.675 128.060 68.120 128.200 ;
        RECT 40.675 128.015 40.965 128.060 ;
        RECT 42.975 128.015 43.265 128.060 ;
        RECT 45.720 128.000 46.040 128.060 ;
        RECT 48.035 128.015 48.325 128.060 ;
        RECT 67.800 128.000 68.120 128.060 ;
        RECT 68.690 128.200 68.980 128.245 ;
        RECT 71.010 128.200 71.225 128.355 ;
        RECT 68.690 128.060 71.225 128.200 ;
        RECT 68.690 128.015 68.980 128.060 ;
        RECT 71.940 128.000 72.260 128.260 ;
        RECT 74.700 128.200 75.020 128.260 ;
        RECT 77.550 128.245 77.690 128.740 ;
        RECT 78.395 128.540 78.685 128.585 ;
        RECT 80.220 128.540 80.540 128.600 ;
        RECT 78.395 128.400 80.540 128.540 ;
        RECT 81.230 128.540 81.370 128.740 ;
        RECT 82.980 128.680 83.300 128.940 ;
        RECT 88.040 128.680 88.360 128.940 ;
        RECT 89.435 128.695 89.725 128.925 ;
        RECT 81.230 128.400 84.130 128.540 ;
        RECT 78.395 128.355 78.685 128.400 ;
        RECT 80.220 128.340 80.540 128.400 ;
        RECT 83.990 128.245 84.130 128.400 ;
        RECT 84.450 128.400 85.510 128.540 ;
        RECT 75.175 128.200 75.465 128.245 ;
        RECT 77.475 128.200 77.765 128.245 ;
        RECT 80.695 128.200 80.985 128.245 ;
        RECT 74.700 128.060 77.765 128.200 ;
        RECT 74.700 128.000 75.020 128.060 ;
        RECT 75.175 128.015 75.465 128.060 ;
        RECT 77.475 128.015 77.765 128.060 ;
        RECT 78.930 128.060 80.985 128.200 ;
        RECT 23.640 127.860 23.960 127.920 ;
        RECT 24.575 127.860 24.865 127.905 ;
        RECT 23.640 127.720 24.865 127.860 ;
        RECT 23.640 127.660 23.960 127.720 ;
        RECT 24.575 127.675 24.865 127.720 ;
        RECT 42.055 127.675 42.345 127.905 ;
        RECT 42.500 127.860 42.820 127.920 ;
        RECT 47.115 127.860 47.405 127.905 ;
        RECT 42.500 127.720 47.405 127.860 ;
        RECT 21.310 127.520 21.600 127.565 ;
        RECT 24.090 127.520 24.380 127.565 ;
        RECT 25.950 127.520 26.240 127.565 ;
        RECT 21.310 127.380 26.240 127.520 ;
        RECT 21.310 127.335 21.600 127.380 ;
        RECT 24.090 127.335 24.380 127.380 ;
        RECT 25.950 127.335 26.240 127.380 ;
        RECT 22.260 127.180 22.580 127.240 ;
        RECT 42.130 127.180 42.270 127.675 ;
        RECT 42.500 127.660 42.820 127.720 ;
        RECT 47.115 127.675 47.405 127.720 ;
        RECT 54.460 127.860 54.780 127.920 ;
        RECT 54.935 127.860 55.225 127.905 ;
        RECT 54.460 127.720 55.225 127.860 ;
        RECT 54.460 127.660 54.780 127.720 ;
        RECT 54.935 127.675 55.225 127.720 ;
        RECT 63.660 127.860 63.980 127.920 ;
        RECT 73.795 127.860 74.085 127.905 ;
        RECT 63.660 127.720 74.085 127.860 ;
        RECT 63.660 127.660 63.980 127.720 ;
        RECT 73.795 127.675 74.085 127.720 ;
        RECT 74.255 127.675 74.545 127.905 ;
        RECT 76.555 127.860 76.845 127.905 ;
        RECT 78.380 127.860 78.700 127.920 ;
        RECT 78.930 127.860 79.070 128.060 ;
        RECT 80.695 128.015 80.985 128.060 ;
        RECT 83.915 128.015 84.205 128.245 ;
        RECT 76.555 127.720 79.070 127.860 ;
        RECT 76.555 127.675 76.845 127.720 ;
        RECT 68.690 127.520 68.980 127.565 ;
        RECT 71.470 127.520 71.760 127.565 ;
        RECT 73.330 127.520 73.620 127.565 ;
        RECT 68.690 127.380 73.620 127.520 ;
        RECT 74.330 127.520 74.470 127.675 ;
        RECT 78.380 127.660 78.700 127.720 ;
        RECT 79.775 127.675 80.065 127.905 ;
        RECT 78.840 127.520 79.160 127.580 ;
        RECT 74.330 127.380 79.160 127.520 ;
        RECT 79.850 127.520 79.990 127.675 ;
        RECT 80.220 127.660 80.540 127.920 ;
        RECT 80.770 127.860 80.910 128.015 ;
        RECT 84.450 127.860 84.590 128.400 ;
        RECT 84.835 128.015 85.125 128.245 ;
        RECT 80.770 127.720 84.590 127.860 ;
        RECT 84.910 127.520 85.050 128.015 ;
        RECT 85.370 127.860 85.510 128.400 ;
        RECT 87.135 128.200 87.425 128.245 ;
        RECT 89.510 128.200 89.650 128.695 ;
        RECT 94.940 128.680 95.260 128.940 ;
        RECT 98.160 128.880 98.480 128.940 ;
        RECT 101.855 128.880 102.145 128.925 ;
        RECT 98.160 128.740 102.145 128.880 ;
        RECT 98.160 128.680 98.480 128.740 ;
        RECT 101.855 128.695 102.145 128.740 ;
        RECT 104.600 128.680 104.920 128.940 ;
        RECT 105.980 128.880 106.300 128.940 ;
        RECT 106.915 128.880 107.205 128.925 ;
        RECT 105.980 128.740 107.205 128.880 ;
        RECT 105.980 128.680 106.300 128.740 ;
        RECT 106.915 128.695 107.205 128.740 ;
        RECT 111.040 128.680 111.360 128.940 ;
        RECT 95.400 128.340 95.720 128.600 ;
        RECT 105.610 128.400 108.050 128.540 ;
        RECT 87.135 128.060 89.650 128.200 ;
        RECT 91.275 128.200 91.565 128.245 ;
        RECT 93.560 128.200 93.880 128.260 ;
        RECT 94.035 128.200 94.325 128.245 ;
        RECT 91.275 128.060 93.330 128.200 ;
        RECT 87.135 128.015 87.425 128.060 ;
        RECT 91.275 128.015 91.565 128.060 ;
        RECT 91.735 127.860 92.025 127.905 ;
        RECT 85.370 127.720 92.025 127.860 ;
        RECT 91.735 127.675 92.025 127.720 ;
        RECT 92.195 127.675 92.485 127.905 ;
        RECT 93.190 127.860 93.330 128.060 ;
        RECT 93.560 128.060 94.325 128.200 ;
        RECT 93.560 128.000 93.880 128.060 ;
        RECT 94.035 128.015 94.325 128.060 ;
        RECT 100.000 128.200 100.320 128.260 ;
        RECT 105.610 128.245 105.750 128.400 ;
        RECT 105.535 128.200 105.825 128.245 ;
        RECT 100.000 128.060 105.825 128.200 ;
        RECT 100.000 128.000 100.320 128.060 ;
        RECT 105.535 128.015 105.825 128.060 ;
        RECT 105.980 128.000 106.300 128.260 ;
        RECT 107.910 128.245 108.050 128.400 ;
        RECT 107.835 128.200 108.125 128.245 ;
        RECT 110.135 128.200 110.425 128.245 ;
        RECT 110.580 128.200 110.900 128.260 ;
        RECT 112.435 128.200 112.725 128.245 ;
        RECT 107.835 128.060 112.725 128.200 ;
        RECT 107.835 128.015 108.125 128.060 ;
        RECT 110.135 128.015 110.425 128.060 ;
        RECT 110.580 128.000 110.900 128.060 ;
        RECT 112.435 128.015 112.725 128.060 ;
        RECT 112.880 128.000 113.200 128.260 ;
        RECT 117.940 128.000 118.260 128.260 ;
        RECT 119.335 128.015 119.625 128.245 ;
        RECT 98.620 127.860 98.940 127.920 ;
        RECT 105.060 127.860 105.380 127.920 ;
        RECT 108.755 127.860 109.045 127.905 ;
        RECT 93.190 127.720 109.045 127.860 ;
        RECT 91.260 127.520 91.580 127.580 ;
        RECT 79.850 127.380 84.590 127.520 ;
        RECT 84.910 127.380 91.580 127.520 ;
        RECT 68.690 127.335 68.980 127.380 ;
        RECT 71.470 127.335 71.760 127.380 ;
        RECT 73.330 127.335 73.620 127.380 ;
        RECT 78.840 127.320 79.160 127.380 ;
        RECT 84.450 127.240 84.590 127.380 ;
        RECT 91.260 127.320 91.580 127.380 ;
        RECT 22.260 127.040 42.270 127.180 ;
        RECT 57.680 127.180 58.000 127.240 ;
        RECT 58.155 127.180 58.445 127.225 ;
        RECT 57.680 127.040 58.445 127.180 ;
        RECT 22.260 126.980 22.580 127.040 ;
        RECT 57.680 126.980 58.000 127.040 ;
        RECT 58.155 126.995 58.445 127.040 ;
        RECT 76.095 127.180 76.385 127.225 ;
        RECT 81.600 127.180 81.920 127.240 ;
        RECT 76.095 127.040 81.920 127.180 ;
        RECT 76.095 126.995 76.385 127.040 ;
        RECT 81.600 126.980 81.920 127.040 ;
        RECT 82.535 127.180 82.825 127.225 ;
        RECT 83.440 127.180 83.760 127.240 ;
        RECT 82.535 127.040 83.760 127.180 ;
        RECT 82.535 126.995 82.825 127.040 ;
        RECT 83.440 126.980 83.760 127.040 ;
        RECT 84.360 127.180 84.680 127.240 ;
        RECT 92.270 127.180 92.410 127.675 ;
        RECT 98.620 127.660 98.940 127.720 ;
        RECT 105.060 127.660 105.380 127.720 ;
        RECT 108.755 127.675 109.045 127.720 ;
        RECT 109.200 127.660 109.520 127.920 ;
        RECT 114.720 127.860 115.040 127.920 ;
        RECT 119.410 127.860 119.550 128.015 ;
        RECT 114.720 127.720 119.550 127.860 ;
        RECT 114.720 127.660 115.040 127.720 ;
        RECT 102.760 127.520 103.080 127.580 ;
        RECT 111.515 127.520 111.805 127.565 ;
        RECT 102.760 127.380 111.805 127.520 ;
        RECT 102.760 127.320 103.080 127.380 ;
        RECT 111.515 127.335 111.805 127.380 ;
        RECT 84.360 127.040 92.410 127.180 ;
        RECT 84.360 126.980 84.680 127.040 ;
        RECT 118.400 126.980 118.720 127.240 ;
        RECT 120.240 126.980 120.560 127.240 ;
        RECT 14.370 126.360 127.530 126.840 ;
        RECT 23.640 125.960 23.960 126.220 ;
        RECT 71.035 126.160 71.325 126.205 ;
        RECT 71.940 126.160 72.260 126.220 ;
        RECT 78.380 126.205 78.700 126.220 ;
        RECT 71.035 126.020 72.260 126.160 ;
        RECT 71.035 125.975 71.325 126.020 ;
        RECT 71.940 125.960 72.260 126.020 ;
        RECT 78.165 125.975 78.700 126.205 ;
        RECT 78.380 125.960 78.700 125.975 ;
        RECT 78.840 126.160 79.160 126.220 ;
        RECT 80.220 126.160 80.540 126.220 ;
        RECT 98.620 126.205 98.940 126.220 ;
        RECT 78.840 126.020 80.540 126.160 ;
        RECT 78.840 125.960 79.160 126.020 ;
        RECT 80.220 125.960 80.540 126.020 ;
        RECT 98.405 125.975 98.940 126.205 ;
        RECT 98.620 125.960 98.940 125.975 ;
        RECT 114.720 125.960 115.040 126.220 ;
        RECT 55.380 125.820 55.700 125.880 ;
        RECT 82.030 125.820 82.320 125.865 ;
        RECT 84.810 125.820 85.100 125.865 ;
        RECT 86.670 125.820 86.960 125.865 ;
        RECT 55.380 125.680 60.670 125.820 ;
        RECT 55.380 125.620 55.700 125.680 ;
        RECT 19.500 125.480 19.820 125.540 ;
        RECT 30.080 125.480 30.400 125.540 ;
        RECT 19.500 125.340 30.400 125.480 ;
        RECT 19.500 125.280 19.820 125.340 ;
        RECT 20.880 125.140 21.200 125.200 ;
        RECT 21.890 125.185 22.030 125.340 ;
        RECT 30.080 125.280 30.400 125.340 ;
        RECT 35.600 125.480 35.920 125.540 ;
        RECT 42.515 125.480 42.805 125.525 ;
        RECT 54.460 125.480 54.780 125.540 ;
        RECT 59.535 125.480 59.825 125.525 ;
        RECT 35.600 125.340 42.805 125.480 ;
        RECT 35.600 125.280 35.920 125.340 ;
        RECT 42.515 125.295 42.805 125.340 ;
        RECT 43.510 125.340 45.950 125.480 ;
        RECT 21.355 125.140 21.645 125.185 ;
        RECT 20.880 125.000 21.645 125.140 ;
        RECT 20.880 124.940 21.200 125.000 ;
        RECT 21.355 124.955 21.645 125.000 ;
        RECT 21.815 124.955 22.105 125.185 ;
        RECT 22.720 124.940 23.040 125.200 ;
        RECT 36.520 124.940 36.840 125.200 ;
        RECT 37.455 124.955 37.745 125.185 ;
        RECT 37.900 125.140 38.220 125.200 ;
        RECT 38.375 125.140 38.665 125.185 ;
        RECT 37.900 125.000 38.665 125.140 ;
        RECT 37.530 124.800 37.670 124.955 ;
        RECT 37.900 124.940 38.220 125.000 ;
        RECT 38.375 124.955 38.665 125.000 ;
        RECT 40.200 124.940 40.520 125.200 ;
        RECT 41.135 124.955 41.425 125.185 ;
        RECT 39.740 124.800 40.060 124.860 ;
        RECT 37.530 124.660 40.060 124.800 ;
        RECT 41.210 124.800 41.350 124.955 ;
        RECT 42.040 124.940 42.360 125.200 ;
        RECT 43.510 125.185 43.650 125.340 ;
        RECT 45.810 125.200 45.950 125.340 ;
        RECT 54.460 125.340 59.825 125.480 ;
        RECT 60.530 125.480 60.670 125.680 ;
        RECT 82.030 125.680 86.960 125.820 ;
        RECT 82.030 125.635 82.320 125.680 ;
        RECT 84.810 125.635 85.100 125.680 ;
        RECT 86.670 125.635 86.960 125.680 ;
        RECT 89.900 125.820 90.190 125.865 ;
        RECT 91.760 125.820 92.050 125.865 ;
        RECT 94.540 125.820 94.830 125.865 ;
        RECT 89.900 125.680 94.830 125.820 ;
        RECT 89.900 125.635 90.190 125.680 ;
        RECT 91.760 125.635 92.050 125.680 ;
        RECT 94.540 125.635 94.830 125.680 ;
        RECT 119.290 125.820 119.580 125.865 ;
        RECT 122.070 125.820 122.360 125.865 ;
        RECT 123.930 125.820 124.220 125.865 ;
        RECT 119.290 125.680 124.220 125.820 ;
        RECT 119.290 125.635 119.580 125.680 ;
        RECT 122.070 125.635 122.360 125.680 ;
        RECT 123.930 125.635 124.220 125.680 ;
        RECT 74.255 125.480 74.545 125.525 ;
        RECT 79.300 125.480 79.620 125.540 ;
        RECT 84.360 125.480 84.680 125.540 ;
        RECT 60.530 125.340 61.130 125.480 ;
        RECT 54.460 125.280 54.780 125.340 ;
        RECT 59.535 125.295 59.825 125.340 ;
        RECT 43.435 125.140 43.725 125.185 ;
        RECT 42.590 125.000 43.725 125.140 ;
        RECT 42.590 124.800 42.730 125.000 ;
        RECT 43.435 124.955 43.725 125.000 ;
        RECT 44.340 124.940 44.660 125.200 ;
        RECT 45.720 124.940 46.040 125.200 ;
        RECT 46.180 124.940 46.500 125.200 ;
        RECT 57.680 124.940 58.000 125.200 ;
        RECT 60.440 124.940 60.760 125.200 ;
        RECT 60.990 125.185 61.130 125.340 ;
        RECT 74.255 125.340 84.680 125.480 ;
        RECT 74.255 125.295 74.545 125.340 ;
        RECT 79.300 125.280 79.620 125.340 ;
        RECT 84.360 125.280 84.680 125.340 ;
        RECT 88.040 125.480 88.360 125.540 ;
        RECT 91.275 125.480 91.565 125.525 ;
        RECT 98.160 125.480 98.480 125.540 ;
        RECT 88.040 125.340 91.565 125.480 ;
        RECT 88.040 125.280 88.360 125.340 ;
        RECT 91.275 125.295 91.565 125.340 ;
        RECT 91.810 125.340 98.480 125.480 ;
        RECT 60.915 124.955 61.205 125.185 ;
        RECT 68.260 125.140 68.580 125.200 ;
        RECT 68.735 125.140 69.025 125.185 ;
        RECT 68.260 125.000 69.025 125.140 ;
        RECT 68.260 124.940 68.580 125.000 ;
        RECT 68.735 124.955 69.025 125.000 ;
        RECT 69.195 125.140 69.485 125.185 ;
        RECT 69.640 125.140 69.960 125.200 ;
        RECT 69.195 125.000 69.960 125.140 ;
        RECT 69.195 124.955 69.485 125.000 ;
        RECT 69.640 124.940 69.960 125.000 ;
        RECT 70.100 124.940 70.420 125.200 ;
        RECT 71.480 125.140 71.800 125.200 ;
        RECT 72.875 125.140 73.165 125.185 ;
        RECT 70.880 125.000 73.165 125.140 ;
        RECT 41.210 124.660 42.730 124.800 ;
        RECT 42.960 124.800 43.280 124.860 ;
        RECT 44.815 124.800 45.105 124.845 ;
        RECT 42.960 124.660 45.105 124.800 ;
        RECT 39.740 124.600 40.060 124.660 ;
        RECT 42.960 124.600 43.280 124.660 ;
        RECT 44.815 124.615 45.105 124.660 ;
        RECT 48.955 124.800 49.245 124.845 ;
        RECT 70.880 124.800 71.020 125.000 ;
        RECT 71.480 124.940 71.800 125.000 ;
        RECT 72.875 124.955 73.165 125.000 ;
        RECT 82.030 125.140 82.320 125.185 ;
        RECT 82.030 125.000 84.565 125.140 ;
        RECT 82.030 124.955 82.320 125.000 ;
        RECT 48.955 124.660 71.020 124.800 ;
        RECT 80.170 124.800 80.460 124.845 ;
        RECT 82.520 124.800 82.840 124.860 ;
        RECT 84.350 124.845 84.565 125.000 ;
        RECT 85.280 124.940 85.600 125.200 ;
        RECT 87.135 125.140 87.425 125.185 ;
        RECT 89.435 125.140 89.725 125.185 ;
        RECT 91.810 125.140 91.950 125.340 ;
        RECT 98.160 125.280 98.480 125.340 ;
        RECT 111.975 125.480 112.265 125.525 ;
        RECT 113.340 125.480 113.660 125.540 ;
        RECT 111.975 125.340 113.660 125.480 ;
        RECT 111.975 125.295 112.265 125.340 ;
        RECT 113.340 125.280 113.660 125.340 ;
        RECT 120.240 125.480 120.560 125.540 ;
        RECT 122.555 125.480 122.845 125.525 ;
        RECT 120.240 125.340 122.845 125.480 ;
        RECT 120.240 125.280 120.560 125.340 ;
        RECT 122.555 125.295 122.845 125.340 ;
        RECT 94.540 125.140 94.830 125.185 ;
        RECT 87.135 125.000 91.950 125.140 ;
        RECT 92.295 125.000 94.830 125.140 ;
        RECT 87.135 124.955 87.425 125.000 ;
        RECT 89.435 124.955 89.725 125.000 ;
        RECT 92.295 124.845 92.510 125.000 ;
        RECT 94.540 124.955 94.830 125.000 ;
        RECT 99.080 124.940 99.400 125.200 ;
        RECT 100.000 124.940 100.320 125.200 ;
        RECT 100.920 124.940 101.240 125.200 ;
        RECT 105.060 125.140 105.380 125.200 ;
        RECT 112.435 125.140 112.725 125.185 ;
        RECT 105.060 125.000 112.725 125.140 ;
        RECT 105.060 124.940 105.380 125.000 ;
        RECT 112.435 124.955 112.725 125.000 ;
        RECT 119.290 125.140 119.580 125.185 ;
        RECT 119.290 125.000 121.825 125.140 ;
        RECT 119.290 124.955 119.580 125.000 ;
        RECT 83.430 124.800 83.720 124.845 ;
        RECT 80.170 124.660 83.720 124.800 ;
        RECT 48.955 124.615 49.245 124.660 ;
        RECT 80.170 124.615 80.460 124.660 ;
        RECT 82.520 124.600 82.840 124.660 ;
        RECT 83.430 124.615 83.720 124.660 ;
        RECT 84.350 124.800 84.640 124.845 ;
        RECT 86.210 124.800 86.500 124.845 ;
        RECT 84.350 124.660 86.500 124.800 ;
        RECT 84.350 124.615 84.640 124.660 ;
        RECT 86.210 124.615 86.500 124.660 ;
        RECT 90.360 124.800 90.650 124.845 ;
        RECT 92.220 124.800 92.510 124.845 ;
        RECT 90.360 124.660 92.510 124.800 ;
        RECT 90.360 124.615 90.650 124.660 ;
        RECT 92.220 124.615 92.510 124.660 ;
        RECT 93.100 124.845 93.420 124.860 ;
        RECT 93.100 124.800 93.430 124.845 ;
        RECT 96.400 124.800 96.690 124.845 ;
        RECT 93.100 124.660 96.690 124.800 ;
        RECT 93.100 124.615 93.430 124.660 ;
        RECT 96.400 124.615 96.690 124.660 ;
        RECT 117.430 124.800 117.720 124.845 ;
        RECT 118.400 124.800 118.720 124.860 ;
        RECT 121.610 124.845 121.825 125.000 ;
        RECT 124.380 124.940 124.700 125.200 ;
        RECT 120.690 124.800 120.980 124.845 ;
        RECT 117.430 124.660 120.980 124.800 ;
        RECT 117.430 124.615 117.720 124.660 ;
        RECT 93.100 124.600 93.420 124.615 ;
        RECT 118.400 124.600 118.720 124.660 ;
        RECT 120.690 124.615 120.980 124.660 ;
        RECT 121.610 124.800 121.900 124.845 ;
        RECT 123.470 124.800 123.760 124.845 ;
        RECT 121.610 124.660 123.760 124.800 ;
        RECT 121.610 124.615 121.900 124.660 ;
        RECT 123.470 124.615 123.760 124.660 ;
        RECT 45.720 124.460 46.040 124.520 ;
        RECT 47.575 124.460 47.865 124.505 ;
        RECT 45.720 124.320 47.865 124.460 ;
        RECT 45.720 124.260 46.040 124.320 ;
        RECT 47.575 124.275 47.865 124.320 ;
        RECT 58.615 124.460 58.905 124.505 ;
        RECT 59.980 124.460 60.300 124.520 ;
        RECT 58.615 124.320 60.300 124.460 ;
        RECT 58.615 124.275 58.905 124.320 ;
        RECT 59.980 124.260 60.300 124.320 ;
        RECT 62.755 124.460 63.045 124.505 ;
        RECT 69.640 124.460 69.960 124.520 ;
        RECT 62.755 124.320 69.960 124.460 ;
        RECT 62.755 124.275 63.045 124.320 ;
        RECT 69.640 124.260 69.960 124.320 ;
        RECT 112.880 124.460 113.200 124.520 ;
        RECT 115.425 124.460 115.715 124.505 ;
        RECT 112.880 124.320 115.715 124.460 ;
        RECT 112.880 124.260 113.200 124.320 ;
        RECT 115.425 124.275 115.715 124.320 ;
        RECT 14.370 123.640 127.530 124.120 ;
        RECT 22.260 123.440 22.580 123.500 ;
        RECT 23.180 123.440 23.500 123.500 ;
        RECT 24.115 123.440 24.405 123.485 ;
        RECT 22.260 123.240 22.720 123.440 ;
        RECT 23.180 123.300 24.405 123.440 ;
        RECT 23.180 123.240 23.500 123.300 ;
        RECT 24.115 123.255 24.405 123.300 ;
        RECT 24.575 123.440 24.865 123.485 ;
        RECT 42.500 123.440 42.820 123.500 ;
        RECT 24.575 123.300 42.820 123.440 ;
        RECT 24.575 123.255 24.865 123.300 ;
        RECT 22.580 123.100 22.720 123.240 ;
        RECT 24.650 123.100 24.790 123.255 ;
        RECT 42.500 123.240 42.820 123.300 ;
        RECT 52.865 123.440 53.155 123.485 ;
        RECT 55.380 123.440 55.700 123.500 ;
        RECT 52.865 123.300 55.700 123.440 ;
        RECT 52.865 123.255 53.155 123.300 ;
        RECT 55.380 123.240 55.700 123.300 ;
        RECT 60.440 123.440 60.760 123.500 ;
        RECT 65.515 123.440 65.805 123.485 ;
        RECT 60.440 123.300 65.805 123.440 ;
        RECT 60.440 123.240 60.760 123.300 ;
        RECT 65.515 123.255 65.805 123.300 ;
        RECT 82.075 123.440 82.365 123.485 ;
        RECT 82.520 123.440 82.840 123.500 ;
        RECT 82.075 123.300 82.840 123.440 ;
        RECT 82.075 123.255 82.365 123.300 ;
        RECT 82.520 123.240 82.840 123.300 ;
        RECT 84.375 123.440 84.665 123.485 ;
        RECT 85.280 123.440 85.600 123.500 ;
        RECT 84.375 123.300 85.600 123.440 ;
        RECT 84.375 123.255 84.665 123.300 ;
        RECT 85.280 123.240 85.600 123.300 ;
        RECT 93.100 123.240 93.420 123.500 ;
        RECT 22.580 122.960 24.790 123.100 ;
        RECT 54.870 123.100 55.160 123.145 ;
        RECT 57.220 123.100 57.540 123.160 ;
        RECT 58.130 123.100 58.420 123.145 ;
        RECT 54.870 122.960 58.420 123.100 ;
        RECT 54.870 122.915 55.160 122.960 ;
        RECT 57.220 122.900 57.540 122.960 ;
        RECT 58.130 122.915 58.420 122.960 ;
        RECT 59.050 123.100 59.340 123.145 ;
        RECT 60.910 123.100 61.200 123.145 ;
        RECT 59.050 122.960 61.200 123.100 ;
        RECT 59.050 122.915 59.340 122.960 ;
        RECT 60.910 122.915 61.200 122.960 ;
        RECT 111.515 123.100 111.805 123.145 ;
        RECT 112.880 123.100 113.200 123.160 ;
        RECT 111.515 122.960 113.200 123.100 ;
        RECT 111.515 122.915 111.805 122.960 ;
        RECT 34.680 122.560 35.000 122.820 ;
        RECT 56.730 122.760 57.020 122.805 ;
        RECT 59.050 122.760 59.265 122.915 ;
        RECT 112.880 122.900 113.200 122.960 ;
        RECT 117.430 123.100 117.720 123.145 ;
        RECT 118.860 123.100 119.180 123.160 ;
        RECT 120.690 123.100 120.980 123.145 ;
        RECT 117.430 122.960 120.980 123.100 ;
        RECT 117.430 122.915 117.720 122.960 ;
        RECT 118.860 122.900 119.180 122.960 ;
        RECT 120.690 122.915 120.980 122.960 ;
        RECT 121.610 123.100 121.900 123.145 ;
        RECT 123.470 123.100 123.760 123.145 ;
        RECT 121.610 122.960 123.760 123.100 ;
        RECT 121.610 122.915 121.900 122.960 ;
        RECT 123.470 122.915 123.760 122.960 ;
        RECT 56.730 122.620 59.265 122.760 ;
        RECT 56.730 122.575 57.020 122.620 ;
        RECT 59.980 122.560 60.300 122.820 ;
        RECT 61.835 122.760 62.125 122.805 ;
        RECT 63.660 122.760 63.980 122.820 ;
        RECT 61.835 122.620 63.980 122.760 ;
        RECT 61.835 122.575 62.125 122.620 ;
        RECT 63.660 122.560 63.980 122.620 ;
        RECT 64.120 122.760 64.440 122.820 ;
        RECT 65.055 122.760 65.345 122.805 ;
        RECT 64.120 122.620 65.345 122.760 ;
        RECT 64.120 122.560 64.440 122.620 ;
        RECT 65.055 122.575 65.345 122.620 ;
        RECT 72.860 122.760 73.180 122.820 ;
        RECT 82.535 122.760 82.825 122.805 ;
        RECT 82.980 122.760 83.300 122.820 ;
        RECT 72.860 122.620 83.300 122.760 ;
        RECT 72.860 122.560 73.180 122.620 ;
        RECT 82.535 122.575 82.825 122.620 ;
        RECT 82.980 122.560 83.300 122.620 ;
        RECT 83.440 122.560 83.760 122.820 ;
        RECT 90.800 122.760 91.120 122.820 ;
        RECT 92.655 122.760 92.945 122.805 ;
        RECT 100.000 122.760 100.320 122.820 ;
        RECT 90.800 122.620 100.320 122.760 ;
        RECT 90.800 122.560 91.120 122.620 ;
        RECT 92.655 122.575 92.945 122.620 ;
        RECT 100.000 122.560 100.320 122.620 ;
        RECT 111.975 122.760 112.265 122.805 ;
        RECT 112.420 122.760 112.740 122.820 ;
        RECT 115.425 122.760 115.715 122.805 ;
        RECT 111.975 122.620 115.715 122.760 ;
        RECT 111.975 122.575 112.265 122.620 ;
        RECT 112.420 122.560 112.740 122.620 ;
        RECT 115.425 122.575 115.715 122.620 ;
        RECT 119.290 122.760 119.580 122.805 ;
        RECT 121.610 122.760 121.825 122.915 ;
        RECT 119.290 122.620 121.825 122.760 ;
        RECT 119.290 122.575 119.580 122.620 ;
        RECT 124.380 122.560 124.700 122.820 ;
        RECT 21.800 122.420 22.120 122.480 ;
        RECT 23.195 122.420 23.485 122.465 ;
        RECT 33.315 122.420 33.605 122.465 ;
        RECT 21.800 122.280 33.605 122.420 ;
        RECT 21.800 122.220 22.120 122.280 ;
        RECT 23.195 122.235 23.485 122.280 ;
        RECT 33.315 122.235 33.605 122.280 ;
        RECT 34.235 122.420 34.525 122.465 ;
        RECT 36.520 122.420 36.840 122.480 ;
        RECT 41.580 122.420 41.900 122.480 ;
        RECT 34.235 122.280 41.900 122.420 ;
        RECT 34.235 122.235 34.525 122.280 ;
        RECT 33.390 122.080 33.530 122.235 ;
        RECT 36.520 122.220 36.840 122.280 ;
        RECT 41.580 122.220 41.900 122.280 ;
        RECT 64.580 122.220 64.900 122.480 ;
        RECT 105.060 122.420 105.380 122.480 ;
        RECT 110.595 122.420 110.885 122.465 ;
        RECT 113.340 122.420 113.660 122.480 ;
        RECT 105.060 122.280 113.660 122.420 ;
        RECT 105.060 122.220 105.380 122.280 ;
        RECT 110.595 122.235 110.885 122.280 ;
        RECT 113.340 122.220 113.660 122.280 ;
        RECT 121.160 122.420 121.480 122.480 ;
        RECT 122.555 122.420 122.845 122.465 ;
        RECT 121.160 122.280 122.845 122.420 ;
        RECT 121.160 122.220 121.480 122.280 ;
        RECT 122.555 122.235 122.845 122.280 ;
        RECT 43.420 122.080 43.740 122.140 ;
        RECT 45.720 122.080 46.040 122.140 ;
        RECT 46.640 122.080 46.960 122.140 ;
        RECT 33.390 121.940 46.960 122.080 ;
        RECT 43.420 121.880 43.740 121.940 ;
        RECT 45.720 121.880 46.040 121.940 ;
        RECT 46.640 121.880 46.960 121.940 ;
        RECT 56.730 122.080 57.020 122.125 ;
        RECT 59.510 122.080 59.800 122.125 ;
        RECT 61.370 122.080 61.660 122.125 ;
        RECT 56.730 121.940 61.660 122.080 ;
        RECT 56.730 121.895 57.020 121.940 ;
        RECT 59.510 121.895 59.800 121.940 ;
        RECT 61.370 121.895 61.660 121.940 ;
        RECT 119.290 122.080 119.580 122.125 ;
        RECT 122.070 122.080 122.360 122.125 ;
        RECT 123.930 122.080 124.220 122.125 ;
        RECT 119.290 121.940 124.220 122.080 ;
        RECT 119.290 121.895 119.580 121.940 ;
        RECT 122.070 121.895 122.360 121.940 ;
        RECT 123.930 121.895 124.220 121.940 ;
        RECT 26.400 121.540 26.720 121.800 ;
        RECT 36.520 121.540 36.840 121.800 ;
        RECT 67.355 121.740 67.645 121.785 ;
        RECT 67.800 121.740 68.120 121.800 ;
        RECT 67.355 121.600 68.120 121.740 ;
        RECT 67.355 121.555 67.645 121.600 ;
        RECT 67.800 121.540 68.120 121.600 ;
        RECT 113.815 121.740 114.105 121.785 ;
        RECT 120.240 121.740 120.560 121.800 ;
        RECT 113.815 121.600 120.560 121.740 ;
        RECT 113.815 121.555 114.105 121.600 ;
        RECT 120.240 121.540 120.560 121.600 ;
        RECT 14.370 120.920 127.530 121.400 ;
        RECT 30.325 120.720 30.615 120.765 ;
        RECT 34.680 120.720 35.000 120.780 ;
        RECT 30.325 120.580 35.000 120.720 ;
        RECT 30.325 120.535 30.615 120.580 ;
        RECT 34.680 120.520 35.000 120.580 ;
        RECT 57.220 120.520 57.540 120.780 ;
        RECT 59.305 120.720 59.595 120.765 ;
        RECT 60.440 120.720 60.760 120.780 ;
        RECT 59.305 120.580 60.760 120.720 ;
        RECT 59.305 120.535 59.595 120.580 ;
        RECT 60.440 120.520 60.760 120.580 ;
        RECT 118.860 120.520 119.180 120.780 ;
        RECT 121.160 120.520 121.480 120.780 ;
        RECT 21.800 120.380 22.120 120.440 ;
        RECT 34.190 120.380 34.480 120.425 ;
        RECT 36.970 120.380 37.260 120.425 ;
        RECT 38.830 120.380 39.120 120.425 ;
        RECT 63.170 120.380 63.460 120.425 ;
        RECT 65.950 120.380 66.240 120.425 ;
        RECT 67.810 120.380 68.100 120.425 ;
        RECT 21.800 120.240 22.950 120.380 ;
        RECT 21.800 120.180 22.120 120.240 ;
        RECT 22.260 119.840 22.580 120.100 ;
        RECT 22.810 120.085 22.950 120.240 ;
        RECT 34.190 120.240 39.120 120.380 ;
        RECT 34.190 120.195 34.480 120.240 ;
        RECT 36.970 120.195 37.260 120.240 ;
        RECT 38.830 120.195 39.120 120.240 ;
        RECT 42.590 120.240 47.330 120.380 ;
        RECT 22.735 119.855 23.025 120.085 ;
        RECT 35.600 120.040 35.920 120.100 ;
        RECT 42.590 120.040 42.730 120.240 ;
        RECT 30.630 119.900 42.730 120.040 ;
        RECT 42.975 120.040 43.265 120.085 ;
        RECT 43.420 120.040 43.740 120.100 ;
        RECT 42.975 119.900 43.740 120.040 ;
        RECT 26.400 119.700 26.720 119.760 ;
        RECT 26.875 119.700 27.165 119.745 ;
        RECT 26.400 119.560 27.165 119.700 ;
        RECT 26.400 119.500 26.720 119.560 ;
        RECT 26.875 119.515 27.165 119.560 ;
        RECT 30.630 119.420 30.770 119.900 ;
        RECT 35.600 119.840 35.920 119.900 ;
        RECT 42.975 119.855 43.265 119.900 ;
        RECT 43.420 119.840 43.740 119.900 ;
        RECT 46.180 119.840 46.500 120.100 ;
        RECT 46.640 119.840 46.960 120.100 ;
        RECT 47.190 120.085 47.330 120.240 ;
        RECT 63.170 120.240 68.100 120.380 ;
        RECT 63.170 120.195 63.460 120.240 ;
        RECT 65.950 120.195 66.240 120.240 ;
        RECT 67.810 120.195 68.100 120.240 ;
        RECT 68.735 120.195 69.025 120.425 ;
        RECT 112.850 120.380 113.140 120.425 ;
        RECT 115.630 120.380 115.920 120.425 ;
        RECT 117.490 120.380 117.780 120.425 ;
        RECT 112.850 120.240 117.780 120.380 ;
        RECT 112.850 120.195 113.140 120.240 ;
        RECT 115.630 120.195 115.920 120.240 ;
        RECT 117.490 120.195 117.780 120.240 ;
        RECT 47.115 119.855 47.405 120.085 ;
        RECT 66.435 120.040 66.725 120.085 ;
        RECT 68.810 120.040 68.950 120.195 ;
        RECT 66.435 119.900 68.950 120.040 ;
        RECT 77.475 120.040 77.765 120.085 ;
        RECT 79.300 120.040 79.620 120.100 ;
        RECT 83.440 120.040 83.760 120.100 ;
        RECT 93.575 120.040 93.865 120.085 ;
        RECT 97.715 120.040 98.005 120.085 ;
        RECT 105.060 120.040 105.380 120.100 ;
        RECT 109.200 120.085 109.520 120.100 ;
        RECT 77.475 119.900 105.380 120.040 ;
        RECT 66.435 119.855 66.725 119.900 ;
        RECT 77.475 119.855 77.765 119.900 ;
        RECT 79.300 119.840 79.620 119.900 ;
        RECT 83.440 119.840 83.760 119.900 ;
        RECT 93.575 119.855 93.865 119.900 ;
        RECT 97.715 119.855 98.005 119.900 ;
        RECT 105.060 119.840 105.380 119.900 ;
        RECT 105.995 120.040 106.285 120.085 ;
        RECT 108.985 120.040 109.520 120.085 ;
        RECT 105.995 119.900 109.520 120.040 ;
        RECT 105.995 119.855 106.285 119.900 ;
        RECT 108.985 119.855 109.520 119.900 ;
        RECT 109.200 119.840 109.520 119.855 ;
        RECT 109.750 119.900 118.630 120.040 ;
        RECT 34.190 119.700 34.480 119.745 ;
        RECT 34.190 119.560 36.725 119.700 ;
        RECT 34.190 119.515 34.480 119.560 ;
        RECT 21.815 119.360 22.105 119.405 ;
        RECT 30.540 119.360 30.860 119.420 ;
        RECT 21.815 119.220 30.860 119.360 ;
        RECT 21.815 119.175 22.105 119.220 ;
        RECT 30.540 119.160 30.860 119.220 ;
        RECT 32.330 119.360 32.620 119.405 ;
        RECT 34.680 119.360 35.000 119.420 ;
        RECT 36.510 119.405 36.725 119.560 ;
        RECT 37.440 119.500 37.760 119.760 ;
        RECT 39.295 119.515 39.585 119.745 ;
        RECT 35.590 119.360 35.880 119.405 ;
        RECT 32.330 119.220 35.880 119.360 ;
        RECT 32.330 119.175 32.620 119.220 ;
        RECT 34.680 119.160 35.000 119.220 ;
        RECT 35.590 119.175 35.880 119.220 ;
        RECT 36.510 119.360 36.800 119.405 ;
        RECT 38.370 119.360 38.660 119.405 ;
        RECT 36.510 119.220 38.660 119.360 ;
        RECT 39.370 119.360 39.510 119.515 ;
        RECT 41.580 119.500 41.900 119.760 ;
        RECT 45.260 119.500 45.580 119.760 ;
        RECT 46.270 119.700 46.410 119.840 ;
        RECT 47.575 119.700 47.865 119.745 ;
        RECT 46.270 119.560 47.865 119.700 ;
        RECT 47.575 119.515 47.865 119.560 ;
        RECT 49.860 119.700 50.180 119.760 ;
        RECT 50.335 119.700 50.625 119.745 ;
        RECT 54.015 119.700 54.305 119.745 ;
        RECT 49.860 119.560 54.305 119.700 ;
        RECT 49.860 119.500 50.180 119.560 ;
        RECT 50.335 119.515 50.625 119.560 ;
        RECT 54.015 119.515 54.305 119.560 ;
        RECT 55.395 119.700 55.685 119.745 ;
        RECT 57.680 119.700 58.000 119.760 ;
        RECT 55.395 119.560 58.000 119.700 ;
        RECT 55.395 119.515 55.685 119.560 ;
        RECT 57.680 119.500 58.000 119.560 ;
        RECT 63.170 119.700 63.460 119.745 ;
        RECT 63.170 119.560 65.705 119.700 ;
        RECT 63.170 119.515 63.460 119.560 ;
        RECT 46.180 119.360 46.500 119.420 ;
        RECT 39.370 119.220 46.500 119.360 ;
        RECT 36.510 119.175 36.800 119.220 ;
        RECT 38.370 119.175 38.660 119.220 ;
        RECT 46.180 119.160 46.500 119.220 ;
        RECT 61.310 119.360 61.600 119.405 ;
        RECT 61.820 119.360 62.140 119.420 ;
        RECT 65.490 119.405 65.705 119.560 ;
        RECT 68.275 119.515 68.565 119.745 ;
        RECT 64.570 119.360 64.860 119.405 ;
        RECT 61.310 119.220 64.860 119.360 ;
        RECT 61.310 119.175 61.600 119.220 ;
        RECT 61.820 119.160 62.140 119.220 ;
        RECT 64.570 119.175 64.860 119.220 ;
        RECT 65.490 119.360 65.780 119.405 ;
        RECT 67.350 119.360 67.640 119.405 ;
        RECT 65.490 119.220 67.640 119.360 ;
        RECT 68.350 119.360 68.490 119.515 ;
        RECT 69.640 119.500 69.960 119.760 ;
        RECT 72.860 119.700 73.180 119.760 ;
        RECT 74.255 119.700 74.545 119.745 ;
        RECT 81.615 119.700 81.905 119.745 ;
        RECT 72.860 119.560 74.545 119.700 ;
        RECT 72.860 119.500 73.180 119.560 ;
        RECT 74.255 119.515 74.545 119.560 ;
        RECT 80.310 119.560 81.905 119.700 ;
        RECT 70.560 119.360 70.880 119.420 ;
        RECT 68.350 119.220 70.880 119.360 ;
        RECT 65.490 119.175 65.780 119.220 ;
        RECT 67.350 119.175 67.640 119.220 ;
        RECT 70.560 119.160 70.880 119.220 ;
        RECT 77.935 119.360 78.225 119.405 ;
        RECT 79.300 119.360 79.620 119.420 ;
        RECT 77.935 119.220 79.620 119.360 ;
        RECT 77.935 119.175 78.225 119.220 ;
        RECT 79.300 119.160 79.620 119.220 ;
        RECT 19.975 119.020 20.265 119.065 ;
        RECT 20.880 119.020 21.200 119.080 ;
        RECT 19.975 118.880 21.200 119.020 ;
        RECT 19.975 118.835 20.265 118.880 ;
        RECT 20.880 118.820 21.200 118.880 ;
        RECT 25.020 119.020 25.340 119.080 ;
        RECT 25.955 119.020 26.245 119.065 ;
        RECT 25.020 118.880 26.245 119.020 ;
        RECT 25.020 118.820 25.340 118.880 ;
        RECT 25.955 118.835 26.245 118.880 ;
        RECT 39.740 118.820 40.060 119.080 ;
        RECT 42.040 118.820 42.360 119.080 ;
        RECT 44.355 119.020 44.645 119.065 ;
        RECT 44.800 119.020 45.120 119.080 ;
        RECT 44.355 118.880 45.120 119.020 ;
        RECT 44.355 118.835 44.645 118.880 ;
        RECT 44.800 118.820 45.120 118.880 ;
        RECT 49.400 118.820 49.720 119.080 ;
        RECT 50.780 118.820 51.100 119.080 ;
        RECT 74.715 119.020 75.005 119.065 ;
        RECT 75.160 119.020 75.480 119.080 ;
        RECT 74.715 118.880 75.480 119.020 ;
        RECT 74.715 118.835 75.005 118.880 ;
        RECT 75.160 118.820 75.480 118.880 ;
        RECT 78.395 119.020 78.685 119.065 ;
        RECT 78.840 119.020 79.160 119.080 ;
        RECT 80.310 119.065 80.450 119.560 ;
        RECT 81.615 119.515 81.905 119.560 ;
        RECT 82.980 119.500 83.300 119.760 ;
        RECT 83.900 119.500 84.220 119.760 ;
        RECT 93.100 119.700 93.420 119.760 ;
        RECT 99.080 119.700 99.400 119.760 ;
        RECT 93.100 119.560 99.400 119.700 ;
        RECT 93.100 119.500 93.420 119.560 ;
        RECT 99.080 119.500 99.400 119.560 ;
        RECT 100.000 119.700 100.320 119.760 ;
        RECT 103.235 119.700 103.525 119.745 ;
        RECT 109.750 119.700 109.890 119.900 ;
        RECT 118.490 119.760 118.630 119.900 ;
        RECT 100.000 119.560 109.890 119.700 ;
        RECT 112.850 119.700 113.140 119.745 ;
        RECT 112.850 119.560 115.385 119.700 ;
        RECT 100.000 119.500 100.320 119.560 ;
        RECT 103.235 119.515 103.525 119.560 ;
        RECT 112.850 119.515 113.140 119.560 ;
        RECT 98.635 119.360 98.925 119.405 ;
        RECT 102.300 119.360 102.620 119.420 ;
        RECT 105.980 119.360 106.300 119.420 ;
        RECT 106.455 119.360 106.745 119.405 ;
        RECT 98.635 119.220 106.745 119.360 ;
        RECT 98.635 119.175 98.925 119.220 ;
        RECT 102.300 119.160 102.620 119.220 ;
        RECT 105.980 119.160 106.300 119.220 ;
        RECT 106.455 119.175 106.745 119.220 ;
        RECT 110.990 119.360 111.280 119.405 ;
        RECT 113.340 119.360 113.660 119.420 ;
        RECT 115.170 119.405 115.385 119.560 ;
        RECT 116.100 119.500 116.420 119.760 ;
        RECT 117.955 119.515 118.245 119.745 ;
        RECT 114.250 119.360 114.540 119.405 ;
        RECT 110.990 119.220 114.540 119.360 ;
        RECT 110.990 119.175 111.280 119.220 ;
        RECT 113.340 119.160 113.660 119.220 ;
        RECT 114.250 119.175 114.540 119.220 ;
        RECT 115.170 119.360 115.460 119.405 ;
        RECT 117.030 119.360 117.320 119.405 ;
        RECT 115.170 119.220 117.320 119.360 ;
        RECT 115.170 119.175 115.460 119.220 ;
        RECT 117.030 119.175 117.320 119.220 ;
        RECT 78.395 118.880 79.160 119.020 ;
        RECT 78.395 118.835 78.685 118.880 ;
        RECT 78.840 118.820 79.160 118.880 ;
        RECT 80.235 118.835 80.525 119.065 ;
        RECT 80.680 118.820 81.000 119.080 ;
        RECT 82.520 118.820 82.840 119.080 ;
        RECT 84.360 119.020 84.680 119.080 ;
        RECT 84.835 119.020 85.125 119.065 ;
        RECT 84.360 118.880 85.125 119.020 ;
        RECT 84.360 118.820 84.680 118.880 ;
        RECT 84.835 118.835 85.125 118.880 ;
        RECT 87.120 119.020 87.440 119.080 ;
        RECT 90.815 119.020 91.105 119.065 ;
        RECT 87.120 118.880 91.105 119.020 ;
        RECT 87.120 118.820 87.440 118.880 ;
        RECT 90.815 118.835 91.105 118.880 ;
        RECT 92.655 119.020 92.945 119.065 ;
        RECT 93.560 119.020 93.880 119.080 ;
        RECT 92.655 118.880 93.880 119.020 ;
        RECT 92.655 118.835 92.945 118.880 ;
        RECT 93.560 118.820 93.880 118.880 ;
        RECT 100.920 118.820 101.240 119.080 ;
        RECT 103.695 119.020 103.985 119.065 ;
        RECT 105.520 119.020 105.840 119.080 ;
        RECT 103.695 118.880 105.840 119.020 ;
        RECT 103.695 118.835 103.985 118.880 ;
        RECT 105.520 118.820 105.840 118.880 ;
        RECT 108.295 119.020 108.585 119.065 ;
        RECT 108.740 119.020 109.060 119.080 ;
        RECT 108.295 118.880 109.060 119.020 ;
        RECT 108.295 118.835 108.585 118.880 ;
        RECT 108.740 118.820 109.060 118.880 ;
        RECT 111.500 119.020 111.820 119.080 ;
        RECT 118.030 119.020 118.170 119.515 ;
        RECT 118.400 119.500 118.720 119.760 ;
        RECT 120.240 119.500 120.560 119.760 ;
        RECT 111.500 118.880 118.170 119.020 ;
        RECT 111.500 118.820 111.820 118.880 ;
        RECT 14.370 118.200 127.530 118.680 ;
        RECT 17.905 118.000 18.195 118.045 ;
        RECT 22.260 118.000 22.580 118.060 ;
        RECT 17.905 117.860 22.580 118.000 ;
        RECT 17.905 117.815 18.195 117.860 ;
        RECT 22.260 117.800 22.580 117.860 ;
        RECT 36.060 118.045 36.380 118.060 ;
        RECT 36.060 117.815 36.595 118.045 ;
        RECT 37.685 118.000 37.975 118.045 ;
        RECT 42.040 118.000 42.360 118.060 ;
        RECT 37.685 117.860 42.360 118.000 ;
        RECT 37.685 117.815 37.975 117.860 ;
        RECT 36.060 117.800 36.380 117.815 ;
        RECT 42.040 117.800 42.360 117.860 ;
        RECT 61.820 117.800 62.140 118.060 ;
        RECT 63.445 118.000 63.735 118.045 ;
        RECT 64.120 118.000 64.440 118.060 ;
        RECT 63.445 117.860 64.440 118.000 ;
        RECT 63.445 117.815 63.735 117.860 ;
        RECT 64.120 117.800 64.440 117.860 ;
        RECT 73.105 118.000 73.395 118.045 ;
        RECT 78.840 118.000 79.160 118.060 ;
        RECT 73.105 117.860 79.160 118.000 ;
        RECT 73.105 117.815 73.395 117.860 ;
        RECT 78.840 117.800 79.160 117.860 ;
        RECT 82.535 118.000 82.825 118.045 ;
        RECT 83.900 118.000 84.220 118.060 ;
        RECT 93.100 118.045 93.420 118.060 ;
        RECT 82.535 117.860 84.220 118.000 ;
        RECT 82.535 117.815 82.825 117.860 ;
        RECT 83.900 117.800 84.220 117.860 ;
        RECT 92.885 117.815 93.420 118.045 ;
        RECT 93.100 117.800 93.420 117.815 ;
        RECT 102.300 118.045 102.620 118.060 ;
        RECT 102.300 117.815 102.835 118.045 ;
        RECT 102.300 117.800 102.620 117.815 ;
        RECT 113.340 117.800 113.660 118.060 ;
        RECT 116.100 117.800 116.420 118.060 ;
        RECT 23.180 117.705 23.500 117.720 ;
        RECT 19.910 117.660 20.200 117.705 ;
        RECT 23.170 117.660 23.500 117.705 ;
        RECT 19.910 117.520 23.500 117.660 ;
        RECT 19.910 117.475 20.200 117.520 ;
        RECT 23.170 117.475 23.500 117.520 ;
        RECT 23.180 117.460 23.500 117.475 ;
        RECT 24.090 117.660 24.380 117.705 ;
        RECT 25.950 117.660 26.240 117.705 ;
        RECT 24.090 117.520 26.240 117.660 ;
        RECT 24.090 117.475 24.380 117.520 ;
        RECT 25.950 117.475 26.240 117.520 ;
        RECT 28.260 117.660 28.550 117.705 ;
        RECT 30.120 117.660 30.410 117.705 ;
        RECT 28.260 117.520 30.410 117.660 ;
        RECT 28.260 117.475 28.550 117.520 ;
        RECT 30.120 117.475 30.410 117.520 ;
        RECT 31.040 117.660 31.330 117.705 ;
        RECT 34.300 117.660 34.590 117.705 ;
        RECT 35.140 117.660 35.460 117.720 ;
        RECT 42.960 117.705 43.280 117.720 ;
        RECT 31.040 117.520 35.460 117.660 ;
        RECT 31.040 117.475 31.330 117.520 ;
        RECT 34.300 117.475 34.590 117.520 ;
        RECT 17.215 117.320 17.505 117.365 ;
        RECT 19.040 117.320 19.360 117.380 ;
        RECT 17.215 117.180 19.360 117.320 ;
        RECT 17.215 117.135 17.505 117.180 ;
        RECT 19.040 117.120 19.360 117.180 ;
        RECT 21.770 117.320 22.060 117.365 ;
        RECT 24.090 117.320 24.305 117.475 ;
        RECT 21.770 117.180 24.305 117.320 ;
        RECT 21.770 117.135 22.060 117.180 ;
        RECT 25.020 117.120 25.340 117.380 ;
        RECT 30.195 117.320 30.410 117.475 ;
        RECT 35.140 117.460 35.460 117.520 ;
        RECT 39.690 117.660 39.980 117.705 ;
        RECT 42.950 117.660 43.280 117.705 ;
        RECT 39.690 117.520 43.280 117.660 ;
        RECT 39.690 117.475 39.980 117.520 ;
        RECT 42.950 117.475 43.280 117.520 ;
        RECT 42.960 117.460 43.280 117.475 ;
        RECT 43.870 117.660 44.160 117.705 ;
        RECT 45.730 117.660 46.020 117.705 ;
        RECT 43.870 117.520 46.020 117.660 ;
        RECT 43.870 117.475 44.160 117.520 ;
        RECT 45.730 117.475 46.020 117.520 ;
        RECT 49.350 117.660 49.640 117.705 ;
        RECT 50.780 117.660 51.100 117.720 ;
        RECT 52.610 117.660 52.900 117.705 ;
        RECT 49.350 117.520 52.900 117.660 ;
        RECT 49.350 117.475 49.640 117.520 ;
        RECT 32.440 117.320 32.730 117.365 ;
        RECT 30.195 117.180 32.730 117.320 ;
        RECT 32.440 117.135 32.730 117.180 ;
        RECT 41.550 117.320 41.840 117.365 ;
        RECT 43.870 117.320 44.085 117.475 ;
        RECT 50.780 117.460 51.100 117.520 ;
        RECT 52.610 117.475 52.900 117.520 ;
        RECT 53.530 117.660 53.820 117.705 ;
        RECT 55.390 117.660 55.680 117.705 ;
        RECT 53.530 117.520 55.680 117.660 ;
        RECT 53.530 117.475 53.820 117.520 ;
        RECT 55.390 117.475 55.680 117.520 ;
        RECT 65.450 117.660 65.740 117.705 ;
        RECT 66.420 117.660 66.740 117.720 ;
        RECT 75.160 117.705 75.480 117.720 ;
        RECT 68.710 117.660 69.000 117.705 ;
        RECT 65.450 117.520 69.000 117.660 ;
        RECT 65.450 117.475 65.740 117.520 ;
        RECT 41.550 117.180 44.085 117.320 ;
        RECT 41.550 117.135 41.840 117.180 ;
        RECT 44.800 117.120 45.120 117.380 ;
        RECT 46.180 117.320 46.500 117.380 ;
        RECT 46.655 117.320 46.945 117.365 ;
        RECT 46.180 117.180 46.945 117.320 ;
        RECT 46.180 117.120 46.500 117.180 ;
        RECT 46.655 117.135 46.945 117.180 ;
        RECT 51.210 117.320 51.500 117.365 ;
        RECT 53.530 117.320 53.745 117.475 ;
        RECT 66.420 117.460 66.740 117.520 ;
        RECT 68.710 117.475 69.000 117.520 ;
        RECT 69.630 117.660 69.920 117.705 ;
        RECT 71.490 117.660 71.780 117.705 ;
        RECT 69.630 117.520 71.780 117.660 ;
        RECT 69.630 117.475 69.920 117.520 ;
        RECT 71.490 117.475 71.780 117.520 ;
        RECT 75.110 117.660 75.480 117.705 ;
        RECT 78.370 117.660 78.660 117.705 ;
        RECT 75.110 117.520 78.660 117.660 ;
        RECT 75.110 117.475 75.480 117.520 ;
        RECT 78.370 117.475 78.660 117.520 ;
        RECT 79.290 117.660 79.580 117.705 ;
        RECT 81.150 117.660 81.440 117.705 ;
        RECT 79.290 117.520 81.440 117.660 ;
        RECT 79.290 117.475 79.580 117.520 ;
        RECT 81.150 117.475 81.440 117.520 ;
        RECT 82.980 117.660 83.300 117.720 ;
        RECT 89.435 117.660 89.725 117.705 ;
        RECT 94.890 117.660 95.180 117.705 ;
        RECT 98.150 117.660 98.440 117.705 ;
        RECT 82.980 117.520 89.190 117.660 ;
        RECT 51.210 117.180 53.745 117.320 ;
        RECT 51.210 117.135 51.500 117.180 ;
        RECT 25.480 116.980 25.800 117.040 ;
        RECT 26.875 116.980 27.165 117.025 ;
        RECT 27.335 116.980 27.625 117.025 ;
        RECT 25.480 116.840 27.625 116.980 ;
        RECT 25.480 116.780 25.800 116.840 ;
        RECT 26.875 116.795 27.165 116.840 ;
        RECT 27.335 116.795 27.625 116.840 ;
        RECT 29.175 116.980 29.465 117.025 ;
        RECT 38.820 116.980 39.140 117.040 ;
        RECT 29.175 116.840 39.140 116.980 ;
        RECT 46.730 116.980 46.870 117.135 ;
        RECT 54.460 117.120 54.780 117.380 ;
        RECT 57.680 117.320 58.000 117.380 ;
        RECT 59.520 117.320 59.840 117.380 ;
        RECT 61.375 117.320 61.665 117.365 ;
        RECT 57.680 117.180 61.665 117.320 ;
        RECT 57.680 117.120 58.000 117.180 ;
        RECT 59.520 117.120 59.840 117.180 ;
        RECT 61.375 117.135 61.665 117.180 ;
        RECT 67.310 117.320 67.600 117.365 ;
        RECT 69.630 117.320 69.845 117.475 ;
        RECT 75.160 117.460 75.480 117.475 ;
        RECT 67.310 117.180 69.845 117.320 ;
        RECT 76.970 117.320 77.260 117.365 ;
        RECT 79.290 117.320 79.505 117.475 ;
        RECT 82.980 117.460 83.300 117.520 ;
        RECT 76.970 117.180 79.505 117.320 ;
        RECT 80.235 117.320 80.525 117.365 ;
        RECT 80.680 117.320 81.000 117.380 ;
        RECT 84.375 117.320 84.665 117.365 ;
        RECT 80.235 117.180 81.000 117.320 ;
        RECT 67.310 117.135 67.600 117.180 ;
        RECT 76.970 117.135 77.260 117.180 ;
        RECT 80.235 117.135 80.525 117.180 ;
        RECT 56.300 116.980 56.620 117.040 ;
        RECT 46.730 116.840 56.620 116.980 ;
        RECT 61.450 116.980 61.590 117.135 ;
        RECT 80.680 117.120 81.000 117.180 ;
        RECT 81.230 117.180 84.665 117.320 ;
        RECT 69.180 116.980 69.500 117.040 ;
        RECT 61.450 116.840 69.500 116.980 ;
        RECT 29.175 116.795 29.465 116.840 ;
        RECT 38.820 116.780 39.140 116.840 ;
        RECT 56.300 116.780 56.620 116.840 ;
        RECT 69.180 116.780 69.500 116.840 ;
        RECT 70.560 116.780 70.880 117.040 ;
        RECT 71.020 116.980 71.340 117.040 ;
        RECT 72.415 116.980 72.705 117.025 ;
        RECT 71.020 116.840 72.705 116.980 ;
        RECT 71.020 116.780 71.340 116.840 ;
        RECT 72.415 116.795 72.705 116.840 ;
        RECT 79.300 116.980 79.620 117.040 ;
        RECT 81.230 116.980 81.370 117.180 ;
        RECT 84.375 117.135 84.665 117.180 ;
        RECT 84.835 117.320 85.125 117.365 ;
        RECT 84.835 117.180 86.890 117.320 ;
        RECT 84.835 117.135 85.125 117.180 ;
        RECT 79.300 116.840 81.370 116.980 ;
        RECT 82.075 116.980 82.365 117.025 ;
        RECT 85.280 116.980 85.600 117.040 ;
        RECT 82.075 116.840 85.600 116.980 ;
        RECT 79.300 116.780 79.620 116.840 ;
        RECT 82.075 116.795 82.365 116.840 ;
        RECT 85.280 116.780 85.600 116.840 ;
        RECT 85.755 116.795 86.045 117.025 ;
        RECT 86.750 116.980 86.890 117.180 ;
        RECT 87.120 117.120 87.440 117.380 ;
        RECT 89.050 117.365 89.190 117.520 ;
        RECT 89.435 117.520 98.440 117.660 ;
        RECT 89.435 117.475 89.725 117.520 ;
        RECT 94.890 117.475 95.180 117.520 ;
        RECT 98.150 117.475 98.440 117.520 ;
        RECT 99.070 117.660 99.360 117.705 ;
        RECT 100.930 117.660 101.220 117.705 ;
        RECT 99.070 117.520 101.220 117.660 ;
        RECT 99.070 117.475 99.360 117.520 ;
        RECT 100.930 117.475 101.220 117.520 ;
        RECT 104.550 117.660 104.840 117.705 ;
        RECT 105.520 117.660 105.840 117.720 ;
        RECT 107.810 117.660 108.100 117.705 ;
        RECT 104.550 117.520 108.100 117.660 ;
        RECT 104.550 117.475 104.840 117.520 ;
        RECT 88.975 117.320 89.265 117.365 ;
        RECT 90.355 117.320 90.645 117.365 ;
        RECT 88.975 117.180 90.645 117.320 ;
        RECT 88.975 117.135 89.265 117.180 ;
        RECT 90.355 117.135 90.645 117.180 ;
        RECT 96.750 117.320 97.040 117.365 ;
        RECT 99.070 117.320 99.285 117.475 ;
        RECT 105.520 117.460 105.840 117.520 ;
        RECT 107.810 117.475 108.100 117.520 ;
        RECT 108.730 117.660 109.020 117.705 ;
        RECT 110.590 117.660 110.880 117.705 ;
        RECT 117.940 117.660 118.260 117.720 ;
        RECT 108.730 117.520 110.880 117.660 ;
        RECT 108.730 117.475 109.020 117.520 ;
        RECT 110.590 117.475 110.880 117.520 ;
        RECT 113.890 117.520 118.260 117.660 ;
        RECT 96.750 117.180 99.285 117.320 ;
        RECT 106.410 117.320 106.700 117.365 ;
        RECT 108.730 117.320 108.945 117.475 ;
        RECT 106.410 117.180 108.945 117.320 ;
        RECT 96.750 117.135 97.040 117.180 ;
        RECT 106.410 117.135 106.700 117.180 ;
        RECT 109.660 117.120 109.980 117.380 ;
        RECT 111.500 117.120 111.820 117.380 ;
        RECT 113.890 117.365 114.030 117.520 ;
        RECT 117.940 117.460 118.260 117.520 ;
        RECT 113.815 117.135 114.105 117.365 ;
        RECT 115.180 117.120 115.500 117.380 ;
        RECT 93.560 116.980 93.880 117.040 ;
        RECT 86.750 116.840 93.880 116.980 ;
        RECT 21.770 116.640 22.060 116.685 ;
        RECT 24.550 116.640 24.840 116.685 ;
        RECT 26.410 116.640 26.700 116.685 ;
        RECT 21.770 116.500 26.700 116.640 ;
        RECT 21.770 116.455 22.060 116.500 ;
        RECT 24.550 116.455 24.840 116.500 ;
        RECT 26.410 116.455 26.700 116.500 ;
        RECT 27.800 116.640 28.090 116.685 ;
        RECT 29.660 116.640 29.950 116.685 ;
        RECT 32.440 116.640 32.730 116.685 ;
        RECT 27.800 116.500 32.730 116.640 ;
        RECT 27.800 116.455 28.090 116.500 ;
        RECT 29.660 116.455 29.950 116.500 ;
        RECT 32.440 116.455 32.730 116.500 ;
        RECT 41.550 116.640 41.840 116.685 ;
        RECT 44.330 116.640 44.620 116.685 ;
        RECT 46.190 116.640 46.480 116.685 ;
        RECT 41.550 116.500 46.480 116.640 ;
        RECT 41.550 116.455 41.840 116.500 ;
        RECT 44.330 116.455 44.620 116.500 ;
        RECT 46.190 116.455 46.480 116.500 ;
        RECT 51.210 116.640 51.500 116.685 ;
        RECT 53.990 116.640 54.280 116.685 ;
        RECT 55.850 116.640 56.140 116.685 ;
        RECT 51.210 116.500 56.140 116.640 ;
        RECT 51.210 116.455 51.500 116.500 ;
        RECT 53.990 116.455 54.280 116.500 ;
        RECT 55.850 116.455 56.140 116.500 ;
        RECT 67.310 116.640 67.600 116.685 ;
        RECT 70.090 116.640 70.380 116.685 ;
        RECT 71.950 116.640 72.240 116.685 ;
        RECT 67.310 116.500 72.240 116.640 ;
        RECT 67.310 116.455 67.600 116.500 ;
        RECT 70.090 116.455 70.380 116.500 ;
        RECT 71.950 116.455 72.240 116.500 ;
        RECT 76.970 116.640 77.260 116.685 ;
        RECT 79.750 116.640 80.040 116.685 ;
        RECT 81.610 116.640 81.900 116.685 ;
        RECT 76.970 116.500 81.900 116.640 ;
        RECT 76.970 116.455 77.260 116.500 ;
        RECT 79.750 116.455 80.040 116.500 ;
        RECT 81.610 116.455 81.900 116.500 ;
        RECT 83.440 116.640 83.760 116.700 ;
        RECT 85.830 116.640 85.970 116.795 ;
        RECT 93.560 116.780 93.880 116.840 ;
        RECT 100.000 116.780 100.320 117.040 ;
        RECT 101.855 116.980 102.145 117.025 ;
        RECT 111.590 116.980 111.730 117.120 ;
        RECT 101.855 116.840 111.730 116.980 ;
        RECT 101.855 116.795 102.145 116.840 ;
        RECT 83.440 116.500 85.970 116.640 ;
        RECT 96.750 116.640 97.040 116.685 ;
        RECT 99.530 116.640 99.820 116.685 ;
        RECT 101.390 116.640 101.680 116.685 ;
        RECT 96.750 116.500 101.680 116.640 ;
        RECT 83.440 116.440 83.760 116.500 ;
        RECT 96.750 116.455 97.040 116.500 ;
        RECT 99.530 116.455 99.820 116.500 ;
        RECT 101.390 116.455 101.680 116.500 ;
        RECT 106.410 116.640 106.700 116.685 ;
        RECT 109.190 116.640 109.480 116.685 ;
        RECT 111.050 116.640 111.340 116.685 ;
        RECT 106.410 116.500 111.340 116.640 ;
        RECT 106.410 116.455 106.700 116.500 ;
        RECT 109.190 116.455 109.480 116.500 ;
        RECT 111.050 116.455 111.340 116.500 ;
        RECT 16.755 116.300 17.045 116.345 ;
        RECT 28.240 116.300 28.560 116.360 ;
        RECT 16.755 116.160 28.560 116.300 ;
        RECT 16.755 116.115 17.045 116.160 ;
        RECT 28.240 116.100 28.560 116.160 ;
        RECT 45.720 116.300 46.040 116.360 ;
        RECT 47.345 116.300 47.635 116.345 ;
        RECT 45.720 116.160 47.635 116.300 ;
        RECT 45.720 116.100 46.040 116.160 ;
        RECT 47.345 116.115 47.635 116.160 ;
        RECT 88.040 116.100 88.360 116.360 ;
        RECT 90.800 116.100 91.120 116.360 ;
        RECT 14.370 115.480 127.530 115.960 ;
        RECT 22.735 115.280 23.025 115.325 ;
        RECT 23.180 115.280 23.500 115.340 ;
        RECT 22.735 115.140 23.500 115.280 ;
        RECT 22.735 115.095 23.025 115.140 ;
        RECT 23.180 115.080 23.500 115.140 ;
        RECT 30.540 115.280 30.860 115.340 ;
        RECT 33.545 115.280 33.835 115.325 ;
        RECT 30.540 115.140 33.835 115.280 ;
        RECT 30.540 115.080 30.860 115.140 ;
        RECT 33.545 115.095 33.835 115.140 ;
        RECT 35.140 115.080 35.460 115.340 ;
        RECT 37.440 115.080 37.760 115.340 ;
        RECT 38.820 115.080 39.140 115.340 ;
        RECT 42.960 115.280 43.280 115.340 ;
        RECT 44.355 115.280 44.645 115.325 ;
        RECT 42.960 115.140 44.645 115.280 ;
        RECT 42.960 115.080 43.280 115.140 ;
        RECT 44.355 115.095 44.645 115.140 ;
        RECT 45.260 115.080 45.580 115.340 ;
        RECT 53.095 115.280 53.385 115.325 ;
        RECT 54.460 115.280 54.780 115.340 ;
        RECT 53.095 115.140 54.780 115.280 ;
        RECT 53.095 115.095 53.385 115.140 ;
        RECT 54.460 115.080 54.780 115.140 ;
        RECT 66.420 115.080 66.740 115.340 ;
        RECT 68.735 115.280 69.025 115.325 ;
        RECT 70.560 115.280 70.880 115.340 ;
        RECT 68.735 115.140 70.880 115.280 ;
        RECT 68.735 115.095 69.025 115.140 ;
        RECT 70.560 115.080 70.880 115.140 ;
        RECT 71.020 115.280 71.340 115.340 ;
        RECT 73.320 115.280 73.640 115.340 ;
        RECT 71.020 115.140 73.640 115.280 ;
        RECT 71.020 115.080 71.340 115.140 ;
        RECT 73.320 115.080 73.640 115.140 ;
        RECT 77.245 115.280 77.535 115.325 ;
        RECT 79.300 115.280 79.620 115.340 ;
        RECT 77.245 115.140 79.620 115.280 ;
        RECT 77.245 115.095 77.535 115.140 ;
        RECT 79.300 115.080 79.620 115.140 ;
        RECT 93.560 115.280 93.880 115.340 ;
        RECT 96.105 115.280 96.395 115.325 ;
        RECT 93.560 115.140 96.395 115.280 ;
        RECT 93.560 115.080 93.880 115.140 ;
        RECT 96.105 115.095 96.395 115.140 ;
        RECT 100.000 115.080 100.320 115.340 ;
        RECT 108.755 115.280 109.045 115.325 ;
        RECT 109.660 115.280 109.980 115.340 ;
        RECT 108.755 115.140 109.980 115.280 ;
        RECT 108.755 115.095 109.045 115.140 ;
        RECT 109.660 115.080 109.980 115.140 ;
        RECT 114.735 115.280 115.025 115.325 ;
        RECT 115.180 115.280 115.500 115.340 ;
        RECT 114.735 115.140 115.500 115.280 ;
        RECT 114.735 115.095 115.025 115.140 ;
        RECT 115.180 115.080 115.500 115.140 ;
        RECT 21.815 114.755 22.105 114.985 ;
        RECT 25.040 114.940 25.330 114.985 ;
        RECT 26.900 114.940 27.190 114.985 ;
        RECT 29.680 114.940 29.970 114.985 ;
        RECT 25.040 114.800 29.970 114.940 ;
        RECT 25.040 114.755 25.330 114.800 ;
        RECT 26.900 114.755 27.190 114.800 ;
        RECT 29.680 114.755 29.970 114.800 ;
        RECT 43.420 114.940 43.740 115.000 ;
        RECT 81.110 114.940 81.400 114.985 ;
        RECT 83.890 114.940 84.180 114.985 ;
        RECT 85.750 114.940 86.040 114.985 ;
        RECT 43.420 114.800 48.250 114.940 ;
        RECT 19.500 114.600 19.820 114.660 ;
        RECT 21.890 114.600 22.030 114.755 ;
        RECT 43.420 114.740 43.740 114.800 ;
        RECT 24.575 114.600 24.865 114.645 ;
        RECT 25.480 114.600 25.800 114.660 ;
        RECT 45.720 114.600 46.040 114.660 ;
        RECT 48.110 114.645 48.250 114.800 ;
        RECT 81.110 114.800 86.040 114.940 ;
        RECT 81.110 114.755 81.400 114.800 ;
        RECT 83.890 114.755 84.180 114.800 ;
        RECT 85.750 114.755 86.040 114.800 ;
        RECT 87.600 114.940 87.890 114.985 ;
        RECT 89.460 114.940 89.750 114.985 ;
        RECT 92.240 114.940 92.530 114.985 ;
        RECT 112.880 114.940 113.200 115.000 ;
        RECT 87.600 114.800 92.530 114.940 ;
        RECT 87.600 114.755 87.890 114.800 ;
        RECT 89.460 114.755 89.750 114.800 ;
        RECT 92.240 114.755 92.530 114.800 ;
        RECT 112.050 114.800 113.200 114.940 ;
        RECT 47.575 114.600 47.865 114.645 ;
        RECT 19.500 114.460 21.570 114.600 ;
        RECT 21.890 114.460 24.330 114.600 ;
        RECT 19.500 114.400 19.820 114.460 ;
        RECT 20.880 114.060 21.200 114.320 ;
        RECT 21.430 114.260 21.570 114.460 ;
        RECT 23.195 114.260 23.485 114.305 ;
        RECT 24.190 114.260 24.330 114.460 ;
        RECT 24.575 114.460 25.800 114.600 ;
        RECT 24.575 114.415 24.865 114.460 ;
        RECT 25.480 114.400 25.800 114.460 ;
        RECT 35.690 114.460 45.030 114.600 ;
        RECT 35.690 114.320 35.830 114.460 ;
        RECT 26.415 114.260 26.705 114.305 ;
        RECT 29.680 114.260 29.970 114.305 ;
        RECT 21.430 114.120 23.870 114.260 ;
        RECT 24.190 114.120 26.705 114.260 ;
        RECT 23.195 114.075 23.485 114.120 ;
        RECT 23.730 113.580 23.870 114.120 ;
        RECT 26.415 114.075 26.705 114.120 ;
        RECT 27.435 114.120 29.970 114.260 ;
        RECT 27.435 113.965 27.650 114.120 ;
        RECT 29.680 114.075 29.970 114.120 ;
        RECT 35.600 114.060 35.920 114.320 ;
        RECT 36.520 114.060 36.840 114.320 ;
        RECT 39.740 114.060 40.060 114.320 ;
        RECT 44.890 114.305 45.030 114.460 ;
        RECT 45.720 114.460 47.865 114.600 ;
        RECT 45.720 114.400 46.040 114.460 ;
        RECT 47.575 114.415 47.865 114.460 ;
        RECT 48.035 114.415 48.325 114.645 ;
        RECT 49.860 114.600 50.180 114.660 ;
        RECT 69.180 114.600 69.500 114.660 ;
        RECT 49.030 114.460 50.180 114.600 ;
        RECT 44.815 114.260 45.105 114.305 ;
        RECT 49.030 114.260 49.170 114.460 ;
        RECT 49.860 114.400 50.180 114.460 ;
        RECT 66.050 114.460 69.500 114.600 ;
        RECT 44.815 114.120 49.170 114.260 ;
        RECT 49.400 114.260 49.720 114.320 ;
        RECT 66.050 114.305 66.190 114.460 ;
        RECT 69.180 114.400 69.500 114.460 ;
        RECT 84.360 114.400 84.680 114.660 ;
        RECT 85.280 114.600 85.600 114.660 ;
        RECT 86.200 114.600 86.520 114.660 ;
        RECT 87.135 114.600 87.425 114.645 ;
        RECT 85.280 114.460 87.425 114.600 ;
        RECT 85.280 114.400 85.600 114.460 ;
        RECT 86.200 114.400 86.520 114.460 ;
        RECT 87.135 114.415 87.425 114.460 ;
        RECT 88.040 114.600 88.360 114.660 ;
        RECT 112.050 114.645 112.190 114.800 ;
        RECT 112.880 114.740 113.200 114.800 ;
        RECT 88.975 114.600 89.265 114.645 ;
        RECT 88.040 114.460 89.265 114.600 ;
        RECT 88.040 114.400 88.360 114.460 ;
        RECT 88.975 114.415 89.265 114.460 ;
        RECT 111.975 114.415 112.265 114.645 ;
        RECT 112.420 114.400 112.740 114.660 ;
        RECT 52.175 114.260 52.465 114.305 ;
        RECT 49.400 114.120 52.465 114.260 ;
        RECT 44.815 114.075 45.105 114.120 ;
        RECT 49.400 114.060 49.720 114.120 ;
        RECT 52.175 114.075 52.465 114.120 ;
        RECT 65.975 114.075 66.265 114.305 ;
        RECT 67.800 114.060 68.120 114.320 ;
        RECT 81.110 114.260 81.400 114.305 ;
        RECT 92.240 114.260 92.530 114.305 ;
        RECT 81.110 114.120 83.645 114.260 ;
        RECT 81.110 114.075 81.400 114.120 ;
        RECT 25.500 113.920 25.790 113.965 ;
        RECT 27.360 113.920 27.650 113.965 ;
        RECT 25.500 113.780 27.650 113.920 ;
        RECT 25.500 113.735 25.790 113.780 ;
        RECT 27.360 113.735 27.650 113.780 ;
        RECT 28.240 113.965 28.560 113.980 ;
        RECT 28.240 113.920 28.570 113.965 ;
        RECT 31.540 113.920 31.830 113.965 ;
        RECT 28.240 113.780 31.830 113.920 ;
        RECT 28.240 113.735 28.570 113.780 ;
        RECT 31.540 113.735 31.830 113.780 ;
        RECT 42.040 113.920 42.360 113.980 ;
        RECT 82.520 113.965 82.840 113.980 ;
        RECT 47.115 113.920 47.405 113.965 ;
        RECT 42.040 113.780 47.405 113.920 ;
        RECT 28.240 113.720 28.560 113.735 ;
        RECT 42.040 113.720 42.360 113.780 ;
        RECT 47.115 113.735 47.405 113.780 ;
        RECT 79.250 113.920 79.540 113.965 ;
        RECT 82.510 113.920 82.840 113.965 ;
        RECT 79.250 113.780 82.840 113.920 ;
        RECT 79.250 113.735 79.540 113.780 ;
        RECT 82.510 113.735 82.840 113.780 ;
        RECT 83.430 113.965 83.645 114.120 ;
        RECT 89.995 114.120 92.530 114.260 ;
        RECT 89.995 113.965 90.210 114.120 ;
        RECT 92.240 114.075 92.530 114.120 ;
        RECT 100.920 114.060 101.240 114.320 ;
        RECT 107.835 114.260 108.125 114.305 ;
        RECT 108.740 114.260 109.060 114.320 ;
        RECT 107.835 114.120 109.060 114.260 ;
        RECT 107.835 114.075 108.125 114.120 ;
        RECT 108.740 114.060 109.060 114.120 ;
        RECT 109.200 114.260 109.520 114.320 ;
        RECT 112.895 114.260 113.185 114.305 ;
        RECT 109.200 114.120 113.185 114.260 ;
        RECT 109.200 114.060 109.520 114.120 ;
        RECT 112.895 114.075 113.185 114.120 ;
        RECT 83.430 113.920 83.720 113.965 ;
        RECT 85.290 113.920 85.580 113.965 ;
        RECT 83.430 113.780 85.580 113.920 ;
        RECT 83.430 113.735 83.720 113.780 ;
        RECT 85.290 113.735 85.580 113.780 ;
        RECT 88.060 113.920 88.350 113.965 ;
        RECT 89.920 113.920 90.210 113.965 ;
        RECT 88.060 113.780 90.210 113.920 ;
        RECT 88.060 113.735 88.350 113.780 ;
        RECT 89.920 113.735 90.210 113.780 ;
        RECT 90.800 113.965 91.120 113.980 ;
        RECT 90.800 113.920 91.130 113.965 ;
        RECT 94.100 113.920 94.390 113.965 ;
        RECT 90.800 113.780 94.390 113.920 ;
        RECT 90.800 113.735 91.130 113.780 ;
        RECT 94.100 113.735 94.390 113.780 ;
        RECT 82.520 113.720 82.840 113.735 ;
        RECT 90.800 113.720 91.120 113.735 ;
        RECT 35.600 113.580 35.920 113.640 ;
        RECT 23.730 113.440 35.920 113.580 ;
        RECT 35.600 113.380 35.920 113.440 ;
        RECT 101.380 113.580 101.700 113.640 ;
        RECT 121.620 113.580 121.940 113.640 ;
        RECT 101.380 113.440 121.940 113.580 ;
        RECT 101.380 113.380 101.700 113.440 ;
        RECT 121.620 113.380 121.940 113.440 ;
        RECT 14.370 112.760 127.530 113.240 ;
        RECT 34.235 112.560 34.525 112.605 ;
        RECT 34.680 112.560 35.000 112.620 ;
        RECT 34.235 112.420 35.000 112.560 ;
        RECT 34.235 112.375 34.525 112.420 ;
        RECT 34.680 112.360 35.000 112.420 ;
        RECT 102.775 112.560 103.065 112.605 ;
        RECT 111.500 112.560 111.820 112.620 ;
        RECT 102.775 112.420 111.820 112.560 ;
        RECT 102.775 112.375 103.065 112.420 ;
        RECT 18.695 112.220 18.985 112.265 ;
        RECT 20.880 112.220 21.200 112.280 ;
        RECT 21.935 112.220 22.585 112.265 ;
        RECT 18.695 112.080 22.585 112.220 ;
        RECT 18.695 112.035 19.285 112.080 ;
        RECT 18.995 111.720 19.285 112.035 ;
        RECT 20.880 112.020 21.200 112.080 ;
        RECT 21.935 112.035 22.585 112.080 ;
        RECT 46.655 112.220 46.945 112.265 ;
        RECT 48.940 112.220 49.260 112.280 ;
        RECT 46.655 112.080 49.260 112.220 ;
        RECT 46.655 112.035 46.945 112.080 ;
        RECT 48.940 112.020 49.260 112.080 ;
        RECT 92.640 112.020 92.960 112.280 ;
        RECT 101.395 112.220 101.685 112.265 ;
        RECT 102.850 112.220 102.990 112.375 ;
        RECT 111.500 112.360 111.820 112.420 ;
        RECT 117.020 112.560 117.340 112.620 ;
        RECT 120.715 112.560 121.005 112.605 ;
        RECT 117.020 112.420 121.005 112.560 ;
        RECT 117.020 112.360 117.340 112.420 ;
        RECT 120.715 112.375 121.005 112.420 ;
        RECT 122.095 112.375 122.385 112.605 ;
        RECT 101.395 112.080 102.990 112.220 ;
        RECT 118.860 112.220 119.180 112.280 ;
        RECT 122.170 112.220 122.310 112.375 ;
        RECT 118.860 112.080 122.310 112.220 ;
        RECT 101.395 112.035 101.685 112.080 ;
        RECT 118.860 112.020 119.180 112.080 ;
        RECT 20.075 111.880 20.365 111.925 ;
        RECT 23.655 111.880 23.945 111.925 ;
        RECT 25.490 111.880 25.780 111.925 ;
        RECT 20.075 111.740 25.780 111.880 ;
        RECT 20.075 111.695 20.365 111.740 ;
        RECT 23.655 111.695 23.945 111.740 ;
        RECT 25.490 111.695 25.780 111.740 ;
        RECT 25.940 111.680 26.260 111.940 ;
        RECT 34.695 111.880 34.985 111.925 ;
        RECT 35.600 111.880 35.920 111.940 ;
        RECT 34.695 111.740 35.920 111.880 ;
        RECT 34.695 111.695 34.985 111.740 ;
        RECT 35.600 111.680 35.920 111.740 ;
        RECT 77.920 111.880 78.240 111.940 ;
        RECT 81.140 111.880 81.460 111.940 ;
        RECT 77.920 111.740 81.460 111.880 ;
        RECT 77.920 111.680 78.240 111.740 ;
        RECT 81.140 111.680 81.460 111.740 ;
        RECT 119.320 111.680 119.640 111.940 ;
        RECT 121.620 111.680 121.940 111.940 ;
        RECT 123.015 111.695 123.305 111.925 ;
        RECT 13.980 111.540 14.300 111.600 ;
        RECT 15.835 111.540 16.125 111.585 ;
        RECT 13.980 111.400 16.125 111.540 ;
        RECT 13.980 111.340 14.300 111.400 ;
        RECT 15.835 111.355 16.125 111.400 ;
        RECT 20.075 111.200 20.365 111.245 ;
        RECT 23.195 111.200 23.485 111.245 ;
        RECT 25.085 111.200 25.375 111.245 ;
        RECT 20.075 111.060 25.375 111.200 ;
        RECT 26.030 111.200 26.170 111.680 ;
        RECT 50.320 111.540 50.640 111.600 ;
        RECT 43.050 111.400 50.640 111.540 ;
        RECT 36.520 111.200 36.840 111.260 ;
        RECT 40.215 111.200 40.505 111.245 ;
        RECT 43.050 111.200 43.190 111.400 ;
        RECT 50.320 111.340 50.640 111.400 ;
        RECT 80.695 111.540 80.985 111.585 ;
        RECT 81.600 111.540 81.920 111.600 ;
        RECT 80.695 111.400 81.920 111.540 ;
        RECT 80.695 111.355 80.985 111.400 ;
        RECT 81.600 111.340 81.920 111.400 ;
        RECT 104.140 111.540 104.460 111.600 ;
        RECT 104.140 111.400 119.550 111.540 ;
        RECT 104.140 111.340 104.460 111.400 ;
        RECT 26.030 111.060 43.190 111.200 ;
        RECT 119.410 111.200 119.550 111.400 ;
        RECT 119.780 111.340 120.100 111.600 ;
        RECT 123.090 111.540 123.230 111.695 ;
        RECT 120.330 111.400 123.230 111.540 ;
        RECT 120.330 111.200 120.470 111.400 ;
        RECT 119.410 111.060 120.470 111.200 ;
        RECT 20.075 111.015 20.365 111.060 ;
        RECT 23.195 111.015 23.485 111.060 ;
        RECT 25.085 111.015 25.375 111.060 ;
        RECT 36.520 111.000 36.840 111.060 ;
        RECT 40.215 111.015 40.505 111.060 ;
        RECT 24.670 110.860 24.960 110.905 ;
        RECT 27.320 110.860 27.640 110.920 ;
        RECT 24.670 110.720 27.640 110.860 ;
        RECT 24.670 110.675 24.960 110.720 ;
        RECT 27.320 110.660 27.640 110.720 ;
        RECT 14.370 110.040 127.530 110.520 ;
        RECT 20.880 109.640 21.200 109.900 ;
        RECT 27.320 109.640 27.640 109.900 ;
        RECT 73.780 109.840 74.100 109.900 ;
        RECT 77.935 109.840 78.225 109.885 ;
        RECT 73.780 109.700 78.225 109.840 ;
        RECT 73.780 109.640 74.100 109.700 ;
        RECT 77.935 109.655 78.225 109.700 ;
        RECT 106.915 109.500 107.205 109.545 ;
        RECT 110.580 109.500 110.900 109.560 ;
        RECT 106.915 109.360 110.900 109.500 ;
        RECT 106.915 109.315 107.205 109.360 ;
        RECT 110.580 109.300 110.900 109.360 ;
        RECT 111.500 109.300 111.820 109.560 ;
        RECT 116.525 109.500 116.815 109.545 ;
        RECT 118.415 109.500 118.705 109.545 ;
        RECT 121.535 109.500 121.825 109.545 ;
        RECT 116.525 109.360 121.825 109.500 ;
        RECT 116.525 109.315 116.815 109.360 ;
        RECT 118.415 109.315 118.705 109.360 ;
        RECT 121.535 109.315 121.825 109.360 ;
        RECT 31.000 109.160 31.320 109.220 ;
        RECT 81.140 109.160 81.460 109.220 ;
        RECT 111.590 109.160 111.730 109.300 ;
        RECT 115.655 109.160 115.945 109.205 ;
        RECT 31.000 109.020 33.070 109.160 ;
        RECT 31.000 108.960 31.320 109.020 ;
        RECT 21.355 108.820 21.645 108.865 ;
        RECT 23.655 108.820 23.945 108.865 ;
        RECT 21.355 108.680 23.945 108.820 ;
        RECT 21.355 108.635 21.645 108.680 ;
        RECT 23.655 108.635 23.945 108.680 ;
        RECT 28.255 108.820 28.545 108.865 ;
        RECT 29.160 108.820 29.480 108.880 ;
        RECT 32.930 108.865 33.070 109.020 ;
        RECT 59.610 109.020 79.530 109.160 ;
        RECT 59.610 108.880 59.750 109.020 ;
        RECT 28.255 108.680 29.480 108.820 ;
        RECT 28.255 108.635 28.545 108.680 ;
        RECT 23.730 108.480 23.870 108.635 ;
        RECT 29.160 108.620 29.480 108.680 ;
        RECT 31.475 108.635 31.765 108.865 ;
        RECT 32.855 108.635 33.145 108.865 ;
        RECT 34.220 108.820 34.540 108.880 ;
        RECT 35.155 108.820 35.445 108.865 ;
        RECT 34.220 108.680 35.445 108.820 ;
        RECT 27.320 108.480 27.640 108.540 ;
        RECT 31.550 108.480 31.690 108.635 ;
        RECT 34.220 108.620 34.540 108.680 ;
        RECT 35.155 108.635 35.445 108.680 ;
        RECT 50.795 108.820 51.085 108.865 ;
        RECT 51.700 108.820 52.020 108.880 ;
        RECT 50.795 108.680 52.020 108.820 ;
        RECT 50.795 108.635 51.085 108.680 ;
        RECT 51.700 108.620 52.020 108.680 ;
        RECT 56.760 108.620 57.080 108.880 ;
        RECT 59.520 108.620 59.840 108.880 ;
        RECT 59.980 108.820 60.300 108.880 ;
        RECT 60.915 108.820 61.205 108.865 ;
        RECT 64.595 108.820 64.885 108.865 ;
        RECT 59.980 108.680 64.885 108.820 ;
        RECT 59.980 108.620 60.300 108.680 ;
        RECT 60.915 108.635 61.205 108.680 ;
        RECT 64.595 108.635 64.885 108.680 ;
        RECT 68.275 108.820 68.565 108.865 ;
        RECT 68.720 108.820 69.040 108.880 ;
        RECT 68.275 108.680 69.040 108.820 ;
        RECT 68.275 108.635 68.565 108.680 ;
        RECT 68.720 108.620 69.040 108.680 ;
        RECT 77.015 108.820 77.305 108.865 ;
        RECT 77.920 108.820 78.240 108.880 ;
        RECT 77.015 108.680 78.240 108.820 ;
        RECT 77.015 108.635 77.305 108.680 ;
        RECT 77.920 108.620 78.240 108.680 ;
        RECT 78.395 108.820 78.685 108.865 ;
        RECT 78.840 108.820 79.160 108.880 ;
        RECT 78.395 108.680 79.160 108.820 ;
        RECT 79.390 108.820 79.530 109.020 ;
        RECT 81.140 109.020 87.350 109.160 ;
        RECT 111.590 109.020 115.945 109.160 ;
        RECT 81.140 108.960 81.460 109.020 ;
        RECT 87.210 108.865 87.350 109.020 ;
        RECT 115.655 108.975 115.945 109.020 ;
        RECT 117.035 109.160 117.325 109.205 ;
        RECT 118.860 109.160 119.180 109.220 ;
        RECT 117.035 109.020 119.180 109.160 ;
        RECT 117.035 108.975 117.325 109.020 ;
        RECT 118.860 108.960 119.180 109.020 ;
        RECT 79.775 108.820 80.065 108.865 ;
        RECT 79.390 108.680 80.065 108.820 ;
        RECT 78.395 108.635 78.685 108.680 ;
        RECT 78.840 108.620 79.160 108.680 ;
        RECT 79.775 108.635 80.065 108.680 ;
        RECT 82.535 108.635 82.825 108.865 ;
        RECT 87.135 108.820 87.425 108.865 ;
        RECT 92.195 108.820 92.485 108.865 ;
        RECT 87.135 108.680 92.485 108.820 ;
        RECT 87.135 108.635 87.425 108.680 ;
        RECT 92.195 108.635 92.485 108.680 ;
        RECT 93.575 108.820 93.865 108.865 ;
        RECT 94.480 108.820 94.800 108.880 ;
        RECT 93.575 108.680 94.800 108.820 ;
        RECT 93.575 108.635 93.865 108.680 ;
        RECT 40.660 108.480 40.980 108.540 ;
        RECT 23.730 108.340 40.980 108.480 ;
        RECT 27.320 108.280 27.640 108.340 ;
        RECT 40.660 108.280 40.980 108.340 ;
        RECT 75.620 108.480 75.940 108.540 ;
        RECT 82.610 108.480 82.750 108.635 ;
        RECT 75.620 108.340 82.750 108.480 ;
        RECT 92.270 108.480 92.410 108.635 ;
        RECT 94.480 108.620 94.800 108.680 ;
        RECT 99.540 108.820 99.860 108.880 ;
        RECT 100.935 108.820 101.225 108.865 ;
        RECT 99.540 108.680 101.225 108.820 ;
        RECT 99.540 108.620 99.860 108.680 ;
        RECT 100.935 108.635 101.225 108.680 ;
        RECT 103.220 108.820 103.540 108.880 ;
        RECT 105.995 108.820 106.285 108.865 ;
        RECT 103.220 108.680 106.285 108.820 ;
        RECT 103.220 108.620 103.540 108.680 ;
        RECT 105.995 108.635 106.285 108.680 ;
        RECT 109.675 108.635 109.965 108.865 ;
        RECT 102.300 108.480 102.620 108.540 ;
        RECT 109.750 108.480 109.890 108.635 ;
        RECT 110.120 108.620 110.440 108.880 ;
        RECT 111.040 108.820 111.360 108.880 ;
        RECT 111.515 108.820 111.805 108.865 ;
        RECT 111.040 108.680 111.805 108.820 ;
        RECT 111.040 108.620 111.360 108.680 ;
        RECT 111.515 108.635 111.805 108.680 ;
        RECT 114.275 108.635 114.565 108.865 ;
        RECT 116.120 108.820 116.410 108.865 ;
        RECT 117.955 108.820 118.245 108.865 ;
        RECT 121.535 108.820 121.825 108.865 ;
        RECT 116.120 108.680 121.825 108.820 ;
        RECT 116.120 108.635 116.410 108.680 ;
        RECT 117.955 108.635 118.245 108.680 ;
        RECT 121.535 108.635 121.825 108.680 ;
        RECT 114.350 108.480 114.490 108.635 ;
        RECT 119.780 108.525 120.100 108.540 ;
        RECT 119.315 108.480 120.100 108.525 ;
        RECT 122.615 108.525 122.905 108.840 ;
        RECT 122.615 108.480 123.205 108.525 ;
        RECT 92.270 108.340 119.090 108.480 ;
        RECT 75.620 108.280 75.940 108.340 ;
        RECT 102.300 108.280 102.620 108.340 ;
        RECT 118.950 108.200 119.090 108.340 ;
        RECT 119.315 108.340 123.205 108.480 ;
        RECT 119.315 108.295 120.100 108.340 ;
        RECT 122.915 108.295 123.205 108.340 ;
        RECT 125.775 108.480 126.065 108.525 ;
        RECT 127.600 108.480 127.920 108.540 ;
        RECT 125.775 108.340 127.920 108.480 ;
        RECT 125.775 108.295 126.065 108.340 ;
        RECT 119.780 108.280 120.100 108.295 ;
        RECT 127.600 108.280 127.920 108.340 ;
        RECT 23.180 107.940 23.500 108.200 ;
        RECT 31.015 108.140 31.305 108.185 ;
        RECT 31.460 108.140 31.780 108.200 ;
        RECT 31.015 108.000 31.780 108.140 ;
        RECT 31.015 107.955 31.305 108.000 ;
        RECT 31.460 107.940 31.780 108.000 ;
        RECT 31.920 107.940 32.240 108.200 ;
        RECT 33.760 108.140 34.080 108.200 ;
        RECT 34.235 108.140 34.525 108.185 ;
        RECT 33.760 108.000 34.525 108.140 ;
        RECT 33.760 107.940 34.080 108.000 ;
        RECT 34.235 107.955 34.525 108.000 ;
        RECT 51.715 108.140 52.005 108.185 ;
        RECT 55.380 108.140 55.700 108.200 ;
        RECT 51.715 108.000 55.700 108.140 ;
        RECT 51.715 107.955 52.005 108.000 ;
        RECT 55.380 107.940 55.700 108.000 ;
        RECT 57.680 107.940 58.000 108.200 ;
        RECT 65.040 107.940 65.360 108.200 ;
        RECT 69.195 108.140 69.485 108.185 ;
        RECT 71.940 108.140 72.260 108.200 ;
        RECT 69.195 108.000 72.260 108.140 ;
        RECT 69.195 107.955 69.485 108.000 ;
        RECT 71.940 107.940 72.260 108.000 ;
        RECT 76.555 108.140 76.845 108.185 ;
        RECT 79.300 108.140 79.620 108.200 ;
        RECT 76.555 108.000 79.620 108.140 ;
        RECT 76.555 107.955 76.845 108.000 ;
        RECT 79.300 107.940 79.620 108.000 ;
        RECT 83.440 107.940 83.760 108.200 ;
        RECT 87.580 107.940 87.900 108.200 ;
        RECT 92.640 107.940 92.960 108.200 ;
        RECT 94.495 108.140 94.785 108.185 ;
        RECT 97.700 108.140 98.020 108.200 ;
        RECT 94.495 108.000 98.020 108.140 ;
        RECT 94.495 107.955 94.785 108.000 ;
        RECT 97.700 107.940 98.020 108.000 ;
        RECT 99.540 108.140 99.860 108.200 ;
        RECT 100.015 108.140 100.305 108.185 ;
        RECT 99.540 108.000 100.305 108.140 ;
        RECT 99.540 107.940 99.860 108.000 ;
        RECT 100.015 107.955 100.305 108.000 ;
        RECT 109.200 107.940 109.520 108.200 ;
        RECT 111.040 107.940 111.360 108.200 ;
        RECT 112.435 108.140 112.725 108.185 ;
        RECT 113.800 108.140 114.120 108.200 ;
        RECT 112.435 108.000 114.120 108.140 ;
        RECT 112.435 107.955 112.725 108.000 ;
        RECT 113.800 107.940 114.120 108.000 ;
        RECT 114.735 108.140 115.025 108.185 ;
        RECT 116.100 108.140 116.420 108.200 ;
        RECT 114.735 108.000 116.420 108.140 ;
        RECT 114.735 107.955 115.025 108.000 ;
        RECT 116.100 107.940 116.420 108.000 ;
        RECT 118.860 107.940 119.180 108.200 ;
        RECT 14.370 107.320 127.530 107.800 ;
        RECT 31.920 107.120 32.240 107.180 ;
        RECT 24.650 106.980 32.240 107.120 ;
        RECT 18.695 106.780 18.985 106.825 ;
        RECT 21.935 106.780 22.585 106.825 ;
        RECT 23.180 106.780 23.500 106.840 ;
        RECT 24.650 106.825 24.790 106.980 ;
        RECT 31.920 106.920 32.240 106.980 ;
        RECT 37.455 106.935 37.745 107.165 ;
        RECT 93.560 107.120 93.880 107.180 ;
        RECT 108.740 107.120 109.060 107.180 ;
        RECT 89.050 106.980 93.880 107.120 ;
        RECT 18.695 106.640 23.500 106.780 ;
        RECT 18.695 106.595 19.285 106.640 ;
        RECT 21.935 106.595 22.585 106.640 ;
        RECT 18.995 106.280 19.285 106.595 ;
        RECT 23.180 106.580 23.500 106.640 ;
        RECT 24.575 106.595 24.865 106.825 ;
        RECT 29.275 106.780 29.565 106.825 ;
        RECT 31.460 106.780 31.780 106.840 ;
        RECT 32.515 106.780 33.165 106.825 ;
        RECT 29.275 106.640 33.165 106.780 ;
        RECT 29.275 106.595 29.865 106.640 ;
        RECT 20.075 106.440 20.365 106.485 ;
        RECT 23.655 106.440 23.945 106.485 ;
        RECT 25.490 106.440 25.780 106.485 ;
        RECT 20.075 106.300 25.780 106.440 ;
        RECT 20.075 106.255 20.365 106.300 ;
        RECT 23.655 106.255 23.945 106.300 ;
        RECT 25.490 106.255 25.780 106.300 ;
        RECT 26.415 106.440 26.705 106.485 ;
        RECT 26.415 106.300 29.390 106.440 ;
        RECT 26.415 106.255 26.705 106.300 ;
        RECT 15.835 106.100 16.125 106.145 ;
        RECT 18.580 106.100 18.900 106.160 ;
        RECT 15.835 105.960 18.900 106.100 ;
        RECT 15.835 105.915 16.125 105.960 ;
        RECT 18.580 105.900 18.900 105.960 ;
        RECT 25.955 106.100 26.245 106.145 ;
        RECT 28.700 106.100 29.020 106.160 ;
        RECT 25.955 105.960 29.020 106.100 ;
        RECT 29.250 106.100 29.390 106.300 ;
        RECT 29.575 106.280 29.865 106.595 ;
        RECT 31.460 106.580 31.780 106.640 ;
        RECT 32.515 106.595 33.165 106.640 ;
        RECT 35.155 106.780 35.445 106.825 ;
        RECT 37.530 106.780 37.670 106.935 ;
        RECT 35.155 106.640 37.670 106.780 ;
        RECT 40.660 106.780 40.980 106.840 ;
        RECT 49.515 106.780 49.805 106.825 ;
        RECT 52.755 106.780 53.405 106.825 ;
        RECT 40.660 106.640 45.030 106.780 ;
        RECT 35.155 106.595 35.445 106.640 ;
        RECT 40.660 106.580 40.980 106.640 ;
        RECT 30.655 106.440 30.945 106.485 ;
        RECT 34.235 106.440 34.525 106.485 ;
        RECT 36.070 106.440 36.360 106.485 ;
        RECT 30.655 106.300 36.360 106.440 ;
        RECT 30.655 106.255 30.945 106.300 ;
        RECT 34.235 106.255 34.525 106.300 ;
        RECT 36.070 106.255 36.360 106.300 ;
        RECT 36.520 106.240 36.840 106.500 ;
        RECT 38.360 106.240 38.680 106.500 ;
        RECT 40.215 106.440 40.505 106.485 ;
        RECT 40.750 106.440 40.890 106.580 ;
        RECT 40.215 106.300 40.890 106.440 ;
        RECT 41.120 106.440 41.440 106.500 ;
        RECT 44.890 106.485 45.030 106.640 ;
        RECT 49.515 106.640 53.405 106.780 ;
        RECT 49.515 106.595 50.105 106.640 ;
        RECT 52.755 106.595 53.405 106.640 ;
        RECT 49.815 106.500 50.105 106.595 ;
        RECT 55.380 106.580 55.700 106.840 ;
        RECT 65.040 106.780 65.360 106.840 ;
        RECT 66.075 106.780 66.365 106.825 ;
        RECT 69.315 106.780 69.965 106.825 ;
        RECT 65.040 106.640 69.965 106.780 ;
        RECT 65.040 106.580 65.360 106.640 ;
        RECT 66.075 106.595 66.665 106.640 ;
        RECT 69.315 106.595 69.965 106.640 ;
        RECT 42.975 106.440 43.265 106.485 ;
        RECT 41.120 106.300 43.265 106.440 ;
        RECT 40.215 106.255 40.505 106.300 ;
        RECT 41.120 106.240 41.440 106.300 ;
        RECT 42.975 106.255 43.265 106.300 ;
        RECT 44.815 106.255 45.105 106.485 ;
        RECT 45.275 106.440 45.565 106.485 ;
        RECT 45.720 106.440 46.040 106.500 ;
        RECT 45.275 106.300 46.040 106.440 ;
        RECT 45.275 106.255 45.565 106.300 ;
        RECT 30.080 106.100 30.400 106.160 ;
        RECT 29.250 105.960 30.400 106.100 ;
        RECT 25.955 105.915 26.245 105.960 ;
        RECT 28.700 105.900 29.020 105.960 ;
        RECT 30.080 105.900 30.400 105.960 ;
        RECT 35.140 106.100 35.460 106.160 ;
        RECT 35.140 105.960 42.270 106.100 ;
        RECT 35.140 105.900 35.460 105.960 ;
        RECT 42.130 105.805 42.270 105.960 ;
        RECT 20.075 105.760 20.365 105.805 ;
        RECT 23.195 105.760 23.485 105.805 ;
        RECT 25.085 105.760 25.375 105.805 ;
        RECT 20.075 105.620 25.375 105.760 ;
        RECT 20.075 105.575 20.365 105.620 ;
        RECT 23.195 105.575 23.485 105.620 ;
        RECT 25.085 105.575 25.375 105.620 ;
        RECT 30.655 105.760 30.945 105.805 ;
        RECT 33.775 105.760 34.065 105.805 ;
        RECT 35.665 105.760 35.955 105.805 ;
        RECT 30.655 105.620 35.955 105.760 ;
        RECT 30.655 105.575 30.945 105.620 ;
        RECT 33.775 105.575 34.065 105.620 ;
        RECT 35.665 105.575 35.955 105.620 ;
        RECT 42.055 105.575 42.345 105.805 ;
        RECT 44.890 105.760 45.030 106.255 ;
        RECT 45.720 106.240 46.040 106.300 ;
        RECT 49.815 106.280 50.180 106.500 ;
        RECT 49.860 106.240 50.180 106.280 ;
        RECT 50.895 106.440 51.185 106.485 ;
        RECT 54.475 106.440 54.765 106.485 ;
        RECT 56.310 106.440 56.600 106.485 ;
        RECT 50.895 106.300 56.600 106.440 ;
        RECT 50.895 106.255 51.185 106.300 ;
        RECT 54.475 106.255 54.765 106.300 ;
        RECT 56.310 106.255 56.600 106.300 ;
        RECT 58.155 106.440 58.445 106.485 ;
        RECT 59.980 106.440 60.300 106.500 ;
        RECT 58.155 106.300 60.300 106.440 ;
        RECT 58.155 106.255 58.445 106.300 ;
        RECT 46.655 106.100 46.945 106.145 ;
        RECT 49.400 106.100 49.720 106.160 ;
        RECT 52.160 106.100 52.480 106.160 ;
        RECT 46.655 105.960 49.720 106.100 ;
        RECT 46.655 105.915 46.945 105.960 ;
        RECT 49.400 105.900 49.720 105.960 ;
        RECT 50.180 105.960 56.530 106.100 ;
        RECT 50.180 105.760 50.320 105.960 ;
        RECT 52.160 105.900 52.480 105.960 ;
        RECT 44.890 105.620 50.320 105.760 ;
        RECT 50.895 105.760 51.185 105.805 ;
        RECT 54.015 105.760 54.305 105.805 ;
        RECT 55.905 105.760 56.195 105.805 ;
        RECT 50.895 105.620 56.195 105.760 ;
        RECT 56.390 105.760 56.530 105.960 ;
        RECT 56.760 105.900 57.080 106.160 ;
        RECT 58.230 105.760 58.370 106.255 ;
        RECT 59.980 106.240 60.300 106.300 ;
        RECT 60.440 106.440 60.760 106.500 ;
        RECT 61.375 106.440 61.665 106.485 ;
        RECT 60.440 106.300 61.665 106.440 ;
        RECT 60.440 106.240 60.760 106.300 ;
        RECT 61.375 106.255 61.665 106.300 ;
        RECT 66.375 106.280 66.665 106.595 ;
        RECT 71.940 106.580 72.260 106.840 ;
        RECT 78.955 106.780 79.245 106.825 ;
        RECT 81.600 106.780 81.920 106.840 ;
        RECT 82.195 106.780 82.845 106.825 ;
        RECT 78.955 106.640 82.845 106.780 ;
        RECT 78.955 106.595 79.545 106.640 ;
        RECT 67.455 106.440 67.745 106.485 ;
        RECT 71.035 106.440 71.325 106.485 ;
        RECT 72.870 106.440 73.160 106.485 ;
        RECT 67.455 106.300 73.160 106.440 ;
        RECT 67.455 106.255 67.745 106.300 ;
        RECT 71.035 106.255 71.325 106.300 ;
        RECT 72.870 106.255 73.160 106.300 ;
        RECT 74.700 106.240 75.020 106.500 ;
        RECT 79.255 106.280 79.545 106.595 ;
        RECT 81.600 106.580 81.920 106.640 ;
        RECT 82.195 106.595 82.845 106.640 ;
        RECT 83.440 106.780 83.760 106.840 ;
        RECT 89.050 106.825 89.190 106.980 ;
        RECT 93.560 106.920 93.880 106.980 ;
        RECT 103.770 106.980 109.060 107.120 ;
        RECT 84.835 106.780 85.125 106.825 ;
        RECT 83.440 106.640 85.125 106.780 ;
        RECT 83.440 106.580 83.760 106.640 ;
        RECT 84.835 106.595 85.125 106.640 ;
        RECT 88.975 106.595 89.265 106.825 ;
        RECT 91.835 106.780 92.125 106.825 ;
        RECT 92.640 106.780 92.960 106.840 ;
        RECT 95.075 106.780 95.725 106.825 ;
        RECT 91.835 106.640 95.725 106.780 ;
        RECT 91.835 106.595 92.425 106.640 ;
        RECT 80.335 106.440 80.625 106.485 ;
        RECT 83.915 106.440 84.205 106.485 ;
        RECT 85.750 106.440 86.040 106.485 ;
        RECT 80.335 106.300 86.040 106.440 ;
        RECT 80.335 106.255 80.625 106.300 ;
        RECT 83.915 106.255 84.205 106.300 ;
        RECT 85.750 106.255 86.040 106.300 ;
        RECT 86.660 106.440 86.980 106.500 ;
        RECT 87.135 106.440 87.425 106.485 ;
        RECT 86.660 106.300 87.425 106.440 ;
        RECT 86.660 106.240 86.980 106.300 ;
        RECT 87.135 106.255 87.425 106.300 ;
        RECT 92.135 106.280 92.425 106.595 ;
        RECT 92.640 106.580 92.960 106.640 ;
        RECT 95.075 106.595 95.725 106.640 ;
        RECT 97.700 106.580 98.020 106.840 ;
        RECT 103.770 106.825 103.910 106.980 ;
        RECT 108.740 106.920 109.060 106.980 ;
        RECT 103.695 106.595 103.985 106.825 ;
        RECT 106.555 106.780 106.845 106.825 ;
        RECT 109.200 106.780 109.520 106.840 ;
        RECT 109.795 106.780 110.445 106.825 ;
        RECT 106.555 106.640 110.445 106.780 ;
        RECT 106.555 106.595 107.145 106.640 ;
        RECT 93.215 106.440 93.505 106.485 ;
        RECT 96.795 106.440 97.085 106.485 ;
        RECT 98.630 106.440 98.920 106.485 ;
        RECT 93.215 106.300 98.920 106.440 ;
        RECT 93.215 106.255 93.505 106.300 ;
        RECT 96.795 106.255 97.085 106.300 ;
        RECT 98.630 106.255 98.920 106.300 ;
        RECT 100.475 106.440 100.765 106.485 ;
        RECT 102.300 106.440 102.620 106.500 ;
        RECT 100.475 106.300 102.620 106.440 ;
        RECT 100.475 106.255 100.765 106.300 ;
        RECT 102.300 106.240 102.620 106.300 ;
        RECT 106.855 106.280 107.145 106.595 ;
        RECT 109.200 106.580 109.520 106.640 ;
        RECT 109.795 106.595 110.445 106.640 ;
        RECT 111.040 106.780 111.360 106.840 ;
        RECT 112.435 106.780 112.725 106.825 ;
        RECT 111.040 106.640 112.725 106.780 ;
        RECT 111.040 106.580 111.360 106.640 ;
        RECT 112.435 106.595 112.725 106.640 ;
        RECT 117.020 106.580 117.340 106.840 ;
        RECT 119.780 106.825 120.100 106.840 ;
        RECT 119.315 106.780 120.100 106.825 ;
        RECT 122.915 106.780 123.205 106.825 ;
        RECT 119.315 106.640 123.205 106.780 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 119.315 106.595 120.100 106.640 ;
        RECT 119.780 106.580 120.100 106.595 ;
        RECT 122.615 106.595 123.205 106.640 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 107.935 106.440 108.225 106.485 ;
        RECT 111.515 106.440 111.805 106.485 ;
        RECT 113.350 106.440 113.640 106.485 ;
        RECT 107.935 106.300 113.640 106.440 ;
        RECT 107.935 106.255 108.225 106.300 ;
        RECT 111.515 106.255 111.805 106.300 ;
        RECT 113.350 106.255 113.640 106.300 ;
        RECT 116.120 106.440 116.410 106.485 ;
        RECT 117.955 106.440 118.245 106.485 ;
        RECT 121.535 106.440 121.825 106.485 ;
        RECT 116.120 106.300 121.825 106.440 ;
        RECT 116.120 106.255 116.410 106.300 ;
        RECT 117.955 106.255 118.245 106.300 ;
        RECT 121.535 106.255 121.825 106.300 ;
        RECT 122.615 106.280 122.905 106.595 ;
        RECT 63.215 106.100 63.505 106.145 ;
        RECT 68.260 106.100 68.580 106.160 ;
        RECT 63.215 105.960 68.580 106.100 ;
        RECT 63.215 105.915 63.505 105.960 ;
        RECT 68.260 105.900 68.580 105.960 ;
        RECT 73.320 105.900 73.640 106.160 ;
        RECT 76.095 106.100 76.385 106.145 ;
        RECT 79.760 106.100 80.080 106.160 ;
        RECT 76.095 105.960 80.080 106.100 ;
        RECT 76.095 105.915 76.385 105.960 ;
        RECT 79.760 105.900 80.080 105.960 ;
        RECT 86.200 106.100 86.520 106.160 ;
        RECT 99.080 106.100 99.400 106.160 ;
        RECT 111.960 106.100 112.280 106.160 ;
        RECT 113.815 106.100 114.105 106.145 ;
        RECT 115.655 106.100 115.945 106.145 ;
        RECT 86.200 105.960 115.945 106.100 ;
        RECT 86.200 105.900 86.520 105.960 ;
        RECT 99.080 105.900 99.400 105.960 ;
        RECT 111.960 105.900 112.280 105.960 ;
        RECT 113.815 105.915 114.105 105.960 ;
        RECT 115.655 105.915 115.945 105.960 ;
        RECT 120.700 106.100 121.020 106.160 ;
        RECT 125.775 106.100 126.065 106.145 ;
        RECT 120.700 105.960 126.065 106.100 ;
        RECT 120.700 105.900 121.020 105.960 ;
        RECT 125.775 105.915 126.065 105.960 ;
        RECT 56.390 105.620 58.370 105.760 ;
        RECT 60.455 105.760 60.745 105.805 ;
        RECT 64.120 105.760 64.440 105.820 ;
        RECT 60.455 105.620 64.440 105.760 ;
        RECT 50.895 105.575 51.185 105.620 ;
        RECT 54.015 105.575 54.305 105.620 ;
        RECT 55.905 105.575 56.195 105.620 ;
        RECT 60.455 105.575 60.745 105.620 ;
        RECT 64.120 105.560 64.440 105.620 ;
        RECT 67.455 105.760 67.745 105.805 ;
        RECT 70.575 105.760 70.865 105.805 ;
        RECT 72.465 105.760 72.755 105.805 ;
        RECT 67.455 105.620 72.755 105.760 ;
        RECT 67.455 105.575 67.745 105.620 ;
        RECT 70.575 105.575 70.865 105.620 ;
        RECT 72.465 105.575 72.755 105.620 ;
        RECT 80.335 105.760 80.625 105.805 ;
        RECT 83.455 105.760 83.745 105.805 ;
        RECT 85.345 105.760 85.635 105.805 ;
        RECT 80.335 105.620 85.635 105.760 ;
        RECT 80.335 105.575 80.625 105.620 ;
        RECT 83.455 105.575 83.745 105.620 ;
        RECT 85.345 105.575 85.635 105.620 ;
        RECT 93.215 105.760 93.505 105.805 ;
        RECT 96.335 105.760 96.625 105.805 ;
        RECT 98.225 105.760 98.515 105.805 ;
        RECT 93.215 105.620 98.515 105.760 ;
        RECT 93.215 105.575 93.505 105.620 ;
        RECT 96.335 105.575 96.625 105.620 ;
        RECT 98.225 105.575 98.515 105.620 ;
        RECT 107.935 105.760 108.225 105.805 ;
        RECT 111.055 105.760 111.345 105.805 ;
        RECT 112.945 105.760 113.235 105.805 ;
        RECT 107.935 105.620 113.235 105.760 ;
        RECT 107.935 105.575 108.225 105.620 ;
        RECT 111.055 105.575 111.345 105.620 ;
        RECT 112.945 105.575 113.235 105.620 ;
        RECT 116.525 105.760 116.815 105.805 ;
        RECT 118.415 105.760 118.705 105.805 ;
        RECT 121.535 105.760 121.825 105.805 ;
        RECT 116.525 105.620 121.825 105.760 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 116.525 105.575 116.815 105.620 ;
        RECT 118.415 105.575 118.705 105.620 ;
        RECT 121.535 105.575 121.825 105.620 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 36.060 105.420 36.380 105.480 ;
        RECT 39.755 105.420 40.045 105.465 ;
        RECT 36.060 105.280 40.045 105.420 ;
        RECT 36.060 105.220 36.380 105.280 ;
        RECT 39.755 105.235 40.045 105.280 ;
        RECT 42.960 105.420 43.280 105.480 ;
        RECT 44.355 105.420 44.645 105.465 ;
        RECT 42.960 105.280 44.645 105.420 ;
        RECT 42.960 105.220 43.280 105.280 ;
        RECT 44.355 105.235 44.645 105.280 ;
        RECT 46.195 105.420 46.485 105.465 ;
        RECT 48.020 105.420 48.340 105.480 ;
        RECT 46.195 105.280 48.340 105.420 ;
        RECT 46.195 105.235 46.485 105.280 ;
        RECT 48.020 105.220 48.340 105.280 ;
        RECT 56.760 105.420 57.080 105.480 ;
        RECT 57.695 105.420 57.985 105.465 ;
        RECT 56.760 105.280 57.985 105.420 ;
        RECT 56.760 105.220 57.080 105.280 ;
        RECT 57.695 105.235 57.985 105.280 ;
        RECT 62.295 105.420 62.585 105.465 ;
        RECT 63.660 105.420 63.980 105.480 ;
        RECT 62.295 105.280 63.980 105.420 ;
        RECT 62.295 105.235 62.585 105.280 ;
        RECT 63.660 105.220 63.980 105.280 ;
        RECT 75.620 105.220 75.940 105.480 ;
        RECT 88.040 105.220 88.360 105.480 ;
        RECT 97.240 105.420 97.560 105.480 ;
        RECT 100.015 105.420 100.305 105.465 ;
        RECT 97.240 105.280 100.305 105.420 ;
        RECT 97.240 105.220 97.560 105.280 ;
        RECT 100.015 105.235 100.305 105.280 ;
        RECT 102.775 105.420 103.065 105.465 ;
        RECT 104.140 105.420 104.460 105.480 ;
        RECT 102.775 105.280 104.460 105.420 ;
        RECT 102.775 105.235 103.065 105.280 ;
        RECT 104.140 105.220 104.460 105.280 ;
        RECT 14.370 104.600 127.530 105.080 ;
        RECT 28.700 104.400 29.020 104.460 ;
        RECT 36.520 104.400 36.840 104.460 ;
        RECT 28.700 104.260 36.840 104.400 ;
        RECT 28.700 104.200 29.020 104.260 ;
        RECT 36.520 104.200 36.840 104.260 ;
        RECT 49.860 104.400 50.180 104.460 ;
        RECT 51.715 104.400 52.005 104.445 ;
        RECT 49.860 104.260 52.005 104.400 ;
        RECT 49.860 104.200 50.180 104.260 ;
        RECT 51.715 104.215 52.005 104.260 ;
        RECT 56.300 104.400 56.620 104.460 ;
        RECT 73.320 104.400 73.640 104.460 ;
        RECT 56.300 104.260 73.640 104.400 ;
        RECT 56.300 104.200 56.620 104.260 ;
        RECT 28.790 103.765 28.930 104.200 ;
        RECT 29.585 104.060 29.875 104.105 ;
        RECT 31.475 104.060 31.765 104.105 ;
        RECT 34.595 104.060 34.885 104.105 ;
        RECT 29.585 103.920 34.885 104.060 ;
        RECT 29.585 103.875 29.875 103.920 ;
        RECT 31.475 103.875 31.765 103.920 ;
        RECT 34.595 103.875 34.885 103.920 ;
        RECT 43.535 104.060 43.825 104.105 ;
        RECT 46.655 104.060 46.945 104.105 ;
        RECT 48.545 104.060 48.835 104.105 ;
        RECT 50.320 104.060 50.640 104.120 ;
        RECT 56.390 104.060 56.530 104.200 ;
        RECT 43.535 103.920 48.835 104.060 ;
        RECT 43.535 103.875 43.825 103.920 ;
        RECT 46.655 103.875 46.945 103.920 ;
        RECT 48.545 103.875 48.835 103.920 ;
        RECT 50.180 103.920 56.530 104.060 ;
        RECT 56.875 104.060 57.165 104.105 ;
        RECT 59.995 104.060 60.285 104.105 ;
        RECT 61.885 104.060 62.175 104.105 ;
        RECT 56.875 103.920 62.175 104.060 ;
        RECT 50.180 103.860 50.640 103.920 ;
        RECT 56.875 103.875 57.165 103.920 ;
        RECT 59.995 103.875 60.285 103.920 ;
        RECT 61.885 103.875 62.175 103.920 ;
        RECT 28.715 103.535 29.005 103.765 ;
        RECT 30.095 103.720 30.385 103.765 ;
        RECT 35.140 103.720 35.460 103.780 ;
        RECT 36.060 103.720 36.380 103.780 ;
        RECT 30.095 103.580 35.460 103.720 ;
        RECT 30.095 103.535 30.385 103.580 ;
        RECT 35.140 103.520 35.460 103.580 ;
        RECT 35.690 103.580 36.380 103.720 ;
        RECT 27.320 103.180 27.640 103.440 ;
        RECT 29.180 103.380 29.470 103.425 ;
        RECT 31.015 103.380 31.305 103.425 ;
        RECT 34.595 103.380 34.885 103.425 ;
        RECT 35.690 103.400 35.830 103.580 ;
        RECT 36.060 103.520 36.380 103.580 ;
        RECT 48.020 103.520 48.340 103.780 ;
        RECT 49.415 103.720 49.705 103.765 ;
        RECT 50.180 103.720 50.320 103.860 ;
        RECT 49.415 103.580 50.320 103.720 ;
        RECT 57.680 103.720 58.000 103.780 ;
        RECT 62.830 103.765 62.970 104.260 ;
        RECT 73.320 104.200 73.640 104.260 ;
        RECT 78.840 104.400 79.160 104.460 ;
        RECT 124.855 104.400 125.145 104.445 ;
        RECT 78.840 104.260 125.145 104.400 ;
        RECT 78.840 104.200 79.160 104.260 ;
        RECT 124.855 104.215 125.145 104.260 ;
        RECT 67.455 104.060 67.745 104.105 ;
        RECT 70.575 104.060 70.865 104.105 ;
        RECT 72.465 104.060 72.755 104.105 ;
        RECT 67.455 103.920 72.755 104.060 ;
        RECT 67.455 103.875 67.745 103.920 ;
        RECT 70.575 103.875 70.865 103.920 ;
        RECT 72.465 103.875 72.755 103.920 ;
        RECT 80.335 104.060 80.625 104.105 ;
        RECT 83.455 104.060 83.745 104.105 ;
        RECT 85.345 104.060 85.635 104.105 ;
        RECT 80.335 103.920 85.635 104.060 ;
        RECT 80.335 103.875 80.625 103.920 ;
        RECT 83.455 103.875 83.745 103.920 ;
        RECT 85.345 103.875 85.635 103.920 ;
        RECT 90.915 104.060 91.205 104.105 ;
        RECT 94.035 104.060 94.325 104.105 ;
        RECT 95.925 104.060 96.215 104.105 ;
        RECT 90.915 103.920 96.215 104.060 ;
        RECT 90.915 103.875 91.205 103.920 ;
        RECT 94.035 103.875 94.325 103.920 ;
        RECT 95.925 103.875 96.215 103.920 ;
        RECT 106.095 104.060 106.385 104.105 ;
        RECT 109.215 104.060 109.505 104.105 ;
        RECT 111.105 104.060 111.395 104.105 ;
        RECT 106.095 103.920 111.395 104.060 ;
        RECT 106.095 103.875 106.385 103.920 ;
        RECT 109.215 103.875 109.505 103.920 ;
        RECT 111.105 103.875 111.395 103.920 ;
        RECT 113.305 104.060 113.595 104.105 ;
        RECT 115.195 104.060 115.485 104.105 ;
        RECT 118.315 104.060 118.605 104.105 ;
        RECT 113.305 103.920 118.605 104.060 ;
        RECT 113.305 103.875 113.595 103.920 ;
        RECT 115.195 103.875 115.485 103.920 ;
        RECT 118.315 103.875 118.605 103.920 ;
        RECT 61.375 103.720 61.665 103.765 ;
        RECT 57.680 103.580 61.665 103.720 ;
        RECT 49.415 103.535 49.705 103.580 ;
        RECT 57.680 103.520 58.000 103.580 ;
        RECT 61.375 103.535 61.665 103.580 ;
        RECT 62.755 103.535 63.045 103.765 ;
        RECT 63.660 103.720 63.980 103.780 ;
        RECT 71.955 103.720 72.245 103.765 ;
        RECT 63.660 103.580 72.245 103.720 ;
        RECT 63.660 103.520 63.980 103.580 ;
        RECT 71.955 103.535 72.245 103.580 ;
        RECT 73.320 103.520 73.640 103.780 ;
        RECT 75.620 103.720 75.940 103.780 ;
        RECT 84.835 103.720 85.125 103.765 ;
        RECT 75.620 103.580 85.125 103.720 ;
        RECT 75.620 103.520 75.940 103.580 ;
        RECT 84.835 103.535 85.125 103.580 ;
        RECT 86.200 103.520 86.520 103.780 ;
        RECT 88.040 103.720 88.360 103.780 ;
        RECT 95.415 103.720 95.705 103.765 ;
        RECT 88.040 103.580 95.705 103.720 ;
        RECT 88.040 103.520 88.360 103.580 ;
        RECT 95.415 103.535 95.705 103.580 ;
        RECT 96.795 103.720 97.085 103.765 ;
        RECT 99.080 103.720 99.400 103.780 ;
        RECT 96.795 103.580 99.400 103.720 ;
        RECT 96.795 103.535 97.085 103.580 ;
        RECT 99.080 103.520 99.400 103.580 ;
        RECT 110.580 103.520 110.900 103.780 ;
        RECT 111.960 103.720 112.280 103.780 ;
        RECT 112.435 103.720 112.725 103.765 ;
        RECT 111.960 103.580 112.725 103.720 ;
        RECT 111.960 103.520 112.280 103.580 ;
        RECT 112.435 103.535 112.725 103.580 ;
        RECT 113.800 103.520 114.120 103.780 ;
        RECT 115.640 103.720 115.960 103.780 ;
        RECT 122.555 103.720 122.845 103.765 ;
        RECT 115.640 103.580 122.845 103.720 ;
        RECT 115.640 103.520 115.960 103.580 ;
        RECT 122.555 103.535 122.845 103.580 ;
        RECT 29.180 103.240 34.885 103.380 ;
        RECT 29.180 103.195 29.470 103.240 ;
        RECT 31.015 103.195 31.305 103.240 ;
        RECT 34.595 103.195 34.885 103.240 ;
        RECT 35.675 103.085 35.965 103.400 ;
        RECT 32.375 103.040 33.025 103.085 ;
        RECT 35.675 103.040 36.265 103.085 ;
        RECT 32.375 102.900 36.265 103.040 ;
        RECT 32.375 102.855 33.025 102.900 ;
        RECT 35.975 102.855 36.265 102.900 ;
        RECT 38.820 102.840 39.140 103.100 ;
        RECT 42.455 103.085 42.745 103.400 ;
        RECT 43.535 103.380 43.825 103.425 ;
        RECT 47.115 103.380 47.405 103.425 ;
        RECT 48.950 103.380 49.240 103.425 ;
        RECT 43.535 103.240 49.240 103.380 ;
        RECT 43.535 103.195 43.825 103.240 ;
        RECT 47.115 103.195 47.405 103.240 ;
        RECT 48.950 103.195 49.240 103.240 ;
        RECT 52.160 103.180 52.480 103.440 ;
        RECT 39.295 102.855 39.585 103.085 ;
        RECT 42.155 103.040 42.745 103.085 ;
        RECT 42.960 103.040 43.280 103.100 ;
        RECT 45.395 103.040 46.045 103.085 ;
        RECT 42.155 102.900 46.045 103.040 ;
        RECT 42.155 102.855 42.445 102.900 ;
        RECT 27.780 102.500 28.100 102.760 ;
        RECT 39.370 102.700 39.510 102.855 ;
        RECT 42.960 102.840 43.280 102.900 ;
        RECT 45.395 102.855 46.045 102.900 ;
        RECT 52.635 103.040 52.925 103.085 ;
        RECT 54.460 103.040 54.780 103.100 ;
        RECT 55.795 103.085 56.085 103.400 ;
        RECT 56.875 103.380 57.165 103.425 ;
        RECT 60.455 103.380 60.745 103.425 ;
        RECT 62.290 103.380 62.580 103.425 ;
        RECT 56.875 103.240 62.580 103.380 ;
        RECT 56.875 103.195 57.165 103.240 ;
        RECT 60.455 103.195 60.745 103.240 ;
        RECT 62.290 103.195 62.580 103.240 ;
        RECT 52.635 102.900 54.780 103.040 ;
        RECT 52.635 102.855 52.925 102.900 ;
        RECT 54.460 102.840 54.780 102.900 ;
        RECT 55.495 103.040 56.085 103.085 ;
        RECT 56.300 103.040 56.620 103.100 ;
        RECT 58.735 103.040 59.385 103.085 ;
        RECT 55.495 102.900 59.385 103.040 ;
        RECT 55.495 102.855 55.785 102.900 ;
        RECT 56.300 102.840 56.620 102.900 ;
        RECT 58.735 102.855 59.385 102.900 ;
        RECT 60.900 103.040 61.220 103.100 ;
        RECT 63.215 103.040 63.505 103.085 ;
        RECT 60.900 102.900 63.505 103.040 ;
        RECT 60.900 102.840 61.220 102.900 ;
        RECT 63.215 102.855 63.505 102.900 ;
        RECT 64.120 103.040 64.440 103.100 ;
        RECT 66.375 103.085 66.665 103.400 ;
        RECT 67.455 103.380 67.745 103.425 ;
        RECT 71.035 103.380 71.325 103.425 ;
        RECT 72.870 103.380 73.160 103.425 ;
        RECT 79.300 103.400 79.620 103.440 ;
        RECT 67.455 103.240 73.160 103.380 ;
        RECT 67.455 103.195 67.745 103.240 ;
        RECT 71.035 103.195 71.325 103.240 ;
        RECT 72.870 103.195 73.160 103.240 ;
        RECT 79.255 103.180 79.620 103.400 ;
        RECT 80.335 103.380 80.625 103.425 ;
        RECT 83.915 103.380 84.205 103.425 ;
        RECT 85.750 103.380 86.040 103.425 ;
        RECT 80.335 103.240 86.040 103.380 ;
        RECT 80.335 103.195 80.625 103.240 ;
        RECT 83.915 103.195 84.205 103.240 ;
        RECT 85.750 103.195 86.040 103.240 ;
        RECT 66.075 103.040 66.665 103.085 ;
        RECT 69.315 103.040 69.965 103.085 ;
        RECT 64.120 102.900 69.965 103.040 ;
        RECT 64.120 102.840 64.440 102.900 ;
        RECT 66.075 102.855 66.365 102.900 ;
        RECT 69.315 102.855 69.965 102.900 ;
        RECT 73.780 103.040 74.100 103.100 ;
        RECT 79.255 103.085 79.545 103.180 ;
        RECT 76.095 103.040 76.385 103.085 ;
        RECT 73.780 102.900 76.385 103.040 ;
        RECT 73.780 102.840 74.100 102.900 ;
        RECT 76.095 102.855 76.385 102.900 ;
        RECT 78.955 103.040 79.545 103.085 ;
        RECT 82.195 103.040 82.845 103.085 ;
        RECT 78.955 102.900 82.845 103.040 ;
        RECT 78.955 102.855 79.245 102.900 ;
        RECT 82.195 102.855 82.845 102.900 ;
        RECT 86.660 102.840 86.980 103.100 ;
        RECT 87.580 103.040 87.900 103.100 ;
        RECT 89.835 103.085 90.125 103.400 ;
        RECT 90.915 103.380 91.205 103.425 ;
        RECT 94.495 103.380 94.785 103.425 ;
        RECT 96.330 103.380 96.620 103.425 ;
        RECT 90.915 103.240 96.620 103.380 ;
        RECT 90.915 103.195 91.205 103.240 ;
        RECT 94.495 103.195 94.785 103.240 ;
        RECT 96.330 103.195 96.620 103.240 ;
        RECT 89.535 103.040 90.125 103.085 ;
        RECT 92.775 103.040 93.425 103.085 ;
        RECT 87.580 102.900 93.425 103.040 ;
        RECT 87.580 102.840 87.900 102.900 ;
        RECT 89.535 102.855 89.825 102.900 ;
        RECT 92.775 102.855 93.425 102.900 ;
        RECT 101.855 103.040 102.145 103.085 ;
        RECT 103.680 103.040 104.000 103.100 ;
        RECT 101.855 102.900 104.000 103.040 ;
        RECT 101.855 102.855 102.145 102.900 ;
        RECT 103.680 102.840 104.000 102.900 ;
        RECT 104.140 103.040 104.460 103.100 ;
        RECT 105.015 103.085 105.305 103.400 ;
        RECT 106.095 103.380 106.385 103.425 ;
        RECT 109.675 103.380 109.965 103.425 ;
        RECT 111.510 103.380 111.800 103.425 ;
        RECT 106.095 103.240 111.800 103.380 ;
        RECT 106.095 103.195 106.385 103.240 ;
        RECT 109.675 103.195 109.965 103.240 ;
        RECT 111.510 103.195 111.800 103.240 ;
        RECT 112.900 103.380 113.190 103.425 ;
        RECT 114.735 103.380 115.025 103.425 ;
        RECT 118.315 103.380 118.605 103.425 ;
        RECT 112.900 103.240 118.605 103.380 ;
        RECT 112.900 103.195 113.190 103.240 ;
        RECT 114.735 103.195 115.025 103.240 ;
        RECT 118.315 103.195 118.605 103.240 ;
        RECT 116.100 103.085 116.420 103.100 ;
        RECT 119.395 103.085 119.685 103.400 ;
        RECT 125.760 103.180 126.080 103.440 ;
        RECT 104.715 103.040 105.305 103.085 ;
        RECT 107.955 103.040 108.605 103.085 ;
        RECT 104.140 102.900 108.605 103.040 ;
        RECT 104.140 102.840 104.460 102.900 ;
        RECT 104.715 102.855 105.005 102.900 ;
        RECT 107.955 102.855 108.605 102.900 ;
        RECT 116.095 103.040 116.745 103.085 ;
        RECT 119.395 103.040 119.985 103.085 ;
        RECT 116.095 102.900 119.985 103.040 ;
        RECT 116.095 102.855 116.745 102.900 ;
        RECT 119.695 102.855 119.985 102.900 ;
        RECT 116.100 102.840 116.420 102.855 ;
        RECT 43.880 102.700 44.200 102.760 ;
        RECT 39.370 102.560 44.200 102.700 ;
        RECT 43.880 102.500 44.200 102.560 ;
        RECT 14.370 101.880 127.530 102.360 ;
        RECT 119.780 101.480 120.100 101.740 ;
        RECT 27.435 101.340 27.725 101.385 ;
        RECT 30.675 101.340 31.325 101.385 ;
        RECT 27.435 101.200 31.325 101.340 ;
        RECT 27.435 101.155 28.025 101.200 ;
        RECT 30.675 101.155 31.325 101.200 ;
        RECT 33.315 101.340 33.605 101.385 ;
        RECT 33.760 101.340 34.080 101.400 ;
        RECT 97.240 101.385 97.560 101.400 ;
        RECT 33.315 101.200 34.080 101.340 ;
        RECT 33.315 101.155 33.605 101.200 ;
        RECT 27.735 101.060 28.025 101.155 ;
        RECT 33.760 101.140 34.080 101.200 ;
        RECT 93.675 101.340 93.965 101.385 ;
        RECT 96.915 101.340 97.565 101.385 ;
        RECT 93.675 101.200 97.565 101.340 ;
        RECT 93.675 101.155 94.265 101.200 ;
        RECT 96.915 101.155 97.565 101.200 ;
        RECT 27.735 100.840 28.100 101.060 ;
        RECT 27.780 100.800 28.100 100.840 ;
        RECT 28.815 101.000 29.105 101.045 ;
        RECT 32.395 101.000 32.685 101.045 ;
        RECT 34.230 101.000 34.520 101.045 ;
        RECT 28.815 100.860 34.520 101.000 ;
        RECT 28.815 100.815 29.105 100.860 ;
        RECT 32.395 100.815 32.685 100.860 ;
        RECT 34.230 100.815 34.520 100.860 ;
        RECT 34.695 101.000 34.985 101.045 ;
        RECT 36.520 101.000 36.840 101.060 ;
        RECT 34.695 100.860 36.840 101.000 ;
        RECT 34.695 100.815 34.985 100.860 ;
        RECT 36.520 100.800 36.840 100.860 ;
        RECT 93.975 100.840 94.265 101.155 ;
        RECT 97.240 101.140 97.560 101.155 ;
        RECT 99.540 101.140 99.860 101.400 ;
        RECT 95.055 101.000 95.345 101.045 ;
        RECT 98.635 101.000 98.925 101.045 ;
        RECT 100.470 101.000 100.760 101.045 ;
        RECT 95.055 100.860 100.760 101.000 ;
        RECT 95.055 100.815 95.345 100.860 ;
        RECT 98.635 100.815 98.925 100.860 ;
        RECT 100.470 100.815 100.760 100.860 ;
        RECT 119.320 100.800 119.640 101.060 ;
        RECT 24.575 100.660 24.865 100.705 ;
        RECT 25.940 100.660 26.260 100.720 ;
        RECT 24.575 100.520 26.260 100.660 ;
        RECT 24.575 100.475 24.865 100.520 ;
        RECT 25.940 100.460 26.260 100.520 ;
        RECT 90.815 100.660 91.105 100.705 ;
        RECT 97.700 100.660 98.020 100.720 ;
        RECT 90.815 100.520 98.020 100.660 ;
        RECT 90.815 100.475 91.105 100.520 ;
        RECT 97.700 100.460 98.020 100.520 ;
        RECT 99.080 100.660 99.400 100.720 ;
        RECT 100.935 100.660 101.225 100.705 ;
        RECT 99.080 100.520 101.225 100.660 ;
        RECT 99.080 100.460 99.400 100.520 ;
        RECT 100.935 100.475 101.225 100.520 ;
        RECT 28.815 100.320 29.105 100.365 ;
        RECT 31.935 100.320 32.225 100.365 ;
        RECT 33.825 100.320 34.115 100.365 ;
        RECT 28.815 100.180 34.115 100.320 ;
        RECT 28.815 100.135 29.105 100.180 ;
        RECT 31.935 100.135 32.225 100.180 ;
        RECT 33.825 100.135 34.115 100.180 ;
        RECT 95.055 100.320 95.345 100.365 ;
        RECT 98.175 100.320 98.465 100.365 ;
        RECT 100.065 100.320 100.355 100.365 ;
        RECT 95.055 100.180 100.355 100.320 ;
        RECT 95.055 100.135 95.345 100.180 ;
        RECT 98.175 100.135 98.465 100.180 ;
        RECT 100.065 100.135 100.355 100.180 ;
        RECT 14.370 99.160 127.530 99.640 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 16.590 210.735 18.470 211.105 ;
        RECT 46.590 210.735 48.470 211.105 ;
        RECT 76.590 210.735 78.470 211.105 ;
        RECT 106.590 210.735 108.470 211.105 ;
        RECT 31.590 208.015 33.470 208.385 ;
        RECT 61.590 208.015 63.470 208.385 ;
        RECT 91.590 208.015 93.470 208.385 ;
        RECT 121.590 208.015 123.470 208.385 ;
        RECT 73.350 207.190 73.610 207.510 ;
        RECT 65.990 206.510 66.250 206.830 ;
        RECT 72.890 206.510 73.150 206.830 ;
        RECT 16.590 205.295 18.470 205.665 ;
        RECT 46.590 205.295 48.470 205.665 ;
        RECT 66.050 204.450 66.190 206.510 ;
        RECT 65.990 204.130 66.250 204.450 ;
        RECT 63.690 203.790 63.950 204.110 ;
        RECT 31.590 202.575 33.470 202.945 ;
        RECT 61.590 202.575 63.470 202.945 ;
        RECT 63.750 202.410 63.890 203.790 ;
        RECT 64.610 203.110 64.870 203.430 ;
        RECT 63.690 202.090 63.950 202.410 ;
        RECT 60.930 201.410 61.190 201.730 ;
        RECT 16.590 199.855 18.470 200.225 ;
        RECT 46.590 199.855 48.470 200.225 ;
        RECT 60.990 199.690 61.130 201.410 ;
        RECT 60.930 199.370 61.190 199.690 ;
        RECT 31.590 197.135 33.470 197.505 ;
        RECT 61.590 197.135 63.470 197.505 ;
        RECT 50.350 195.970 50.610 196.290 ;
        RECT 48.970 195.630 49.230 195.950 ;
        RECT 16.590 194.415 18.470 194.785 ;
        RECT 46.590 194.415 48.470 194.785 ;
        RECT 49.030 193.910 49.170 195.630 ;
        RECT 50.410 194.250 50.550 195.970 ;
        RECT 53.110 194.950 53.370 195.270 ;
        RECT 57.710 194.950 57.970 195.270 ;
        RECT 50.350 194.160 50.610 194.250 ;
        RECT 49.490 194.020 50.610 194.160 ;
        RECT 48.970 193.590 49.230 193.910 ;
        RECT 45.750 193.250 46.010 193.570 ;
        RECT 31.590 191.695 33.470 192.065 ;
        RECT 41.150 190.530 41.410 190.850 ;
        RECT 38.850 189.850 39.110 190.170 ;
        RECT 16.590 188.975 18.470 189.345 ;
        RECT 28.270 187.470 28.530 187.790 ;
        RECT 36.090 187.470 36.350 187.790 ;
        RECT 22.750 185.090 23.010 185.410 ;
        RECT 16.590 183.535 18.470 183.905 ;
        RECT 22.810 183.370 22.950 185.090 ;
        RECT 28.330 184.730 28.470 187.470 ;
        RECT 31.590 186.255 33.470 186.625 ;
        RECT 36.150 185.070 36.290 187.470 ;
        RECT 37.470 186.790 37.730 187.110 ;
        RECT 36.090 184.750 36.350 185.070 ;
        RECT 28.270 184.410 28.530 184.730 ;
        RECT 29.650 184.070 29.910 184.390 ;
        RECT 30.110 184.070 30.370 184.390 ;
        RECT 22.750 183.050 23.010 183.370 ;
        RECT 29.710 182.690 29.850 184.070 ;
        RECT 30.170 183.370 30.310 184.070 ;
        RECT 30.110 183.050 30.370 183.370 ;
        RECT 33.790 182.710 34.050 183.030 ;
        RECT 29.650 182.370 29.910 182.690 ;
        RECT 31.590 180.815 33.470 181.185 ;
        RECT 33.850 179.290 33.990 182.710 ;
        RECT 35.630 182.370 35.890 182.690 ;
        RECT 25.970 178.970 26.230 179.290 ;
        RECT 27.350 178.970 27.610 179.290 ;
        RECT 33.790 178.970 34.050 179.290 ;
        RECT 34.710 178.970 34.970 179.290 ;
        RECT 16.590 178.095 18.470 178.465 ;
        RECT 26.030 175.210 26.170 178.970 ;
        RECT 27.410 177.930 27.550 178.970 ;
        RECT 27.350 177.610 27.610 177.930 ;
        RECT 30.110 176.590 30.370 176.910 ;
        RECT 27.810 175.910 28.070 176.230 ;
        RECT 25.970 174.890 26.230 175.210 ;
        RECT 27.870 173.850 28.010 175.910 ;
        RECT 27.810 173.530 28.070 173.850 ;
        RECT 16.590 172.655 18.470 173.025 ;
        RECT 30.170 168.750 30.310 176.590 ;
        RECT 31.590 175.375 33.470 175.745 ;
        RECT 33.850 173.850 33.990 178.970 ;
        RECT 34.250 175.910 34.510 176.230 ;
        RECT 34.310 174.190 34.450 175.910 ;
        RECT 34.250 173.870 34.510 174.190 ;
        RECT 33.790 173.530 34.050 173.850 ;
        RECT 31.590 169.935 33.470 170.305 ;
        RECT 30.110 168.430 30.370 168.750 ;
        RECT 29.650 167.750 29.910 168.070 ;
        RECT 33.790 167.750 34.050 168.070 ;
        RECT 16.590 167.215 18.470 167.585 ;
        RECT 29.710 166.710 29.850 167.750 ;
        RECT 24.590 166.390 24.850 166.710 ;
        RECT 29.650 166.390 29.910 166.710 ;
        RECT 24.650 164.330 24.790 166.390 ;
        RECT 26.890 165.710 27.150 166.030 ;
        RECT 24.590 164.010 24.850 164.330 ;
        RECT 26.950 163.310 27.090 165.710 ;
        RECT 29.650 165.370 29.910 165.690 ;
        RECT 28.270 165.030 28.530 165.350 ;
        RECT 28.330 163.650 28.470 165.030 ;
        RECT 28.270 163.330 28.530 163.650 ;
        RECT 28.730 163.330 28.990 163.650 ;
        RECT 26.430 162.990 26.690 163.310 ;
        RECT 26.890 162.990 27.150 163.310 ;
        RECT 16.590 161.775 18.470 162.145 ;
        RECT 26.490 161.610 26.630 162.990 ;
        RECT 28.790 162.970 28.930 163.330 ;
        RECT 28.730 162.650 28.990 162.970 ;
        RECT 26.430 161.290 26.690 161.610 ;
        RECT 18.610 160.950 18.870 161.270 ;
        RECT 18.670 158.890 18.810 160.950 ;
        RECT 28.790 160.930 28.930 162.650 ;
        RECT 29.710 161.610 29.850 165.370 ;
        RECT 31.590 164.495 33.470 164.865 ;
        RECT 33.850 163.310 33.990 167.750 ;
        RECT 34.250 166.050 34.510 166.370 ;
        RECT 33.790 162.990 34.050 163.310 ;
        RECT 34.310 161.610 34.450 166.050 ;
        RECT 29.650 161.290 29.910 161.610 ;
        RECT 34.250 161.290 34.510 161.610 ;
        RECT 31.030 160.950 31.290 161.270 ;
        RECT 34.770 161.010 34.910 178.970 ;
        RECT 35.170 176.590 35.430 176.910 ;
        RECT 35.230 172.490 35.370 176.590 ;
        RECT 35.170 172.170 35.430 172.490 ;
        RECT 35.690 171.470 35.830 182.370 ;
        RECT 35.630 171.150 35.890 171.470 ;
        RECT 35.170 170.470 35.430 170.790 ;
        RECT 36.150 170.530 36.290 184.750 ;
        RECT 37.530 184.730 37.670 186.790 ;
        RECT 38.910 186.090 39.050 189.850 ;
        RECT 38.850 185.770 39.110 186.090 ;
        RECT 41.210 185.410 41.350 190.530 ;
        RECT 44.830 190.190 45.090 190.510 ;
        RECT 44.370 187.470 44.630 187.790 ;
        RECT 44.430 185.750 44.570 187.470 ;
        RECT 44.370 185.430 44.630 185.750 ;
        RECT 37.930 185.090 38.190 185.410 ;
        RECT 41.150 185.090 41.410 185.410 ;
        RECT 37.470 184.410 37.730 184.730 ;
        RECT 37.530 182.690 37.670 184.410 ;
        RECT 37.470 182.370 37.730 182.690 ;
        RECT 37.010 179.310 37.270 179.630 ;
        RECT 36.550 178.630 36.810 178.950 ;
        RECT 36.610 176.910 36.750 178.630 ;
        RECT 36.550 176.590 36.810 176.910 ;
        RECT 26.890 160.610 27.150 160.930 ;
        RECT 28.730 160.610 28.990 160.930 ;
        RECT 25.510 160.270 25.770 160.590 ;
        RECT 21.370 159.590 21.630 159.910 ;
        RECT 18.610 158.570 18.870 158.890 ;
        RECT 21.430 158.210 21.570 159.590 ;
        RECT 25.570 158.890 25.710 160.270 ;
        RECT 25.510 158.570 25.770 158.890 ;
        RECT 20.910 157.890 21.170 158.210 ;
        RECT 21.370 157.890 21.630 158.210 ;
        RECT 19.070 156.870 19.330 157.190 ;
        RECT 16.590 156.335 18.470 156.705 ;
        RECT 19.130 155.830 19.270 156.870 ;
        RECT 19.070 155.510 19.330 155.830 ;
        RECT 20.970 152.770 21.110 157.890 ;
        RECT 21.830 156.870 22.090 157.190 ;
        RECT 21.890 156.170 22.030 156.870 ;
        RECT 21.830 155.850 22.090 156.170 ;
        RECT 21.890 152.770 22.030 155.850 ;
        RECT 26.950 155.490 27.090 160.610 ;
        RECT 30.570 160.270 30.830 160.590 ;
        RECT 30.630 158.550 30.770 160.270 ;
        RECT 31.090 158.890 31.230 160.950 ;
        RECT 33.790 160.610 34.050 160.930 ;
        RECT 34.310 160.870 34.910 161.010 ;
        RECT 33.850 159.910 33.990 160.610 ;
        RECT 33.790 159.590 34.050 159.910 ;
        RECT 31.590 159.055 33.470 159.425 ;
        RECT 31.030 158.570 31.290 158.890 ;
        RECT 30.570 158.230 30.830 158.550 ;
        RECT 29.650 157.890 29.910 158.210 ;
        RECT 26.890 155.170 27.150 155.490 ;
        RECT 27.350 155.170 27.610 155.490 ;
        RECT 27.410 153.450 27.550 155.170 ;
        RECT 27.350 153.130 27.610 153.450 ;
        RECT 20.910 152.450 21.170 152.770 ;
        RECT 21.830 152.450 22.090 152.770 ;
        RECT 16.590 150.895 18.470 151.265 ;
        RECT 19.990 150.070 20.250 150.390 ;
        RECT 16.590 145.455 18.470 145.825 ;
        RECT 20.050 145.290 20.190 150.070 ;
        RECT 20.970 147.330 21.110 152.450 ;
        RECT 22.290 151.430 22.550 151.750 ;
        RECT 22.350 149.710 22.490 151.430 ;
        RECT 29.710 150.050 29.850 157.890 ;
        RECT 30.630 155.150 30.770 158.230 ;
        RECT 31.950 157.550 32.210 157.870 ;
        RECT 31.030 155.170 31.290 155.490 ;
        RECT 30.570 154.830 30.830 155.150 ;
        RECT 31.090 151.750 31.230 155.170 ;
        RECT 32.010 154.810 32.150 157.550 ;
        RECT 33.330 155.850 33.590 156.170 ;
        RECT 33.390 155.490 33.530 155.850 ;
        RECT 33.330 155.170 33.590 155.490 ;
        RECT 33.790 154.830 34.050 155.150 ;
        RECT 31.950 154.490 32.210 154.810 ;
        RECT 31.590 153.615 33.470 153.985 ;
        RECT 33.330 151.770 33.590 152.090 ;
        RECT 31.030 151.430 31.290 151.750 ;
        RECT 31.090 150.390 31.230 151.430 ;
        RECT 33.390 150.730 33.530 151.770 ;
        RECT 33.330 150.410 33.590 150.730 ;
        RECT 31.030 150.070 31.290 150.390 ;
        RECT 29.650 149.730 29.910 150.050 ;
        RECT 22.290 149.390 22.550 149.710 ;
        RECT 24.590 149.390 24.850 149.710 ;
        RECT 20.910 147.010 21.170 147.330 ;
        RECT 22.350 146.310 22.490 149.390 ;
        RECT 24.650 148.010 24.790 149.390 ;
        RECT 24.590 147.690 24.850 148.010 ;
        RECT 28.270 147.350 28.530 147.670 ;
        RECT 22.750 146.330 23.010 146.650 ;
        RECT 22.290 145.990 22.550 146.310 ;
        RECT 22.810 145.290 22.950 146.330 ;
        RECT 28.330 146.310 28.470 147.350 ;
        RECT 28.270 145.990 28.530 146.310 ;
        RECT 28.730 145.990 28.990 146.310 ;
        RECT 19.990 144.970 20.250 145.290 ;
        RECT 22.750 144.970 23.010 145.290 ;
        RECT 28.790 144.270 28.930 145.990 ;
        RECT 29.710 144.690 29.850 149.730 ;
        RECT 31.090 146.990 31.230 150.070 ;
        RECT 31.590 148.175 33.470 148.545 ;
        RECT 33.850 147.330 33.990 154.830 ;
        RECT 33.790 147.010 34.050 147.330 ;
        RECT 31.030 146.670 31.290 146.990 ;
        RECT 29.710 144.610 30.310 144.690 ;
        RECT 29.710 144.550 30.370 144.610 ;
        RECT 28.730 143.950 28.990 144.270 ;
        RECT 29.710 143.590 29.850 144.550 ;
        RECT 30.110 144.290 30.370 144.550 ;
        RECT 29.650 143.270 29.910 143.590 ;
        RECT 31.590 142.735 33.470 143.105 ;
        RECT 34.310 141.890 34.450 160.870 ;
        RECT 34.710 159.590 34.970 159.910 ;
        RECT 34.770 157.190 34.910 159.590 ;
        RECT 34.710 156.870 34.970 157.190 ;
        RECT 34.770 156.170 34.910 156.870 ;
        RECT 34.710 155.850 34.970 156.170 ;
        RECT 34.710 151.430 34.970 151.750 ;
        RECT 34.250 141.570 34.510 141.890 ;
        RECT 34.770 141.550 34.910 151.430 ;
        RECT 34.710 141.230 34.970 141.550 ;
        RECT 29.190 140.550 29.450 140.870 ;
        RECT 16.590 140.015 18.470 140.385 ;
        RECT 19.070 139.190 19.330 139.510 ;
        RECT 18.610 135.110 18.870 135.430 ;
        RECT 16.590 134.575 18.470 134.945 ;
        RECT 18.670 133.730 18.810 135.110 ;
        RECT 19.130 134.410 19.270 139.190 ;
        RECT 23.210 138.510 23.470 138.830 ;
        RECT 22.290 137.830 22.550 138.150 ;
        RECT 21.370 136.130 21.630 136.450 ;
        RECT 19.070 134.090 19.330 134.410 ;
        RECT 21.430 133.810 21.570 136.130 ;
        RECT 22.350 136.110 22.490 137.830 ;
        RECT 22.290 135.790 22.550 136.110 ;
        RECT 21.830 135.110 22.090 135.430 ;
        RECT 21.890 134.410 22.030 135.110 ;
        RECT 21.830 134.090 22.090 134.410 ;
        RECT 18.610 133.410 18.870 133.730 ;
        RECT 21.430 133.670 22.030 133.810 ;
        RECT 21.890 133.390 22.030 133.670 ;
        RECT 19.530 133.070 19.790 133.390 ;
        RECT 21.830 133.070 22.090 133.390 ;
        RECT 16.590 129.135 18.470 129.505 ;
        RECT 19.590 125.570 19.730 133.070 ;
        RECT 21.890 131.010 22.030 133.070 ;
        RECT 21.830 130.690 22.090 131.010 ;
        RECT 20.910 128.310 21.170 128.630 ;
        RECT 19.530 125.250 19.790 125.570 ;
        RECT 16.590 123.695 18.470 124.065 ;
        RECT 16.590 118.255 18.470 118.625 ;
        RECT 19.590 117.490 19.730 125.250 ;
        RECT 20.970 125.230 21.110 128.310 ;
        RECT 20.910 124.910 21.170 125.230 ;
        RECT 21.890 122.510 22.030 130.690 ;
        RECT 22.350 129.990 22.490 135.790 ;
        RECT 23.270 133.050 23.410 138.510 ;
        RECT 28.270 135.110 28.530 135.430 ;
        RECT 23.210 132.730 23.470 133.050 ;
        RECT 28.330 130.670 28.470 135.110 ;
        RECT 28.730 133.070 28.990 133.390 ;
        RECT 28.790 131.690 28.930 133.070 ;
        RECT 28.730 131.370 28.990 131.690 ;
        RECT 28.270 130.350 28.530 130.670 ;
        RECT 23.210 130.010 23.470 130.330 ;
        RECT 22.290 129.670 22.550 129.990 ;
        RECT 22.750 129.670 23.010 129.990 ;
        RECT 22.350 127.270 22.490 129.670 ;
        RECT 22.290 126.950 22.550 127.270 ;
        RECT 22.810 125.230 22.950 129.670 ;
        RECT 23.270 128.970 23.410 130.010 ;
        RECT 23.210 128.650 23.470 128.970 ;
        RECT 22.750 124.910 23.010 125.230 ;
        RECT 23.270 123.530 23.410 128.650 ;
        RECT 23.670 127.630 23.930 127.950 ;
        RECT 23.730 126.250 23.870 127.630 ;
        RECT 23.670 125.930 23.930 126.250 ;
        RECT 22.290 123.210 22.550 123.530 ;
        RECT 23.210 123.210 23.470 123.530 ;
        RECT 21.830 122.190 22.090 122.510 ;
        RECT 21.890 120.470 22.030 122.190 ;
        RECT 21.830 120.150 22.090 120.470 ;
        RECT 22.350 120.130 22.490 123.210 ;
        RECT 26.430 121.510 26.690 121.830 ;
        RECT 22.290 119.810 22.550 120.130 ;
        RECT 20.910 118.790 21.170 119.110 ;
        RECT 19.130 117.410 19.730 117.490 ;
        RECT 19.070 117.350 19.730 117.410 ;
        RECT 19.070 117.090 19.330 117.350 ;
        RECT 19.590 114.690 19.730 117.350 ;
        RECT 19.530 114.370 19.790 114.690 ;
        RECT 20.970 114.350 21.110 118.790 ;
        RECT 22.350 118.090 22.490 119.810 ;
        RECT 26.490 119.790 26.630 121.510 ;
        RECT 26.430 119.470 26.690 119.790 ;
        RECT 25.050 118.790 25.310 119.110 ;
        RECT 22.290 117.770 22.550 118.090 ;
        RECT 23.210 117.430 23.470 117.750 ;
        RECT 23.270 115.370 23.410 117.430 ;
        RECT 25.110 117.410 25.250 118.790 ;
        RECT 25.050 117.090 25.310 117.410 ;
        RECT 25.510 116.750 25.770 117.070 ;
        RECT 23.210 115.050 23.470 115.370 ;
        RECT 25.570 114.770 25.710 116.750 ;
        RECT 28.270 116.070 28.530 116.390 ;
        RECT 25.570 114.690 26.170 114.770 ;
        RECT 25.510 114.630 26.170 114.690 ;
        RECT 25.510 114.370 25.770 114.630 ;
        RECT 20.910 114.030 21.170 114.350 ;
        RECT 16.590 112.815 18.470 113.185 ;
        RECT 20.910 111.990 21.170 112.310 ;
        RECT 14.010 111.310 14.270 111.630 ;
        RECT 14.070 89.420 14.210 111.310 ;
        RECT 20.970 109.930 21.110 111.990 ;
        RECT 26.030 111.970 26.170 114.630 ;
        RECT 28.330 114.010 28.470 116.070 ;
        RECT 28.270 113.690 28.530 114.010 ;
        RECT 25.970 111.650 26.230 111.970 ;
        RECT 27.350 110.630 27.610 110.950 ;
        RECT 27.410 109.930 27.550 110.630 ;
        RECT 20.910 109.610 21.170 109.930 ;
        RECT 27.350 109.610 27.610 109.930 ;
        RECT 29.250 108.910 29.390 140.550 ;
        RECT 34.710 138.850 34.970 139.170 ;
        RECT 29.650 138.510 29.910 138.830 ;
        RECT 30.110 138.510 30.370 138.830 ;
        RECT 29.710 133.730 29.850 138.510 ;
        RECT 30.170 135.770 30.310 138.510 ;
        RECT 34.250 137.830 34.510 138.150 ;
        RECT 31.590 137.295 33.470 137.665 ;
        RECT 34.310 137.130 34.450 137.830 ;
        RECT 34.250 136.810 34.510 137.130 ;
        RECT 33.790 136.470 34.050 136.790 ;
        RECT 31.030 136.130 31.290 136.450 ;
        RECT 30.110 135.450 30.370 135.770 ;
        RECT 30.570 135.110 30.830 135.430 ;
        RECT 29.650 133.410 29.910 133.730 ;
        RECT 29.710 128.290 29.850 133.410 ;
        RECT 30.630 131.690 30.770 135.110 ;
        RECT 31.090 133.730 31.230 136.130 ;
        RECT 33.330 135.790 33.590 136.110 ;
        RECT 32.410 135.110 32.670 135.430 ;
        RECT 32.470 133.730 32.610 135.110 ;
        RECT 31.030 133.410 31.290 133.730 ;
        RECT 31.950 133.410 32.210 133.730 ;
        RECT 32.410 133.410 32.670 133.730 ;
        RECT 32.010 133.130 32.150 133.410 ;
        RECT 33.390 133.130 33.530 135.790 ;
        RECT 33.850 134.410 33.990 136.470 ;
        RECT 34.770 136.110 34.910 138.850 ;
        RECT 35.230 136.450 35.370 170.470 ;
        RECT 35.690 170.390 36.290 170.530 ;
        RECT 35.690 168.750 35.830 170.390 ;
        RECT 35.630 168.430 35.890 168.750 ;
        RECT 35.690 166.710 35.830 168.430 ;
        RECT 36.610 168.070 36.750 176.590 ;
        RECT 37.070 172.150 37.210 179.310 ;
        RECT 37.530 174.530 37.670 182.370 ;
        RECT 37.990 182.350 38.130 185.090 ;
        RECT 37.930 182.030 38.190 182.350 ;
        RECT 37.990 176.910 38.130 182.030 ;
        RECT 39.310 181.350 39.570 181.670 ;
        RECT 39.370 177.930 39.510 181.350 ;
        RECT 40.690 179.540 40.950 179.630 ;
        RECT 41.210 179.540 41.350 185.090 ;
        RECT 43.450 184.070 43.710 184.390 ;
        RECT 43.910 184.070 44.170 184.390 ;
        RECT 43.510 182.350 43.650 184.070 ;
        RECT 43.970 182.690 44.110 184.070 ;
        RECT 44.890 183.370 45.030 190.190 ;
        RECT 45.810 186.090 45.950 193.250 ;
        RECT 48.970 192.910 49.230 193.230 ;
        RECT 46.210 190.530 46.470 190.850 ;
        RECT 46.270 187.530 46.410 190.530 ;
        RECT 49.030 190.170 49.170 192.910 ;
        RECT 48.970 189.850 49.230 190.170 ;
        RECT 46.590 188.975 48.470 189.345 ;
        RECT 46.670 187.530 46.930 187.790 ;
        RECT 46.270 187.470 46.930 187.530 ;
        RECT 46.270 187.390 46.870 187.470 ;
        RECT 49.030 187.450 49.170 189.850 ;
        RECT 45.750 185.770 46.010 186.090 ;
        RECT 46.270 185.750 46.410 187.390 ;
        RECT 48.970 187.130 49.230 187.450 ;
        RECT 46.210 185.430 46.470 185.750 ;
        RECT 45.290 184.750 45.550 185.070 ;
        RECT 44.830 183.050 45.090 183.370 ;
        RECT 43.910 182.370 44.170 182.690 ;
        RECT 43.450 182.030 43.710 182.350 ;
        RECT 45.350 180.650 45.490 184.750 ;
        RECT 45.750 184.070 46.010 184.390 ;
        RECT 46.210 184.070 46.470 184.390 ;
        RECT 45.810 181.670 45.950 184.070 ;
        RECT 46.270 182.690 46.410 184.070 ;
        RECT 46.590 183.535 48.470 183.905 ;
        RECT 46.210 182.370 46.470 182.690 ;
        RECT 45.750 181.350 46.010 181.670 ;
        RECT 45.290 180.330 45.550 180.650 ;
        RECT 46.270 179.970 46.410 182.370 ;
        RECT 47.130 181.350 47.390 181.670 ;
        RECT 46.670 180.330 46.930 180.650 ;
        RECT 46.730 179.970 46.870 180.330 ;
        RECT 47.190 179.970 47.330 181.350 ;
        RECT 46.210 179.650 46.470 179.970 ;
        RECT 46.670 179.650 46.930 179.970 ;
        RECT 47.130 179.650 47.390 179.970 ;
        RECT 40.220 179.115 40.500 179.485 ;
        RECT 40.690 179.400 41.350 179.540 ;
        RECT 40.690 179.310 40.950 179.400 ;
        RECT 41.600 179.115 41.880 179.485 ;
        RECT 43.910 179.310 44.170 179.630 ;
        RECT 45.290 179.310 45.550 179.630 ;
        RECT 40.290 178.950 40.430 179.115 ;
        RECT 39.770 178.630 40.030 178.950 ;
        RECT 40.230 178.630 40.490 178.950 ;
        RECT 40.690 178.630 40.950 178.950 ;
        RECT 39.310 177.610 39.570 177.930 ;
        RECT 37.930 176.590 38.190 176.910 ;
        RECT 37.990 175.210 38.130 176.590 ;
        RECT 37.930 174.890 38.190 175.210 ;
        RECT 39.830 174.725 39.970 178.630 ;
        RECT 40.750 175.210 40.890 178.630 ;
        RECT 40.690 174.890 40.950 175.210 ;
        RECT 37.470 174.210 37.730 174.530 ;
        RECT 39.760 174.355 40.040 174.725 ;
        RECT 40.230 174.550 40.490 174.870 ;
        RECT 39.830 174.190 39.970 174.355 ;
        RECT 37.930 173.870 38.190 174.190 ;
        RECT 39.770 173.870 40.030 174.190 ;
        RECT 37.010 171.830 37.270 172.150 ;
        RECT 37.990 171.810 38.130 173.870 ;
        RECT 38.850 173.530 39.110 173.850 ;
        RECT 39.310 173.530 39.570 173.850 ;
        RECT 37.930 171.490 38.190 171.810 ;
        RECT 36.550 167.750 36.810 168.070 ;
        RECT 35.630 166.390 35.890 166.710 ;
        RECT 36.610 166.370 36.750 167.750 ;
        RECT 36.550 166.050 36.810 166.370 ;
        RECT 36.610 163.650 36.750 166.050 ;
        RECT 37.930 165.030 38.190 165.350 ;
        RECT 36.550 163.330 36.810 163.650 ;
        RECT 37.990 163.310 38.130 165.030 ;
        RECT 37.930 162.990 38.190 163.310 ;
        RECT 35.630 162.310 35.890 162.630 ;
        RECT 36.090 162.310 36.350 162.630 ;
        RECT 35.690 157.870 35.830 162.310 ;
        RECT 36.150 161.270 36.290 162.310 ;
        RECT 36.090 160.950 36.350 161.270 ;
        RECT 35.630 157.550 35.890 157.870 ;
        RECT 36.150 157.530 36.290 160.950 ;
        RECT 37.470 159.930 37.730 160.250 ;
        RECT 36.090 157.210 36.350 157.530 ;
        RECT 35.630 154.150 35.890 154.470 ;
        RECT 35.690 150.050 35.830 154.150 ;
        RECT 37.530 152.770 37.670 159.930 ;
        RECT 37.010 152.450 37.270 152.770 ;
        RECT 37.470 152.450 37.730 152.770 ;
        RECT 36.550 152.340 36.810 152.430 ;
        RECT 36.150 152.200 36.810 152.340 ;
        RECT 35.630 149.730 35.890 150.050 ;
        RECT 36.150 149.710 36.290 152.200 ;
        RECT 36.550 152.110 36.810 152.200 ;
        RECT 37.070 150.730 37.210 152.450 ;
        RECT 37.010 150.410 37.270 150.730 ;
        RECT 36.090 149.390 36.350 149.710 ;
        RECT 35.630 147.690 35.890 148.010 ;
        RECT 35.690 146.990 35.830 147.690 ;
        RECT 35.630 146.670 35.890 146.990 ;
        RECT 36.150 144.270 36.290 149.390 ;
        RECT 36.550 145.990 36.810 146.310 ;
        RECT 38.390 145.990 38.650 146.310 ;
        RECT 36.090 143.950 36.350 144.270 ;
        RECT 35.630 142.250 35.890 142.570 ;
        RECT 35.690 139.850 35.830 142.250 ;
        RECT 35.630 139.530 35.890 139.850 ;
        RECT 35.630 138.850 35.890 139.170 ;
        RECT 35.170 136.130 35.430 136.450 ;
        RECT 34.710 135.790 34.970 136.110 ;
        RECT 34.250 135.110 34.510 135.430 ;
        RECT 33.790 134.090 34.050 134.410 ;
        RECT 32.010 132.990 33.990 133.130 ;
        RECT 31.030 132.390 31.290 132.710 ;
        RECT 30.570 131.370 30.830 131.690 ;
        RECT 29.650 127.970 29.910 128.290 ;
        RECT 30.110 127.970 30.370 128.290 ;
        RECT 30.170 125.570 30.310 127.970 ;
        RECT 30.110 125.250 30.370 125.570 ;
        RECT 30.570 119.130 30.830 119.450 ;
        RECT 30.630 115.370 30.770 119.130 ;
        RECT 30.570 115.050 30.830 115.370 ;
        RECT 31.090 109.250 31.230 132.390 ;
        RECT 31.590 131.855 33.470 132.225 ;
        RECT 33.850 131.690 33.990 132.990 ;
        RECT 33.790 131.370 34.050 131.690 ;
        RECT 33.790 130.010 34.050 130.330 ;
        RECT 33.850 128.970 33.990 130.010 ;
        RECT 33.790 128.650 34.050 128.970 ;
        RECT 31.590 126.415 33.470 126.785 ;
        RECT 31.590 120.975 33.470 121.345 ;
        RECT 31.590 115.535 33.470 115.905 ;
        RECT 31.590 110.095 33.470 110.465 ;
        RECT 31.030 108.930 31.290 109.250 ;
        RECT 34.310 108.910 34.450 135.110 ;
        RECT 34.710 132.730 34.970 133.050 ;
        RECT 34.770 122.850 34.910 132.730 ;
        RECT 35.690 132.710 35.830 138.850 ;
        RECT 36.150 134.070 36.290 143.950 ;
        RECT 36.610 136.110 36.750 145.990 ;
        RECT 37.930 136.810 38.190 137.130 ;
        RECT 36.550 135.790 36.810 136.110 ;
        RECT 36.090 133.750 36.350 134.070 ;
        RECT 35.630 132.390 35.890 132.710 ;
        RECT 36.150 131.010 36.290 133.750 ;
        RECT 36.090 130.690 36.350 131.010 ;
        RECT 37.470 130.690 37.730 131.010 ;
        RECT 37.530 128.970 37.670 130.690 ;
        RECT 37.470 128.650 37.730 128.970 ;
        RECT 35.630 125.250 35.890 125.570 ;
        RECT 34.710 122.530 34.970 122.850 ;
        RECT 34.770 120.810 34.910 122.530 ;
        RECT 34.710 120.490 34.970 120.810 ;
        RECT 35.690 120.130 35.830 125.250 ;
        RECT 37.990 125.230 38.130 136.810 ;
        RECT 38.450 136.110 38.590 145.990 ;
        RECT 38.910 136.450 39.050 173.530 ;
        RECT 39.370 171.810 39.510 173.530 ;
        RECT 39.310 171.490 39.570 171.810 ;
        RECT 39.770 154.150 40.030 154.470 ;
        RECT 39.310 140.890 39.570 141.210 ;
        RECT 39.370 139.850 39.510 140.890 ;
        RECT 39.310 139.530 39.570 139.850 ;
        RECT 39.830 138.830 39.970 154.150 ;
        RECT 39.770 138.510 40.030 138.830 ;
        RECT 38.850 136.130 39.110 136.450 ;
        RECT 38.390 135.790 38.650 136.110 ;
        RECT 38.390 135.110 38.650 135.430 ;
        RECT 36.550 124.910 36.810 125.230 ;
        RECT 37.930 124.910 38.190 125.230 ;
        RECT 36.610 122.510 36.750 124.910 ;
        RECT 36.550 122.420 36.810 122.510 ;
        RECT 36.150 122.280 36.810 122.420 ;
        RECT 35.630 119.810 35.890 120.130 ;
        RECT 34.710 119.130 34.970 119.450 ;
        RECT 34.770 112.650 34.910 119.130 ;
        RECT 36.150 118.090 36.290 122.280 ;
        RECT 36.550 122.190 36.810 122.280 ;
        RECT 36.550 121.510 36.810 121.830 ;
        RECT 36.090 117.770 36.350 118.090 ;
        RECT 35.170 117.430 35.430 117.750 ;
        RECT 35.230 115.370 35.370 117.430 ;
        RECT 35.170 115.050 35.430 115.370 ;
        RECT 36.610 114.350 36.750 121.510 ;
        RECT 37.470 119.470 37.730 119.790 ;
        RECT 37.530 115.370 37.670 119.470 ;
        RECT 37.470 115.050 37.730 115.370 ;
        RECT 35.630 114.030 35.890 114.350 ;
        RECT 36.550 114.030 36.810 114.350 ;
        RECT 35.690 113.670 35.830 114.030 ;
        RECT 35.630 113.350 35.890 113.670 ;
        RECT 34.710 112.330 34.970 112.650 ;
        RECT 35.690 111.970 35.830 113.350 ;
        RECT 35.630 111.650 35.890 111.970 ;
        RECT 36.550 110.970 36.810 111.290 ;
        RECT 29.190 108.590 29.450 108.910 ;
        RECT 34.250 108.590 34.510 108.910 ;
        RECT 27.350 108.250 27.610 108.570 ;
        RECT 23.210 107.910 23.470 108.230 ;
        RECT 16.590 107.375 18.470 107.745 ;
        RECT 23.270 106.870 23.410 107.910 ;
        RECT 23.210 106.550 23.470 106.870 ;
        RECT 18.610 105.870 18.870 106.190 ;
        RECT 16.590 101.935 18.470 102.305 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 18.670 88.250 18.810 105.870 ;
        RECT 27.410 103.470 27.550 108.250 ;
        RECT 31.490 107.910 31.750 108.230 ;
        RECT 31.950 107.910 32.210 108.230 ;
        RECT 33.790 107.910 34.050 108.230 ;
        RECT 31.550 106.870 31.690 107.910 ;
        RECT 32.010 107.210 32.150 107.910 ;
        RECT 31.950 106.890 32.210 107.210 ;
        RECT 31.490 106.550 31.750 106.870 ;
        RECT 28.730 105.870 28.990 106.190 ;
        RECT 30.110 105.870 30.370 106.190 ;
        RECT 28.790 104.490 28.930 105.870 ;
        RECT 28.730 104.170 28.990 104.490 ;
        RECT 27.350 103.150 27.610 103.470 ;
        RECT 27.810 102.470 28.070 102.790 ;
        RECT 27.870 101.090 28.010 102.470 ;
        RECT 27.810 100.770 28.070 101.090 ;
        RECT 25.970 100.430 26.230 100.750 ;
        RECT 19.910 88.250 21.130 89.850 ;
        RECT 26.030 88.990 26.170 100.430 ;
        RECT 18.670 88.110 21.130 88.250 ;
        RECT 19.910 85.980 21.130 88.110 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 30.170 88.250 30.310 105.870 ;
        RECT 31.590 104.655 33.470 105.025 ;
        RECT 33.850 101.430 33.990 107.910 ;
        RECT 36.610 106.530 36.750 110.970 ;
        RECT 38.450 106.530 38.590 135.110 ;
        RECT 40.290 133.730 40.430 174.550 ;
        RECT 40.750 171.810 40.890 174.890 ;
        RECT 41.670 173.850 41.810 179.115 ;
        RECT 42.070 178.630 42.330 178.950 ;
        RECT 41.610 173.530 41.870 173.850 ;
        RECT 40.690 171.490 40.950 171.810 ;
        RECT 40.750 169.430 40.890 171.490 ;
        RECT 41.150 170.470 41.410 170.790 ;
        RECT 40.690 169.110 40.950 169.430 ;
        RECT 40.750 155.830 40.890 169.110 ;
        RECT 40.690 155.510 40.950 155.830 ;
        RECT 40.690 148.710 40.950 149.030 ;
        RECT 40.750 133.730 40.890 148.710 ;
        RECT 41.210 139.510 41.350 170.470 ;
        RECT 42.130 159.770 42.270 178.630 ;
        RECT 43.450 176.930 43.710 177.250 ;
        RECT 42.530 175.910 42.790 176.230 ;
        RECT 42.590 171.810 42.730 175.910 ;
        RECT 43.510 174.190 43.650 176.930 ;
        RECT 43.970 174.190 44.110 179.310 ;
        RECT 44.370 178.630 44.630 178.950 ;
        RECT 44.430 174.190 44.570 178.630 ;
        RECT 45.350 177.250 45.490 179.310 ;
        RECT 46.730 179.200 46.870 179.650 ;
        RECT 46.270 179.060 46.870 179.200 ;
        RECT 45.750 178.630 46.010 178.950 ;
        RECT 45.810 177.930 45.950 178.630 ;
        RECT 45.750 177.610 46.010 177.930 ;
        RECT 45.290 176.930 45.550 177.250 ;
        RECT 45.350 174.530 45.490 176.930 ;
        RECT 46.270 175.210 46.410 179.060 ;
        RECT 46.590 178.095 48.470 178.465 ;
        RECT 47.590 176.930 47.850 177.250 ;
        RECT 48.970 176.930 49.230 177.250 ;
        RECT 46.210 174.890 46.470 175.210 ;
        RECT 45.290 174.210 45.550 174.530 ;
        RECT 43.450 173.870 43.710 174.190 ;
        RECT 43.910 173.870 44.170 174.190 ;
        RECT 44.370 173.870 44.630 174.190 ;
        RECT 44.430 172.490 44.570 173.870 ;
        RECT 47.650 173.850 47.790 176.930 ;
        RECT 45.290 173.530 45.550 173.850 ;
        RECT 47.590 173.530 47.850 173.850 ;
        RECT 44.370 172.170 44.630 172.490 ;
        RECT 42.530 171.490 42.790 171.810 ;
        RECT 43.900 168.915 44.180 169.285 ;
        RECT 43.970 168.750 44.110 168.915 ;
        RECT 43.910 168.430 44.170 168.750 ;
        RECT 42.990 165.710 43.250 166.030 ;
        RECT 42.530 165.030 42.790 165.350 ;
        RECT 42.590 161.610 42.730 165.030 ;
        RECT 42.530 161.290 42.790 161.610 ;
        RECT 42.130 159.630 42.730 159.770 ;
        RECT 41.610 157.550 41.870 157.870 ;
        RECT 41.670 156.170 41.810 157.550 ;
        RECT 42.070 156.870 42.330 157.190 ;
        RECT 41.610 155.850 41.870 156.170 ;
        RECT 41.600 155.315 41.880 155.685 ;
        RECT 41.610 155.170 41.870 155.315 ;
        RECT 41.610 151.430 41.870 151.750 ;
        RECT 41.670 150.050 41.810 151.430 ;
        RECT 41.610 149.730 41.870 150.050 ;
        RECT 41.670 146.310 41.810 149.730 ;
        RECT 41.610 145.990 41.870 146.310 ;
        RECT 41.150 139.190 41.410 139.510 ;
        RECT 42.130 136.110 42.270 156.870 ;
        RECT 42.070 135.790 42.330 136.110 ;
        RECT 42.590 133.730 42.730 159.630 ;
        RECT 43.050 157.870 43.190 165.710 ;
        RECT 42.990 157.550 43.250 157.870 ;
        RECT 44.830 157.550 45.090 157.870 ;
        RECT 42.990 156.870 43.250 157.190 ;
        RECT 43.050 155.685 43.190 156.870 ;
        RECT 44.890 156.170 45.030 157.550 ;
        RECT 44.830 155.850 45.090 156.170 ;
        RECT 42.980 155.315 43.260 155.685 ;
        RECT 43.050 155.060 43.190 155.315 ;
        RECT 43.450 155.060 43.710 155.150 ;
        RECT 43.050 154.920 43.710 155.060 ;
        RECT 43.450 154.830 43.710 154.920 ;
        RECT 43.450 154.150 43.710 154.470 ;
        RECT 44.830 154.150 45.090 154.470 ;
        RECT 42.990 151.770 43.250 152.090 ;
        RECT 43.050 150.050 43.190 151.770 ;
        RECT 42.990 149.730 43.250 150.050 ;
        RECT 43.050 146.650 43.190 149.730 ;
        RECT 42.990 146.330 43.250 146.650 ;
        RECT 43.510 133.730 43.650 154.150 ;
        RECT 44.370 152.285 44.630 152.430 ;
        RECT 44.360 151.915 44.640 152.285 ;
        RECT 43.910 148.710 44.170 149.030 ;
        RECT 40.230 133.410 40.490 133.730 ;
        RECT 40.690 133.410 40.950 133.730 ;
        RECT 42.530 133.410 42.790 133.730 ;
        RECT 43.450 133.410 43.710 133.730 ;
        RECT 43.970 133.130 44.110 148.710 ;
        RECT 44.430 146.990 44.570 151.915 ;
        RECT 44.890 150.050 45.030 154.150 ;
        RECT 44.830 149.730 45.090 150.050 ;
        RECT 44.370 146.670 44.630 146.990 ;
        RECT 44.830 141.910 45.090 142.230 ;
        RECT 44.370 136.810 44.630 137.130 ;
        RECT 43.510 132.990 44.110 133.130 ;
        RECT 39.310 132.390 39.570 132.710 ;
        RECT 40.230 132.390 40.490 132.710 ;
        RECT 41.150 132.390 41.410 132.710 ;
        RECT 42.990 132.390 43.250 132.710 ;
        RECT 39.370 128.290 39.510 132.390 ;
        RECT 39.770 131.030 40.030 131.350 ;
        RECT 39.310 127.970 39.570 128.290 ;
        RECT 39.830 124.890 39.970 131.030 ;
        RECT 40.290 125.230 40.430 132.390 ;
        RECT 40.230 124.910 40.490 125.230 ;
        RECT 39.770 124.570 40.030 124.890 ;
        RECT 39.770 118.790 40.030 119.110 ;
        RECT 38.850 116.750 39.110 117.070 ;
        RECT 38.910 115.370 39.050 116.750 ;
        RECT 38.850 115.050 39.110 115.370 ;
        RECT 39.830 114.350 39.970 118.790 ;
        RECT 39.770 114.030 40.030 114.350 ;
        RECT 40.690 108.250 40.950 108.570 ;
        RECT 40.750 106.870 40.890 108.250 ;
        RECT 40.690 106.550 40.950 106.870 ;
        RECT 41.210 106.530 41.350 132.390 ;
        RECT 42.530 129.670 42.790 129.990 ;
        RECT 42.590 128.630 42.730 129.670 ;
        RECT 42.530 128.310 42.790 128.630 ;
        RECT 42.530 127.630 42.790 127.950 ;
        RECT 42.070 124.910 42.330 125.230 ;
        RECT 41.610 122.190 41.870 122.510 ;
        RECT 41.670 119.790 41.810 122.190 ;
        RECT 41.610 119.470 41.870 119.790 ;
        RECT 42.130 119.110 42.270 124.910 ;
        RECT 42.590 123.530 42.730 127.630 ;
        RECT 43.050 124.890 43.190 132.390 ;
        RECT 43.510 128.970 43.650 132.990 ;
        RECT 43.910 132.390 44.170 132.710 ;
        RECT 43.450 128.650 43.710 128.970 ;
        RECT 42.990 124.570 43.250 124.890 ;
        RECT 42.530 123.210 42.790 123.530 ;
        RECT 43.450 121.850 43.710 122.170 ;
        RECT 43.510 120.130 43.650 121.850 ;
        RECT 43.450 119.810 43.710 120.130 ;
        RECT 42.070 118.790 42.330 119.110 ;
        RECT 42.130 118.090 42.270 118.790 ;
        RECT 42.070 117.770 42.330 118.090 ;
        RECT 42.130 114.010 42.270 117.770 ;
        RECT 42.990 117.430 43.250 117.750 ;
        RECT 43.050 115.370 43.190 117.430 ;
        RECT 42.990 115.050 43.250 115.370 ;
        RECT 43.510 115.030 43.650 119.810 ;
        RECT 43.450 114.710 43.710 115.030 ;
        RECT 42.070 113.690 42.330 114.010 ;
        RECT 43.970 111.470 44.110 132.390 ;
        RECT 44.430 125.230 44.570 136.810 ;
        RECT 44.890 128.970 45.030 141.910 ;
        RECT 45.350 136.450 45.490 173.530 ;
        RECT 46.590 172.655 48.470 173.025 ;
        RECT 49.030 172.490 49.170 176.930 ;
        RECT 49.490 172.490 49.630 194.020 ;
        RECT 50.350 193.930 50.610 194.020 ;
        RECT 53.170 193.910 53.310 194.950 ;
        RECT 53.110 193.590 53.370 193.910 ;
        RECT 50.350 192.910 50.610 193.230 ;
        RECT 50.410 191.530 50.550 192.910 ;
        RECT 54.030 192.230 54.290 192.550 ;
        RECT 50.350 191.210 50.610 191.530 ;
        RECT 52.190 190.530 52.450 190.850 ;
        RECT 49.890 186.790 50.150 187.110 ;
        RECT 49.950 183.370 50.090 186.790 ;
        RECT 49.890 183.050 50.150 183.370 ;
        RECT 49.890 182.030 50.150 182.350 ;
        RECT 49.950 180.650 50.090 182.030 ;
        RECT 49.890 180.330 50.150 180.650 ;
        RECT 52.250 179.970 52.390 190.530 ;
        RECT 54.090 190.510 54.230 192.230 ;
        RECT 54.030 190.190 54.290 190.510 ;
        RECT 57.770 189.830 57.910 194.950 ;
        RECT 61.590 191.695 63.470 192.065 ;
        RECT 63.750 191.190 63.890 202.090 ;
        RECT 64.670 201.050 64.810 203.110 ;
        RECT 64.610 200.730 64.870 201.050 ;
        RECT 64.610 197.670 64.870 197.990 ;
        RECT 63.690 190.870 63.950 191.190 ;
        RECT 59.090 190.530 59.350 190.850 ;
        RECT 57.710 189.510 57.970 189.830 ;
        RECT 57.770 188.810 57.910 189.510 ;
        RECT 57.710 188.490 57.970 188.810 ;
        RECT 55.410 187.810 55.670 188.130 ;
        RECT 56.330 187.810 56.590 188.130 ;
        RECT 55.470 187.645 55.610 187.810 ;
        RECT 55.400 187.275 55.680 187.645 ;
        RECT 55.870 181.350 56.130 181.670 ;
        RECT 52.190 179.650 52.450 179.970 ;
        RECT 54.030 179.650 54.290 179.970 ;
        RECT 50.350 178.630 50.610 178.950 ;
        RECT 50.410 177.250 50.550 178.630 ;
        RECT 52.250 177.590 52.390 179.650 ;
        RECT 53.570 178.970 53.830 179.290 ;
        RECT 53.630 177.930 53.770 178.970 ;
        RECT 53.570 177.610 53.830 177.930 ;
        RECT 52.190 177.270 52.450 177.590 ;
        RECT 50.350 176.930 50.610 177.250 ;
        RECT 50.810 176.250 51.070 176.570 ;
        RECT 49.890 175.910 50.150 176.230 ;
        RECT 48.970 172.170 49.230 172.490 ;
        RECT 49.430 172.170 49.690 172.490 ;
        RECT 49.030 171.810 49.170 172.170 ;
        RECT 47.130 171.490 47.390 171.810 ;
        RECT 48.970 171.490 49.230 171.810 ;
        RECT 49.430 171.490 49.690 171.810 ;
        RECT 45.750 170.470 46.010 170.790 ;
        RECT 45.810 159.770 45.950 170.470 ;
        RECT 47.190 169.770 47.330 171.490 ;
        RECT 49.490 171.130 49.630 171.490 ;
        RECT 49.430 170.810 49.690 171.130 ;
        RECT 47.130 169.450 47.390 169.770 ;
        RECT 46.590 167.215 48.470 167.585 ;
        RECT 49.430 165.030 49.690 165.350 ;
        RECT 48.970 162.990 49.230 163.310 ;
        RECT 46.210 162.650 46.470 162.970 ;
        RECT 46.270 161.610 46.410 162.650 ;
        RECT 46.590 161.775 48.470 162.145 ;
        RECT 49.030 161.610 49.170 162.990 ;
        RECT 49.490 161.610 49.630 165.030 ;
        RECT 46.210 161.290 46.470 161.610 ;
        RECT 48.970 161.290 49.230 161.610 ;
        RECT 49.430 161.290 49.690 161.610 ;
        RECT 49.430 160.610 49.690 160.930 ;
        RECT 48.970 160.270 49.230 160.590 ;
        RECT 45.810 159.630 46.410 159.770 ;
        RECT 45.750 156.870 46.010 157.190 ;
        RECT 45.810 141.550 45.950 156.870 ;
        RECT 46.270 141.890 46.410 159.630 ;
        RECT 46.590 156.335 48.470 156.705 ;
        RECT 49.030 156.170 49.170 160.270 ;
        RECT 49.490 158.890 49.630 160.610 ;
        RECT 49.430 158.570 49.690 158.890 ;
        RECT 49.950 157.610 50.090 175.910 ;
        RECT 50.870 172.490 51.010 176.250 ;
        RECT 54.090 175.210 54.230 179.650 ;
        RECT 55.930 177.590 56.070 181.350 ;
        RECT 56.390 180.310 56.530 187.810 ;
        RECT 59.150 187.450 59.290 190.530 ;
        RECT 60.010 189.850 60.270 190.170 ;
        RECT 60.070 188.810 60.210 189.850 ;
        RECT 61.850 189.510 62.110 189.830 ;
        RECT 60.010 188.490 60.270 188.810 ;
        RECT 61.910 187.790 62.050 189.510 ;
        RECT 61.850 187.470 62.110 187.790 ;
        RECT 59.090 187.130 59.350 187.450 ;
        RECT 59.150 185.410 59.290 187.130 ;
        RECT 64.670 186.850 64.810 197.670 ;
        RECT 66.050 193.570 66.190 204.130 ;
        RECT 72.950 203.430 73.090 206.510 ;
        RECT 72.890 203.110 73.150 203.430 ;
        RECT 66.450 202.090 66.710 202.410 ;
        RECT 65.990 193.250 66.250 193.570 ;
        RECT 65.530 192.230 65.790 192.550 ;
        RECT 65.590 190.170 65.730 192.230 ;
        RECT 65.530 189.850 65.790 190.170 ;
        RECT 66.050 189.830 66.190 193.250 ;
        RECT 65.990 189.510 66.250 189.830 ;
        RECT 65.530 187.470 65.790 187.790 ;
        RECT 64.210 186.710 64.810 186.850 ;
        RECT 61.590 186.255 63.470 186.625 ;
        RECT 60.470 185.430 60.730 185.750 ;
        RECT 59.090 185.090 59.350 185.410 ;
        RECT 57.710 184.410 57.970 184.730 ;
        RECT 57.770 183.370 57.910 184.410 ;
        RECT 57.710 183.050 57.970 183.370 ;
        RECT 59.150 182.690 59.290 185.090 ;
        RECT 60.530 182.690 60.670 185.430 ;
        RECT 59.090 182.370 59.350 182.690 ;
        RECT 60.470 182.370 60.730 182.690 ;
        RECT 56.330 179.990 56.590 180.310 ;
        RECT 55.870 177.270 56.130 177.590 ;
        RECT 54.030 174.890 54.290 175.210 ;
        RECT 54.090 174.530 54.230 174.890 ;
        RECT 53.570 174.210 53.830 174.530 ;
        RECT 54.030 174.210 54.290 174.530 ;
        RECT 53.110 173.530 53.370 173.850 ;
        RECT 50.810 172.170 51.070 172.490 ;
        RECT 50.870 171.810 51.010 172.170 ;
        RECT 53.170 171.810 53.310 173.530 ;
        RECT 53.630 171.810 53.770 174.210 ;
        RECT 56.390 174.190 56.530 179.990 ;
        RECT 57.710 178.630 57.970 178.950 ;
        RECT 57.770 174.530 57.910 178.630 ;
        RECT 59.150 176.910 59.290 182.370 ;
        RECT 59.090 176.590 59.350 176.910 ;
        RECT 57.710 174.210 57.970 174.530 ;
        RECT 54.480 173.675 54.760 174.045 ;
        RECT 56.330 173.870 56.590 174.190 ;
        RECT 54.550 172.490 54.690 173.675 ;
        RECT 56.790 173.190 57.050 173.510 ;
        RECT 54.490 172.170 54.750 172.490 ;
        RECT 54.550 171.810 54.690 172.170 ;
        RECT 56.850 172.150 56.990 173.190 ;
        RECT 56.790 171.830 57.050 172.150 ;
        RECT 60.530 171.810 60.670 182.370 ;
        RECT 61.590 180.815 63.470 181.185 ;
        RECT 60.990 177.930 62.050 178.010 ;
        RECT 60.990 177.870 62.110 177.930 ;
        RECT 60.990 177.590 61.130 177.870 ;
        RECT 61.850 177.610 62.110 177.870 ;
        RECT 60.930 177.270 61.190 177.590 ;
        RECT 63.690 176.590 63.950 176.910 ;
        RECT 61.590 175.375 63.470 175.745 ;
        RECT 63.750 175.210 63.890 176.590 ;
        RECT 63.690 174.890 63.950 175.210 ;
        RECT 60.930 173.530 61.190 173.850 ;
        RECT 62.760 173.675 63.040 174.045 ;
        RECT 60.990 172.490 61.130 173.530 ;
        RECT 62.830 173.510 62.970 173.675 ;
        RECT 62.770 173.190 63.030 173.510 ;
        RECT 60.930 172.170 61.190 172.490 ;
        RECT 50.810 171.490 51.070 171.810 ;
        RECT 53.110 171.490 53.370 171.810 ;
        RECT 53.570 171.490 53.830 171.810 ;
        RECT 54.490 171.490 54.750 171.810 ;
        RECT 60.470 171.490 60.730 171.810 ;
        RECT 52.190 170.470 52.450 170.790 ;
        RECT 50.810 166.390 51.070 166.710 ;
        RECT 50.870 164.330 51.010 166.390 ;
        RECT 50.810 164.010 51.070 164.330 ;
        RECT 50.350 158.570 50.610 158.890 ;
        RECT 50.410 158.210 50.550 158.570 ;
        RECT 50.350 157.890 50.610 158.210 ;
        RECT 49.490 157.470 50.090 157.610 ;
        RECT 48.970 155.850 49.230 156.170 ;
        RECT 46.670 155.170 46.930 155.490 ;
        RECT 46.730 154.810 46.870 155.170 ;
        RECT 46.670 154.490 46.930 154.810 ;
        RECT 48.970 154.150 49.230 154.470 ;
        RECT 46.590 150.895 48.470 151.265 ;
        RECT 49.030 150.130 49.170 154.150 ;
        RECT 48.570 149.990 49.170 150.130 ;
        RECT 49.490 150.050 49.630 157.470 ;
        RECT 49.890 156.870 50.150 157.190 ;
        RECT 49.950 150.050 50.090 156.870 ;
        RECT 50.350 155.850 50.610 156.170 ;
        RECT 50.410 151.750 50.550 155.850 ;
        RECT 50.810 152.110 51.070 152.430 ;
        RECT 50.350 151.430 50.610 151.750 ;
        RECT 48.570 146.990 48.710 149.990 ;
        RECT 49.430 149.730 49.690 150.050 ;
        RECT 49.890 149.730 50.150 150.050 ;
        RECT 50.350 149.390 50.610 149.710 ;
        RECT 50.410 148.010 50.550 149.390 ;
        RECT 48.970 147.690 49.230 148.010 ;
        RECT 50.350 147.690 50.610 148.010 ;
        RECT 48.510 146.670 48.770 146.990 ;
        RECT 46.590 145.455 48.470 145.825 ;
        RECT 49.030 144.010 49.170 147.690 ;
        RECT 49.430 145.990 49.690 146.310 ;
        RECT 49.490 144.610 49.630 145.990 ;
        RECT 50.870 145.290 51.010 152.110 ;
        RECT 51.270 148.710 51.530 149.030 ;
        RECT 51.330 146.650 51.470 148.710 ;
        RECT 52.250 147.330 52.390 170.470 ;
        RECT 53.110 166.390 53.370 166.710 ;
        RECT 53.170 163.310 53.310 166.390 ;
        RECT 54.030 165.710 54.290 166.030 ;
        RECT 54.490 165.710 54.750 166.030 ;
        RECT 57.250 165.710 57.510 166.030 ;
        RECT 53.110 162.990 53.370 163.310 ;
        RECT 52.650 162.310 52.910 162.630 ;
        RECT 52.710 158.890 52.850 162.310 ;
        RECT 54.090 161.610 54.230 165.710 ;
        RECT 54.550 164.330 54.690 165.710 ;
        RECT 54.490 164.010 54.750 164.330 ;
        RECT 57.310 163.990 57.450 165.710 ;
        RECT 58.630 165.030 58.890 165.350 ;
        RECT 57.250 163.670 57.510 163.990 ;
        RECT 58.690 162.970 58.830 165.030 ;
        RECT 60.530 163.650 60.670 171.490 ;
        RECT 61.590 169.935 63.470 170.305 ;
        RECT 61.390 166.050 61.650 166.370 ;
        RECT 61.450 165.770 61.590 166.050 ;
        RECT 60.990 165.630 61.590 165.770 ;
        RECT 63.690 165.710 63.950 166.030 ;
        RECT 60.990 163.730 61.130 165.630 ;
        RECT 61.590 164.495 63.470 164.865 ;
        RECT 61.390 164.010 61.650 164.330 ;
        RECT 61.450 163.730 61.590 164.010 ;
        RECT 60.470 163.330 60.730 163.650 ;
        RECT 60.990 163.590 61.590 163.730 ;
        RECT 58.630 162.650 58.890 162.970 ;
        RECT 54.030 161.290 54.290 161.610 ;
        RECT 53.110 159.930 53.370 160.250 ;
        RECT 52.650 158.570 52.910 158.890 ;
        RECT 52.710 157.870 52.850 158.570 ;
        RECT 52.650 157.550 52.910 157.870 ;
        RECT 53.170 157.190 53.310 159.930 ;
        RECT 53.570 157.550 53.830 157.870 ;
        RECT 56.790 157.550 57.050 157.870 ;
        RECT 60.990 157.780 61.130 163.590 ;
        RECT 63.750 163.310 63.890 165.710 ;
        RECT 63.690 162.990 63.950 163.310 ;
        RECT 62.310 162.650 62.570 162.970 ;
        RECT 62.370 161.610 62.510 162.650 ;
        RECT 62.310 161.290 62.570 161.610 ;
        RECT 61.590 159.055 63.470 159.425 ;
        RECT 62.770 157.780 63.030 157.870 ;
        RECT 60.990 157.640 63.030 157.780 ;
        RECT 62.770 157.550 63.030 157.640 ;
        RECT 53.110 156.870 53.370 157.190 ;
        RECT 53.170 155.830 53.310 156.870 ;
        RECT 53.110 155.510 53.370 155.830 ;
        RECT 53.630 155.490 53.770 157.550 ;
        RECT 53.570 155.170 53.830 155.490 ;
        RECT 53.570 154.150 53.830 154.470 ;
        RECT 54.030 154.150 54.290 154.470 ;
        RECT 53.630 150.050 53.770 154.150 ;
        RECT 54.090 153.110 54.230 154.150 ;
        RECT 54.030 152.790 54.290 153.110 ;
        RECT 56.850 152.430 56.990 157.550 ;
        RECT 58.630 156.870 58.890 157.190 ;
        RECT 58.690 155.830 58.830 156.870 ;
        RECT 58.630 155.510 58.890 155.830 ;
        RECT 63.750 155.490 63.890 162.990 ;
        RECT 63.690 155.170 63.950 155.490 ;
        RECT 60.930 154.830 61.190 155.150 ;
        RECT 56.790 152.110 57.050 152.430 ;
        RECT 58.630 151.430 58.890 151.750 ;
        RECT 58.690 150.050 58.830 151.430 ;
        RECT 60.990 150.730 61.130 154.830 ;
        RECT 61.590 153.615 63.470 153.985 ;
        RECT 64.210 152.770 64.350 186.710 ;
        RECT 65.590 179.630 65.730 187.470 ;
        RECT 65.530 179.310 65.790 179.630 ;
        RECT 65.990 178.630 66.250 178.950 ;
        RECT 66.050 177.445 66.190 178.630 ;
        RECT 65.980 177.075 66.260 177.445 ;
        RECT 65.070 176.250 65.330 176.570 ;
        RECT 64.610 175.910 64.870 176.230 ;
        RECT 64.670 174.530 64.810 175.910 ;
        RECT 65.130 174.725 65.270 176.250 ;
        RECT 65.990 174.890 66.250 175.210 ;
        RECT 64.610 174.210 64.870 174.530 ;
        RECT 65.060 174.355 65.340 174.725 ;
        RECT 66.050 174.530 66.190 174.890 ;
        RECT 65.990 174.210 66.250 174.530 ;
        RECT 64.610 173.530 64.870 173.850 ;
        RECT 64.670 172.490 64.810 173.530 ;
        RECT 64.610 172.170 64.870 172.490 ;
        RECT 66.510 166.030 66.650 202.090 ;
        RECT 72.950 201.730 73.090 203.110 ;
        RECT 72.890 201.410 73.150 201.730 ;
        RECT 71.510 200.390 71.770 200.710 ;
        RECT 72.430 200.390 72.690 200.710 ;
        RECT 71.570 199.010 71.710 200.390 ;
        RECT 68.290 198.690 68.550 199.010 ;
        RECT 71.510 198.690 71.770 199.010 ;
        RECT 68.350 196.970 68.490 198.690 ;
        RECT 72.490 197.990 72.630 200.390 ;
        RECT 73.410 198.330 73.550 207.190 ;
        RECT 79.330 206.850 79.590 207.170 ;
        RECT 73.810 205.830 74.070 206.150 ;
        RECT 75.650 205.830 75.910 206.150 ;
        RECT 73.870 205.130 74.010 205.830 ;
        RECT 73.810 204.810 74.070 205.130 ;
        RECT 75.710 204.790 75.850 205.830 ;
        RECT 76.590 205.295 78.470 205.665 ;
        RECT 75.650 204.470 75.910 204.790 ;
        RECT 73.810 203.110 74.070 203.430 ;
        RECT 73.870 201.390 74.010 203.110 ;
        RECT 76.110 201.750 76.370 202.070 ;
        RECT 74.270 201.410 74.530 201.730 ;
        RECT 73.810 201.070 74.070 201.390 ;
        RECT 73.870 199.690 74.010 201.070 ;
        RECT 73.810 199.370 74.070 199.690 ;
        RECT 74.330 199.350 74.470 201.410 ;
        RECT 74.730 200.730 74.990 201.050 ;
        RECT 75.190 200.730 75.450 201.050 ;
        RECT 74.790 199.690 74.930 200.730 ;
        RECT 74.730 199.370 74.990 199.690 ;
        RECT 74.270 199.030 74.530 199.350 ;
        RECT 72.890 198.010 73.150 198.330 ;
        RECT 73.350 198.010 73.610 198.330 ;
        RECT 72.430 197.670 72.690 197.990 ;
        RECT 68.290 196.650 68.550 196.970 ;
        RECT 69.670 196.650 69.930 196.970 ;
        RECT 68.750 195.630 69.010 195.950 ;
        RECT 68.810 193.570 68.950 195.630 ;
        RECT 68.750 193.250 69.010 193.570 ;
        RECT 69.730 190.250 69.870 196.650 ;
        RECT 72.490 196.290 72.630 197.670 ;
        RECT 72.950 196.290 73.090 198.010 ;
        RECT 73.410 196.970 73.550 198.010 ;
        RECT 73.350 196.650 73.610 196.970 ;
        RECT 70.130 195.970 70.390 196.290 ;
        RECT 72.430 195.970 72.690 196.290 ;
        RECT 72.890 195.970 73.150 196.290 ;
        RECT 70.190 192.550 70.330 195.970 ;
        RECT 71.510 195.290 71.770 195.610 ;
        RECT 71.570 194.250 71.710 195.290 ;
        RECT 71.510 193.930 71.770 194.250 ;
        RECT 72.490 193.910 72.630 195.970 ;
        RECT 72.430 193.590 72.690 193.910 ;
        RECT 72.950 193.570 73.090 195.970 ;
        RECT 72.890 193.250 73.150 193.570 ;
        RECT 70.130 192.230 70.390 192.550 ;
        RECT 72.430 192.460 72.690 192.550 ;
        RECT 72.030 192.320 72.690 192.460 ;
        RECT 71.050 190.530 71.310 190.850 ;
        RECT 71.110 190.250 71.250 190.530 ;
        RECT 69.730 190.110 71.250 190.250 ;
        RECT 69.670 189.510 69.930 189.830 ;
        RECT 67.830 185.090 68.090 185.410 ;
        RECT 67.890 182.690 68.030 185.090 ;
        RECT 67.830 182.370 68.090 182.690 ;
        RECT 69.210 181.350 69.470 181.670 ;
        RECT 67.370 179.990 67.630 180.310 ;
        RECT 67.430 179.485 67.570 179.990 ;
        RECT 67.360 179.115 67.640 179.485 ;
        RECT 68.290 179.370 68.550 179.630 ;
        RECT 68.290 179.310 68.950 179.370 ;
        RECT 68.350 179.230 68.950 179.310 ;
        RECT 68.810 177.250 68.950 179.230 ;
        RECT 69.270 177.250 69.410 181.350 ;
        RECT 68.750 176.930 69.010 177.250 ;
        RECT 69.210 176.930 69.470 177.250 ;
        RECT 68.810 176.230 68.950 176.930 ;
        RECT 67.830 175.910 68.090 176.230 ;
        RECT 68.750 175.910 69.010 176.230 ;
        RECT 67.890 175.210 68.030 175.910 ;
        RECT 67.830 174.890 68.090 175.210 ;
        RECT 69.730 174.530 69.870 189.510 ;
        RECT 72.030 187.790 72.170 192.320 ;
        RECT 72.430 192.230 72.690 192.320 ;
        RECT 72.950 190.930 73.090 193.250 ;
        RECT 72.490 190.790 73.090 190.930 ;
        RECT 71.970 187.470 72.230 187.790 ;
        RECT 71.050 185.430 71.310 185.750 ;
        RECT 71.110 183.370 71.250 185.430 ;
        RECT 71.050 183.050 71.310 183.370 ;
        RECT 71.510 183.050 71.770 183.370 ;
        RECT 71.570 182.690 71.710 183.050 ;
        RECT 71.510 182.370 71.770 182.690 ;
        RECT 72.030 182.600 72.170 187.470 ;
        RECT 72.490 184.730 72.630 190.790 ;
        RECT 72.890 190.190 73.150 190.510 ;
        RECT 72.950 188.810 73.090 190.190 ;
        RECT 73.410 190.170 73.550 196.650 ;
        RECT 74.330 195.950 74.470 199.030 ;
        RECT 74.270 195.630 74.530 195.950 ;
        RECT 74.330 190.510 74.470 195.630 ;
        RECT 75.250 195.610 75.390 200.730 ;
        RECT 75.650 200.390 75.910 200.710 ;
        RECT 75.710 198.670 75.850 200.390 ;
        RECT 76.170 199.690 76.310 201.750 ;
        RECT 78.870 201.410 79.130 201.730 ;
        RECT 76.590 199.855 78.470 200.225 ;
        RECT 76.110 199.370 76.370 199.690 ;
        RECT 78.930 199.010 79.070 201.410 ;
        RECT 79.390 201.050 79.530 206.850 ;
        RECT 106.590 205.295 108.470 205.665 ;
        RECT 83.470 204.470 83.730 204.790 ;
        RECT 79.330 200.730 79.590 201.050 ;
        RECT 79.390 199.690 79.530 200.730 ;
        RECT 83.530 199.690 83.670 204.470 ;
        RECT 88.070 203.790 88.330 204.110 ;
        RECT 84.390 201.410 84.650 201.730 ;
        RECT 84.450 199.690 84.590 201.410 ;
        RECT 88.130 201.390 88.270 203.790 ;
        RECT 91.590 202.575 93.470 202.945 ;
        RECT 121.590 202.575 123.470 202.945 ;
        RECT 88.070 201.070 88.330 201.390 ;
        RECT 96.350 201.070 96.610 201.390 ;
        RECT 85.310 200.730 85.570 201.050 ;
        RECT 85.370 199.690 85.510 200.730 ;
        RECT 79.330 199.370 79.590 199.690 ;
        RECT 83.470 199.370 83.730 199.690 ;
        RECT 84.390 199.370 84.650 199.690 ;
        RECT 85.310 199.370 85.570 199.690 ;
        RECT 80.710 199.030 80.970 199.350 ;
        RECT 78.870 198.690 79.130 199.010 ;
        RECT 79.790 198.690 80.050 199.010 ;
        RECT 75.650 198.350 75.910 198.670 ;
        RECT 79.850 196.630 79.990 198.690 ;
        RECT 80.770 197.990 80.910 199.030 ;
        RECT 86.690 198.690 86.950 199.010 ;
        RECT 80.710 197.670 80.970 197.990 ;
        RECT 79.790 196.310 80.050 196.630 ;
        RECT 75.190 195.290 75.450 195.610 ;
        RECT 76.590 194.415 78.470 194.785 ;
        RECT 76.110 193.250 76.370 193.570 ;
        RECT 74.270 190.190 74.530 190.510 ;
        RECT 73.350 189.850 73.610 190.170 ;
        RECT 72.890 188.490 73.150 188.810 ;
        RECT 73.410 185.410 73.550 189.850 ;
        RECT 73.350 185.090 73.610 185.410 ;
        RECT 72.430 184.410 72.690 184.730 ;
        RECT 72.490 183.370 72.630 184.410 ;
        RECT 72.430 183.050 72.690 183.370 ;
        RECT 73.410 183.030 73.550 185.090 ;
        RECT 74.330 185.070 74.470 190.190 ;
        RECT 76.170 189.830 76.310 193.250 ;
        RECT 79.850 190.850 79.990 196.310 ;
        RECT 85.310 194.950 85.570 195.270 ;
        RECT 85.370 194.250 85.510 194.950 ;
        RECT 85.310 193.930 85.570 194.250 ;
        RECT 84.850 192.910 85.110 193.230 ;
        RECT 79.790 190.530 80.050 190.850 ;
        RECT 76.110 189.510 76.370 189.830 ;
        RECT 76.170 185.750 76.310 189.510 ;
        RECT 76.590 188.975 78.470 189.345 ;
        RECT 76.110 185.430 76.370 185.750 ;
        RECT 74.270 184.750 74.530 185.070 ;
        RECT 75.650 184.410 75.910 184.730 ;
        RECT 74.270 184.070 74.530 184.390 ;
        RECT 73.810 183.050 74.070 183.370 ;
        RECT 73.350 182.940 73.610 183.030 ;
        RECT 72.950 182.800 73.610 182.940 ;
        RECT 72.430 182.600 72.690 182.690 ;
        RECT 72.030 182.460 72.690 182.600 ;
        RECT 72.430 182.370 72.690 182.460 ;
        RECT 72.430 181.690 72.690 182.010 ;
        RECT 72.490 179.970 72.630 181.690 ;
        RECT 72.950 179.970 73.090 182.800 ;
        RECT 73.350 182.710 73.610 182.800 ;
        RECT 73.350 182.030 73.610 182.350 ;
        RECT 72.430 179.650 72.690 179.970 ;
        RECT 72.890 179.650 73.150 179.970 ;
        RECT 71.050 179.310 71.310 179.630 ;
        RECT 70.120 177.075 70.400 177.445 ;
        RECT 69.670 174.210 69.930 174.530 ;
        RECT 68.750 173.870 69.010 174.190 ;
        RECT 68.810 171.810 68.950 173.870 ;
        RECT 68.750 171.490 69.010 171.810 ;
        RECT 67.370 169.450 67.630 169.770 ;
        RECT 66.450 165.710 66.710 166.030 ;
        RECT 66.510 160.930 66.650 165.710 ;
        RECT 66.910 162.310 67.170 162.630 ;
        RECT 66.450 160.610 66.710 160.930 ;
        RECT 66.970 160.590 67.110 162.310 ;
        RECT 66.910 160.270 67.170 160.590 ;
        RECT 66.910 159.590 67.170 159.910 ;
        RECT 66.970 156.170 67.110 159.590 ;
        RECT 66.910 155.850 67.170 156.170 ;
        RECT 65.530 155.005 65.790 155.150 ;
        RECT 65.520 154.635 65.800 155.005 ;
        RECT 64.150 152.450 64.410 152.770 ;
        RECT 65.530 152.110 65.790 152.430 ;
        RECT 65.590 150.730 65.730 152.110 ;
        RECT 60.930 150.410 61.190 150.730 ;
        RECT 65.530 150.410 65.790 150.730 ;
        RECT 53.110 149.730 53.370 150.050 ;
        RECT 53.570 149.730 53.830 150.050 ;
        RECT 56.330 149.730 56.590 150.050 ;
        RECT 58.630 149.730 58.890 150.050 ;
        RECT 63.690 149.730 63.950 150.050 ;
        RECT 53.170 147.330 53.310 149.730 ;
        RECT 52.190 147.010 52.450 147.330 ;
        RECT 53.110 147.010 53.370 147.330 ;
        RECT 51.730 146.670 51.990 146.990 ;
        RECT 51.270 146.330 51.530 146.650 ;
        RECT 51.790 145.290 51.930 146.670 ;
        RECT 50.810 144.970 51.070 145.290 ;
        RECT 51.730 144.970 51.990 145.290 ;
        RECT 49.430 144.290 49.690 144.610 ;
        RECT 49.030 143.870 49.630 144.010 ;
        RECT 50.350 143.950 50.610 144.270 ;
        RECT 46.210 141.570 46.470 141.890 ;
        RECT 45.750 141.230 46.010 141.550 ;
        RECT 46.590 140.015 48.470 140.385 ;
        RECT 47.590 137.830 47.850 138.150 ;
        RECT 45.290 136.130 45.550 136.450 ;
        RECT 47.650 136.110 47.790 137.830 ;
        RECT 48.050 136.810 48.310 137.130 ;
        RECT 48.110 136.110 48.250 136.810 ;
        RECT 47.590 136.020 47.850 136.110 ;
        RECT 46.270 135.880 47.850 136.020 ;
        RECT 46.270 133.730 46.410 135.880 ;
        RECT 47.590 135.790 47.850 135.880 ;
        RECT 48.050 135.790 48.310 136.110 ;
        RECT 48.970 135.450 49.230 135.770 ;
        RECT 46.590 134.575 48.470 134.945 ;
        RECT 46.210 133.410 46.470 133.730 ;
        RECT 49.030 133.390 49.170 135.450 ;
        RECT 48.970 133.070 49.230 133.390 ;
        RECT 48.960 131.515 49.240 131.885 ;
        RECT 49.030 130.330 49.170 131.515 ;
        RECT 48.970 130.010 49.230 130.330 ;
        RECT 46.590 129.135 48.470 129.505 ;
        RECT 44.830 128.650 45.090 128.970 ;
        RECT 45.750 127.970 46.010 128.290 ;
        RECT 45.810 125.230 45.950 127.970 ;
        RECT 44.370 124.910 44.630 125.230 ;
        RECT 45.750 124.910 46.010 125.230 ;
        RECT 46.210 124.910 46.470 125.230 ;
        RECT 45.750 124.230 46.010 124.550 ;
        RECT 45.810 122.170 45.950 124.230 ;
        RECT 45.750 121.850 46.010 122.170 ;
        RECT 46.270 120.130 46.410 124.910 ;
        RECT 46.590 123.695 48.470 124.065 ;
        RECT 46.670 121.850 46.930 122.170 ;
        RECT 46.730 120.130 46.870 121.850 ;
        RECT 46.210 120.040 46.470 120.130 ;
        RECT 45.810 119.900 46.470 120.040 ;
        RECT 45.290 119.470 45.550 119.790 ;
        RECT 44.830 118.790 45.090 119.110 ;
        RECT 44.890 117.410 45.030 118.790 ;
        RECT 44.830 117.090 45.090 117.410 ;
        RECT 45.350 115.370 45.490 119.470 ;
        RECT 45.810 116.390 45.950 119.900 ;
        RECT 46.210 119.810 46.470 119.900 ;
        RECT 46.670 119.810 46.930 120.130 ;
        RECT 46.210 119.130 46.470 119.450 ;
        RECT 46.270 117.410 46.410 119.130 ;
        RECT 46.590 118.255 48.470 118.625 ;
        RECT 46.210 117.090 46.470 117.410 ;
        RECT 45.750 116.070 46.010 116.390 ;
        RECT 45.290 115.050 45.550 115.370 ;
        RECT 45.810 114.690 45.950 116.070 ;
        RECT 45.750 114.370 46.010 114.690 ;
        RECT 46.590 112.815 48.470 113.185 ;
        RECT 49.030 112.310 49.170 130.010 ;
        RECT 49.490 128.970 49.630 143.870 ;
        RECT 49.890 137.830 50.150 138.150 ;
        RECT 49.950 133.730 50.090 137.830 ;
        RECT 50.410 136.450 50.550 143.950 ;
        RECT 53.170 141.890 53.310 147.010 ;
        RECT 53.630 145.290 53.770 149.730 ;
        RECT 54.030 149.450 54.290 149.710 ;
        RECT 54.030 149.390 54.690 149.450 ;
        RECT 54.090 149.310 54.690 149.390 ;
        RECT 54.550 148.010 54.690 149.310 ;
        RECT 54.490 147.690 54.750 148.010 ;
        RECT 54.550 146.990 54.690 147.690 ;
        RECT 56.390 146.990 56.530 149.730 ;
        RECT 56.790 147.350 57.050 147.670 ;
        RECT 54.490 146.900 54.750 146.990 ;
        RECT 56.330 146.900 56.590 146.990 ;
        RECT 54.090 146.760 54.750 146.900 ;
        RECT 53.570 144.970 53.830 145.290 ;
        RECT 54.090 141.970 54.230 146.760 ;
        RECT 54.490 146.670 54.750 146.760 ;
        RECT 55.930 146.760 56.590 146.900 ;
        RECT 54.950 144.630 55.210 144.950 ;
        RECT 54.490 143.950 54.750 144.270 ;
        RECT 53.110 141.570 53.370 141.890 ;
        RECT 53.630 141.830 54.230 141.970 ;
        RECT 53.170 137.130 53.310 141.570 ;
        RECT 53.630 141.550 53.770 141.830 ;
        RECT 53.570 141.230 53.830 141.550 ;
        RECT 53.630 138.150 53.770 141.230 ;
        RECT 53.570 137.830 53.830 138.150 ;
        RECT 50.810 136.810 51.070 137.130 ;
        RECT 53.110 136.810 53.370 137.130 ;
        RECT 50.350 136.130 50.610 136.450 ;
        RECT 50.350 135.450 50.610 135.770 ;
        RECT 50.410 134.410 50.550 135.450 ;
        RECT 50.350 134.090 50.610 134.410 ;
        RECT 50.870 133.810 51.010 136.810 ;
        RECT 54.550 136.450 54.690 143.950 ;
        RECT 55.010 138.830 55.150 144.630 ;
        RECT 55.930 141.550 56.070 146.760 ;
        RECT 56.330 146.670 56.590 146.760 ;
        RECT 55.870 141.230 56.130 141.550 ;
        RECT 55.930 139.930 56.070 141.230 ;
        RECT 55.470 139.790 56.070 139.930 ;
        RECT 54.950 138.510 55.210 138.830 ;
        RECT 54.490 136.130 54.750 136.450 ;
        RECT 52.190 135.450 52.450 135.770 ;
        RECT 51.730 135.110 51.990 135.430 ;
        RECT 50.410 133.730 51.010 133.810 ;
        RECT 49.890 133.410 50.150 133.730 ;
        RECT 50.350 133.670 51.010 133.730 ;
        RECT 50.350 133.410 50.610 133.670 ;
        RECT 50.410 132.710 50.550 133.410 ;
        RECT 50.350 132.390 50.610 132.710 ;
        RECT 49.430 128.650 49.690 128.970 ;
        RECT 49.890 119.470 50.150 119.790 ;
        RECT 49.430 118.790 49.690 119.110 ;
        RECT 49.490 114.350 49.630 118.790 ;
        RECT 49.950 114.690 50.090 119.470 ;
        RECT 50.810 118.790 51.070 119.110 ;
        RECT 50.870 117.750 51.010 118.790 ;
        RECT 50.810 117.430 51.070 117.750 ;
        RECT 49.890 114.370 50.150 114.690 ;
        RECT 49.430 114.030 49.690 114.350 ;
        RECT 48.970 111.990 49.230 112.310 ;
        RECT 43.970 111.330 45.950 111.470 ;
        RECT 45.810 106.530 45.950 111.330 ;
        RECT 50.350 111.310 50.610 111.630 ;
        RECT 46.590 107.375 48.470 107.745 ;
        RECT 36.550 106.210 36.810 106.530 ;
        RECT 38.390 106.210 38.650 106.530 ;
        RECT 41.150 106.210 41.410 106.530 ;
        RECT 45.750 106.210 46.010 106.530 ;
        RECT 49.890 106.210 50.150 106.530 ;
        RECT 35.170 105.870 35.430 106.190 ;
        RECT 35.230 103.810 35.370 105.870 ;
        RECT 36.090 105.190 36.350 105.510 ;
        RECT 36.150 103.810 36.290 105.190 ;
        RECT 36.610 104.490 36.750 106.210 ;
        RECT 49.430 105.870 49.690 106.190 ;
        RECT 42.990 105.190 43.250 105.510 ;
        RECT 48.050 105.190 48.310 105.510 ;
        RECT 36.550 104.170 36.810 104.490 ;
        RECT 35.170 103.490 35.430 103.810 ;
        RECT 36.090 103.490 36.350 103.810 ;
        RECT 33.790 101.110 34.050 101.430 ;
        RECT 36.610 101.090 36.750 104.170 ;
        RECT 43.050 103.130 43.190 105.190 ;
        RECT 48.110 103.810 48.250 105.190 ;
        RECT 49.490 103.890 49.630 105.870 ;
        RECT 49.950 104.490 50.090 106.210 ;
        RECT 49.890 104.170 50.150 104.490 ;
        RECT 50.410 104.150 50.550 111.310 ;
        RECT 51.790 108.910 51.930 135.110 ;
        RECT 52.250 133.730 52.390 135.450 ;
        RECT 52.190 133.410 52.450 133.730 ;
        RECT 54.550 127.950 54.690 136.130 ;
        RECT 55.470 135.770 55.610 139.790 ;
        RECT 55.870 138.850 56.130 139.170 ;
        RECT 55.410 135.450 55.670 135.770 ;
        RECT 55.930 134.070 56.070 138.850 ;
        RECT 56.330 135.110 56.590 135.430 ;
        RECT 56.390 134.410 56.530 135.110 ;
        RECT 56.330 134.090 56.590 134.410 ;
        RECT 55.870 133.750 56.130 134.070 ;
        RECT 55.410 132.730 55.670 133.050 ;
        RECT 55.470 128.970 55.610 132.730 ;
        RECT 56.390 128.970 56.530 134.090 ;
        RECT 55.410 128.650 55.670 128.970 ;
        RECT 56.330 128.650 56.590 128.970 ;
        RECT 54.490 127.630 54.750 127.950 ;
        RECT 54.550 125.570 54.690 127.630 ;
        RECT 55.470 125.910 55.610 128.650 ;
        RECT 55.410 125.590 55.670 125.910 ;
        RECT 54.490 125.250 54.750 125.570 ;
        RECT 55.470 123.530 55.610 125.590 ;
        RECT 55.410 123.210 55.670 123.530 ;
        RECT 54.490 117.090 54.750 117.410 ;
        RECT 54.550 115.370 54.690 117.090 ;
        RECT 56.330 116.750 56.590 117.070 ;
        RECT 54.490 115.050 54.750 115.370 ;
        RECT 51.730 108.590 51.990 108.910 ;
        RECT 55.410 107.910 55.670 108.230 ;
        RECT 55.470 106.870 55.610 107.910 ;
        RECT 55.410 106.550 55.670 106.870 ;
        RECT 52.190 105.870 52.450 106.190 ;
        RECT 56.390 106.100 56.530 116.750 ;
        RECT 56.850 108.910 56.990 147.350 ;
        RECT 58.690 146.650 58.830 149.730 ;
        RECT 60.010 149.050 60.270 149.370 ;
        RECT 58.630 146.330 58.890 146.650 ;
        RECT 59.090 145.990 59.350 146.310 ;
        RECT 59.150 144.950 59.290 145.990 ;
        RECT 59.090 144.630 59.350 144.950 ;
        RECT 58.630 143.270 58.890 143.590 ;
        RECT 58.690 141.210 58.830 143.270 ;
        RECT 59.150 142.570 59.290 144.630 ;
        RECT 59.090 142.250 59.350 142.570 ;
        RECT 58.630 140.890 58.890 141.210 ;
        RECT 59.550 135.110 59.810 135.430 ;
        RECT 59.610 133.730 59.750 135.110 ;
        RECT 59.550 133.410 59.810 133.730 ;
        RECT 60.070 133.130 60.210 149.050 ;
        RECT 61.590 148.175 63.470 148.545 ;
        RECT 63.750 146.310 63.890 149.730 ;
        RECT 65.530 149.390 65.790 149.710 ;
        RECT 64.610 149.050 64.870 149.370 ;
        RECT 64.670 147.330 64.810 149.050 ;
        RECT 65.070 148.710 65.330 149.030 ;
        RECT 64.610 147.010 64.870 147.330 ;
        RECT 63.690 145.990 63.950 146.310 ;
        RECT 64.670 144.270 64.810 147.010 ;
        RECT 64.610 143.950 64.870 144.270 ;
        RECT 63.690 143.610 63.950 143.930 ;
        RECT 61.590 142.735 63.470 143.105 ;
        RECT 63.750 140.870 63.890 143.610 ;
        RECT 63.690 140.550 63.950 140.870 ;
        RECT 60.930 139.530 61.190 139.850 ;
        RECT 60.470 138.850 60.730 139.170 ;
        RECT 60.530 137.130 60.670 138.850 ;
        RECT 60.470 136.810 60.730 137.130 ;
        RECT 60.470 135.450 60.730 135.770 ;
        RECT 59.610 132.990 60.210 133.130 ;
        RECT 57.710 126.950 57.970 127.270 ;
        RECT 57.770 125.230 57.910 126.950 ;
        RECT 57.710 124.910 57.970 125.230 ;
        RECT 57.250 122.870 57.510 123.190 ;
        RECT 57.310 120.810 57.450 122.870 ;
        RECT 59.610 122.250 59.750 132.990 ;
        RECT 60.530 125.230 60.670 135.450 ;
        RECT 60.990 135.430 61.130 139.530 ;
        RECT 61.590 137.295 63.470 137.665 ;
        RECT 60.930 135.110 61.190 135.430 ;
        RECT 63.750 133.730 63.890 140.550 ;
        RECT 65.130 139.170 65.270 148.710 ;
        RECT 65.590 146.990 65.730 149.390 ;
        RECT 65.530 146.670 65.790 146.990 ;
        RECT 65.530 144.290 65.790 144.610 ;
        RECT 65.590 139.850 65.730 144.290 ;
        RECT 65.530 139.530 65.790 139.850 ;
        RECT 65.070 138.850 65.330 139.170 ;
        RECT 64.150 138.170 64.410 138.490 ;
        RECT 64.210 136.110 64.350 138.170 ;
        RECT 65.130 137.130 65.270 138.850 ;
        RECT 65.070 136.810 65.330 137.130 ;
        RECT 65.130 136.530 65.270 136.810 ;
        RECT 64.670 136.390 65.270 136.530 ;
        RECT 65.590 136.450 65.730 139.530 ;
        RECT 65.990 138.850 66.250 139.170 ;
        RECT 64.150 135.790 64.410 136.110 ;
        RECT 64.210 134.070 64.350 135.790 ;
        RECT 64.150 133.750 64.410 134.070 ;
        RECT 64.670 133.730 64.810 136.390 ;
        RECT 65.530 136.130 65.790 136.450 ;
        RECT 65.070 135.450 65.330 135.770 ;
        RECT 65.130 133.730 65.270 135.450 ;
        RECT 63.690 133.410 63.950 133.730 ;
        RECT 64.610 133.410 64.870 133.730 ;
        RECT 65.070 133.410 65.330 133.730 ;
        RECT 65.530 133.410 65.790 133.730 ;
        RECT 61.590 131.855 63.470 132.225 ;
        RECT 63.750 128.630 63.890 133.410 ;
        RECT 64.610 130.690 64.870 131.010 ;
        RECT 64.150 130.010 64.410 130.330 ;
        RECT 63.690 128.310 63.950 128.630 ;
        RECT 63.750 127.950 63.890 128.310 ;
        RECT 63.690 127.630 63.950 127.950 ;
        RECT 61.590 126.415 63.470 126.785 ;
        RECT 60.470 124.910 60.730 125.230 ;
        RECT 60.010 124.230 60.270 124.550 ;
        RECT 60.070 122.850 60.210 124.230 ;
        RECT 60.530 123.530 60.670 124.910 ;
        RECT 60.470 123.210 60.730 123.530 ;
        RECT 60.010 122.530 60.270 122.850 ;
        RECT 59.610 122.110 60.210 122.250 ;
        RECT 57.250 120.490 57.510 120.810 ;
        RECT 57.710 119.470 57.970 119.790 ;
        RECT 57.770 117.410 57.910 119.470 ;
        RECT 57.710 117.090 57.970 117.410 ;
        RECT 59.550 117.090 59.810 117.410 ;
        RECT 59.610 108.910 59.750 117.090 ;
        RECT 60.070 111.470 60.210 122.110 ;
        RECT 60.530 120.810 60.670 123.210 ;
        RECT 63.750 122.850 63.890 127.630 ;
        RECT 64.210 122.850 64.350 130.010 ;
        RECT 63.690 122.530 63.950 122.850 ;
        RECT 64.150 122.530 64.410 122.850 ;
        RECT 61.590 120.975 63.470 121.345 ;
        RECT 60.470 120.490 60.730 120.810 ;
        RECT 61.850 119.130 62.110 119.450 ;
        RECT 61.910 118.090 62.050 119.130 ;
        RECT 64.210 118.090 64.350 122.530 ;
        RECT 64.670 122.510 64.810 130.690 ;
        RECT 65.590 130.330 65.730 133.410 ;
        RECT 65.530 130.010 65.790 130.330 ;
        RECT 66.050 129.990 66.190 138.850 ;
        RECT 67.430 138.490 67.570 169.450 ;
        RECT 68.290 166.050 68.550 166.370 ;
        RECT 68.350 163.310 68.490 166.050 ;
        RECT 68.810 165.350 68.950 171.490 ;
        RECT 70.190 168.750 70.330 177.075 ;
        RECT 70.590 173.190 70.850 173.510 ;
        RECT 70.650 169.770 70.790 173.190 ;
        RECT 70.590 169.450 70.850 169.770 ;
        RECT 70.130 168.430 70.390 168.750 ;
        RECT 70.190 167.050 70.330 168.430 ;
        RECT 70.130 166.730 70.390 167.050 ;
        RECT 68.750 165.030 69.010 165.350 ;
        RECT 68.290 162.990 68.550 163.310 ;
        RECT 67.820 158.035 68.100 158.405 ;
        RECT 67.890 152.285 68.030 158.035 ;
        RECT 67.820 151.915 68.100 152.285 ;
        RECT 68.290 152.110 68.550 152.430 ;
        RECT 67.890 139.170 68.030 151.915 ;
        RECT 68.350 141.890 68.490 152.110 ;
        RECT 68.810 143.930 68.950 165.030 ;
        RECT 69.670 159.590 69.930 159.910 ;
        RECT 69.210 157.550 69.470 157.870 ;
        RECT 69.270 152.770 69.410 157.550 ;
        RECT 69.730 154.470 69.870 159.590 ;
        RECT 70.190 157.870 70.330 166.730 ;
        RECT 71.110 166.450 71.250 179.310 ;
        RECT 72.890 178.970 73.150 179.290 ;
        RECT 72.950 177.930 73.090 178.970 ;
        RECT 71.510 177.610 71.770 177.930 ;
        RECT 72.890 177.610 73.150 177.930 ;
        RECT 71.570 176.765 71.710 177.610 ;
        RECT 72.420 177.075 72.700 177.445 ;
        RECT 72.430 176.930 72.690 177.075 ;
        RECT 71.500 176.395 71.780 176.765 ;
        RECT 72.490 174.190 72.630 176.930 ;
        RECT 72.430 173.870 72.690 174.190 ;
        RECT 73.410 171.210 73.550 182.030 ;
        RECT 73.870 179.630 74.010 183.050 ;
        RECT 73.810 179.310 74.070 179.630 ;
        RECT 73.810 176.930 74.070 177.250 ;
        RECT 70.650 166.370 71.250 166.450 ;
        RECT 70.590 166.310 71.250 166.370 ;
        RECT 70.590 166.050 70.850 166.310 ;
        RECT 71.110 160.930 71.250 166.310 ;
        RECT 72.490 171.070 73.550 171.210 ;
        RECT 71.050 160.610 71.310 160.930 ;
        RECT 70.590 159.930 70.850 160.250 ;
        RECT 70.650 158.550 70.790 159.930 ;
        RECT 71.510 158.570 71.770 158.890 ;
        RECT 70.590 158.230 70.850 158.550 ;
        RECT 71.570 158.405 71.710 158.570 ;
        RECT 71.500 158.035 71.780 158.405 ;
        RECT 70.130 157.550 70.390 157.870 ;
        RECT 69.670 154.150 69.930 154.470 ;
        RECT 69.730 153.110 69.870 154.150 ;
        RECT 70.130 153.130 70.390 153.450 ;
        RECT 69.670 152.790 69.930 153.110 ;
        RECT 69.210 152.450 69.470 152.770 ;
        RECT 69.270 150.050 69.410 152.450 ;
        RECT 70.190 151.750 70.330 153.130 ;
        RECT 70.590 152.170 70.850 152.430 ;
        RECT 71.510 152.170 71.770 152.430 ;
        RECT 70.590 152.110 71.770 152.170 ;
        RECT 70.650 152.030 71.710 152.110 ;
        RECT 70.130 151.430 70.390 151.750 ;
        RECT 69.210 149.730 69.470 150.050 ;
        RECT 69.210 143.950 69.470 144.270 ;
        RECT 68.750 143.610 69.010 143.930 ;
        RECT 68.750 141.910 69.010 142.230 ;
        RECT 68.290 141.570 68.550 141.890 ;
        RECT 68.350 140.870 68.490 141.570 ;
        RECT 68.290 140.550 68.550 140.870 ;
        RECT 67.830 138.850 68.090 139.170 ;
        RECT 67.370 138.170 67.630 138.490 ;
        RECT 66.450 137.830 66.710 138.150 ;
        RECT 66.510 135.770 66.650 137.830 ;
        RECT 66.450 135.450 66.710 135.770 ;
        RECT 67.830 130.010 68.090 130.330 ;
        RECT 65.990 129.670 66.250 129.990 ;
        RECT 66.050 128.970 66.190 129.670 ;
        RECT 65.990 128.650 66.250 128.970 ;
        RECT 67.890 128.290 68.030 130.010 ;
        RECT 68.290 128.310 68.550 128.630 ;
        RECT 67.830 127.970 68.090 128.290 ;
        RECT 68.350 125.230 68.490 128.310 ;
        RECT 68.290 124.910 68.550 125.230 ;
        RECT 64.610 122.190 64.870 122.510 ;
        RECT 67.830 121.510 68.090 121.830 ;
        RECT 61.850 117.770 62.110 118.090 ;
        RECT 64.150 117.770 64.410 118.090 ;
        RECT 66.450 117.430 66.710 117.750 ;
        RECT 61.590 115.535 63.470 115.905 ;
        RECT 66.510 115.370 66.650 117.430 ;
        RECT 66.450 115.050 66.710 115.370 ;
        RECT 67.890 114.350 68.030 121.510 ;
        RECT 67.830 114.030 68.090 114.350 ;
        RECT 60.070 111.330 60.670 111.470 ;
        RECT 56.790 108.590 57.050 108.910 ;
        RECT 59.550 108.590 59.810 108.910 ;
        RECT 60.010 108.590 60.270 108.910 ;
        RECT 57.710 107.910 57.970 108.230 ;
        RECT 56.790 106.100 57.050 106.190 ;
        RECT 56.390 105.960 57.050 106.100 ;
        RECT 48.050 103.490 48.310 103.810 ;
        RECT 49.490 103.750 50.090 103.890 ;
        RECT 50.350 103.830 50.610 104.150 ;
        RECT 38.850 102.810 39.110 103.130 ;
        RECT 42.990 102.810 43.250 103.130 ;
        RECT 36.550 100.770 36.810 101.090 ;
        RECT 31.590 99.215 33.470 99.585 ;
        RECT 31.780 88.250 33.000 89.380 ;
        RECT 38.910 89.290 39.050 102.810 ;
        RECT 43.910 102.470 44.170 102.790 ;
        RECT 43.970 89.530 44.110 102.470 ;
        RECT 46.590 101.935 48.470 102.305 ;
        RECT 37.750 88.780 39.050 89.290 ;
        RECT 30.170 88.110 33.000 88.250 ;
        RECT 31.780 85.510 33.000 88.110 ;
        RECT 37.680 88.620 39.050 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.950 89.040 50.090 103.750 ;
        RECT 52.250 103.470 52.390 105.870 ;
        RECT 56.390 104.490 56.530 105.960 ;
        RECT 56.790 105.870 57.050 105.960 ;
        RECT 56.790 105.190 57.050 105.510 ;
        RECT 56.330 104.170 56.590 104.490 ;
        RECT 56.850 103.890 56.990 105.190 ;
        RECT 56.390 103.750 56.990 103.890 ;
        RECT 57.770 103.810 57.910 107.910 ;
        RECT 60.070 106.530 60.210 108.590 ;
        RECT 60.530 106.530 60.670 111.330 ;
        RECT 61.590 110.095 63.470 110.465 ;
        RECT 68.810 108.910 68.950 141.910 ;
        RECT 69.270 136.110 69.410 143.950 ;
        RECT 69.670 143.270 69.930 143.590 ;
        RECT 69.730 141.550 69.870 143.270 ;
        RECT 69.670 141.230 69.930 141.550 ;
        RECT 70.190 138.830 70.330 151.430 ;
        RECT 70.650 150.050 70.790 152.030 ;
        RECT 71.970 151.770 72.230 152.090 ;
        RECT 70.590 149.730 70.850 150.050 ;
        RECT 70.650 147.330 70.790 149.730 ;
        RECT 70.590 147.010 70.850 147.330 ;
        RECT 72.030 146.990 72.170 151.770 ;
        RECT 71.970 146.670 72.230 146.990 ;
        RECT 70.590 143.610 70.850 143.930 ;
        RECT 70.650 141.550 70.790 143.610 ;
        RECT 70.590 141.230 70.850 141.550 ;
        RECT 70.130 138.510 70.390 138.830 ;
        RECT 69.210 135.790 69.470 136.110 ;
        RECT 69.270 131.010 69.410 135.790 ;
        RECT 69.210 130.690 69.470 131.010 ;
        RECT 70.650 130.410 70.790 141.230 ;
        RECT 71.970 140.550 72.230 140.870 ;
        RECT 72.030 139.510 72.170 140.550 ;
        RECT 71.970 139.190 72.230 139.510 ;
        RECT 72.490 130.670 72.630 171.070 ;
        RECT 73.870 166.030 74.010 176.930 ;
        RECT 73.810 165.710 74.070 166.030 ;
        RECT 72.890 165.030 73.150 165.350 ;
        RECT 72.950 163.310 73.090 165.030 ;
        RECT 72.890 162.990 73.150 163.310 ;
        RECT 72.950 157.870 73.090 162.990 ;
        RECT 74.330 160.840 74.470 184.070 ;
        RECT 75.710 182.690 75.850 184.410 ;
        RECT 75.650 182.370 75.910 182.690 ;
        RECT 75.710 182.010 75.850 182.370 ;
        RECT 75.650 181.690 75.910 182.010 ;
        RECT 74.730 181.350 74.990 181.670 ;
        RECT 76.170 181.410 76.310 185.430 ;
        RECT 84.910 185.410 85.050 192.910 ;
        RECT 85.370 191.530 85.510 193.930 ;
        RECT 86.750 193.910 86.890 198.690 ;
        RECT 91.590 197.135 93.470 197.505 ;
        RECT 93.590 195.970 93.850 196.290 ;
        RECT 89.910 195.290 90.170 195.610 ;
        RECT 89.970 194.250 90.110 195.290 ;
        RECT 89.910 193.930 90.170 194.250 ;
        RECT 86.690 193.590 86.950 193.910 ;
        RECT 85.770 193.250 86.030 193.570 ;
        RECT 89.910 193.250 90.170 193.570 ;
        RECT 85.310 191.210 85.570 191.530 ;
        RECT 84.850 185.090 85.110 185.410 ;
        RECT 76.590 183.535 78.470 183.905 ;
        RECT 76.570 182.370 76.830 182.690 ;
        RECT 76.630 181.410 76.770 182.370 ;
        RECT 84.910 181.670 85.050 185.090 ;
        RECT 74.790 177.250 74.930 181.350 ;
        RECT 75.710 181.270 76.770 181.410 ;
        RECT 79.330 181.350 79.590 181.670 ;
        RECT 84.850 181.350 85.110 181.670 ;
        RECT 75.710 179.970 75.850 181.270 ;
        RECT 78.870 179.990 79.130 180.310 ;
        RECT 75.650 179.650 75.910 179.970 ;
        RECT 76.110 179.310 76.370 179.630 ;
        RECT 76.170 177.250 76.310 179.310 ;
        RECT 78.400 179.115 78.680 179.485 ;
        RECT 78.470 178.950 78.610 179.115 ;
        RECT 78.410 178.630 78.670 178.950 ;
        RECT 76.590 178.095 78.470 178.465 ;
        RECT 74.730 176.930 74.990 177.250 ;
        RECT 76.110 176.930 76.370 177.250 ;
        RECT 77.490 176.930 77.750 177.250 ;
        RECT 77.950 176.930 78.210 177.250 ;
        RECT 74.790 176.230 74.930 176.930 ;
        RECT 74.730 175.910 74.990 176.230 ;
        RECT 76.170 174.870 76.310 176.930 ;
        RECT 77.550 175.210 77.690 176.930 ;
        RECT 78.010 176.765 78.150 176.930 ;
        RECT 78.930 176.910 79.070 179.990 ;
        RECT 79.390 179.970 79.530 181.350 ;
        RECT 82.090 180.330 82.350 180.650 ;
        RECT 79.330 179.650 79.590 179.970 ;
        RECT 81.170 179.310 81.430 179.630 ;
        RECT 81.630 179.310 81.890 179.630 ;
        RECT 79.330 177.270 79.590 177.590 ;
        RECT 77.940 176.395 78.220 176.765 ;
        RECT 78.870 176.590 79.130 176.910 ;
        RECT 77.490 174.890 77.750 175.210 ;
        RECT 76.110 174.550 76.370 174.870 ;
        RECT 78.010 174.190 78.150 176.395 ;
        RECT 77.950 173.870 78.210 174.190 ;
        RECT 76.590 172.655 78.470 173.025 ;
        RECT 76.110 167.750 76.370 168.070 ;
        RECT 78.870 167.750 79.130 168.070 ;
        RECT 74.730 165.710 74.990 166.030 ;
        RECT 73.410 160.700 74.470 160.840 ;
        RECT 72.890 157.550 73.150 157.870 ;
        RECT 72.880 155.995 73.160 156.365 ;
        RECT 69.730 130.270 70.790 130.410 ;
        RECT 72.430 130.350 72.690 130.670 ;
        RECT 69.730 125.230 69.870 130.270 ;
        RECT 70.130 129.670 70.390 129.990 ;
        RECT 71.510 129.670 71.770 129.990 ;
        RECT 70.190 125.230 70.330 129.670 ;
        RECT 71.570 125.230 71.710 129.670 ;
        RECT 71.970 127.970 72.230 128.290 ;
        RECT 72.030 126.250 72.170 127.970 ;
        RECT 71.970 125.930 72.230 126.250 ;
        RECT 69.670 125.140 69.930 125.230 ;
        RECT 69.270 125.000 69.930 125.140 ;
        RECT 69.270 117.070 69.410 125.000 ;
        RECT 69.670 124.910 69.930 125.000 ;
        RECT 70.130 124.910 70.390 125.230 ;
        RECT 71.510 124.910 71.770 125.230 ;
        RECT 69.670 124.230 69.930 124.550 ;
        RECT 69.730 119.790 69.870 124.230 ;
        RECT 72.950 122.850 73.090 155.995 ;
        RECT 73.410 153.450 73.550 160.700 ;
        RECT 73.810 159.590 74.070 159.910 ;
        RECT 73.870 157.870 74.010 159.590 ;
        RECT 73.810 157.550 74.070 157.870 ;
        RECT 73.870 157.190 74.010 157.550 ;
        RECT 73.810 156.870 74.070 157.190 ;
        RECT 73.870 155.830 74.010 156.870 ;
        RECT 73.810 155.510 74.070 155.830 ;
        RECT 74.270 155.170 74.530 155.490 ;
        RECT 74.330 155.005 74.470 155.170 ;
        RECT 74.260 154.635 74.540 155.005 ;
        RECT 73.350 153.130 73.610 153.450 ;
        RECT 73.410 152.090 73.550 153.130 ;
        RECT 73.810 152.680 74.070 152.770 ;
        RECT 74.790 152.680 74.930 165.710 ;
        RECT 75.190 162.650 75.450 162.970 ;
        RECT 75.250 156.365 75.390 162.650 ;
        RECT 76.170 158.210 76.310 167.750 ;
        RECT 76.590 167.215 78.470 167.585 ;
        RECT 78.410 165.370 78.670 165.690 ;
        RECT 78.470 163.650 78.610 165.370 ;
        RECT 78.410 163.330 78.670 163.650 ;
        RECT 78.930 162.970 79.070 167.750 ;
        RECT 78.870 162.650 79.130 162.970 ;
        RECT 76.590 161.775 78.470 162.145 ;
        RECT 76.110 157.890 76.370 158.210 ;
        RECT 78.870 157.550 79.130 157.870 ;
        RECT 76.110 157.210 76.370 157.530 ;
        RECT 75.650 156.870 75.910 157.190 ;
        RECT 75.180 155.995 75.460 156.365 ;
        RECT 73.810 152.540 74.930 152.680 ;
        RECT 73.810 152.450 74.070 152.540 ;
        RECT 73.350 151.770 73.610 152.090 ;
        RECT 73.350 147.690 73.610 148.010 ;
        RECT 73.410 146.310 73.550 147.690 ;
        RECT 73.350 145.990 73.610 146.310 ;
        RECT 73.870 136.450 74.010 152.450 ;
        RECT 74.730 151.430 74.990 151.750 ;
        RECT 74.790 150.390 74.930 151.430 ;
        RECT 74.730 150.070 74.990 150.390 ;
        RECT 75.710 150.050 75.850 156.870 ;
        RECT 76.170 155.150 76.310 157.210 ;
        RECT 76.590 156.335 78.470 156.705 ;
        RECT 78.930 156.080 79.070 157.550 ;
        RECT 78.010 155.940 79.070 156.080 ;
        RECT 78.010 155.490 78.150 155.940 ;
        RECT 77.950 155.170 78.210 155.490 ;
        RECT 78.410 155.170 78.670 155.490 ;
        RECT 76.110 154.830 76.370 155.150 ;
        RECT 78.470 154.810 78.610 155.170 ;
        RECT 78.410 154.490 78.670 154.810 ;
        RECT 76.110 154.150 76.370 154.470 ;
        RECT 75.650 149.730 75.910 150.050 ;
        RECT 75.650 148.710 75.910 149.030 ;
        RECT 75.190 143.610 75.450 143.930 ;
        RECT 74.730 138.510 74.990 138.830 ;
        RECT 74.790 137.130 74.930 138.510 ;
        RECT 74.730 136.810 74.990 137.130 ;
        RECT 74.270 136.470 74.530 136.790 ;
        RECT 73.810 136.130 74.070 136.450 ;
        RECT 73.870 131.010 74.010 136.130 ;
        RECT 74.330 134.410 74.470 136.470 ;
        RECT 74.270 134.090 74.530 134.410 ;
        RECT 73.810 130.690 74.070 131.010 ;
        RECT 72.890 122.530 73.150 122.850 ;
        RECT 72.950 119.790 73.090 122.530 ;
        RECT 69.670 119.470 69.930 119.790 ;
        RECT 72.890 119.470 73.150 119.790 ;
        RECT 70.590 119.130 70.850 119.450 ;
        RECT 70.650 118.170 70.790 119.130 ;
        RECT 70.650 118.030 71.250 118.170 ;
        RECT 71.110 117.070 71.250 118.030 ;
        RECT 69.210 116.750 69.470 117.070 ;
        RECT 70.590 116.750 70.850 117.070 ;
        RECT 71.050 116.750 71.310 117.070 ;
        RECT 69.270 114.690 69.410 116.750 ;
        RECT 70.650 115.370 70.790 116.750 ;
        RECT 71.110 115.370 71.250 116.750 ;
        RECT 70.590 115.050 70.850 115.370 ;
        RECT 71.050 115.050 71.310 115.370 ;
        RECT 73.350 115.050 73.610 115.370 ;
        RECT 69.210 114.370 69.470 114.690 ;
        RECT 68.750 108.590 69.010 108.910 ;
        RECT 65.070 107.910 65.330 108.230 ;
        RECT 71.970 107.910 72.230 108.230 ;
        RECT 65.130 106.870 65.270 107.910 ;
        RECT 72.030 106.870 72.170 107.910 ;
        RECT 65.070 106.550 65.330 106.870 ;
        RECT 71.970 106.550 72.230 106.870 ;
        RECT 60.010 106.210 60.270 106.530 ;
        RECT 60.470 106.210 60.730 106.530 ;
        RECT 73.410 106.190 73.550 115.050 ;
        RECT 73.870 109.930 74.010 130.690 ;
        RECT 74.730 129.670 74.990 129.990 ;
        RECT 74.790 128.290 74.930 129.670 ;
        RECT 74.730 127.970 74.990 128.290 ;
        RECT 75.250 127.690 75.390 143.610 ;
        RECT 74.790 127.550 75.390 127.690 ;
        RECT 73.810 109.610 74.070 109.930 ;
        RECT 74.790 106.530 74.930 127.550 ;
        RECT 75.190 118.790 75.450 119.110 ;
        RECT 75.250 117.750 75.390 118.790 ;
        RECT 75.190 117.430 75.450 117.750 ;
        RECT 75.710 108.570 75.850 148.710 ;
        RECT 76.170 136.110 76.310 154.150 ;
        RECT 76.590 150.895 78.470 151.265 ;
        RECT 79.390 149.710 79.530 177.270 ;
        RECT 81.230 177.160 81.370 179.310 ;
        RECT 81.690 177.930 81.830 179.310 ;
        RECT 82.150 177.930 82.290 180.330 ;
        RECT 84.910 179.970 85.050 181.350 ;
        RECT 85.370 180.310 85.510 191.210 ;
        RECT 85.830 189.830 85.970 193.250 ;
        RECT 87.610 189.850 87.870 190.170 ;
        RECT 85.770 189.510 86.030 189.830 ;
        RECT 85.830 184.390 85.970 189.510 ;
        RECT 87.670 188.810 87.810 189.850 ;
        RECT 87.610 188.490 87.870 188.810 ;
        RECT 88.990 187.810 89.250 188.130 ;
        RECT 89.050 186.090 89.190 187.810 ;
        RECT 89.970 187.790 90.110 193.250 ;
        RECT 90.830 192.230 91.090 192.550 ;
        RECT 90.890 190.510 91.030 192.230 ;
        RECT 91.590 191.695 93.470 192.065 ;
        RECT 93.650 191.530 93.790 195.970 ;
        RECT 96.410 195.950 96.550 201.070 ;
        RECT 106.590 199.855 108.470 200.225 ;
        RECT 97.730 199.030 97.990 199.350 ;
        RECT 96.350 195.630 96.610 195.950 ;
        RECT 96.410 193.910 96.550 195.630 ;
        RECT 97.790 194.250 97.930 199.030 ;
        RECT 104.170 198.350 104.430 198.670 ;
        RECT 105.550 198.350 105.810 198.670 ;
        RECT 98.190 197.670 98.450 197.990 ;
        RECT 98.250 195.950 98.390 197.670 ;
        RECT 98.190 195.630 98.450 195.950 ;
        RECT 97.730 193.930 97.990 194.250 ;
        RECT 96.350 193.590 96.610 193.910 ;
        RECT 94.510 193.250 94.770 193.570 ;
        RECT 93.590 191.210 93.850 191.530 ;
        RECT 93.590 190.530 93.850 190.850 ;
        RECT 90.370 190.190 90.630 190.510 ;
        RECT 90.830 190.190 91.090 190.510 ;
        RECT 90.430 188.810 90.570 190.190 ;
        RECT 90.370 188.490 90.630 188.810 ;
        RECT 89.910 187.470 90.170 187.790 ;
        RECT 90.830 187.470 91.090 187.790 ;
        RECT 88.990 185.770 89.250 186.090 ;
        RECT 90.890 185.750 91.030 187.470 ;
        RECT 91.590 186.255 93.470 186.625 ;
        RECT 90.830 185.430 91.090 185.750 ;
        RECT 85.770 184.070 86.030 184.390 ;
        RECT 86.230 184.070 86.490 184.390 ;
        RECT 85.310 179.990 85.570 180.310 ;
        RECT 84.850 179.650 85.110 179.970 ;
        RECT 84.910 179.485 85.050 179.650 ;
        RECT 84.840 179.115 85.120 179.485 ;
        RECT 82.550 178.630 82.810 178.950 ;
        RECT 83.470 178.630 83.730 178.950 ;
        RECT 81.630 177.610 81.890 177.930 ;
        RECT 82.090 177.610 82.350 177.930 ;
        RECT 82.610 177.250 82.750 178.630 ;
        RECT 81.630 177.160 81.890 177.250 ;
        RECT 81.230 177.020 81.890 177.160 ;
        RECT 81.630 176.930 81.890 177.020 ;
        RECT 82.550 176.930 82.810 177.250 ;
        RECT 80.250 176.590 80.510 176.910 ;
        RECT 79.790 168.770 80.050 169.090 ;
        RECT 79.850 165.350 79.990 168.770 ;
        RECT 79.790 165.030 80.050 165.350 ;
        RECT 79.850 160.590 79.990 165.030 ;
        RECT 79.790 160.270 80.050 160.590 ;
        RECT 79.780 158.715 80.060 159.085 ;
        RECT 79.790 158.570 80.050 158.715 ;
        RECT 80.310 154.890 80.450 176.590 ;
        RECT 81.690 175.210 81.830 176.930 ;
        RECT 81.630 174.890 81.890 175.210 ;
        RECT 81.630 173.530 81.890 173.850 ;
        RECT 80.710 162.310 80.970 162.630 ;
        RECT 81.690 162.370 81.830 173.530 ;
        RECT 83.010 167.750 83.270 168.070 ;
        RECT 82.550 165.710 82.810 166.030 ;
        RECT 82.610 164.330 82.750 165.710 ;
        RECT 82.550 164.010 82.810 164.330 ;
        RECT 83.070 163.310 83.210 167.750 ;
        RECT 83.530 165.770 83.670 178.630 ;
        RECT 85.830 177.590 85.970 184.070 ;
        RECT 86.290 179.290 86.430 184.070 ;
        RECT 90.890 182.690 91.030 185.430 ;
        RECT 90.830 182.370 91.090 182.690 ;
        RECT 89.450 181.690 89.710 182.010 ;
        RECT 89.510 180.650 89.650 181.690 ;
        RECT 89.450 180.330 89.710 180.650 ;
        RECT 90.890 179.630 91.030 182.370 ;
        RECT 93.650 182.350 93.790 190.530 ;
        RECT 94.570 187.645 94.710 193.250 ;
        RECT 96.410 190.510 96.550 193.590 ;
        RECT 97.730 190.530 97.990 190.850 ;
        RECT 96.350 190.190 96.610 190.510 ;
        RECT 94.500 187.275 94.780 187.645 ;
        RECT 97.270 184.070 97.530 184.390 ;
        RECT 97.330 183.370 97.470 184.070 ;
        RECT 97.270 183.050 97.530 183.370 ;
        RECT 95.890 182.370 96.150 182.690 ;
        RECT 93.590 182.030 93.850 182.350 ;
        RECT 91.590 180.815 93.470 181.185 ;
        RECT 90.370 179.310 90.630 179.630 ;
        RECT 90.830 179.310 91.090 179.630 ;
        RECT 86.230 178.970 86.490 179.290 ;
        RECT 87.150 178.630 87.410 178.950 ;
        RECT 88.990 178.630 89.250 178.950 ;
        RECT 85.770 177.270 86.030 177.590 ;
        RECT 83.930 176.930 84.190 177.250 ;
        RECT 83.990 174.190 84.130 176.930 ;
        RECT 87.210 174.530 87.350 178.630 ;
        RECT 89.050 177.250 89.190 178.630 ;
        RECT 90.430 177.930 90.570 179.310 ;
        RECT 90.370 177.610 90.630 177.930 ;
        RECT 88.990 176.930 89.250 177.250 ;
        RECT 87.150 174.210 87.410 174.530 ;
        RECT 83.930 173.870 84.190 174.190 ;
        RECT 90.890 172.490 91.030 179.310 ;
        RECT 95.950 178.950 96.090 182.370 ;
        RECT 97.790 182.350 97.930 190.530 ;
        RECT 97.730 182.030 97.990 182.350 ;
        RECT 98.250 182.010 98.390 195.630 ;
        RECT 100.950 194.950 101.210 195.270 ;
        RECT 101.010 190.850 101.150 194.950 ;
        RECT 104.230 191.530 104.370 198.350 ;
        RECT 105.610 193.910 105.750 198.350 ;
        RECT 121.590 197.135 123.470 197.505 ;
        RECT 115.210 195.290 115.470 195.610 ;
        RECT 117.510 195.290 117.770 195.610 ;
        RECT 117.970 195.290 118.230 195.610 ;
        RECT 108.770 194.950 109.030 195.270 ;
        RECT 106.590 194.415 108.470 194.785 ;
        RECT 105.550 193.590 105.810 193.910 ;
        RECT 107.850 192.910 108.110 193.230 ;
        RECT 104.170 191.210 104.430 191.530 ;
        RECT 107.910 191.190 108.050 192.910 ;
        RECT 107.850 190.870 108.110 191.190 ;
        RECT 100.950 190.530 101.210 190.850 ;
        RECT 106.010 190.530 106.270 190.850 ;
        RECT 106.070 188.810 106.210 190.530 ;
        RECT 106.590 188.975 108.470 189.345 ;
        RECT 106.010 188.490 106.270 188.810 ;
        RECT 100.030 188.150 100.290 188.470 ;
        RECT 99.110 186.790 99.370 187.110 ;
        RECT 99.570 186.790 99.830 187.110 ;
        RECT 99.170 185.410 99.310 186.790 ;
        RECT 99.630 186.090 99.770 186.790 ;
        RECT 100.090 186.090 100.230 188.150 ;
        RECT 99.570 185.770 99.830 186.090 ;
        RECT 100.030 185.770 100.290 186.090 ;
        RECT 108.830 185.410 108.970 194.950 ;
        RECT 115.270 194.250 115.410 195.290 ;
        RECT 112.450 193.930 112.710 194.250 ;
        RECT 115.210 193.930 115.470 194.250 ;
        RECT 110.610 192.910 110.870 193.230 ;
        RECT 109.230 192.230 109.490 192.550 ;
        RECT 109.290 190.170 109.430 192.230 ;
        RECT 109.690 190.530 109.950 190.850 ;
        RECT 109.230 189.850 109.490 190.170 ;
        RECT 109.750 188.130 109.890 190.530 ;
        RECT 109.690 187.810 109.950 188.130 ;
        RECT 99.110 185.090 99.370 185.410 ;
        RECT 105.090 185.090 105.350 185.410 ;
        RECT 108.770 185.090 109.030 185.410 ;
        RECT 99.170 182.690 99.310 185.090 ;
        RECT 99.110 182.370 99.370 182.690 ;
        RECT 98.190 181.690 98.450 182.010 ;
        RECT 95.890 178.630 96.150 178.950 ;
        RECT 99.170 177.250 99.310 182.370 ;
        RECT 104.170 182.090 104.430 182.350 ;
        RECT 103.310 182.030 104.430 182.090 ;
        RECT 103.310 181.950 104.370 182.030 ;
        RECT 99.570 178.970 99.830 179.290 ;
        RECT 101.870 178.970 102.130 179.290 ;
        RECT 99.630 177.930 99.770 178.970 ;
        RECT 99.570 177.610 99.830 177.930 ;
        RECT 101.930 177.250 102.070 178.970 ;
        RECT 98.190 176.930 98.450 177.250 ;
        RECT 99.110 176.930 99.370 177.250 ;
        RECT 101.870 176.930 102.130 177.250 ;
        RECT 91.590 175.375 93.470 175.745 ;
        RECT 98.250 174.190 98.390 176.930 ;
        RECT 100.490 175.910 100.750 176.230 ;
        RECT 101.870 175.910 102.130 176.230 ;
        RECT 98.190 173.870 98.450 174.190 ;
        RECT 98.250 173.510 98.390 173.870 ;
        RECT 98.190 173.190 98.450 173.510 ;
        RECT 90.830 172.170 91.090 172.490 ;
        RECT 98.190 171.150 98.450 171.470 ;
        RECT 89.450 170.470 89.710 170.790 ;
        RECT 89.510 169.430 89.650 170.470 ;
        RECT 91.590 169.935 93.470 170.305 ;
        RECT 98.250 169.770 98.390 171.150 ;
        RECT 98.190 169.450 98.450 169.770 ;
        RECT 89.450 169.110 89.710 169.430 ;
        RECT 91.750 168.770 92.010 169.090 ;
        RECT 87.610 168.430 87.870 168.750 ;
        RECT 90.830 168.430 91.090 168.750 ;
        RECT 83.930 168.090 84.190 168.410 ;
        RECT 83.990 166.710 84.130 168.090 ;
        RECT 83.930 166.390 84.190 166.710 ;
        RECT 83.530 165.630 84.130 165.770 ;
        RECT 83.010 162.990 83.270 163.310 ;
        RECT 80.770 160.250 80.910 162.310 ;
        RECT 81.690 162.230 83.670 162.370 ;
        RECT 82.550 161.290 82.810 161.610 ;
        RECT 80.710 159.930 80.970 160.250 ;
        RECT 80.770 158.890 80.910 159.930 ;
        RECT 80.710 158.570 80.970 158.890 ;
        RECT 81.160 158.715 81.440 159.085 ;
        RECT 80.770 155.830 80.910 158.570 ;
        RECT 80.710 155.510 80.970 155.830 ;
        RECT 80.310 154.750 80.910 154.890 ;
        RECT 80.250 154.150 80.510 154.470 ;
        RECT 79.790 149.730 80.050 150.050 ;
        RECT 79.330 149.390 79.590 149.710 ;
        RECT 77.950 149.050 78.210 149.370 ;
        RECT 78.010 147.670 78.150 149.050 ;
        RECT 79.850 148.010 79.990 149.730 ;
        RECT 79.790 147.690 80.050 148.010 ;
        RECT 77.950 147.350 78.210 147.670 ;
        RECT 77.950 146.670 78.210 146.990 ;
        RECT 79.790 146.670 80.050 146.990 ;
        RECT 78.010 146.310 78.150 146.670 ;
        RECT 77.950 145.990 78.210 146.310 ;
        RECT 79.330 145.990 79.590 146.310 ;
        RECT 76.590 145.455 78.470 145.825 ;
        RECT 79.390 144.950 79.530 145.990 ;
        RECT 79.330 144.630 79.590 144.950 ;
        RECT 76.590 140.015 78.470 140.385 ;
        RECT 79.850 139.510 79.990 146.670 ;
        RECT 79.790 139.190 80.050 139.510 ;
        RECT 79.330 137.830 79.590 138.150 ;
        RECT 79.390 136.110 79.530 137.830 ;
        RECT 79.790 136.810 80.050 137.130 ;
        RECT 76.110 135.790 76.370 136.110 ;
        RECT 79.330 135.790 79.590 136.110 ;
        RECT 78.870 135.110 79.130 135.430 ;
        RECT 76.590 134.575 78.470 134.945 ;
        RECT 78.930 134.070 79.070 135.110 ;
        RECT 78.870 133.750 79.130 134.070 ;
        RECT 79.850 131.690 79.990 136.810 ;
        RECT 80.310 133.730 80.450 154.150 ;
        RECT 80.770 145.290 80.910 154.750 ;
        RECT 80.710 144.970 80.970 145.290 ;
        RECT 81.230 144.610 81.370 158.715 ;
        RECT 81.630 157.550 81.890 157.870 ;
        RECT 81.690 155.490 81.830 157.550 ;
        RECT 82.090 157.210 82.350 157.530 ;
        RECT 82.150 155.490 82.290 157.210 ;
        RECT 82.610 155.490 82.750 161.290 ;
        RECT 83.010 159.590 83.270 159.910 ;
        RECT 83.070 157.530 83.210 159.590 ;
        RECT 83.010 157.210 83.270 157.530 ;
        RECT 81.630 155.170 81.890 155.490 ;
        RECT 82.090 155.170 82.350 155.490 ;
        RECT 82.550 155.170 82.810 155.490 ;
        RECT 82.150 154.810 82.290 155.170 ;
        RECT 82.090 154.490 82.350 154.810 ;
        RECT 81.630 148.710 81.890 149.030 ;
        RECT 81.170 144.290 81.430 144.610 ;
        RECT 80.710 143.270 80.970 143.590 ;
        RECT 80.250 133.410 80.510 133.730 ;
        RECT 80.770 133.130 80.910 143.270 ;
        RECT 81.170 139.530 81.430 139.850 ;
        RECT 81.230 136.110 81.370 139.530 ;
        RECT 81.170 135.790 81.430 136.110 ;
        RECT 80.310 132.990 80.910 133.130 ;
        RECT 79.790 131.370 80.050 131.690 ;
        RECT 79.790 130.350 80.050 130.670 ;
        RECT 76.590 129.135 78.470 129.505 ;
        RECT 78.410 127.630 78.670 127.950 ;
        RECT 78.470 126.250 78.610 127.630 ;
        RECT 78.870 127.290 79.130 127.610 ;
        RECT 78.930 126.250 79.070 127.290 ;
        RECT 78.410 125.930 78.670 126.250 ;
        RECT 78.870 125.930 79.130 126.250 ;
        RECT 76.590 123.695 78.470 124.065 ;
        RECT 78.930 119.110 79.070 125.930 ;
        RECT 79.330 125.250 79.590 125.570 ;
        RECT 79.390 120.130 79.530 125.250 ;
        RECT 79.330 119.810 79.590 120.130 ;
        RECT 79.330 119.360 79.590 119.450 ;
        RECT 79.850 119.360 79.990 130.350 ;
        RECT 80.310 128.630 80.450 132.990 ;
        RECT 80.250 128.310 80.510 128.630 ;
        RECT 80.250 127.630 80.510 127.950 ;
        RECT 80.310 126.250 80.450 127.630 ;
        RECT 81.690 127.270 81.830 148.710 ;
        RECT 83.010 147.350 83.270 147.670 ;
        RECT 83.070 146.990 83.210 147.350 ;
        RECT 82.090 146.670 82.350 146.990 ;
        RECT 83.010 146.670 83.270 146.990 ;
        RECT 82.150 146.310 82.290 146.670 ;
        RECT 82.550 146.330 82.810 146.650 ;
        RECT 82.090 145.990 82.350 146.310 ;
        RECT 82.090 138.740 82.350 138.830 ;
        RECT 82.610 138.740 82.750 146.330 ;
        RECT 83.070 138.830 83.210 146.670 ;
        RECT 82.090 138.600 82.750 138.740 ;
        RECT 82.090 138.510 82.350 138.600 ;
        RECT 83.010 138.510 83.270 138.830 ;
        RECT 82.150 136.790 82.290 138.510 ;
        RECT 82.090 136.470 82.350 136.790 ;
        RECT 83.070 136.110 83.210 138.510 ;
        RECT 83.010 135.790 83.270 136.110 ;
        RECT 83.530 133.390 83.670 162.230 ;
        RECT 83.990 135.770 84.130 165.630 ;
        RECT 87.670 164.330 87.810 168.430 ;
        RECT 88.530 166.050 88.790 166.370 ;
        RECT 87.610 164.010 87.870 164.330 ;
        RECT 88.590 160.250 88.730 166.050 ;
        RECT 90.890 166.030 91.030 168.430 ;
        RECT 91.810 166.030 91.950 168.770 ;
        RECT 100.030 166.390 100.290 166.710 ;
        RECT 90.830 165.710 91.090 166.030 ;
        RECT 91.750 165.710 92.010 166.030 ;
        RECT 93.590 165.710 93.850 166.030 ;
        RECT 94.510 165.710 94.770 166.030 ;
        RECT 98.190 165.710 98.450 166.030 ;
        RECT 90.890 162.630 91.030 165.710 ;
        RECT 91.810 165.350 91.950 165.710 ;
        RECT 91.750 165.030 92.010 165.350 ;
        RECT 91.590 164.495 93.470 164.865 ;
        RECT 93.650 163.650 93.790 165.710 ;
        RECT 93.590 163.330 93.850 163.650 ;
        RECT 90.830 162.310 91.090 162.630 ;
        RECT 88.530 159.930 88.790 160.250 ;
        RECT 88.070 159.590 88.330 159.910 ;
        RECT 84.380 158.035 84.660 158.405 ;
        RECT 88.130 158.210 88.270 159.590 ;
        RECT 88.590 158.210 88.730 159.930 ;
        RECT 84.450 155.490 84.590 158.035 ;
        RECT 88.070 157.890 88.330 158.210 ;
        RECT 88.530 157.890 88.790 158.210 ;
        RECT 90.890 157.870 91.030 162.310 ;
        RECT 94.570 161.610 94.710 165.710 ;
        RECT 96.350 165.030 96.610 165.350 ;
        RECT 94.510 161.290 94.770 161.610 ;
        RECT 94.050 160.950 94.310 161.270 ;
        RECT 91.590 159.055 93.470 159.425 ;
        RECT 94.110 158.890 94.250 160.950 ;
        RECT 94.050 158.570 94.310 158.890 ;
        RECT 96.410 157.870 96.550 165.030 ;
        RECT 98.250 162.970 98.390 165.710 ;
        RECT 98.190 162.650 98.450 162.970 ;
        RECT 97.270 162.310 97.530 162.630 ;
        RECT 97.330 160.930 97.470 162.310 ;
        RECT 97.270 160.610 97.530 160.930 ;
        RECT 96.810 160.270 97.070 160.590 ;
        RECT 96.870 158.890 97.010 160.270 ;
        RECT 96.810 158.570 97.070 158.890 ;
        RECT 90.830 157.550 91.090 157.870 ;
        RECT 96.350 157.550 96.610 157.870 ;
        RECT 84.390 155.170 84.650 155.490 ;
        RECT 90.890 153.360 91.030 157.550 ;
        RECT 94.970 157.210 95.230 157.530 ;
        RECT 91.590 153.615 93.470 153.985 ;
        RECT 90.890 153.220 91.950 153.360 ;
        RECT 91.810 152.770 91.950 153.220 ;
        RECT 91.750 152.450 92.010 152.770 ;
        RECT 93.590 152.680 93.850 152.770 ;
        RECT 93.190 152.540 93.850 152.680 ;
        RECT 87.610 151.770 87.870 152.090 ;
        RECT 86.230 151.430 86.490 151.750 ;
        RECT 86.290 150.730 86.430 151.430 ;
        RECT 86.230 150.410 86.490 150.730 ;
        RECT 85.770 149.730 86.030 150.050 ;
        RECT 84.850 149.390 85.110 149.710 ;
        RECT 84.910 148.010 85.050 149.390 ;
        RECT 84.850 147.690 85.110 148.010 ;
        RECT 84.390 144.290 84.650 144.610 ;
        RECT 84.450 139.850 84.590 144.290 ;
        RECT 84.910 144.270 85.050 147.690 ;
        RECT 85.830 146.310 85.970 149.730 ;
        RECT 86.290 147.330 86.430 150.410 ;
        RECT 87.670 150.245 87.810 151.770 ;
        RECT 93.190 150.730 93.330 152.540 ;
        RECT 93.590 152.450 93.850 152.540 ;
        RECT 93.590 151.430 93.850 151.750 ;
        RECT 93.650 150.730 93.790 151.430 ;
        RECT 93.130 150.410 93.390 150.730 ;
        RECT 93.590 150.410 93.850 150.730 ;
        RECT 87.600 149.875 87.880 150.245 ;
        RECT 93.590 149.050 93.850 149.370 ;
        RECT 94.050 149.050 94.310 149.370 ;
        RECT 90.370 148.710 90.630 149.030 ;
        RECT 86.230 147.010 86.490 147.330 ;
        RECT 90.430 146.650 90.570 148.710 ;
        RECT 91.590 148.175 93.470 148.545 ;
        RECT 90.830 147.010 91.090 147.330 ;
        RECT 90.370 146.330 90.630 146.650 ;
        RECT 85.770 145.990 86.030 146.310 ;
        RECT 85.830 145.290 85.970 145.990 ;
        RECT 90.890 145.290 91.030 147.010 ;
        RECT 93.650 146.650 93.790 149.050 ;
        RECT 94.110 146.990 94.250 149.050 ;
        RECT 95.030 146.990 95.170 157.210 ;
        RECT 98.250 155.490 98.390 162.650 ;
        RECT 100.090 158.890 100.230 166.390 ;
        RECT 100.030 158.570 100.290 158.890 ;
        RECT 98.190 155.170 98.450 155.490 ;
        RECT 98.650 155.170 98.910 155.490 ;
        RECT 98.710 153.450 98.850 155.170 ;
        RECT 99.570 154.150 99.830 154.470 ;
        RECT 98.650 153.130 98.910 153.450 ;
        RECT 95.430 150.070 95.690 150.390 ;
        RECT 95.490 148.010 95.630 150.070 ;
        RECT 99.100 149.875 99.380 150.245 ;
        RECT 96.350 148.710 96.610 149.030 ;
        RECT 96.410 148.010 96.550 148.710 ;
        RECT 95.430 147.690 95.690 148.010 ;
        RECT 96.350 147.690 96.610 148.010 ;
        RECT 94.050 146.670 94.310 146.990 ;
        RECT 94.970 146.670 95.230 146.990 ;
        RECT 93.590 146.330 93.850 146.650 ;
        RECT 85.770 144.970 86.030 145.290 ;
        RECT 90.830 144.970 91.090 145.290 ;
        RECT 84.850 143.950 85.110 144.270 ;
        RECT 84.390 139.530 84.650 139.850 ;
        RECT 84.450 137.130 84.590 139.530 ;
        RECT 84.910 138.830 85.050 143.950 ;
        RECT 91.590 142.735 93.470 143.105 ;
        RECT 86.230 138.850 86.490 139.170 ;
        RECT 84.850 138.510 85.110 138.830 ;
        RECT 84.910 137.130 85.050 138.510 ;
        RECT 84.390 136.810 84.650 137.130 ;
        RECT 84.850 136.810 85.110 137.130 ;
        RECT 86.290 136.450 86.430 138.850 ;
        RECT 94.110 138.490 94.250 146.670 ;
        RECT 96.410 144.610 96.550 147.690 ;
        RECT 96.810 145.990 97.070 146.310 ;
        RECT 96.870 145.290 97.010 145.990 ;
        RECT 96.810 144.970 97.070 145.290 ;
        RECT 96.350 144.290 96.610 144.610 ;
        RECT 98.650 138.510 98.910 138.830 ;
        RECT 94.050 138.170 94.310 138.490 ;
        RECT 90.830 137.830 91.090 138.150 ;
        RECT 86.690 136.470 86.950 136.790 ;
        RECT 86.230 136.130 86.490 136.450 ;
        RECT 83.930 135.450 84.190 135.770 ;
        RECT 84.850 135.110 85.110 135.430 ;
        RECT 84.910 134.070 85.050 135.110 ;
        RECT 84.850 133.750 85.110 134.070 ;
        RECT 86.290 133.390 86.430 136.130 ;
        RECT 83.470 133.070 83.730 133.390 ;
        RECT 86.230 133.070 86.490 133.390 ;
        RECT 83.010 132.390 83.270 132.710 ;
        RECT 83.070 128.970 83.210 132.390 ;
        RECT 83.010 128.650 83.270 128.970 ;
        RECT 81.630 126.950 81.890 127.270 ;
        RECT 83.470 126.950 83.730 127.270 ;
        RECT 84.390 126.950 84.650 127.270 ;
        RECT 80.250 125.930 80.510 126.250 ;
        RECT 82.550 124.570 82.810 124.890 ;
        RECT 82.610 123.530 82.750 124.570 ;
        RECT 82.550 123.210 82.810 123.530 ;
        RECT 83.530 122.850 83.670 126.950 ;
        RECT 84.450 125.570 84.590 126.950 ;
        RECT 84.390 125.250 84.650 125.570 ;
        RECT 85.310 124.910 85.570 125.230 ;
        RECT 85.370 123.530 85.510 124.910 ;
        RECT 85.310 123.210 85.570 123.530 ;
        RECT 83.010 122.530 83.270 122.850 ;
        RECT 83.470 122.530 83.730 122.850 ;
        RECT 83.070 119.790 83.210 122.530 ;
        RECT 83.470 119.810 83.730 120.130 ;
        RECT 83.010 119.470 83.270 119.790 ;
        RECT 79.330 119.220 79.990 119.360 ;
        RECT 79.330 119.130 79.590 119.220 ;
        RECT 78.870 118.790 79.130 119.110 ;
        RECT 76.590 118.255 78.470 118.625 ;
        RECT 78.930 118.090 79.070 118.790 ;
        RECT 78.870 117.770 79.130 118.090 ;
        RECT 79.390 117.070 79.530 119.130 ;
        RECT 80.710 118.790 80.970 119.110 ;
        RECT 82.550 118.790 82.810 119.110 ;
        RECT 80.770 117.410 80.910 118.790 ;
        RECT 80.710 117.090 80.970 117.410 ;
        RECT 79.330 116.750 79.590 117.070 ;
        RECT 79.390 115.370 79.530 116.750 ;
        RECT 79.330 115.050 79.590 115.370 ;
        RECT 82.610 114.010 82.750 118.790 ;
        RECT 83.070 117.750 83.210 119.470 ;
        RECT 83.010 117.430 83.270 117.750 ;
        RECT 83.530 116.730 83.670 119.810 ;
        RECT 83.930 119.470 84.190 119.790 ;
        RECT 83.990 118.090 84.130 119.470 ;
        RECT 84.390 118.790 84.650 119.110 ;
        RECT 83.930 117.770 84.190 118.090 ;
        RECT 83.470 116.410 83.730 116.730 ;
        RECT 84.450 114.690 84.590 118.790 ;
        RECT 85.310 116.750 85.570 117.070 ;
        RECT 85.370 114.690 85.510 116.750 ;
        RECT 84.390 114.370 84.650 114.690 ;
        RECT 85.310 114.370 85.570 114.690 ;
        RECT 86.230 114.370 86.490 114.690 ;
        RECT 82.550 113.690 82.810 114.010 ;
        RECT 76.590 112.815 78.470 113.185 ;
        RECT 77.950 111.650 78.210 111.970 ;
        RECT 81.170 111.650 81.430 111.970 ;
        RECT 78.010 108.910 78.150 111.650 ;
        RECT 81.230 109.250 81.370 111.650 ;
        RECT 81.630 111.310 81.890 111.630 ;
        RECT 81.170 108.930 81.430 109.250 ;
        RECT 77.950 108.590 78.210 108.910 ;
        RECT 78.870 108.590 79.130 108.910 ;
        RECT 75.650 108.250 75.910 108.570 ;
        RECT 76.590 107.375 78.470 107.745 ;
        RECT 74.730 106.210 74.990 106.530 ;
        RECT 68.290 106.100 68.550 106.190 ;
        RECT 67.890 105.960 68.550 106.100 ;
        RECT 64.150 105.530 64.410 105.850 ;
        RECT 63.690 105.190 63.950 105.510 ;
        RECT 61.590 104.655 63.470 105.025 ;
        RECT 63.750 103.810 63.890 105.190 ;
        RECT 52.190 103.150 52.450 103.470 ;
        RECT 56.390 103.130 56.530 103.750 ;
        RECT 57.710 103.490 57.970 103.810 ;
        RECT 63.690 103.490 63.950 103.810 ;
        RECT 64.210 103.130 64.350 105.530 ;
        RECT 54.490 102.810 54.750 103.130 ;
        RECT 56.330 102.810 56.590 103.130 ;
        RECT 60.930 102.810 61.190 103.130 ;
        RECT 64.150 102.810 64.410 103.130 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 54.550 88.250 54.690 102.810 ;
        RECT 60.990 98.450 61.130 102.810 ;
        RECT 61.590 99.215 63.470 99.585 ;
        RECT 60.990 98.310 62.050 98.450 ;
        RECT 55.530 88.250 56.750 89.190 ;
        RECT 61.910 88.870 62.050 98.310 ;
        RECT 67.890 89.840 68.030 105.960 ;
        RECT 68.290 105.870 68.550 105.960 ;
        RECT 73.350 105.870 73.610 106.190 ;
        RECT 73.410 104.490 73.550 105.870 ;
        RECT 75.650 105.190 75.910 105.510 ;
        RECT 73.350 104.170 73.610 104.490 ;
        RECT 73.410 103.810 73.550 104.170 ;
        RECT 75.710 103.810 75.850 105.190 ;
        RECT 78.930 104.490 79.070 108.590 ;
        RECT 79.330 107.910 79.590 108.230 ;
        RECT 78.870 104.170 79.130 104.490 ;
        RECT 73.350 103.490 73.610 103.810 ;
        RECT 75.650 103.490 75.910 103.810 ;
        RECT 79.390 103.470 79.530 107.910 ;
        RECT 81.690 106.870 81.830 111.310 ;
        RECT 83.470 107.910 83.730 108.230 ;
        RECT 83.530 106.870 83.670 107.910 ;
        RECT 81.630 106.550 81.890 106.870 ;
        RECT 83.470 106.550 83.730 106.870 ;
        RECT 86.290 106.190 86.430 114.370 ;
        RECT 86.750 106.530 86.890 136.470 ;
        RECT 90.890 136.450 91.030 137.830 ;
        RECT 91.590 137.295 93.470 137.665 ;
        RECT 90.830 136.130 91.090 136.450 ;
        RECT 91.290 136.130 91.550 136.450 ;
        RECT 88.070 135.450 88.330 135.770 ;
        RECT 88.130 134.410 88.270 135.450 ;
        RECT 88.070 134.090 88.330 134.410 ;
        RECT 90.370 133.750 90.630 134.070 ;
        RECT 88.070 133.410 88.330 133.730 ;
        RECT 88.130 130.670 88.270 133.410 ;
        RECT 90.430 131.690 90.570 133.750 ;
        RECT 91.350 133.390 91.490 136.130 ;
        RECT 93.130 136.020 93.390 136.110 ;
        RECT 92.730 135.880 93.390 136.020 ;
        RECT 92.730 135.430 92.870 135.880 ;
        RECT 93.130 135.790 93.390 135.880 ;
        RECT 94.110 135.770 94.250 138.170 ;
        RECT 98.190 137.830 98.450 138.150 ;
        RECT 97.730 135.790 97.990 136.110 ;
        RECT 94.050 135.450 94.310 135.770 ;
        RECT 92.670 135.110 92.930 135.430 ;
        RECT 93.590 135.110 93.850 135.430 ;
        RECT 91.290 133.070 91.550 133.390 ;
        RECT 91.590 131.855 93.470 132.225 ;
        RECT 90.370 131.370 90.630 131.690 ;
        RECT 88.070 130.350 88.330 130.670 ;
        RECT 90.830 130.350 91.090 130.670 ;
        RECT 88.070 128.650 88.330 128.970 ;
        RECT 88.130 125.570 88.270 128.650 ;
        RECT 88.070 125.250 88.330 125.570 ;
        RECT 90.890 122.850 91.030 130.350 ;
        RECT 93.650 128.290 93.790 135.110 ;
        RECT 97.790 133.730 97.930 135.790 ;
        RECT 98.250 135.770 98.390 137.830 ;
        RECT 98.710 136.110 98.850 138.510 ;
        RECT 99.170 136.110 99.310 149.875 ;
        RECT 98.650 135.790 98.910 136.110 ;
        RECT 99.110 135.790 99.370 136.110 ;
        RECT 98.190 135.450 98.450 135.770 ;
        RECT 98.250 133.730 98.390 135.450 ;
        RECT 99.170 133.925 99.310 135.790 ;
        RECT 97.730 133.410 97.990 133.730 ;
        RECT 98.190 133.410 98.450 133.730 ;
        RECT 99.100 133.555 99.380 133.925 ;
        RECT 99.630 133.730 99.770 154.150 ;
        RECT 100.030 135.790 100.290 136.110 ;
        RECT 100.090 134.410 100.230 135.790 ;
        RECT 100.030 134.090 100.290 134.410 ;
        RECT 99.570 133.410 99.830 133.730 ;
        RECT 94.970 133.070 95.230 133.390 ;
        RECT 94.510 132.390 94.770 132.710 ;
        RECT 93.590 127.970 93.850 128.290 ;
        RECT 91.350 127.610 93.790 127.690 ;
        RECT 91.290 127.550 93.790 127.610 ;
        RECT 91.290 127.290 91.550 127.550 ;
        RECT 91.590 126.415 93.470 126.785 ;
        RECT 93.130 124.570 93.390 124.890 ;
        RECT 93.190 123.530 93.330 124.570 ;
        RECT 93.130 123.210 93.390 123.530 ;
        RECT 90.830 122.530 91.090 122.850 ;
        RECT 91.590 120.975 93.470 121.345 ;
        RECT 93.130 119.470 93.390 119.790 ;
        RECT 87.150 118.790 87.410 119.110 ;
        RECT 87.210 117.410 87.350 118.790 ;
        RECT 93.190 118.090 93.330 119.470 ;
        RECT 93.650 119.110 93.790 127.550 ;
        RECT 93.590 118.790 93.850 119.110 ;
        RECT 93.130 117.770 93.390 118.090 ;
        RECT 87.150 117.090 87.410 117.410 ;
        RECT 93.650 117.070 93.790 118.790 ;
        RECT 93.590 116.750 93.850 117.070 ;
        RECT 88.070 116.070 88.330 116.390 ;
        RECT 90.830 116.070 91.090 116.390 ;
        RECT 88.130 114.690 88.270 116.070 ;
        RECT 88.070 114.370 88.330 114.690 ;
        RECT 90.890 114.010 91.030 116.070 ;
        RECT 91.590 115.535 93.470 115.905 ;
        RECT 93.650 115.370 93.790 116.750 ;
        RECT 93.590 115.050 93.850 115.370 ;
        RECT 90.830 113.690 91.090 114.010 ;
        RECT 92.660 112.475 92.940 112.845 ;
        RECT 92.730 112.310 92.870 112.475 ;
        RECT 92.670 111.990 92.930 112.310 ;
        RECT 91.590 110.095 93.470 110.465 ;
        RECT 94.570 108.910 94.710 132.390 ;
        RECT 95.030 128.970 95.170 133.070 ;
        RECT 98.250 130.670 98.390 133.410 ;
        RECT 100.550 133.390 100.690 175.910 ;
        RECT 100.940 163.475 101.220 163.845 ;
        RECT 101.010 163.310 101.150 163.475 ;
        RECT 100.950 162.990 101.210 163.310 ;
        RECT 101.410 151.430 101.670 151.750 ;
        RECT 100.950 135.110 101.210 135.430 ;
        RECT 101.010 134.070 101.150 135.110 ;
        RECT 100.950 133.750 101.210 134.070 ;
        RECT 100.490 133.070 100.750 133.390 ;
        RECT 99.570 132.390 99.830 132.710 ;
        RECT 100.950 132.390 101.210 132.710 ;
        RECT 98.190 130.350 98.450 130.670 ;
        RECT 94.970 128.650 95.230 128.970 ;
        RECT 95.420 128.795 95.700 129.165 ;
        RECT 98.250 128.970 98.390 130.350 ;
        RECT 95.490 128.630 95.630 128.795 ;
        RECT 98.190 128.650 98.450 128.970 ;
        RECT 95.430 128.310 95.690 128.630 ;
        RECT 98.250 125.570 98.390 128.650 ;
        RECT 98.650 127.630 98.910 127.950 ;
        RECT 98.710 126.250 98.850 127.630 ;
        RECT 98.650 125.930 98.910 126.250 ;
        RECT 98.190 125.250 98.450 125.570 ;
        RECT 99.110 124.910 99.370 125.230 ;
        RECT 99.170 119.790 99.310 124.910 ;
        RECT 99.110 119.470 99.370 119.790 ;
        RECT 99.630 108.910 99.770 132.390 ;
        RECT 100.030 131.030 100.290 131.350 ;
        RECT 100.090 128.290 100.230 131.030 ;
        RECT 100.030 127.970 100.290 128.290 ;
        RECT 100.090 125.230 100.230 127.970 ;
        RECT 101.010 125.230 101.150 132.390 ;
        RECT 100.030 124.910 100.290 125.230 ;
        RECT 100.950 124.910 101.210 125.230 ;
        RECT 100.030 122.530 100.290 122.850 ;
        RECT 100.090 119.790 100.230 122.530 ;
        RECT 100.030 119.470 100.290 119.790 ;
        RECT 100.950 118.790 101.210 119.110 ;
        RECT 100.030 116.750 100.290 117.070 ;
        RECT 100.090 115.370 100.230 116.750 ;
        RECT 100.030 115.050 100.290 115.370 ;
        RECT 101.010 114.350 101.150 118.790 ;
        RECT 100.950 114.030 101.210 114.350 ;
        RECT 101.470 113.670 101.610 151.430 ;
        RECT 101.930 133.390 102.070 175.910 ;
        RECT 102.330 167.750 102.590 168.070 ;
        RECT 102.390 160.930 102.530 167.750 ;
        RECT 102.330 160.610 102.590 160.930 ;
        RECT 102.390 159.770 102.530 160.610 ;
        RECT 102.390 159.630 102.990 159.770 ;
        RECT 102.330 155.850 102.590 156.170 ;
        RECT 102.390 154.810 102.530 155.850 ;
        RECT 102.850 155.830 102.990 159.630 ;
        RECT 102.790 155.510 103.050 155.830 ;
        RECT 102.330 154.490 102.590 154.810 ;
        RECT 102.790 153.360 103.050 153.450 ;
        RECT 102.390 153.220 103.050 153.360 ;
        RECT 102.390 146.730 102.530 153.220 ;
        RECT 102.790 153.130 103.050 153.220 ;
        RECT 103.310 150.810 103.450 181.950 ;
        RECT 104.630 181.350 104.890 181.670 ;
        RECT 104.690 179.970 104.830 181.350 ;
        RECT 104.630 179.650 104.890 179.970 ;
        RECT 104.630 174.100 104.890 174.190 ;
        RECT 105.150 174.100 105.290 185.090 ;
        RECT 105.550 184.750 105.810 185.070 ;
        RECT 105.610 183.370 105.750 184.750 ;
        RECT 106.590 183.535 108.470 183.905 ;
        RECT 105.550 183.050 105.810 183.370 ;
        RECT 105.550 182.370 105.810 182.690 ;
        RECT 106.010 182.370 106.270 182.690 ;
        RECT 107.850 182.370 108.110 182.690 ;
        RECT 109.230 182.370 109.490 182.690 ;
        RECT 105.610 180.650 105.750 182.370 ;
        RECT 105.550 180.330 105.810 180.650 ;
        RECT 105.550 179.650 105.810 179.970 ;
        RECT 105.610 176.910 105.750 179.650 ;
        RECT 106.070 177.160 106.210 182.370 ;
        RECT 107.910 179.970 108.050 182.370 ;
        RECT 107.850 179.650 108.110 179.970 ;
        RECT 108.770 179.310 109.030 179.630 ;
        RECT 106.590 178.095 108.470 178.465 ;
        RECT 108.830 177.590 108.970 179.310 ;
        RECT 108.770 177.270 109.030 177.590 ;
        RECT 109.290 177.250 109.430 182.370 ;
        RECT 106.470 177.160 106.730 177.250 ;
        RECT 106.070 177.020 106.730 177.160 ;
        RECT 106.470 176.930 106.730 177.020 ;
        RECT 107.850 176.930 108.110 177.250 ;
        RECT 109.230 176.930 109.490 177.250 ;
        RECT 105.550 176.590 105.810 176.910 ;
        RECT 105.610 174.190 105.750 176.590 ;
        RECT 106.010 174.890 106.270 175.210 ;
        RECT 104.630 173.960 105.290 174.100 ;
        RECT 104.630 173.870 104.890 173.960 ;
        RECT 105.550 173.870 105.810 174.190 ;
        RECT 104.170 173.530 104.430 173.850 ;
        RECT 103.710 154.150 103.970 154.470 ;
        RECT 102.850 150.670 103.450 150.810 ;
        RECT 102.850 147.330 102.990 150.670 ;
        RECT 103.250 150.070 103.510 150.390 ;
        RECT 103.310 148.010 103.450 150.070 ;
        RECT 103.250 147.690 103.510 148.010 ;
        RECT 102.790 147.010 103.050 147.330 ;
        RECT 102.390 146.590 102.990 146.730 ;
        RECT 102.330 139.190 102.590 139.510 ;
        RECT 102.390 134.410 102.530 139.190 ;
        RECT 102.330 134.090 102.590 134.410 ;
        RECT 102.330 133.410 102.590 133.730 ;
        RECT 101.870 133.070 102.130 133.390 ;
        RECT 102.390 131.350 102.530 133.410 ;
        RECT 102.330 131.030 102.590 131.350 ;
        RECT 102.850 127.610 102.990 146.590 ;
        RECT 103.770 133.730 103.910 154.150 ;
        RECT 104.230 152.770 104.370 173.530 ;
        RECT 106.070 172.150 106.210 174.890 ;
        RECT 106.530 174.530 106.670 176.930 ;
        RECT 107.910 175.210 108.050 176.930 ;
        RECT 107.850 174.890 108.110 175.210 ;
        RECT 108.770 174.550 109.030 174.870 ;
        RECT 106.470 174.210 106.730 174.530 ;
        RECT 106.590 172.655 108.470 173.025 ;
        RECT 106.010 171.830 106.270 172.150 ;
        RECT 105.550 171.150 105.810 171.470 ;
        RECT 105.610 166.030 105.750 171.150 ;
        RECT 106.930 170.470 107.190 170.790 ;
        RECT 106.990 168.410 107.130 170.470 ;
        RECT 106.930 168.090 107.190 168.410 ;
        RECT 106.590 167.215 108.470 167.585 ;
        RECT 104.630 165.710 104.890 166.030 ;
        RECT 105.550 165.710 105.810 166.030 ;
        RECT 104.690 158.890 104.830 165.710 ;
        RECT 105.090 162.310 105.350 162.630 ;
        RECT 104.630 158.570 104.890 158.890 ;
        RECT 105.150 157.870 105.290 162.310 ;
        RECT 105.610 160.590 105.750 165.710 ;
        RECT 108.830 165.690 108.970 174.550 ;
        RECT 109.750 174.190 109.890 187.810 ;
        RECT 110.150 184.750 110.410 185.070 ;
        RECT 110.210 182.010 110.350 184.750 ;
        RECT 110.670 182.350 110.810 192.910 ;
        RECT 111.990 192.570 112.250 192.890 ;
        RECT 112.050 184.730 112.190 192.570 ;
        RECT 112.510 191.530 112.650 193.930 ;
        RECT 115.670 193.250 115.930 193.570 ;
        RECT 112.450 191.210 112.710 191.530 ;
        RECT 112.910 189.510 113.170 189.830 ;
        RECT 112.970 188.130 113.110 189.510 ;
        RECT 112.910 187.810 113.170 188.130 ;
        RECT 111.990 184.410 112.250 184.730 ;
        RECT 111.530 184.070 111.790 184.390 ;
        RECT 111.590 182.690 111.730 184.070 ;
        RECT 111.530 182.370 111.790 182.690 ;
        RECT 110.610 182.030 110.870 182.350 ;
        RECT 110.150 181.690 110.410 182.010 ;
        RECT 109.230 173.870 109.490 174.190 ;
        RECT 109.690 173.870 109.950 174.190 ;
        RECT 109.290 171.810 109.430 173.870 ;
        RECT 109.690 173.190 109.950 173.510 ;
        RECT 109.750 171.810 109.890 173.190 ;
        RECT 110.210 172.150 110.350 181.690 ;
        RECT 110.670 176.910 110.810 182.030 ;
        RECT 111.590 177.930 111.730 182.370 ;
        RECT 112.050 177.930 112.190 184.410 ;
        RECT 115.730 179.970 115.870 193.250 ;
        RECT 117.570 191.530 117.710 195.290 ;
        RECT 118.030 193.910 118.170 195.290 ;
        RECT 117.970 193.590 118.230 193.910 ;
        RECT 117.510 191.210 117.770 191.530 ;
        RECT 118.030 190.510 118.170 193.590 ;
        RECT 118.890 192.230 119.150 192.550 ;
        RECT 118.950 190.510 119.090 192.230 ;
        RECT 121.590 191.695 123.470 192.065 ;
        RECT 117.970 190.190 118.230 190.510 ;
        RECT 118.890 190.190 119.150 190.510 ;
        RECT 116.130 189.850 116.390 190.170 ;
        RECT 116.190 188.810 116.330 189.850 ;
        RECT 116.130 188.490 116.390 188.810 ;
        RECT 118.030 187.790 118.170 190.190 ;
        RECT 117.970 187.470 118.230 187.790 ;
        RECT 117.510 182.370 117.770 182.690 ;
        RECT 116.590 181.350 116.850 181.670 ;
        RECT 115.670 179.650 115.930 179.970 ;
        RECT 111.530 177.610 111.790 177.930 ;
        RECT 111.990 177.610 112.250 177.930 ;
        RECT 116.650 177.250 116.790 181.350 ;
        RECT 117.570 180.650 117.710 182.370 ;
        RECT 118.030 182.350 118.170 187.470 ;
        RECT 121.590 186.255 123.470 186.625 ;
        RECT 124.410 182.710 124.670 183.030 ;
        RECT 117.970 182.030 118.230 182.350 ;
        RECT 117.510 180.330 117.770 180.650 ;
        RECT 118.030 178.950 118.170 182.030 ;
        RECT 121.590 180.815 123.470 181.185 ;
        RECT 124.470 180.650 124.610 182.710 ;
        RECT 124.410 180.330 124.670 180.650 ;
        RECT 121.650 179.310 121.910 179.630 ;
        RECT 118.430 178.970 118.690 179.290 ;
        RECT 117.970 178.630 118.230 178.950 ;
        RECT 118.490 177.930 118.630 178.970 ;
        RECT 118.430 177.610 118.690 177.930 ;
        RECT 121.710 177.590 121.850 179.310 ;
        RECT 121.650 177.270 121.910 177.590 ;
        RECT 116.590 176.930 116.850 177.250 ;
        RECT 110.610 176.590 110.870 176.910 ;
        RECT 121.590 175.375 123.470 175.745 ;
        RECT 118.890 173.870 119.150 174.190 ;
        RECT 117.970 173.190 118.230 173.510 ;
        RECT 118.030 172.150 118.170 173.190 ;
        RECT 118.950 172.490 119.090 173.870 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 118.890 172.170 119.150 172.490 ;
        RECT 110.150 171.830 110.410 172.150 ;
        RECT 117.970 171.830 118.230 172.150 ;
        RECT 109.230 171.490 109.490 171.810 ;
        RECT 109.690 171.490 109.950 171.810 ;
        RECT 114.290 170.810 114.550 171.130 ;
        RECT 111.070 170.470 111.330 170.790 ;
        RECT 113.370 170.470 113.630 170.790 ;
        RECT 109.690 168.770 109.950 169.090 ;
        RECT 108.770 165.370 109.030 165.690 ;
        RECT 109.750 164.410 109.890 168.770 ;
        RECT 110.150 168.090 110.410 168.410 ;
        RECT 110.210 167.050 110.350 168.090 ;
        RECT 110.610 167.750 110.870 168.070 ;
        RECT 110.150 166.730 110.410 167.050 ;
        RECT 110.670 166.370 110.810 167.750 ;
        RECT 110.610 166.050 110.870 166.370 ;
        RECT 110.610 165.370 110.870 165.690 ;
        RECT 109.290 164.270 109.890 164.410 ;
        RECT 108.770 163.670 109.030 163.990 ;
        RECT 106.010 162.650 106.270 162.970 ;
        RECT 106.070 161.610 106.210 162.650 ;
        RECT 106.590 161.775 108.470 162.145 ;
        RECT 106.010 161.290 106.270 161.610 ;
        RECT 105.550 160.270 105.810 160.590 ;
        RECT 108.830 157.870 108.970 163.670 ;
        RECT 109.290 158.550 109.430 164.270 ;
        RECT 110.150 163.330 110.410 163.650 ;
        RECT 109.690 162.310 109.950 162.630 ;
        RECT 109.750 161.610 109.890 162.310 ;
        RECT 109.690 161.290 109.950 161.610 ;
        RECT 110.210 160.930 110.350 163.330 ;
        RECT 110.150 160.610 110.410 160.930 ;
        RECT 110.670 160.330 110.810 165.370 ;
        RECT 110.210 160.190 110.810 160.330 ;
        RECT 109.230 158.230 109.490 158.550 ;
        RECT 105.090 157.550 105.350 157.870 ;
        RECT 108.770 157.550 109.030 157.870 ;
        RECT 109.230 157.550 109.490 157.870 ;
        RECT 109.690 157.550 109.950 157.870 ;
        RECT 108.770 156.870 109.030 157.190 ;
        RECT 106.590 156.335 108.470 156.705 ;
        RECT 108.310 155.850 108.570 156.170 ;
        RECT 105.090 155.170 105.350 155.490 ;
        RECT 105.150 153.110 105.290 155.170 ;
        RECT 106.470 154.150 106.730 154.470 ;
        RECT 105.090 152.790 105.350 153.110 ;
        RECT 104.170 152.450 104.430 152.770 ;
        RECT 106.530 152.430 106.670 154.150 ;
        RECT 107.850 152.790 108.110 153.110 ;
        RECT 106.470 152.110 106.730 152.430 ;
        RECT 107.390 152.340 107.650 152.430 ;
        RECT 107.910 152.340 108.050 152.790 ;
        RECT 108.370 152.430 108.510 155.850 ;
        RECT 107.390 152.200 108.050 152.340 ;
        RECT 107.390 152.110 107.650 152.200 ;
        RECT 108.310 152.110 108.570 152.430 ;
        RECT 104.630 151.770 104.890 152.090 ;
        RECT 104.690 150.730 104.830 151.770 ;
        RECT 108.370 151.750 108.510 152.110 ;
        RECT 105.090 151.430 105.350 151.750 ;
        RECT 108.310 151.430 108.570 151.750 ;
        RECT 104.630 150.410 104.890 150.730 ;
        RECT 104.170 147.690 104.430 148.010 ;
        RECT 103.710 133.410 103.970 133.730 ;
        RECT 103.250 132.390 103.510 132.710 ;
        RECT 102.790 127.290 103.050 127.610 ;
        RECT 102.330 119.130 102.590 119.450 ;
        RECT 102.390 118.090 102.530 119.130 ;
        RECT 102.330 117.770 102.590 118.090 ;
        RECT 101.410 113.350 101.670 113.670 ;
        RECT 103.310 108.910 103.450 132.390 ;
        RECT 104.230 111.630 104.370 147.690 ;
        RECT 105.150 146.990 105.290 151.430 ;
        RECT 106.590 150.895 108.470 151.265 ;
        RECT 107.380 149.875 107.660 150.245 ;
        RECT 107.450 149.710 107.590 149.875 ;
        RECT 107.850 149.730 108.110 150.050 ;
        RECT 107.390 149.390 107.650 149.710 ;
        RECT 106.010 147.690 106.270 148.010 ;
        RECT 105.090 146.670 105.350 146.990 ;
        RECT 105.090 138.510 105.350 138.830 ;
        RECT 105.150 137.130 105.290 138.510 ;
        RECT 105.090 136.810 105.350 137.130 ;
        RECT 104.630 132.390 104.890 132.710 ;
        RECT 104.690 128.970 104.830 132.390 ;
        RECT 106.070 128.970 106.210 147.690 ;
        RECT 107.450 147.330 107.590 149.390 ;
        RECT 107.390 147.010 107.650 147.330 ;
        RECT 107.910 146.990 108.050 149.730 ;
        RECT 107.850 146.670 108.110 146.990 ;
        RECT 107.910 146.310 108.050 146.670 ;
        RECT 107.850 145.990 108.110 146.310 ;
        RECT 106.590 145.455 108.470 145.825 ;
        RECT 108.830 144.610 108.970 156.870 ;
        RECT 109.290 155.490 109.430 157.550 ;
        RECT 109.230 155.170 109.490 155.490 ;
        RECT 109.290 152.430 109.430 155.170 ;
        RECT 109.750 153.450 109.890 157.550 ;
        RECT 109.690 153.130 109.950 153.450 ;
        RECT 109.750 152.770 109.890 153.130 ;
        RECT 109.690 152.450 109.950 152.770 ;
        RECT 109.230 152.110 109.490 152.430 ;
        RECT 109.690 149.730 109.950 150.050 ;
        RECT 109.750 146.990 109.890 149.730 ;
        RECT 109.690 146.670 109.950 146.990 ;
        RECT 109.230 145.990 109.490 146.310 ;
        RECT 109.290 144.610 109.430 145.990 ;
        RECT 108.770 144.290 109.030 144.610 ;
        RECT 109.230 144.290 109.490 144.610 ;
        RECT 109.750 144.010 109.890 146.670 ;
        RECT 110.210 144.270 110.350 160.190 ;
        RECT 110.610 159.590 110.870 159.910 ;
        RECT 110.670 155.830 110.810 159.590 ;
        RECT 110.610 155.510 110.870 155.830 ;
        RECT 110.610 154.150 110.870 154.470 ;
        RECT 108.770 143.610 109.030 143.930 ;
        RECT 109.290 143.870 109.890 144.010 ;
        RECT 110.150 143.950 110.410 144.270 ;
        RECT 108.830 142.570 108.970 143.610 ;
        RECT 108.770 142.250 109.030 142.570 ;
        RECT 106.590 140.015 108.470 140.385 ;
        RECT 109.290 139.170 109.430 143.870 ;
        RECT 109.690 143.270 109.950 143.590 ;
        RECT 110.150 143.270 110.410 143.590 ;
        RECT 109.230 138.850 109.490 139.170 ;
        RECT 108.770 135.450 109.030 135.770 ;
        RECT 106.590 134.575 108.470 134.945 ;
        RECT 107.840 133.555 108.120 133.925 ;
        RECT 108.830 133.730 108.970 135.450 ;
        RECT 109.290 133.730 109.430 138.850 ;
        RECT 107.850 133.410 108.110 133.555 ;
        RECT 108.770 133.410 109.030 133.730 ;
        RECT 109.230 133.410 109.490 133.730 ;
        RECT 109.750 131.690 109.890 143.270 ;
        RECT 110.210 139.510 110.350 143.270 ;
        RECT 110.150 139.190 110.410 139.510 ;
        RECT 110.210 134.070 110.350 139.190 ;
        RECT 110.150 133.750 110.410 134.070 ;
        RECT 110.670 133.730 110.810 154.150 ;
        RECT 111.130 133.730 111.270 170.470 ;
        RECT 112.450 168.770 112.710 169.090 ;
        RECT 111.530 168.430 111.790 168.750 ;
        RECT 111.590 166.030 111.730 168.430 ;
        RECT 111.990 166.050 112.250 166.370 ;
        RECT 111.530 165.710 111.790 166.030 ;
        RECT 112.050 165.690 112.190 166.050 ;
        RECT 111.990 165.370 112.250 165.690 ;
        RECT 111.530 162.650 111.790 162.970 ;
        RECT 111.590 158.290 111.730 162.650 ;
        RECT 112.050 158.890 112.190 165.370 ;
        RECT 112.510 163.310 112.650 168.770 ;
        RECT 112.910 167.750 113.170 168.070 ;
        RECT 112.970 164.330 113.110 167.750 ;
        RECT 112.910 164.010 113.170 164.330 ;
        RECT 112.970 163.310 113.110 164.010 ;
        RECT 112.450 162.990 112.710 163.310 ;
        RECT 112.910 162.990 113.170 163.310 ;
        RECT 112.510 160.590 112.650 162.990 ;
        RECT 112.450 160.270 112.710 160.590 ;
        RECT 111.990 158.570 112.250 158.890 ;
        RECT 111.590 158.150 112.190 158.290 ;
        RECT 111.530 157.550 111.790 157.870 ;
        RECT 111.590 156.170 111.730 157.550 ;
        RECT 112.050 157.530 112.190 158.150 ;
        RECT 111.990 157.210 112.250 157.530 ;
        RECT 111.530 155.850 111.790 156.170 ;
        RECT 112.050 151.750 112.190 157.210 ;
        RECT 112.970 155.490 113.110 162.990 ;
        RECT 113.430 162.970 113.570 170.470 ;
        RECT 114.350 168.750 114.490 170.810 ;
        RECT 117.050 170.470 117.310 170.790 ;
        RECT 117.110 169.090 117.250 170.470 ;
        RECT 117.050 168.770 117.310 169.090 ;
        RECT 114.290 168.430 114.550 168.750 ;
        RECT 113.830 165.030 114.090 165.350 ;
        RECT 113.370 162.650 113.630 162.970 ;
        RECT 113.890 160.930 114.030 165.030 ;
        RECT 113.830 160.610 114.090 160.930 ;
        RECT 112.910 155.170 113.170 155.490 ;
        RECT 114.350 153.110 114.490 168.430 ;
        RECT 117.110 161.610 117.250 168.770 ;
        RECT 116.130 161.290 116.390 161.610 ;
        RECT 117.050 161.290 117.310 161.610 ;
        RECT 114.290 152.790 114.550 153.110 ;
        RECT 116.190 152.770 116.330 161.290 ;
        RECT 118.950 160.930 119.090 172.170 ;
        RECT 121.190 171.150 121.450 171.470 ;
        RECT 124.410 171.150 124.670 171.470 ;
        RECT 121.250 169.770 121.390 171.150 ;
        RECT 121.590 169.935 123.470 170.305 ;
        RECT 121.190 169.450 121.450 169.770 ;
        RECT 119.350 166.390 119.610 166.710 ;
        RECT 119.410 161.610 119.550 166.390 ;
        RECT 124.470 166.370 124.610 171.150 ;
        RECT 127.620 170.955 127.900 171.325 ;
        RECT 127.690 168.750 127.830 170.955 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 127.630 168.430 127.890 168.750 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 124.410 166.050 124.670 166.370 ;
        RECT 121.190 165.030 121.450 165.350 ;
        RECT 121.250 161.610 121.390 165.030 ;
        RECT 121.590 164.495 123.470 164.865 ;
        RECT 124.470 163.650 124.610 166.050 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 124.410 163.330 124.670 163.650 ;
        RECT 123.490 162.990 123.750 163.310 ;
        RECT 119.350 161.290 119.610 161.610 ;
        RECT 121.190 161.290 121.450 161.610 ;
        RECT 123.550 161.270 123.690 162.990 ;
        RECT 123.490 160.950 123.750 161.270 ;
        RECT 118.890 160.610 119.150 160.930 ;
        RECT 120.730 160.610 120.990 160.930 ;
        RECT 116.590 159.590 116.850 159.910 ;
        RECT 116.650 158.210 116.790 159.590 ;
        RECT 120.790 158.890 120.930 160.610 ;
        RECT 121.590 159.055 123.470 159.425 ;
        RECT 120.730 158.570 120.990 158.890 ;
        RECT 116.590 157.890 116.850 158.210 ;
        RECT 117.510 154.830 117.770 155.150 ;
        RECT 116.130 152.450 116.390 152.770 ;
        RECT 115.670 151.770 115.930 152.090 ;
        RECT 111.990 151.430 112.250 151.750 ;
        RECT 111.530 149.050 111.790 149.370 ;
        RECT 111.590 144.610 111.730 149.050 ;
        RECT 113.830 148.710 114.090 149.030 ;
        RECT 112.910 147.010 113.170 147.330 ;
        RECT 111.990 146.670 112.250 146.990 ;
        RECT 111.530 144.290 111.790 144.610 ;
        RECT 112.050 144.520 112.190 146.670 ;
        RECT 112.450 144.520 112.710 144.610 ;
        RECT 112.050 144.380 112.710 144.520 ;
        RECT 112.450 144.290 112.710 144.380 ;
        RECT 111.590 143.330 111.730 144.290 ;
        RECT 112.970 144.180 113.110 147.010 ;
        RECT 113.890 146.310 114.030 148.710 ;
        RECT 115.730 148.010 115.870 151.770 ;
        RECT 116.590 150.300 116.850 150.390 ;
        RECT 117.570 150.300 117.710 154.830 ;
        RECT 121.590 153.615 123.470 153.985 ;
        RECT 119.350 152.110 119.610 152.430 ;
        RECT 117.970 151.430 118.230 151.750 ;
        RECT 118.030 150.390 118.170 151.430 ;
        RECT 116.590 150.160 117.710 150.300 ;
        RECT 116.590 150.070 116.850 150.160 ;
        RECT 115.670 147.690 115.930 148.010 ;
        RECT 117.570 147.240 117.710 150.160 ;
        RECT 117.970 150.070 118.230 150.390 ;
        RECT 117.570 147.100 118.170 147.240 ;
        RECT 117.510 146.330 117.770 146.650 ;
        RECT 113.830 145.990 114.090 146.310 ;
        RECT 117.050 145.990 117.310 146.310 ;
        RECT 117.110 145.290 117.250 145.990 ;
        RECT 117.050 144.970 117.310 145.290 ;
        RECT 117.570 144.270 117.710 146.330 ;
        RECT 113.370 144.180 113.630 144.270 ;
        RECT 112.970 144.040 113.630 144.180 ;
        RECT 111.590 143.190 112.650 143.330 ;
        RECT 111.530 142.250 111.790 142.570 ;
        RECT 110.610 133.410 110.870 133.730 ;
        RECT 111.070 133.410 111.330 133.730 ;
        RECT 110.150 132.390 110.410 132.710 ;
        RECT 111.070 132.390 111.330 132.710 ;
        RECT 109.690 131.370 109.950 131.690 ;
        RECT 106.590 129.135 108.470 129.505 ;
        RECT 104.630 128.650 104.890 128.970 ;
        RECT 106.010 128.650 106.270 128.970 ;
        RECT 106.010 127.970 106.270 128.290 ;
        RECT 105.090 127.630 105.350 127.950 ;
        RECT 105.150 125.230 105.290 127.630 ;
        RECT 105.090 124.910 105.350 125.230 ;
        RECT 105.090 122.190 105.350 122.510 ;
        RECT 105.150 120.130 105.290 122.190 ;
        RECT 105.090 119.810 105.350 120.130 ;
        RECT 106.070 119.450 106.210 127.970 ;
        RECT 109.230 127.630 109.490 127.950 ;
        RECT 106.590 123.695 108.470 124.065 ;
        RECT 109.290 120.130 109.430 127.630 ;
        RECT 109.230 119.810 109.490 120.130 ;
        RECT 106.010 119.130 106.270 119.450 ;
        RECT 105.550 118.790 105.810 119.110 ;
        RECT 108.770 118.790 109.030 119.110 ;
        RECT 105.610 117.750 105.750 118.790 ;
        RECT 106.590 118.255 108.470 118.625 ;
        RECT 105.550 117.430 105.810 117.750 ;
        RECT 108.830 114.350 108.970 118.790 ;
        RECT 109.290 114.350 109.430 119.810 ;
        RECT 109.690 117.090 109.950 117.410 ;
        RECT 109.750 115.370 109.890 117.090 ;
        RECT 109.690 115.050 109.950 115.370 ;
        RECT 108.770 114.030 109.030 114.350 ;
        RECT 109.230 114.030 109.490 114.350 ;
        RECT 106.590 112.815 108.470 113.185 ;
        RECT 104.170 111.310 104.430 111.630 ;
        RECT 110.210 108.910 110.350 132.390 ;
        RECT 110.610 130.350 110.870 130.670 ;
        RECT 110.670 128.290 110.810 130.350 ;
        RECT 111.130 128.970 111.270 132.390 ;
        RECT 111.070 128.650 111.330 128.970 ;
        RECT 111.590 128.370 111.730 142.250 ;
        RECT 111.990 139.190 112.250 139.510 ;
        RECT 112.050 134.070 112.190 139.190 ;
        RECT 112.510 139.170 112.650 143.190 ;
        RECT 112.970 141.890 113.110 144.040 ;
        RECT 113.370 143.950 113.630 144.040 ;
        RECT 117.510 143.950 117.770 144.270 ;
        RECT 112.910 141.570 113.170 141.890 ;
        RECT 112.450 138.850 112.710 139.170 ;
        RECT 112.450 138.170 112.710 138.490 ;
        RECT 112.510 136.110 112.650 138.170 ;
        RECT 112.970 136.790 113.110 141.570 ;
        RECT 117.570 141.550 117.710 143.950 ;
        RECT 117.510 141.230 117.770 141.550 ;
        RECT 117.050 140.550 117.310 140.870 ;
        RECT 117.110 139.510 117.250 140.550 ;
        RECT 117.050 139.190 117.310 139.510 ;
        RECT 115.670 138.850 115.930 139.170 ;
        RECT 112.910 136.470 113.170 136.790 ;
        RECT 112.450 135.790 112.710 136.110 ;
        RECT 115.730 135.770 115.870 138.850 ;
        RECT 115.670 135.450 115.930 135.770 ;
        RECT 112.910 135.110 113.170 135.430 ;
        RECT 111.990 133.750 112.250 134.070 ;
        RECT 112.970 133.730 113.110 135.110 ;
        RECT 112.910 133.410 113.170 133.730 ;
        RECT 118.030 131.350 118.170 147.100 ;
        RECT 119.410 144.610 119.550 152.110 ;
        RECT 123.030 151.430 123.290 151.750 ;
        RECT 123.090 150.390 123.230 151.430 ;
        RECT 123.030 150.070 123.290 150.390 ;
        RECT 125.790 149.390 126.050 149.710 ;
        RECT 121.590 148.175 123.470 148.545 ;
        RECT 125.850 146.990 125.990 149.390 ;
        RECT 123.490 146.670 123.750 146.990 ;
        RECT 125.790 146.670 126.050 146.990 ;
        RECT 119.810 146.330 120.070 146.650 ;
        RECT 119.870 145.290 120.010 146.330 ;
        RECT 123.550 145.290 123.690 146.670 ;
        RECT 119.810 144.970 120.070 145.290 ;
        RECT 123.490 144.970 123.750 145.290 ;
        RECT 119.350 144.290 119.610 144.610 ;
        RECT 119.410 141.550 119.550 144.290 ;
        RECT 121.590 142.735 123.470 143.105 ;
        RECT 119.350 141.290 119.610 141.550 ;
        RECT 119.350 141.230 120.010 141.290 ;
        RECT 119.410 141.150 120.010 141.230 ;
        RECT 119.350 140.550 119.610 140.870 ;
        RECT 119.410 137.130 119.550 140.550 ;
        RECT 119.870 138.490 120.010 141.150 ;
        RECT 120.270 140.550 120.530 140.870 ;
        RECT 120.330 139.510 120.470 140.550 ;
        RECT 120.270 139.190 120.530 139.510 ;
        RECT 123.950 138.850 124.210 139.170 ;
        RECT 119.810 138.170 120.070 138.490 ;
        RECT 121.190 137.830 121.450 138.150 ;
        RECT 119.350 136.810 119.610 137.130 ;
        RECT 121.250 136.450 121.390 137.830 ;
        RECT 121.590 137.295 123.470 137.665 ;
        RECT 124.010 137.130 124.150 138.850 ;
        RECT 125.850 138.830 125.990 146.670 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 125.790 138.510 126.050 138.830 ;
        RECT 124.410 137.830 124.670 138.150 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 123.950 136.810 124.210 137.130 ;
        RECT 121.190 136.130 121.450 136.450 ;
        RECT 120.730 135.790 120.990 136.110 ;
        RECT 120.790 134.410 120.930 135.790 ;
        RECT 120.730 134.090 120.990 134.410 ;
        RECT 121.590 131.855 123.470 132.225 ;
        RECT 117.970 131.030 118.230 131.350 ;
        RECT 111.990 130.350 112.250 130.670 ;
        RECT 110.610 127.970 110.870 128.290 ;
        RECT 111.130 128.230 111.730 128.370 ;
        RECT 110.610 109.270 110.870 109.590 ;
        RECT 94.510 108.590 94.770 108.910 ;
        RECT 99.570 108.590 99.830 108.910 ;
        RECT 103.250 108.590 103.510 108.910 ;
        RECT 110.150 108.590 110.410 108.910 ;
        RECT 102.330 108.250 102.590 108.570 ;
        RECT 87.610 107.910 87.870 108.230 ;
        RECT 92.670 107.910 92.930 108.230 ;
        RECT 97.730 107.910 97.990 108.230 ;
        RECT 99.570 107.910 99.830 108.230 ;
        RECT 86.690 106.210 86.950 106.530 ;
        RECT 79.790 105.870 80.050 106.190 ;
        RECT 86.230 105.870 86.490 106.190 ;
        RECT 79.330 103.150 79.590 103.470 ;
        RECT 73.810 102.810 74.070 103.130 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 54.550 88.110 56.750 88.250 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 88.110 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.870 88.800 74.010 102.810 ;
        RECT 76.590 101.935 78.470 102.305 ;
        RECT 79.850 88.800 79.990 105.870 ;
        RECT 86.290 103.810 86.430 105.870 ;
        RECT 86.230 103.490 86.490 103.810 ;
        RECT 87.670 103.130 87.810 107.910 ;
        RECT 92.730 106.870 92.870 107.910 ;
        RECT 93.590 106.890 93.850 107.210 ;
        RECT 92.670 106.550 92.930 106.870 ;
        RECT 88.070 105.190 88.330 105.510 ;
        RECT 88.130 103.810 88.270 105.190 ;
        RECT 91.590 104.655 93.470 105.025 ;
        RECT 88.070 103.490 88.330 103.810 ;
        RECT 86.690 102.810 86.950 103.130 ;
        RECT 87.610 102.810 87.870 103.130 ;
        RECT 73.800 88.160 74.080 88.800 ;
        RECT 79.780 88.180 80.060 88.800 ;
        RECT 85.760 88.250 86.040 88.800 ;
        RECT 86.750 88.250 86.890 102.810 ;
        RECT 91.590 99.215 93.470 99.585 ;
        RECT 91.740 88.320 92.020 88.800 ;
        RECT 73.800 86.800 75.070 88.160 ;
        RECT 73.850 84.290 75.070 86.800 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 85.760 88.110 86.890 88.250 ;
        RECT 91.460 88.250 92.680 88.320 ;
        RECT 93.650 88.250 93.790 106.890 ;
        RECT 97.790 106.870 97.930 107.910 ;
        RECT 97.730 106.550 97.990 106.870 ;
        RECT 99.110 105.870 99.370 106.190 ;
        RECT 97.270 105.190 97.530 105.510 ;
        RECT 97.330 101.430 97.470 105.190 ;
        RECT 99.170 103.810 99.310 105.870 ;
        RECT 99.110 103.490 99.370 103.810 ;
        RECT 97.270 101.110 97.530 101.430 ;
        RECT 99.170 100.750 99.310 103.490 ;
        RECT 99.630 101.430 99.770 107.910 ;
        RECT 102.390 106.530 102.530 108.250 ;
        RECT 109.230 107.910 109.490 108.230 ;
        RECT 106.590 107.375 108.470 107.745 ;
        RECT 108.770 106.890 109.030 107.210 ;
        RECT 102.330 106.210 102.590 106.530 ;
        RECT 104.170 105.190 104.430 105.510 ;
        RECT 104.230 103.130 104.370 105.190 ;
        RECT 103.710 102.810 103.970 103.130 ;
        RECT 104.170 102.810 104.430 103.130 ;
        RECT 99.570 101.110 99.830 101.430 ;
        RECT 97.730 100.430 97.990 100.750 ;
        RECT 99.110 100.430 99.370 100.750 ;
        RECT 97.790 88.800 97.930 100.430 ;
        RECT 103.770 88.800 103.910 102.810 ;
        RECT 106.590 101.935 108.470 102.305 ;
        RECT 108.830 97.770 108.970 106.890 ;
        RECT 109.290 106.870 109.430 107.910 ;
        RECT 109.230 106.550 109.490 106.870 ;
        RECT 110.670 103.810 110.810 109.270 ;
        RECT 111.130 108.910 111.270 128.230 ;
        RECT 112.050 125.140 112.190 130.350 ;
        RECT 118.030 128.290 118.170 131.030 ;
        RECT 112.910 127.970 113.170 128.290 ;
        RECT 117.970 127.970 118.230 128.290 ;
        RECT 112.050 125.000 112.650 125.140 ;
        RECT 112.510 122.850 112.650 125.000 ;
        RECT 112.970 124.550 113.110 127.970 ;
        RECT 114.750 127.630 115.010 127.950 ;
        RECT 114.810 126.250 114.950 127.630 ;
        RECT 114.750 125.930 115.010 126.250 ;
        RECT 113.370 125.250 113.630 125.570 ;
        RECT 112.910 124.230 113.170 124.550 ;
        RECT 112.970 123.190 113.110 124.230 ;
        RECT 112.910 122.870 113.170 123.190 ;
        RECT 112.450 122.530 112.710 122.850 ;
        RECT 111.530 118.790 111.790 119.110 ;
        RECT 111.590 117.410 111.730 118.790 ;
        RECT 111.530 117.090 111.790 117.410 ;
        RECT 111.590 112.650 111.730 117.090 ;
        RECT 112.510 114.690 112.650 122.530 ;
        RECT 113.430 122.510 113.570 125.250 ;
        RECT 113.370 122.420 113.630 122.510 ;
        RECT 112.970 122.280 113.630 122.420 ;
        RECT 112.970 115.030 113.110 122.280 ;
        RECT 113.370 122.190 113.630 122.280 ;
        RECT 116.130 119.470 116.390 119.790 ;
        RECT 118.030 119.700 118.170 127.970 ;
        RECT 118.430 126.950 118.690 127.270 ;
        RECT 120.270 126.950 120.530 127.270 ;
        RECT 118.490 124.890 118.630 126.950 ;
        RECT 120.330 125.570 120.470 126.950 ;
        RECT 121.590 126.415 123.470 126.785 ;
        RECT 120.270 125.250 120.530 125.570 ;
        RECT 124.470 125.230 124.610 137.830 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 124.410 124.910 124.670 125.230 ;
        RECT 118.430 124.570 118.690 124.890 ;
        RECT 118.890 122.870 119.150 123.190 ;
        RECT 118.950 120.810 119.090 122.870 ;
        RECT 124.470 122.850 124.610 124.910 ;
        RECT 124.410 122.530 124.670 122.850 ;
        RECT 121.190 122.190 121.450 122.510 ;
        RECT 120.270 121.510 120.530 121.830 ;
        RECT 118.890 120.490 119.150 120.810 ;
        RECT 120.330 119.790 120.470 121.510 ;
        RECT 121.250 120.810 121.390 122.190 ;
        RECT 121.590 120.975 123.470 121.345 ;
        RECT 121.190 120.490 121.450 120.810 ;
        RECT 118.430 119.700 118.690 119.790 ;
        RECT 118.030 119.560 118.690 119.700 ;
        RECT 113.370 119.130 113.630 119.450 ;
        RECT 113.430 118.090 113.570 119.130 ;
        RECT 116.190 118.090 116.330 119.470 ;
        RECT 113.370 117.770 113.630 118.090 ;
        RECT 116.130 117.770 116.390 118.090 ;
        RECT 118.030 117.750 118.170 119.560 ;
        RECT 118.430 119.470 118.690 119.560 ;
        RECT 120.270 119.470 120.530 119.790 ;
        RECT 117.970 117.430 118.230 117.750 ;
        RECT 115.210 117.090 115.470 117.410 ;
        RECT 115.270 115.370 115.410 117.090 ;
        RECT 121.590 115.535 123.470 115.905 ;
        RECT 115.210 115.050 115.470 115.370 ;
        RECT 112.910 114.710 113.170 115.030 ;
        RECT 112.450 114.370 112.710 114.690 ;
        RECT 121.650 113.350 121.910 113.670 ;
        RECT 111.530 112.330 111.790 112.650 ;
        RECT 117.050 112.330 117.310 112.650 ;
        RECT 111.590 109.590 111.730 112.330 ;
        RECT 111.530 109.270 111.790 109.590 ;
        RECT 111.070 108.590 111.330 108.910 ;
        RECT 111.070 107.910 111.330 108.230 ;
        RECT 111.130 106.870 111.270 107.910 ;
        RECT 111.070 106.550 111.330 106.870 ;
        RECT 111.590 106.610 111.730 109.270 ;
        RECT 113.830 107.910 114.090 108.230 ;
        RECT 116.130 107.910 116.390 108.230 ;
        RECT 111.590 106.470 112.190 106.610 ;
        RECT 112.050 106.190 112.190 106.470 ;
        RECT 111.990 105.870 112.250 106.190 ;
        RECT 112.050 103.810 112.190 105.870 ;
        RECT 113.890 103.810 114.030 107.910 ;
        RECT 110.610 103.490 110.870 103.810 ;
        RECT 111.990 103.490 112.250 103.810 ;
        RECT 113.830 103.490 114.090 103.810 ;
        RECT 115.670 103.490 115.930 103.810 ;
        RECT 108.830 97.630 109.890 97.770 ;
        RECT 109.750 89.290 109.890 97.630 ;
        RECT 115.730 89.570 115.870 103.490 ;
        RECT 116.190 103.130 116.330 107.910 ;
        RECT 117.110 106.870 117.250 112.330 ;
        RECT 118.890 111.990 119.150 112.310 ;
        RECT 118.950 109.250 119.090 111.990 ;
        RECT 121.710 111.970 121.850 113.350 ;
        RECT 119.350 111.650 119.610 111.970 ;
        RECT 121.650 111.650 121.910 111.970 ;
        RECT 118.890 108.930 119.150 109.250 ;
        RECT 118.890 108.140 119.150 108.230 ;
        RECT 119.410 108.140 119.550 111.650 ;
        RECT 119.810 111.310 120.070 111.630 ;
        RECT 119.870 108.570 120.010 111.310 ;
        RECT 121.590 110.095 123.470 110.465 ;
        RECT 119.810 108.250 120.070 108.570 ;
        RECT 127.630 108.250 127.890 108.570 ;
        RECT 118.890 108.000 119.550 108.140 ;
        RECT 118.890 107.910 119.150 108.000 ;
        RECT 117.050 106.550 117.310 106.870 ;
        RECT 116.130 102.810 116.390 103.130 ;
        RECT 119.410 101.090 119.550 108.000 ;
        RECT 119.810 106.550 120.070 106.870 ;
        RECT 119.870 101.770 120.010 106.550 ;
        RECT 120.730 105.870 120.990 106.190 ;
        RECT 119.810 101.450 120.070 101.770 ;
        RECT 119.350 100.770 119.610 101.090 ;
        RECT 120.790 98.450 120.930 105.870 ;
        RECT 125.780 105.675 126.060 106.045 ;
        RECT 121.590 104.655 123.470 105.025 ;
        RECT 125.850 103.470 125.990 105.675 ;
        RECT 125.790 103.150 126.050 103.470 ;
        RECT 121.590 99.215 123.470 99.585 ;
        RECT 120.790 98.310 121.850 98.450 ;
        RECT 121.710 89.570 121.850 98.310 ;
        RECT 91.460 88.110 93.790 88.250 ;
        RECT 97.720 88.240 98.000 88.800 ;
        RECT 103.700 88.610 103.980 88.800 ;
        RECT 85.760 87.970 86.040 88.110 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.110 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.730 88.800 116.960 89.570 ;
        RECT 115.660 86.800 116.960 88.800 ;
        RECT 115.740 85.700 116.960 86.800 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 127.690 89.380 127.830 108.250 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 16.540 210.755 18.520 211.085 ;
        RECT 46.540 210.755 48.520 211.085 ;
        RECT 76.540 210.755 78.520 211.085 ;
        RECT 106.540 210.755 108.520 211.085 ;
        RECT 31.540 208.035 33.520 208.365 ;
        RECT 61.540 208.035 63.520 208.365 ;
        RECT 91.540 208.035 93.520 208.365 ;
        RECT 121.540 208.035 123.520 208.365 ;
        RECT 16.540 205.315 18.520 205.645 ;
        RECT 46.540 205.315 48.520 205.645 ;
        RECT 76.540 205.315 78.520 205.645 ;
        RECT 106.540 205.315 108.520 205.645 ;
        RECT 31.540 202.595 33.520 202.925 ;
        RECT 61.540 202.595 63.520 202.925 ;
        RECT 91.540 202.595 93.520 202.925 ;
        RECT 121.540 202.595 123.520 202.925 ;
        RECT 16.540 199.875 18.520 200.205 ;
        RECT 46.540 199.875 48.520 200.205 ;
        RECT 76.540 199.875 78.520 200.205 ;
        RECT 106.540 199.875 108.520 200.205 ;
        RECT 31.540 197.155 33.520 197.485 ;
        RECT 61.540 197.155 63.520 197.485 ;
        RECT 91.540 197.155 93.520 197.485 ;
        RECT 121.540 197.155 123.520 197.485 ;
        RECT 16.540 194.435 18.520 194.765 ;
        RECT 46.540 194.435 48.520 194.765 ;
        RECT 76.540 194.435 78.520 194.765 ;
        RECT 106.540 194.435 108.520 194.765 ;
        RECT 31.540 191.715 33.520 192.045 ;
        RECT 61.540 191.715 63.520 192.045 ;
        RECT 91.540 191.715 93.520 192.045 ;
        RECT 121.540 191.715 123.520 192.045 ;
        RECT 16.540 188.995 18.520 189.325 ;
        RECT 46.540 188.995 48.520 189.325 ;
        RECT 76.540 188.995 78.520 189.325 ;
        RECT 106.540 188.995 108.520 189.325 ;
        RECT 44.080 187.610 44.460 187.620 ;
        RECT 55.375 187.610 55.705 187.625 ;
        RECT 44.080 187.310 55.705 187.610 ;
        RECT 44.080 187.300 44.460 187.310 ;
        RECT 55.375 187.295 55.705 187.310 ;
        RECT 94.475 187.610 94.805 187.625 ;
        RECT 98.360 187.610 98.740 187.620 ;
        RECT 94.475 187.310 98.740 187.610 ;
        RECT 94.475 187.295 94.805 187.310 ;
        RECT 98.360 187.300 98.740 187.310 ;
        RECT 31.540 186.275 33.520 186.605 ;
        RECT 61.540 186.275 63.520 186.605 ;
        RECT 91.540 186.275 93.520 186.605 ;
        RECT 121.540 186.275 123.520 186.605 ;
        RECT 16.540 183.555 18.520 183.885 ;
        RECT 46.540 183.555 48.520 183.885 ;
        RECT 76.540 183.555 78.520 183.885 ;
        RECT 106.540 183.555 108.520 183.885 ;
        RECT 31.540 180.835 33.520 181.165 ;
        RECT 61.540 180.835 63.520 181.165 ;
        RECT 91.540 180.835 93.520 181.165 ;
        RECT 121.540 180.835 123.520 181.165 ;
        RECT 40.195 179.450 40.525 179.465 ;
        RECT 41.575 179.450 41.905 179.465 ;
        RECT 67.335 179.450 67.665 179.465 ;
        RECT 40.195 179.150 67.665 179.450 ;
        RECT 40.195 179.135 40.525 179.150 ;
        RECT 41.575 179.135 41.905 179.150 ;
        RECT 67.335 179.135 67.665 179.150 ;
        RECT 78.375 179.450 78.705 179.465 ;
        RECT 84.815 179.450 85.145 179.465 ;
        RECT 78.375 179.150 85.145 179.450 ;
        RECT 78.375 179.135 78.705 179.150 ;
        RECT 84.815 179.135 85.145 179.150 ;
        RECT 16.540 178.115 18.520 178.445 ;
        RECT 46.540 178.115 48.520 178.445 ;
        RECT 76.540 178.115 78.520 178.445 ;
        RECT 106.540 178.115 108.520 178.445 ;
        RECT 65.955 177.410 66.285 177.425 ;
        RECT 70.095 177.410 70.425 177.425 ;
        RECT 72.395 177.410 72.725 177.425 ;
        RECT 65.955 177.110 72.725 177.410 ;
        RECT 65.955 177.095 66.285 177.110 ;
        RECT 70.095 177.095 70.425 177.110 ;
        RECT 72.395 177.095 72.725 177.110 ;
        RECT 71.475 176.730 71.805 176.745 ;
        RECT 77.915 176.730 78.245 176.745 ;
        RECT 71.475 176.430 78.245 176.730 ;
        RECT 71.475 176.415 71.805 176.430 ;
        RECT 77.915 176.415 78.245 176.430 ;
        RECT 31.540 175.395 33.520 175.725 ;
        RECT 61.540 175.395 63.520 175.725 ;
        RECT 91.540 175.395 93.520 175.725 ;
        RECT 121.540 175.395 123.520 175.725 ;
        RECT 39.735 174.690 40.065 174.705 ;
        RECT 65.035 174.690 65.365 174.705 ;
        RECT 39.735 174.390 65.365 174.690 ;
        RECT 39.735 174.375 40.065 174.390 ;
        RECT 65.035 174.375 65.365 174.390 ;
        RECT 54.455 174.010 54.785 174.025 ;
        RECT 62.735 174.010 63.065 174.025 ;
        RECT 54.455 173.710 63.065 174.010 ;
        RECT 54.455 173.695 54.785 173.710 ;
        RECT 62.735 173.695 63.065 173.710 ;
        RECT 16.540 172.675 18.520 173.005 ;
        RECT 46.540 172.675 48.520 173.005 ;
        RECT 76.540 172.675 78.520 173.005 ;
        RECT 106.540 172.675 108.520 173.005 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 127.595 171.290 127.925 171.305 ;
        RECT 129.030 171.290 134.930 172.500 ;
        RECT 127.595 170.990 134.930 171.290 ;
        RECT 127.595 170.975 127.925 170.990 ;
        RECT 31.540 169.955 33.520 170.285 ;
        RECT 61.540 169.955 63.520 170.285 ;
        RECT 91.540 169.955 93.520 170.285 ;
        RECT 121.540 169.955 123.520 170.285 ;
        RECT 129.030 170.130 134.930 170.990 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 43.875 169.260 44.205 169.265 ;
        RECT 43.875 169.250 44.460 169.260 ;
        RECT 43.650 168.950 44.460 169.250 ;
        RECT 43.875 168.940 44.460 168.950 ;
        RECT 43.875 168.935 44.205 168.940 ;
        RECT 16.540 167.235 18.520 167.565 ;
        RECT 46.540 167.235 48.520 167.565 ;
        RECT 76.540 167.235 78.520 167.565 ;
        RECT 106.540 167.235 108.520 167.565 ;
        RECT 31.540 164.515 33.520 164.845 ;
        RECT 61.540 164.515 63.520 164.845 ;
        RECT 91.540 164.515 93.520 164.845 ;
        RECT 121.540 164.515 123.520 164.845 ;
        RECT 94.680 163.810 95.060 163.820 ;
        RECT 98.360 163.810 98.740 163.820 ;
        RECT 100.915 163.810 101.245 163.825 ;
        RECT 94.680 163.510 101.245 163.810 ;
        RECT 94.680 163.500 95.060 163.510 ;
        RECT 98.360 163.500 98.740 163.510 ;
        RECT 100.915 163.495 101.245 163.510 ;
        RECT 16.540 161.795 18.520 162.125 ;
        RECT 46.540 161.795 48.520 162.125 ;
        RECT 76.540 161.795 78.520 162.125 ;
        RECT 106.540 161.795 108.520 162.125 ;
        RECT 31.540 159.075 33.520 159.405 ;
        RECT 61.540 159.075 63.520 159.405 ;
        RECT 91.540 159.075 93.520 159.405 ;
        RECT 121.540 159.075 123.520 159.405 ;
        RECT 79.755 159.050 80.085 159.065 ;
        RECT 81.135 159.050 81.465 159.065 ;
        RECT 79.755 158.750 81.465 159.050 ;
        RECT 79.755 158.735 80.085 158.750 ;
        RECT 81.135 158.735 81.465 158.750 ;
        RECT 67.795 158.370 68.125 158.385 ;
        RECT 71.475 158.370 71.805 158.385 ;
        RECT 84.355 158.370 84.685 158.385 ;
        RECT 67.795 158.070 84.685 158.370 ;
        RECT 67.795 158.055 68.125 158.070 ;
        RECT 71.475 158.055 71.805 158.070 ;
        RECT 84.355 158.055 84.685 158.070 ;
        RECT 16.540 156.355 18.520 156.685 ;
        RECT 46.540 156.355 48.520 156.685 ;
        RECT 76.540 156.355 78.520 156.685 ;
        RECT 106.540 156.355 108.520 156.685 ;
        RECT 72.855 156.330 73.185 156.345 ;
        RECT 75.155 156.330 75.485 156.345 ;
        RECT 72.855 156.030 75.485 156.330 ;
        RECT 72.855 156.015 73.185 156.030 ;
        RECT 75.155 156.015 75.485 156.030 ;
        RECT 41.575 155.650 41.905 155.665 ;
        RECT 42.955 155.650 43.285 155.665 ;
        RECT 94.680 155.650 95.060 155.660 ;
        RECT 41.575 155.350 43.285 155.650 ;
        RECT 41.575 155.335 41.905 155.350 ;
        RECT 42.955 155.335 43.285 155.350 ;
        RECT 70.800 155.350 95.060 155.650 ;
        RECT 44.080 154.970 44.460 154.980 ;
        RECT 65.495 154.970 65.825 154.985 ;
        RECT 70.800 154.970 71.100 155.350 ;
        RECT 94.680 155.340 95.060 155.350 ;
        RECT 44.080 154.670 71.100 154.970 ;
        RECT 74.235 154.970 74.565 154.985 ;
        RECT 112.160 154.970 112.540 154.980 ;
        RECT 74.235 154.670 112.540 154.970 ;
        RECT 44.080 154.660 44.460 154.670 ;
        RECT 65.495 154.655 65.825 154.670 ;
        RECT 74.235 154.655 74.565 154.670 ;
        RECT 112.160 154.660 112.540 154.670 ;
        RECT 31.540 153.635 33.520 153.965 ;
        RECT 61.540 153.635 63.520 153.965 ;
        RECT 91.540 153.635 93.520 153.965 ;
        RECT 121.540 153.635 123.520 153.965 ;
        RECT 44.335 152.250 44.665 152.265 ;
        RECT 67.795 152.250 68.125 152.265 ;
        RECT 44.335 151.950 68.125 152.250 ;
        RECT 44.335 151.935 44.665 151.950 ;
        RECT 67.795 151.935 68.125 151.950 ;
        RECT 16.540 150.915 18.520 151.245 ;
        RECT 46.540 150.915 48.520 151.245 ;
        RECT 76.540 150.915 78.520 151.245 ;
        RECT 106.540 150.915 108.520 151.245 ;
        RECT 87.575 150.210 87.905 150.225 ;
        RECT 99.075 150.210 99.405 150.225 ;
        RECT 107.355 150.210 107.685 150.225 ;
        RECT 87.575 149.910 107.685 150.210 ;
        RECT 87.575 149.895 87.905 149.910 ;
        RECT 99.075 149.895 99.405 149.910 ;
        RECT 107.355 149.895 107.685 149.910 ;
        RECT 31.540 148.195 33.520 148.525 ;
        RECT 61.540 148.195 63.520 148.525 ;
        RECT 91.540 148.195 93.520 148.525 ;
        RECT 121.540 148.195 123.520 148.525 ;
        RECT 16.540 145.475 18.520 145.805 ;
        RECT 46.540 145.475 48.520 145.805 ;
        RECT 76.540 145.475 78.520 145.805 ;
        RECT 106.540 145.475 108.520 145.805 ;
        RECT 31.540 142.755 33.520 143.085 ;
        RECT 61.540 142.755 63.520 143.085 ;
        RECT 91.540 142.755 93.520 143.085 ;
        RECT 121.540 142.755 123.520 143.085 ;
        RECT 16.540 140.035 18.520 140.365 ;
        RECT 46.540 140.035 48.520 140.365 ;
        RECT 76.540 140.035 78.520 140.365 ;
        RECT 106.540 140.035 108.520 140.365 ;
        RECT 132.510 138.800 135.210 140.035 ;
        RECT 112.160 138.650 112.540 138.660 ;
        RECT 131.050 138.650 135.210 138.800 ;
        RECT 112.160 138.350 135.210 138.650 ;
        RECT 112.160 138.340 112.540 138.350 ;
        RECT 131.050 138.200 135.210 138.350 ;
        RECT 132.510 138.165 135.210 138.200 ;
        RECT 31.540 137.315 33.520 137.645 ;
        RECT 61.540 137.315 63.520 137.645 ;
        RECT 91.540 137.315 93.520 137.645 ;
        RECT 121.540 137.315 123.520 137.645 ;
        RECT 16.540 134.595 18.520 134.925 ;
        RECT 46.540 134.595 48.520 134.925 ;
        RECT 76.540 134.595 78.520 134.925 ;
        RECT 106.540 134.595 108.520 134.925 ;
        RECT 99.075 133.890 99.405 133.905 ;
        RECT 107.815 133.890 108.145 133.905 ;
        RECT 99.075 133.590 108.145 133.890 ;
        RECT 99.075 133.575 99.405 133.590 ;
        RECT 107.815 133.575 108.145 133.590 ;
        RECT 31.540 131.875 33.520 132.205 ;
        RECT 61.540 131.875 63.520 132.205 ;
        RECT 91.540 131.875 93.520 132.205 ;
        RECT 121.540 131.875 123.520 132.205 ;
        RECT 44.080 131.850 44.460 131.860 ;
        RECT 48.935 131.850 49.265 131.865 ;
        RECT 44.080 131.550 49.265 131.850 ;
        RECT 44.080 131.540 44.460 131.550 ;
        RECT 48.935 131.535 49.265 131.550 ;
        RECT 16.540 129.155 18.520 129.485 ;
        RECT 46.540 129.155 48.520 129.485 ;
        RECT 76.540 129.155 78.520 129.485 ;
        RECT 106.540 129.155 108.520 129.485 ;
        RECT 94.680 129.130 95.060 129.140 ;
        RECT 95.395 129.130 95.725 129.145 ;
        RECT 94.680 128.830 95.725 129.130 ;
        RECT 94.680 128.820 95.060 128.830 ;
        RECT 95.395 128.815 95.725 128.830 ;
        RECT 31.540 126.435 33.520 126.765 ;
        RECT 61.540 126.435 63.520 126.765 ;
        RECT 91.540 126.435 93.520 126.765 ;
        RECT 121.540 126.435 123.520 126.765 ;
        RECT 16.540 123.715 18.520 124.045 ;
        RECT 46.540 123.715 48.520 124.045 ;
        RECT 76.540 123.715 78.520 124.045 ;
        RECT 106.540 123.715 108.520 124.045 ;
        RECT 31.540 120.995 33.520 121.325 ;
        RECT 61.540 120.995 63.520 121.325 ;
        RECT 91.540 120.995 93.520 121.325 ;
        RECT 121.540 120.995 123.520 121.325 ;
        RECT 16.540 118.275 18.520 118.605 ;
        RECT 46.540 118.275 48.520 118.605 ;
        RECT 76.540 118.275 78.520 118.605 ;
        RECT 106.540 118.275 108.520 118.605 ;
        RECT 31.540 115.555 33.520 115.885 ;
        RECT 61.540 115.555 63.520 115.885 ;
        RECT 91.540 115.555 93.520 115.885 ;
        RECT 121.540 115.555 123.520 115.885 ;
        RECT 16.540 112.835 18.520 113.165 ;
        RECT 46.540 112.835 48.520 113.165 ;
        RECT 76.540 112.835 78.520 113.165 ;
        RECT 106.540 112.835 108.520 113.165 ;
        RECT 92.635 112.810 92.965 112.825 ;
        RECT 94.680 112.810 95.060 112.820 ;
        RECT 92.635 112.510 95.060 112.810 ;
        RECT 92.635 112.495 92.965 112.510 ;
        RECT 94.680 112.500 95.060 112.510 ;
        RECT 31.540 110.115 33.520 110.445 ;
        RECT 61.540 110.115 63.520 110.445 ;
        RECT 91.540 110.115 93.520 110.445 ;
        RECT 121.540 110.115 123.520 110.445 ;
        RECT 16.540 107.395 18.520 107.725 ;
        RECT 46.540 107.395 48.520 107.725 ;
        RECT 76.540 107.395 78.520 107.725 ;
        RECT 106.540 107.395 108.520 107.725 ;
        RECT 125.755 106.010 126.085 106.025 ;
        RECT 129.700 106.010 133.210 106.625 ;
        RECT 125.755 105.710 133.210 106.010 ;
        RECT 125.755 105.695 126.085 105.710 ;
        RECT 129.700 105.605 133.210 105.710 ;
        RECT 131.050 105.560 133.050 105.605 ;
        RECT 31.540 104.675 33.520 105.005 ;
        RECT 61.540 104.675 63.520 105.005 ;
        RECT 91.540 104.675 93.520 105.005 ;
        RECT 121.540 104.675 123.520 105.005 ;
        RECT 16.540 101.955 18.520 102.285 ;
        RECT 46.540 101.955 48.520 102.285 ;
        RECT 76.540 101.955 78.520 102.285 ;
        RECT 106.540 101.955 108.520 102.285 ;
        RECT 31.540 99.235 33.520 99.565 ;
        RECT 61.540 99.235 63.520 99.565 ;
        RECT 91.540 99.235 93.520 99.565 ;
        RECT 121.540 99.235 123.520 99.565 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 16.530 99.160 18.530 211.160 ;
        RECT 31.530 99.160 33.530 211.160 ;
        RECT 44.105 187.295 44.435 187.625 ;
        RECT 44.120 169.265 44.420 187.295 ;
        RECT 44.105 168.935 44.435 169.265 ;
        RECT 44.120 154.985 44.420 168.935 ;
        RECT 44.105 154.655 44.435 154.985 ;
        RECT 44.120 131.865 44.420 154.655 ;
        RECT 44.105 131.535 44.435 131.865 ;
        RECT 46.530 99.160 48.530 211.160 ;
        RECT 61.530 99.160 63.530 211.160 ;
        RECT 76.530 99.160 78.530 211.160 ;
        RECT 91.530 99.160 93.530 211.160 ;
        RECT 98.385 187.295 98.715 187.625 ;
        RECT 98.400 163.825 98.700 187.295 ;
        RECT 94.705 163.495 95.035 163.825 ;
        RECT 98.385 163.495 98.715 163.825 ;
        RECT 94.720 155.665 95.020 163.495 ;
        RECT 94.705 155.335 95.035 155.665 ;
        RECT 94.720 129.145 95.020 155.335 ;
        RECT 94.705 128.815 95.035 129.145 ;
        RECT 94.720 112.825 95.020 128.815 ;
        RECT 94.705 112.495 95.035 112.825 ;
        RECT 106.530 99.160 108.530 211.160 ;
        RECT 112.185 154.655 112.515 154.985 ;
        RECT 112.200 138.665 112.500 154.655 ;
        RECT 112.185 138.335 112.515 138.665 ;
        RECT 121.530 99.720 123.530 211.160 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.530 99.160 123.830 99.720 ;
        RECT 121.810 97.750 123.830 99.160 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

