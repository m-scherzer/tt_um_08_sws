VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.795 206.170 14.965 206.360 ;
        RECT 19.395 206.170 19.565 206.360 ;
        RECT 24.915 206.170 25.085 206.360 ;
        RECT 26.755 206.170 26.925 206.360 ;
        RECT 32.275 206.170 32.445 206.360 ;
        RECT 37.795 206.170 37.965 206.360 ;
        RECT 39.635 206.170 39.805 206.360 ;
        RECT 45.155 206.170 45.325 206.360 ;
        RECT 50.675 206.170 50.845 206.360 ;
        RECT 52.515 206.170 52.685 206.360 ;
        RECT 58.035 206.170 58.205 206.360 ;
        RECT 63.555 206.170 63.725 206.360 ;
        RECT 65.395 206.170 65.565 206.360 ;
        RECT 70.915 206.170 71.085 206.360 ;
        RECT 76.435 206.170 76.605 206.360 ;
        RECT 78.275 206.170 78.445 206.360 ;
        RECT 83.795 206.170 83.965 206.360 ;
        RECT 89.315 206.170 89.485 206.360 ;
        RECT 91.155 206.170 91.325 206.360 ;
        RECT 96.675 206.170 96.845 206.360 ;
        RECT 102.195 206.170 102.365 206.360 ;
        RECT 103.170 206.220 103.290 206.330 ;
        RECT 108.635 206.170 108.805 206.360 ;
        RECT 114.155 206.170 114.325 206.360 ;
        RECT 115.535 206.170 115.705 206.360 ;
        RECT 14.655 205.360 16.025 206.170 ;
        RECT 16.035 205.360 19.705 206.170 ;
        RECT 19.715 205.360 25.225 206.170 ;
        RECT 25.245 205.300 25.675 206.085 ;
        RECT 25.695 205.360 27.065 206.170 ;
        RECT 27.075 205.360 32.585 206.170 ;
        RECT 32.595 205.360 38.105 206.170 ;
        RECT 38.125 205.300 38.555 206.085 ;
        RECT 38.575 205.360 39.945 206.170 ;
        RECT 39.955 205.360 45.465 206.170 ;
        RECT 45.475 205.360 50.985 206.170 ;
        RECT 51.005 205.300 51.435 206.085 ;
        RECT 51.455 205.360 52.825 206.170 ;
        RECT 52.835 205.360 58.345 206.170 ;
        RECT 58.355 205.360 63.865 206.170 ;
        RECT 63.885 205.300 64.315 206.085 ;
        RECT 64.335 205.360 65.705 206.170 ;
        RECT 65.715 205.360 71.225 206.170 ;
        RECT 71.235 205.360 76.745 206.170 ;
        RECT 76.765 205.300 77.195 206.085 ;
        RECT 77.215 205.360 78.585 206.170 ;
        RECT 78.595 205.360 84.105 206.170 ;
        RECT 84.115 205.360 89.625 206.170 ;
        RECT 89.645 205.300 90.075 206.085 ;
        RECT 90.095 205.360 91.465 206.170 ;
        RECT 91.475 205.360 96.985 206.170 ;
        RECT 96.995 205.360 102.505 206.170 ;
        RECT 102.525 205.300 102.955 206.085 ;
        RECT 103.435 205.360 108.945 206.170 ;
        RECT 108.955 205.360 114.465 206.170 ;
        RECT 114.475 205.360 115.845 206.170 ;
      LAYER nwell ;
        RECT 14.460 202.140 116.040 204.970 ;
      LAYER pwell ;
        RECT 14.655 200.940 16.025 201.750 ;
        RECT 16.035 200.940 21.545 201.750 ;
        RECT 21.555 200.940 27.065 201.750 ;
        RECT 27.075 200.940 32.585 201.750 ;
        RECT 32.595 200.940 38.105 201.750 ;
        RECT 38.125 201.025 38.555 201.810 ;
        RECT 38.575 200.940 44.085 201.750 ;
        RECT 44.095 200.940 49.605 201.750 ;
        RECT 49.615 200.940 55.125 201.750 ;
        RECT 55.135 200.940 60.645 201.750 ;
        RECT 60.665 200.940 62.015 201.850 ;
        RECT 62.520 201.620 63.865 201.850 ;
        RECT 62.035 200.940 63.865 201.620 ;
        RECT 63.885 201.025 64.315 201.810 ;
        RECT 64.335 200.940 65.705 201.720 ;
        RECT 66.175 200.940 68.005 201.620 ;
        RECT 68.475 200.940 70.305 201.750 ;
        RECT 70.315 201.620 71.235 201.850 ;
        RECT 74.065 201.620 74.995 201.840 ;
        RECT 70.315 200.940 79.505 201.620 ;
        RECT 80.435 200.940 84.105 201.750 ;
        RECT 84.115 200.940 89.625 201.750 ;
        RECT 89.645 201.025 90.075 201.810 ;
        RECT 90.555 200.940 92.385 201.750 ;
        RECT 92.395 200.940 97.905 201.750 ;
        RECT 97.915 200.940 103.425 201.750 ;
        RECT 103.435 200.940 108.945 201.750 ;
        RECT 108.955 200.940 114.465 201.750 ;
        RECT 114.475 200.940 115.845 201.750 ;
        RECT 14.795 200.730 14.965 200.940 ;
        RECT 19.395 200.730 19.565 200.920 ;
        RECT 21.235 200.750 21.405 200.940 ;
        RECT 24.915 200.730 25.085 200.920 ;
        RECT 25.890 200.780 26.010 200.890 ;
        RECT 26.755 200.750 26.925 200.940 ;
        RECT 28.595 200.730 28.765 200.920 ;
        RECT 32.275 200.750 32.445 200.940 ;
        RECT 34.115 200.730 34.285 200.920 ;
        RECT 37.795 200.750 37.965 200.940 ;
        RECT 39.635 200.730 39.805 200.920 ;
        RECT 43.775 200.750 43.945 200.940 ;
        RECT 45.155 200.730 45.325 200.920 ;
        RECT 49.295 200.750 49.465 200.940 ;
        RECT 50.675 200.730 50.845 200.920 ;
        RECT 52.055 200.775 52.215 200.885 ;
        RECT 54.815 200.750 54.985 200.940 ;
        RECT 57.575 200.730 57.745 200.920 ;
        RECT 58.955 200.730 59.125 200.920 ;
        RECT 60.335 200.750 60.505 200.940 ;
        RECT 60.795 200.750 60.965 200.940 ;
        RECT 62.175 200.750 62.345 200.940 ;
        RECT 65.395 200.750 65.565 200.940 ;
        RECT 65.910 200.780 66.030 200.890 ;
        RECT 67.695 200.750 67.865 200.940 ;
        RECT 68.155 200.890 68.325 200.920 ;
        RECT 68.155 200.780 68.330 200.890 ;
        RECT 68.155 200.730 68.325 200.780 ;
        RECT 69.075 200.775 69.235 200.885 ;
        RECT 69.995 200.750 70.165 200.940 ;
        RECT 72.295 200.730 72.465 200.920 ;
        RECT 72.755 200.750 72.925 200.920 ;
        RECT 72.760 200.730 72.925 200.750 ;
        RECT 75.055 200.730 75.225 200.920 ;
        RECT 76.490 200.780 76.610 200.890 ;
        RECT 79.195 200.730 79.365 200.940 ;
        RECT 80.115 200.785 80.275 200.895 ;
        RECT 80.575 200.730 80.745 200.920 ;
        RECT 81.035 200.730 81.205 200.920 ;
        RECT 83.335 200.730 83.505 200.920 ;
        RECT 83.795 200.890 83.965 200.940 ;
        RECT 83.795 200.780 83.970 200.890 ;
        RECT 83.795 200.750 83.965 200.780 ;
        RECT 85.635 200.730 85.805 200.920 ;
        RECT 89.315 200.750 89.485 200.940 ;
        RECT 90.290 200.780 90.410 200.890 ;
        RECT 91.155 200.730 91.325 200.920 ;
        RECT 92.075 200.750 92.245 200.940 ;
        RECT 96.675 200.730 96.845 200.920 ;
        RECT 97.595 200.750 97.765 200.940 ;
        RECT 102.195 200.730 102.365 200.920 ;
        RECT 103.115 200.890 103.285 200.940 ;
        RECT 103.115 200.780 103.290 200.890 ;
        RECT 103.115 200.750 103.285 200.780 ;
        RECT 108.635 200.730 108.805 200.940 ;
        RECT 114.155 200.730 114.325 200.940 ;
        RECT 115.535 200.730 115.705 200.940 ;
        RECT 14.655 199.920 16.025 200.730 ;
        RECT 16.035 199.920 19.705 200.730 ;
        RECT 19.715 199.920 25.225 200.730 ;
        RECT 25.245 199.860 25.675 200.645 ;
        RECT 26.155 199.920 28.905 200.730 ;
        RECT 28.915 199.920 34.425 200.730 ;
        RECT 34.435 199.920 39.945 200.730 ;
        RECT 39.955 199.920 45.465 200.730 ;
        RECT 45.475 199.920 50.985 200.730 ;
        RECT 51.005 199.860 51.435 200.645 ;
        RECT 52.375 199.920 57.885 200.730 ;
        RECT 57.905 199.820 59.255 200.730 ;
        RECT 59.275 200.050 68.465 200.730 ;
        RECT 59.275 199.820 60.195 200.050 ;
        RECT 63.025 199.830 63.955 200.050 ;
        RECT 69.395 199.820 72.505 200.730 ;
        RECT 72.760 200.050 74.595 200.730 ;
        RECT 73.665 199.820 74.595 200.050 ;
        RECT 74.915 199.950 76.285 200.730 ;
        RECT 76.765 199.860 77.195 200.645 ;
        RECT 77.215 200.050 79.505 200.730 ;
        RECT 77.215 199.820 78.135 200.050 ;
        RECT 79.525 199.820 80.875 200.730 ;
        RECT 80.905 199.820 82.255 200.730 ;
        RECT 82.285 199.820 83.635 200.730 ;
        RECT 84.115 199.920 85.945 200.730 ;
        RECT 85.955 199.920 91.465 200.730 ;
        RECT 91.475 199.920 96.985 200.730 ;
        RECT 96.995 199.920 102.505 200.730 ;
        RECT 102.525 199.860 102.955 200.645 ;
        RECT 103.435 199.920 108.945 200.730 ;
        RECT 108.955 199.920 114.465 200.730 ;
        RECT 114.475 199.920 115.845 200.730 ;
      LAYER nwell ;
        RECT 14.460 196.700 116.040 199.530 ;
      LAYER pwell ;
        RECT 14.655 195.500 16.025 196.310 ;
        RECT 16.035 195.500 21.545 196.310 ;
        RECT 21.555 195.500 27.065 196.310 ;
        RECT 27.075 195.500 32.585 196.310 ;
        RECT 32.595 195.500 38.105 196.310 ;
        RECT 38.125 195.585 38.555 196.370 ;
        RECT 38.575 195.500 42.245 196.310 ;
        RECT 42.255 195.500 47.765 196.310 ;
        RECT 47.775 195.500 53.285 196.310 ;
        RECT 57.805 196.180 58.735 196.400 ;
        RECT 61.455 196.180 63.665 196.410 ;
        RECT 53.295 195.500 63.665 196.180 ;
        RECT 63.885 195.585 64.315 196.370 ;
        RECT 65.265 196.180 68.265 196.410 ;
        RECT 65.265 196.090 69.845 196.180 ;
        RECT 65.255 195.730 69.845 196.090 ;
        RECT 65.255 195.540 66.185 195.730 ;
        RECT 65.265 195.500 66.185 195.540 ;
        RECT 68.275 195.500 69.845 195.730 ;
        RECT 69.855 195.500 72.145 196.410 ;
        RECT 73.075 196.180 73.995 196.410 ;
        RECT 76.825 196.180 77.755 196.400 ;
        RECT 73.075 195.500 82.265 196.180 ;
        RECT 82.275 195.500 84.105 196.310 ;
        RECT 84.115 195.500 89.625 196.310 ;
        RECT 89.645 195.585 90.075 196.370 ;
        RECT 90.095 195.500 93.765 196.310 ;
        RECT 96.430 196.180 97.350 196.410 ;
        RECT 93.885 195.500 97.350 196.180 ;
        RECT 97.455 196.180 98.375 196.410 ;
        RECT 101.205 196.180 102.135 196.400 ;
        RECT 97.455 195.500 106.645 196.180 ;
        RECT 107.115 195.500 108.945 196.310 ;
        RECT 108.955 195.500 114.465 196.310 ;
        RECT 114.475 195.500 115.845 196.310 ;
        RECT 14.795 195.290 14.965 195.500 ;
        RECT 19.395 195.290 19.565 195.480 ;
        RECT 21.235 195.310 21.405 195.500 ;
        RECT 24.915 195.290 25.085 195.480 ;
        RECT 25.890 195.340 26.010 195.450 ;
        RECT 26.755 195.310 26.925 195.500 ;
        RECT 29.515 195.290 29.685 195.480 ;
        RECT 32.275 195.310 32.445 195.500 ;
        RECT 35.035 195.290 35.205 195.480 ;
        RECT 37.795 195.310 37.965 195.500 ;
        RECT 40.555 195.290 40.725 195.480 ;
        RECT 41.015 195.290 41.185 195.480 ;
        RECT 41.935 195.310 42.105 195.500 ;
        RECT 44.750 195.340 44.870 195.450 ;
        RECT 47.455 195.290 47.625 195.500 ;
        RECT 48.835 195.290 49.005 195.480 ;
        RECT 50.215 195.290 50.385 195.480 ;
        RECT 50.730 195.340 50.850 195.450 ;
        RECT 51.650 195.340 51.770 195.450 ;
        RECT 52.975 195.310 53.145 195.500 ;
        RECT 53.435 195.310 53.605 195.500 ;
        RECT 55.275 195.290 55.445 195.480 ;
        RECT 60.795 195.290 60.965 195.480 ;
        RECT 64.010 195.290 64.180 195.480 ;
        RECT 64.475 195.290 64.645 195.480 ;
        RECT 64.935 195.345 65.095 195.455 ;
        RECT 69.075 195.290 69.245 195.480 ;
        RECT 69.535 195.290 69.705 195.500 ;
        RECT 70.000 195.310 70.170 195.500 ;
        RECT 72.755 195.345 72.915 195.455 ;
        RECT 75.055 195.290 75.225 195.480 ;
        RECT 76.440 195.290 76.610 195.480 ;
        RECT 77.410 195.340 77.530 195.450 ;
        RECT 81.955 195.310 82.125 195.500 ;
        RECT 82.875 195.290 83.045 195.480 ;
        RECT 83.335 195.290 83.505 195.480 ;
        RECT 83.795 195.310 83.965 195.500 ;
        RECT 85.635 195.290 85.805 195.480 ;
        RECT 86.095 195.290 86.265 195.480 ;
        RECT 87.475 195.290 87.645 195.480 ;
        RECT 89.315 195.310 89.485 195.500 ;
        RECT 93.455 195.310 93.625 195.500 ;
        RECT 93.915 195.310 94.085 195.500 ;
        RECT 96.730 195.340 96.850 195.450 ;
        RECT 97.135 195.290 97.305 195.480 ;
        RECT 101.920 195.290 102.090 195.480 ;
        RECT 103.115 195.290 103.285 195.480 ;
        RECT 106.335 195.310 106.505 195.500 ;
        RECT 106.795 195.450 106.965 195.480 ;
        RECT 106.795 195.340 106.970 195.450 ;
        RECT 106.795 195.290 106.965 195.340 ;
        RECT 108.175 195.290 108.345 195.480 ;
        RECT 108.635 195.310 108.805 195.500 ;
        RECT 110.475 195.290 110.645 195.480 ;
        RECT 114.155 195.290 114.325 195.500 ;
        RECT 115.535 195.290 115.705 195.500 ;
        RECT 14.655 194.480 16.025 195.290 ;
        RECT 16.035 194.480 19.705 195.290 ;
        RECT 19.715 194.480 25.225 195.290 ;
        RECT 25.245 194.420 25.675 195.205 ;
        RECT 26.155 194.480 29.825 195.290 ;
        RECT 29.835 194.480 35.345 195.290 ;
        RECT 35.355 194.480 40.865 195.290 ;
        RECT 40.985 194.610 44.450 195.290 ;
        RECT 43.530 194.380 44.450 194.610 ;
        RECT 45.015 194.480 47.765 195.290 ;
        RECT 47.785 194.380 49.135 195.290 ;
        RECT 49.155 194.510 50.525 195.290 ;
        RECT 51.005 194.420 51.435 195.205 ;
        RECT 51.915 194.480 55.585 195.290 ;
        RECT 55.595 194.480 61.105 195.290 ;
        RECT 61.405 194.380 64.325 195.290 ;
        RECT 64.335 194.610 68.005 195.290 ;
        RECT 67.075 194.380 68.005 194.610 ;
        RECT 68.015 194.480 69.385 195.290 ;
        RECT 69.505 194.610 72.970 195.290 ;
        RECT 72.050 194.380 72.970 194.610 ;
        RECT 73.075 194.610 75.365 195.290 ;
        RECT 73.075 194.380 73.995 194.610 ;
        RECT 75.375 194.380 76.725 195.290 ;
        RECT 76.765 194.420 77.195 195.205 ;
        RECT 77.675 194.480 83.185 195.290 ;
        RECT 83.195 194.510 84.565 195.290 ;
        RECT 84.575 194.480 85.945 195.290 ;
        RECT 85.965 194.380 87.315 195.290 ;
        RECT 87.335 194.610 96.525 195.290 ;
        RECT 91.845 194.390 92.775 194.610 ;
        RECT 95.605 194.380 96.525 194.610 ;
        RECT 97.005 194.380 98.355 195.290 ;
        RECT 98.605 194.610 102.505 195.290 ;
        RECT 101.575 194.380 102.505 194.610 ;
        RECT 102.525 194.420 102.955 195.205 ;
        RECT 103.085 194.610 106.550 195.290 ;
        RECT 105.630 194.380 106.550 194.610 ;
        RECT 106.665 194.380 108.015 195.290 ;
        RECT 108.035 194.510 109.405 195.290 ;
        RECT 109.415 194.480 110.785 195.290 ;
        RECT 110.795 194.480 114.465 195.290 ;
        RECT 114.475 194.480 115.845 195.290 ;
      LAYER nwell ;
        RECT 14.460 191.260 116.040 194.090 ;
      LAYER pwell ;
        RECT 14.655 190.060 16.025 190.870 ;
        RECT 16.035 190.060 17.405 190.870 ;
        RECT 17.415 190.060 21.085 190.870 ;
        RECT 21.095 190.060 26.605 190.870 ;
        RECT 29.270 190.740 30.190 190.970 ;
        RECT 26.725 190.060 30.190 190.740 ;
        RECT 30.755 190.060 32.585 190.870 ;
        RECT 32.605 190.060 33.955 190.970 ;
        RECT 37.175 190.740 38.105 190.970 ;
        RECT 34.205 190.060 38.105 190.740 ;
        RECT 38.125 190.145 38.555 190.930 ;
        RECT 38.575 190.060 39.945 190.840 ;
        RECT 40.415 190.740 41.335 190.970 ;
        RECT 44.165 190.740 45.095 190.960 ;
        RECT 49.615 190.740 50.535 190.970 ;
        RECT 53.365 190.740 54.295 190.960 ;
        RECT 40.415 190.060 49.605 190.740 ;
        RECT 49.615 190.060 58.805 190.740 ;
        RECT 58.825 190.060 60.175 190.970 ;
        RECT 62.850 190.740 63.770 190.970 ;
        RECT 60.305 190.060 63.770 190.740 ;
        RECT 63.885 190.145 64.315 190.930 ;
        RECT 64.335 190.060 66.165 190.870 ;
        RECT 66.175 190.770 67.105 190.970 ;
        RECT 68.440 190.770 69.385 190.970 ;
        RECT 66.175 190.290 69.385 190.770 ;
        RECT 69.395 190.770 70.325 190.970 ;
        RECT 71.660 190.770 72.605 190.970 ;
        RECT 69.395 190.290 72.605 190.770 ;
        RECT 66.315 190.090 69.385 190.290 ;
        RECT 14.795 189.850 14.965 190.060 ;
        RECT 17.095 189.870 17.265 190.060 ;
        RECT 19.395 189.850 19.565 190.040 ;
        RECT 20.775 189.870 20.945 190.060 ;
        RECT 24.915 189.850 25.085 190.040 ;
        RECT 26.295 189.870 26.465 190.060 ;
        RECT 26.755 189.870 26.925 190.060 ;
        RECT 27.675 189.850 27.845 190.040 ;
        RECT 28.135 189.850 28.305 190.040 ;
        RECT 30.490 189.900 30.610 190.010 ;
        RECT 32.275 189.870 32.445 190.060 ;
        RECT 32.735 189.870 32.905 190.060 ;
        RECT 37.520 189.870 37.690 190.060 ;
        RECT 38.715 189.870 38.885 190.060 ;
        RECT 40.150 189.900 40.270 190.010 ;
        RECT 41.015 189.850 41.185 190.040 ;
        RECT 42.395 189.850 42.565 190.040 ;
        RECT 46.260 189.850 46.430 190.040 ;
        RECT 49.295 189.870 49.465 190.060 ;
        RECT 50.400 189.850 50.570 190.040 ;
        RECT 52.515 189.850 52.685 190.040 ;
        RECT 53.895 189.850 54.065 190.040 ;
        RECT 54.410 189.900 54.530 190.010 ;
        RECT 54.815 189.850 54.985 190.040 ;
        RECT 56.250 189.900 56.370 190.010 ;
        RECT 58.035 189.850 58.205 190.040 ;
        RECT 58.495 189.870 58.665 190.060 ;
        RECT 58.955 189.870 59.125 190.060 ;
        RECT 60.335 189.870 60.505 190.060 ;
        RECT 65.855 189.870 66.025 190.060 ;
        RECT 66.315 189.870 66.485 190.090 ;
        RECT 68.440 190.060 69.385 190.090 ;
        RECT 69.535 190.090 72.605 190.290 ;
        RECT 67.235 189.850 67.405 190.040 ;
        RECT 69.535 189.870 69.705 190.090 ;
        RECT 71.660 190.060 72.605 190.090 ;
        RECT 72.615 190.060 74.445 190.740 ;
        RECT 74.915 190.060 77.665 190.870 ;
        RECT 78.045 190.860 78.965 190.970 ;
        RECT 78.045 190.740 80.380 190.860 ;
        RECT 85.045 190.740 85.965 190.960 ;
        RECT 78.045 190.060 87.325 190.740 ;
        RECT 88.255 190.060 89.625 190.840 ;
        RECT 89.645 190.145 90.075 190.930 ;
        RECT 90.095 190.740 91.025 190.970 ;
        RECT 90.095 190.060 93.995 190.740 ;
        RECT 94.235 190.060 96.985 190.870 ;
        RECT 96.995 190.740 97.925 190.970 ;
        RECT 101.135 190.740 102.055 190.970 ;
        RECT 104.885 190.740 105.815 190.960 ;
        RECT 96.995 190.060 100.895 190.740 ;
        RECT 101.135 190.060 110.325 190.740 ;
        RECT 110.795 190.060 114.465 190.870 ;
        RECT 114.475 190.060 115.845 190.870 ;
        RECT 70.455 189.850 70.625 190.040 ;
        RECT 70.970 189.900 71.090 190.010 ;
        RECT 72.755 189.870 72.925 190.060 ;
        RECT 74.650 189.900 74.770 190.010 ;
        RECT 76.435 189.850 76.605 190.040 ;
        RECT 77.355 189.870 77.525 190.060 ;
        RECT 78.275 189.850 78.445 190.040 ;
        RECT 82.140 189.850 82.310 190.040 ;
        RECT 83.795 189.850 83.965 190.040 ;
        RECT 85.175 189.850 85.345 190.040 ;
        RECT 87.015 189.870 87.185 190.060 ;
        RECT 87.935 189.905 88.095 190.015 ;
        RECT 88.855 189.850 89.025 190.040 ;
        RECT 89.315 189.850 89.485 190.060 ;
        RECT 90.510 189.870 90.680 190.060 ;
        RECT 93.915 189.850 94.085 190.040 ;
        RECT 94.430 189.900 94.550 190.010 ;
        RECT 94.835 189.850 95.005 190.040 ;
        RECT 96.675 189.870 96.845 190.060 ;
        RECT 97.410 189.870 97.580 190.060 ;
        RECT 99.435 189.850 99.605 190.040 ;
        RECT 99.895 189.850 100.065 190.040 ;
        RECT 101.275 189.850 101.445 190.040 ;
        RECT 106.335 189.850 106.505 190.040 ;
        RECT 106.850 189.900 106.970 190.010 ;
        RECT 108.635 189.850 108.805 190.040 ;
        RECT 110.015 189.870 110.185 190.060 ;
        RECT 110.530 189.900 110.650 190.010 ;
        RECT 114.155 189.850 114.325 190.060 ;
        RECT 115.535 189.850 115.705 190.060 ;
        RECT 14.655 189.040 16.025 189.850 ;
        RECT 16.035 189.040 19.705 189.850 ;
        RECT 19.715 189.040 25.225 189.850 ;
        RECT 25.245 188.980 25.675 189.765 ;
        RECT 26.615 189.070 27.985 189.850 ;
        RECT 28.105 189.170 31.570 189.850 ;
        RECT 30.650 188.940 31.570 189.170 ;
        RECT 32.045 189.170 41.325 189.850 ;
        RECT 32.045 189.050 34.380 189.170 ;
        RECT 32.045 188.940 32.965 189.050 ;
        RECT 39.045 188.950 39.965 189.170 ;
        RECT 41.335 189.070 42.705 189.850 ;
        RECT 42.945 189.170 46.845 189.850 ;
        RECT 47.085 189.170 50.985 189.850 ;
        RECT 45.915 188.940 46.845 189.170 ;
        RECT 50.055 188.940 50.985 189.170 ;
        RECT 51.005 188.980 51.435 189.765 ;
        RECT 51.455 189.040 52.825 189.850 ;
        RECT 52.845 188.940 54.195 189.850 ;
        RECT 54.675 189.070 56.045 189.850 ;
        RECT 56.515 189.040 58.345 189.850 ;
        RECT 58.355 189.170 67.545 189.850 ;
        RECT 58.355 188.940 59.275 189.170 ;
        RECT 62.105 188.950 63.035 189.170 ;
        RECT 67.555 188.940 70.665 189.850 ;
        RECT 71.235 189.040 76.745 189.850 ;
        RECT 76.765 188.980 77.195 189.765 ;
        RECT 77.225 188.940 78.575 189.850 ;
        RECT 78.825 189.170 82.725 189.850 ;
        RECT 81.795 188.940 82.725 189.170 ;
        RECT 82.745 188.940 84.095 189.850 ;
        RECT 84.115 189.040 85.485 189.850 ;
        RECT 85.495 189.040 89.165 189.850 ;
        RECT 89.185 188.940 90.535 189.850 ;
        RECT 90.650 189.170 94.115 189.850 ;
        RECT 90.650 188.940 91.570 189.170 ;
        RECT 94.695 189.070 96.065 189.850 ;
        RECT 96.170 189.170 99.635 189.850 ;
        RECT 96.170 188.940 97.090 189.170 ;
        RECT 99.765 188.940 101.115 189.850 ;
        RECT 101.145 188.940 102.495 189.850 ;
        RECT 102.525 188.980 102.955 189.765 ;
        RECT 103.070 189.170 106.535 189.850 ;
        RECT 103.070 188.940 103.990 189.170 ;
        RECT 107.115 189.040 108.945 189.850 ;
        RECT 108.955 189.040 114.465 189.850 ;
        RECT 114.475 189.040 115.845 189.850 ;
      LAYER nwell ;
        RECT 14.460 185.820 116.040 188.650 ;
      LAYER pwell ;
        RECT 14.655 184.620 16.025 185.430 ;
        RECT 16.495 184.620 19.245 185.430 ;
        RECT 19.265 184.620 20.615 185.530 ;
        RECT 23.290 185.300 24.210 185.530 ;
        RECT 28.825 185.300 29.755 185.520 ;
        RECT 32.585 185.300 33.505 185.530 ;
        RECT 20.745 184.620 24.210 185.300 ;
        RECT 24.315 184.620 33.505 185.300 ;
        RECT 34.630 184.620 38.105 185.530 ;
        RECT 38.125 184.705 38.555 185.490 ;
        RECT 39.035 185.300 39.965 185.530 ;
        RECT 43.175 185.300 44.095 185.530 ;
        RECT 46.925 185.300 47.855 185.520 ;
        RECT 39.035 184.620 42.935 185.300 ;
        RECT 43.175 184.620 52.365 185.300 ;
        RECT 52.835 184.620 58.345 185.430 ;
        RECT 58.355 184.620 63.865 185.430 ;
        RECT 63.885 184.705 64.315 185.490 ;
        RECT 64.335 184.620 69.845 185.430 ;
        RECT 69.855 184.620 75.365 185.430 ;
        RECT 75.745 185.420 76.665 185.530 ;
        RECT 75.745 185.300 78.080 185.420 ;
        RECT 82.745 185.300 83.665 185.520 ;
        RECT 75.745 184.620 85.025 185.300 ;
        RECT 85.035 184.620 86.405 185.400 ;
        RECT 86.415 184.620 87.785 185.430 ;
        RECT 87.805 184.620 89.155 185.530 ;
        RECT 89.645 184.705 90.075 185.490 ;
        RECT 90.095 185.300 91.015 185.530 ;
        RECT 93.845 185.300 94.775 185.520 ;
        RECT 99.390 185.300 100.310 185.530 ;
        RECT 103.895 185.300 104.815 185.530 ;
        RECT 107.645 185.300 108.575 185.520 ;
        RECT 90.095 184.620 99.285 185.300 ;
        RECT 99.390 184.620 102.855 185.300 ;
        RECT 103.895 184.620 113.085 185.300 ;
        RECT 113.095 184.620 114.465 185.430 ;
        RECT 114.475 184.620 115.845 185.430 ;
        RECT 14.795 184.410 14.965 184.620 ;
        RECT 16.230 184.460 16.350 184.570 ;
        RECT 17.555 184.410 17.725 184.600 ;
        RECT 18.015 184.410 18.185 184.600 ;
        RECT 18.935 184.430 19.105 184.620 ;
        RECT 19.395 184.430 19.565 184.620 ;
        RECT 20.775 184.430 20.945 184.620 ;
        RECT 21.695 184.410 21.865 184.600 ;
        RECT 24.455 184.430 24.625 184.620 ;
        RECT 26.755 184.410 26.925 184.600 ;
        RECT 28.135 184.410 28.305 184.600 ;
        RECT 28.870 184.410 29.040 184.600 ;
        RECT 33.195 184.455 33.355 184.565 ;
        RECT 34.115 184.465 34.275 184.575 ;
        RECT 37.790 184.430 37.960 184.620 ;
        RECT 38.770 184.460 38.890 184.570 ;
        RECT 39.450 184.430 39.620 184.620 ;
        RECT 42.395 184.410 42.565 184.600 ;
        RECT 42.910 184.460 43.030 184.570 ;
        RECT 44.235 184.410 44.405 184.600 ;
        RECT 44.695 184.410 44.865 184.600 ;
        RECT 46.075 184.410 46.245 184.600 ;
        RECT 49.755 184.410 49.925 184.600 ;
        RECT 52.055 184.430 52.225 184.620 ;
        RECT 52.570 184.460 52.690 184.570 ;
        RECT 54.815 184.410 54.985 184.600 ;
        RECT 58.035 184.430 58.205 184.620 ;
        RECT 60.335 184.410 60.505 184.600 ;
        RECT 63.555 184.430 63.725 184.620 ;
        RECT 65.855 184.410 66.025 184.600 ;
        RECT 66.315 184.430 66.485 184.600 ;
        RECT 69.535 184.570 69.705 184.620 ;
        RECT 69.535 184.460 69.710 184.570 ;
        RECT 69.535 184.430 69.705 184.460 ;
        RECT 66.415 184.410 66.485 184.430 ;
        RECT 72.295 184.410 72.465 184.600 ;
        RECT 75.055 184.430 75.225 184.620 ;
        RECT 76.160 184.410 76.330 184.600 ;
        RECT 78.275 184.410 78.445 184.600 ;
        RECT 82.140 184.410 82.310 184.600 ;
        RECT 82.875 184.410 83.045 184.600 ;
        RECT 84.715 184.430 84.885 184.620 ;
        RECT 85.175 184.410 85.345 184.600 ;
        RECT 86.095 184.430 86.265 184.620 ;
        RECT 87.475 184.430 87.645 184.620 ;
        RECT 87.935 184.430 88.105 184.620 ;
        RECT 89.370 184.460 89.490 184.570 ;
        RECT 97.780 184.410 97.950 184.600 ;
        RECT 98.975 184.430 99.145 184.620 ;
        RECT 101.920 184.410 102.090 184.600 ;
        RECT 102.655 184.430 102.825 184.620 ;
        RECT 103.575 184.465 103.735 184.575 ;
        RECT 111.855 184.410 112.025 184.600 ;
        RECT 112.370 184.460 112.490 184.570 ;
        RECT 112.775 184.430 112.945 184.620 ;
        RECT 114.155 184.410 114.325 184.620 ;
        RECT 115.535 184.410 115.705 184.620 ;
        RECT 14.655 183.600 16.025 184.410 ;
        RECT 16.035 183.600 17.865 184.410 ;
        RECT 17.985 183.730 21.450 184.410 ;
        RECT 21.665 183.730 25.130 184.410 ;
        RECT 20.530 183.500 21.450 183.730 ;
        RECT 24.210 183.500 25.130 183.730 ;
        RECT 25.245 183.540 25.675 184.325 ;
        RECT 25.705 183.500 27.055 184.410 ;
        RECT 27.075 183.600 28.445 184.410 ;
        RECT 28.455 183.730 32.355 184.410 ;
        RECT 33.515 183.730 42.705 184.410 ;
        RECT 28.455 183.500 29.385 183.730 ;
        RECT 33.515 183.500 34.435 183.730 ;
        RECT 37.265 183.510 38.195 183.730 ;
        RECT 43.185 183.500 44.535 184.410 ;
        RECT 44.555 183.630 45.925 184.410 ;
        RECT 46.045 183.730 49.510 184.410 ;
        RECT 48.590 183.500 49.510 183.730 ;
        RECT 49.625 183.500 50.975 184.410 ;
        RECT 51.005 183.540 51.435 184.325 ;
        RECT 51.550 183.730 55.015 184.410 ;
        RECT 51.550 183.500 52.470 183.730 ;
        RECT 55.135 183.600 60.645 184.410 ;
        RECT 60.655 183.600 66.165 184.410 ;
        RECT 66.415 184.180 68.685 184.410 ;
        RECT 66.415 183.500 69.170 184.180 ;
        RECT 69.855 183.600 72.605 184.410 ;
        RECT 72.845 183.730 76.745 184.410 ;
        RECT 75.815 183.500 76.745 183.730 ;
        RECT 76.765 183.540 77.195 184.325 ;
        RECT 77.225 183.500 78.575 184.410 ;
        RECT 78.825 183.730 82.725 184.410 ;
        RECT 81.795 183.500 82.725 183.730 ;
        RECT 82.735 183.630 84.105 184.410 ;
        RECT 85.035 183.730 94.225 184.410 ;
        RECT 94.465 183.730 98.365 184.410 ;
        RECT 98.605 183.730 102.505 184.410 ;
        RECT 89.545 183.510 90.475 183.730 ;
        RECT 93.305 183.500 94.225 183.730 ;
        RECT 97.435 183.500 98.365 183.730 ;
        RECT 101.575 183.500 102.505 183.730 ;
        RECT 102.525 183.540 102.955 184.325 ;
        RECT 102.975 183.730 112.165 184.410 ;
        RECT 102.975 183.500 103.895 183.730 ;
        RECT 106.725 183.510 107.655 183.730 ;
        RECT 112.635 183.600 114.465 184.410 ;
        RECT 114.475 183.600 115.845 184.410 ;
      LAYER nwell ;
        RECT 14.460 180.380 116.040 183.210 ;
      LAYER pwell ;
        RECT 14.655 179.180 16.025 179.990 ;
        RECT 16.495 179.180 18.325 179.990 ;
        RECT 20.990 179.860 21.910 180.090 ;
        RECT 18.445 179.180 21.910 179.860 ;
        RECT 22.015 179.860 22.935 180.090 ;
        RECT 25.765 179.860 26.695 180.080 ;
        RECT 22.015 179.180 31.205 179.860 ;
        RECT 31.215 179.180 33.045 179.990 ;
        RECT 33.065 179.180 34.415 180.090 ;
        RECT 37.090 179.860 38.010 180.090 ;
        RECT 34.545 179.180 38.010 179.860 ;
        RECT 38.125 179.265 38.555 180.050 ;
        RECT 39.495 179.180 42.970 180.090 ;
        RECT 46.375 179.860 47.305 180.090 ;
        RECT 43.405 179.180 47.305 179.860 ;
        RECT 47.315 179.860 48.235 180.090 ;
        RECT 51.065 179.860 51.995 180.080 ;
        RECT 47.315 179.180 56.505 179.860 ;
        RECT 56.515 179.180 57.885 179.990 ;
        RECT 57.895 179.180 60.505 180.090 ;
        RECT 60.895 179.410 63.650 180.090 ;
        RECT 60.895 179.180 63.165 179.410 ;
        RECT 63.885 179.265 64.315 180.050 ;
        RECT 64.335 179.180 65.705 179.990 ;
        RECT 67.295 179.860 70.295 180.090 ;
        RECT 73.170 179.860 74.090 180.090 ;
        RECT 76.755 179.860 77.675 180.090 ;
        RECT 80.505 179.860 81.435 180.080 ;
        RECT 88.610 179.860 89.530 180.090 ;
        RECT 65.715 179.770 70.295 179.860 ;
        RECT 65.715 179.410 70.305 179.770 ;
        RECT 65.715 179.180 67.285 179.410 ;
        RECT 69.375 179.220 70.305 179.410 ;
        RECT 69.375 179.180 70.295 179.220 ;
        RECT 70.315 179.180 73.055 179.860 ;
        RECT 73.170 179.180 76.635 179.860 ;
        RECT 76.755 179.180 85.945 179.860 ;
        RECT 86.065 179.180 89.530 179.860 ;
        RECT 89.645 179.265 90.075 180.050 ;
        RECT 90.095 179.860 91.025 180.090 ;
        RECT 90.095 179.180 93.995 179.860 ;
        RECT 95.155 179.180 98.630 180.090 ;
        RECT 98.835 179.180 100.205 179.960 ;
        RECT 100.215 179.180 102.045 179.990 ;
        RECT 105.255 179.860 106.185 180.090 ;
        RECT 102.285 179.180 106.185 179.860 ;
        RECT 106.390 179.180 109.865 180.090 ;
        RECT 109.875 179.180 111.245 179.960 ;
        RECT 111.255 179.180 112.625 179.960 ;
        RECT 112.635 179.180 114.465 179.990 ;
        RECT 114.475 179.180 115.845 179.990 ;
        RECT 14.795 178.970 14.965 179.180 ;
        RECT 16.230 179.020 16.350 179.130 ;
        RECT 18.015 178.990 18.185 179.180 ;
        RECT 18.475 178.990 18.645 179.180 ;
        RECT 21.235 178.970 21.405 179.160 ;
        RECT 21.695 178.970 21.865 179.160 ;
        RECT 25.835 178.970 26.005 179.160 ;
        RECT 27.215 178.970 27.385 179.160 ;
        RECT 28.870 178.970 29.040 179.160 ;
        RECT 30.895 178.990 31.065 179.180 ;
        RECT 32.735 179.130 32.905 179.180 ;
        RECT 32.735 179.020 32.910 179.130 ;
        RECT 32.735 178.990 32.905 179.020 ;
        RECT 33.195 178.990 33.365 179.180 ;
        RECT 34.575 178.990 34.745 179.180 ;
        RECT 36.600 178.970 36.770 179.160 ;
        RECT 37.390 179.020 37.510 179.130 ;
        RECT 39.175 179.025 39.335 179.135 ;
        RECT 39.640 178.990 39.810 179.180 ;
        RECT 40.095 178.970 40.265 179.160 ;
        RECT 40.560 178.970 40.730 179.160 ;
        RECT 46.535 178.970 46.705 179.160 ;
        RECT 46.720 178.990 46.890 179.180 ;
        RECT 50.400 178.970 50.570 179.160 ;
        RECT 51.595 178.970 51.765 179.160 ;
        RECT 56.195 178.990 56.365 179.180 ;
        RECT 57.575 178.970 57.745 179.180 ;
        RECT 58.040 178.990 58.210 179.180 ;
        RECT 60.895 179.160 60.965 179.180 ;
        RECT 58.955 178.970 59.125 179.160 ;
        RECT 59.470 179.020 59.590 179.130 ;
        RECT 60.795 178.990 60.965 179.160 ;
        RECT 62.175 178.970 62.345 179.160 ;
        RECT 62.635 178.970 62.805 179.160 ;
        RECT 65.395 178.970 65.565 179.180 ;
        RECT 65.855 178.990 66.025 179.180 ;
        RECT 69.535 179.015 69.695 179.125 ;
        RECT 69.995 178.990 70.165 179.160 ;
        RECT 70.455 178.990 70.625 179.180 ;
        RECT 65.955 178.970 66.025 178.990 ;
        RECT 70.095 178.970 70.165 178.990 ;
        RECT 73.220 178.970 73.390 179.160 ;
        RECT 76.435 178.990 76.605 179.180 ;
        RECT 78.735 178.970 78.905 179.160 ;
        RECT 79.195 178.970 79.365 179.160 ;
        RECT 82.880 178.970 83.050 179.160 ;
        RECT 85.635 178.970 85.805 179.180 ;
        RECT 86.095 178.990 86.265 179.180 ;
        RECT 90.235 178.970 90.405 179.160 ;
        RECT 90.510 178.990 90.680 179.180 ;
        RECT 90.700 178.970 90.870 179.160 ;
        RECT 94.380 178.970 94.550 179.160 ;
        RECT 94.835 179.025 94.995 179.135 ;
        RECT 95.300 178.990 95.470 179.180 ;
        RECT 98.515 179.015 98.675 179.125 ;
        RECT 99.895 178.990 100.065 179.180 ;
        RECT 101.735 178.990 101.905 179.180 ;
        RECT 102.190 178.970 102.360 179.160 ;
        RECT 103.575 179.015 103.735 179.125 ;
        RECT 104.035 178.970 104.205 179.160 ;
        RECT 105.600 178.990 105.770 179.180 ;
        RECT 108.635 178.970 108.805 179.160 ;
        RECT 109.095 178.970 109.265 179.160 ;
        RECT 109.550 178.990 109.720 179.180 ;
        RECT 110.015 178.990 110.185 179.180 ;
        RECT 110.530 179.020 110.650 179.130 ;
        RECT 112.315 178.990 112.485 179.180 ;
        RECT 114.155 178.970 114.325 179.180 ;
        RECT 115.535 178.970 115.705 179.180 ;
        RECT 14.655 178.160 16.025 178.970 ;
        RECT 16.035 178.160 21.545 178.970 ;
        RECT 21.665 178.290 25.130 178.970 ;
        RECT 24.210 178.060 25.130 178.290 ;
        RECT 25.245 178.100 25.675 178.885 ;
        RECT 25.695 178.190 27.065 178.970 ;
        RECT 27.085 178.060 28.435 178.970 ;
        RECT 28.455 178.290 32.355 178.970 ;
        RECT 33.285 178.290 37.185 178.970 ;
        RECT 28.455 178.060 29.385 178.290 ;
        RECT 36.255 178.060 37.185 178.290 ;
        RECT 37.655 178.160 40.405 178.970 ;
        RECT 40.415 178.060 43.890 178.970 ;
        RECT 44.095 178.160 46.845 178.970 ;
        RECT 47.085 178.290 50.985 178.970 ;
        RECT 50.055 178.060 50.985 178.290 ;
        RECT 51.005 178.100 51.435 178.885 ;
        RECT 51.565 178.290 55.030 178.970 ;
        RECT 55.145 178.290 57.885 178.970 ;
        RECT 54.110 178.060 55.030 178.290 ;
        RECT 57.895 178.190 59.265 178.970 ;
        RECT 59.735 178.160 62.485 178.970 ;
        RECT 62.505 178.060 63.855 178.970 ;
        RECT 63.875 178.290 65.705 178.970 ;
        RECT 65.955 178.740 68.225 178.970 ;
        RECT 70.095 178.740 72.365 178.970 ;
        RECT 63.875 178.060 65.220 178.290 ;
        RECT 65.955 178.060 68.710 178.740 ;
        RECT 70.095 178.060 72.850 178.740 ;
        RECT 73.075 178.060 76.550 178.970 ;
        RECT 76.765 178.100 77.195 178.885 ;
        RECT 77.215 178.160 79.045 178.970 ;
        RECT 79.165 178.290 82.630 178.970 ;
        RECT 81.710 178.060 82.630 178.290 ;
        RECT 82.735 178.060 85.345 178.970 ;
        RECT 85.495 178.190 86.865 178.970 ;
        RECT 86.970 178.290 90.435 178.970 ;
        RECT 86.970 178.060 87.890 178.290 ;
        RECT 90.555 178.060 94.030 178.970 ;
        RECT 94.235 178.060 97.710 178.970 ;
        RECT 99.030 178.060 102.505 178.970 ;
        RECT 102.525 178.100 102.955 178.885 ;
        RECT 104.005 178.290 107.470 178.970 ;
        RECT 106.550 178.060 107.470 178.290 ;
        RECT 107.575 178.160 108.945 178.970 ;
        RECT 108.955 178.190 110.325 178.970 ;
        RECT 110.795 178.160 114.465 178.970 ;
        RECT 114.475 178.160 115.845 178.970 ;
      LAYER nwell ;
        RECT 14.460 174.940 116.040 177.770 ;
      LAYER pwell ;
        RECT 14.655 173.740 16.025 174.550 ;
        RECT 16.955 173.740 20.625 174.550 ;
        RECT 20.830 173.740 24.305 174.650 ;
        RECT 26.970 174.420 27.890 174.650 ;
        RECT 24.425 173.740 27.890 174.420 ;
        RECT 27.995 174.420 28.915 174.650 ;
        RECT 31.745 174.420 32.675 174.640 ;
        RECT 27.995 173.740 37.185 174.420 ;
        RECT 38.125 173.825 38.555 174.610 ;
        RECT 38.575 173.740 39.945 174.520 ;
        RECT 40.610 173.740 44.085 174.650 ;
        RECT 46.750 174.420 47.670 174.650 ;
        RECT 50.975 174.420 51.905 174.650 ;
        RECT 44.205 173.740 47.670 174.420 ;
        RECT 48.005 173.740 51.905 174.420 ;
        RECT 51.915 174.420 52.835 174.650 ;
        RECT 55.665 174.420 56.595 174.640 ;
        RECT 62.035 174.420 63.380 174.650 ;
        RECT 51.915 173.740 61.105 174.420 ;
        RECT 62.035 173.740 63.865 174.420 ;
        RECT 63.885 173.825 64.315 174.610 ;
        RECT 64.795 174.420 66.140 174.650 ;
        RECT 64.795 173.740 66.625 174.420 ;
        RECT 66.635 173.740 69.355 174.650 ;
        RECT 69.395 173.740 72.870 174.650 ;
        RECT 73.075 173.740 76.550 174.650 ;
        RECT 76.755 173.740 80.230 174.650 ;
        RECT 80.435 173.740 82.265 174.550 ;
        RECT 82.275 173.740 87.785 174.550 ;
        RECT 87.805 173.740 89.155 174.650 ;
        RECT 89.645 173.825 90.075 174.610 ;
        RECT 93.210 174.420 94.130 174.650 ;
        RECT 90.665 173.740 94.130 174.420 ;
        RECT 94.235 173.740 95.605 174.550 ;
        RECT 95.625 173.740 96.975 174.650 ;
        RECT 97.190 173.740 100.665 174.650 ;
        RECT 103.330 174.420 104.250 174.650 ;
        RECT 100.785 173.740 104.250 174.420 ;
        RECT 104.355 174.420 105.275 174.650 ;
        RECT 108.105 174.420 109.035 174.640 ;
        RECT 104.355 173.740 113.545 174.420 ;
        RECT 114.475 173.740 115.845 174.550 ;
        RECT 14.795 173.530 14.965 173.740 ;
        RECT 16.230 173.580 16.350 173.690 ;
        RECT 16.635 173.585 16.795 173.695 ;
        RECT 19.855 173.530 20.025 173.720 ;
        RECT 20.315 173.550 20.485 173.740 ;
        RECT 23.535 173.530 23.705 173.720 ;
        RECT 23.990 173.550 24.160 173.740 ;
        RECT 24.455 173.550 24.625 173.740 ;
        RECT 24.915 173.530 25.085 173.720 ;
        RECT 26.755 173.530 26.925 173.720 ;
        RECT 30.430 173.530 30.600 173.720 ;
        RECT 34.110 173.530 34.280 173.720 ;
        RECT 36.875 173.550 37.045 173.740 ;
        RECT 37.790 173.530 37.960 173.720 ;
        RECT 38.255 173.530 38.425 173.720 ;
        RECT 39.635 173.550 39.805 173.740 ;
        RECT 43.770 173.720 43.940 173.740 ;
        RECT 40.150 173.580 40.270 173.690 ;
        RECT 43.315 173.530 43.485 173.720 ;
        RECT 43.770 173.550 43.950 173.720 ;
        RECT 44.235 173.550 44.405 173.740 ;
        RECT 43.780 173.530 43.950 173.550 ;
        RECT 47.460 173.530 47.630 173.720 ;
        RECT 51.320 173.550 51.490 173.740 ;
        RECT 54.815 173.530 54.985 173.720 ;
        RECT 56.195 173.530 56.365 173.720 ;
        RECT 56.710 173.580 56.830 173.690 ;
        RECT 57.115 173.530 57.285 173.720 ;
        RECT 58.550 173.580 58.670 173.690 ;
        RECT 60.795 173.550 60.965 173.740 ;
        RECT 61.715 173.585 61.875 173.695 ;
        RECT 62.175 173.530 62.345 173.720 ;
        RECT 63.555 173.550 63.725 173.740 ;
        RECT 64.015 173.530 64.185 173.720 ;
        RECT 64.475 173.690 64.645 173.720 ;
        RECT 64.475 173.580 64.650 173.690 ;
        RECT 64.475 173.530 64.645 173.580 ;
        RECT 66.315 173.550 66.485 173.740 ;
        RECT 66.775 173.550 66.945 173.740 ;
        RECT 67.235 173.530 67.405 173.720 ;
        RECT 69.540 173.550 69.710 173.740 ;
        RECT 70.915 173.530 71.085 173.720 ;
        RECT 73.220 173.550 73.390 173.740 ;
        RECT 76.435 173.530 76.605 173.720 ;
        RECT 76.900 173.550 77.070 173.740 ;
        RECT 81.955 173.550 82.125 173.740 ;
        RECT 86.555 173.530 86.725 173.720 ;
        RECT 87.015 173.530 87.185 173.720 ;
        RECT 87.475 173.550 87.645 173.740 ;
        RECT 87.935 173.550 88.105 173.740 ;
        RECT 89.370 173.580 89.490 173.690 ;
        RECT 90.290 173.580 90.410 173.690 ;
        RECT 90.695 173.550 90.865 173.740 ;
        RECT 95.295 173.550 95.465 173.740 ;
        RECT 95.755 173.550 95.925 173.740 ;
        RECT 96.675 173.575 96.835 173.685 ;
        RECT 97.135 173.530 97.305 173.720 ;
        RECT 100.350 173.550 100.520 173.740 ;
        RECT 100.815 173.550 100.985 173.740 ;
        RECT 101.920 173.530 102.090 173.720 ;
        RECT 103.115 173.530 103.285 173.720 ;
        RECT 113.235 173.530 113.405 173.740 ;
        RECT 114.155 173.575 114.315 173.695 ;
        RECT 115.535 173.530 115.705 173.740 ;
        RECT 14.655 172.720 16.025 173.530 ;
        RECT 16.495 172.720 20.165 173.530 ;
        RECT 20.270 172.850 23.735 173.530 ;
        RECT 20.270 172.620 21.190 172.850 ;
        RECT 23.855 172.720 25.225 173.530 ;
        RECT 25.245 172.660 25.675 173.445 ;
        RECT 25.705 172.620 27.055 173.530 ;
        RECT 27.270 172.620 30.745 173.530 ;
        RECT 30.950 172.620 34.425 173.530 ;
        RECT 34.630 172.620 38.105 173.530 ;
        RECT 38.225 172.850 41.690 173.530 ;
        RECT 40.770 172.620 41.690 172.850 ;
        RECT 41.795 172.720 43.625 173.530 ;
        RECT 43.635 172.620 47.110 173.530 ;
        RECT 47.315 172.620 50.790 173.530 ;
        RECT 51.005 172.660 51.435 173.445 ;
        RECT 51.455 172.720 55.125 173.530 ;
        RECT 55.145 172.620 56.495 173.530 ;
        RECT 56.975 172.750 58.345 173.530 ;
        RECT 58.815 172.720 62.485 173.530 ;
        RECT 62.495 172.850 64.325 173.530 ;
        RECT 64.335 172.850 66.165 173.530 ;
        RECT 62.495 172.620 63.840 172.850 ;
        RECT 64.820 172.620 66.165 172.850 ;
        RECT 66.175 172.720 67.545 173.530 ;
        RECT 67.555 172.720 71.225 173.530 ;
        RECT 71.235 172.720 76.745 173.530 ;
        RECT 76.765 172.660 77.195 173.445 ;
        RECT 77.585 172.850 86.865 173.530 ;
        RECT 86.875 172.850 96.065 173.530 ;
        RECT 77.585 172.730 79.920 172.850 ;
        RECT 77.585 172.620 78.505 172.730 ;
        RECT 84.585 172.630 85.505 172.850 ;
        RECT 91.385 172.630 92.315 172.850 ;
        RECT 95.145 172.620 96.065 172.850 ;
        RECT 97.005 172.620 98.355 173.530 ;
        RECT 98.605 172.850 102.505 173.530 ;
        RECT 101.575 172.620 102.505 172.850 ;
        RECT 102.525 172.660 102.955 173.445 ;
        RECT 102.985 172.620 104.335 173.530 ;
        RECT 104.355 172.850 113.545 173.530 ;
        RECT 104.355 172.620 105.275 172.850 ;
        RECT 108.105 172.630 109.035 172.850 ;
        RECT 114.475 172.720 115.845 173.530 ;
      LAYER nwell ;
        RECT 14.460 169.500 116.040 172.330 ;
      LAYER pwell ;
        RECT 14.655 168.300 16.025 169.110 ;
        RECT 16.505 168.300 17.855 169.210 ;
        RECT 17.875 168.300 19.245 169.080 ;
        RECT 21.910 168.980 22.830 169.210 ;
        RECT 19.365 168.300 22.830 168.980 ;
        RECT 22.935 168.980 23.855 169.210 ;
        RECT 26.685 168.980 27.615 169.200 ;
        RECT 22.935 168.300 32.125 168.980 ;
        RECT 33.065 168.300 34.415 169.210 ;
        RECT 37.090 168.980 38.010 169.210 ;
        RECT 34.545 168.300 38.010 168.980 ;
        RECT 38.125 168.385 38.555 169.170 ;
        RECT 39.035 168.300 41.785 169.110 ;
        RECT 41.795 168.980 42.715 169.210 ;
        RECT 45.545 168.980 46.475 169.200 ;
        RECT 41.795 168.300 50.985 168.980 ;
        RECT 51.005 168.300 52.355 169.210 ;
        RECT 52.385 168.300 53.735 169.210 ;
        RECT 53.895 168.300 56.505 169.210 ;
        RECT 56.515 168.300 58.345 169.110 ;
        RECT 58.355 168.300 63.865 169.110 ;
        RECT 63.885 168.385 64.315 169.170 ;
        RECT 64.335 168.980 65.680 169.210 ;
        RECT 64.335 168.300 66.165 168.980 ;
        RECT 66.175 168.300 68.915 168.980 ;
        RECT 69.395 168.300 72.145 169.110 ;
        RECT 72.525 169.100 73.445 169.210 ;
        RECT 72.525 168.980 74.860 169.100 ;
        RECT 79.525 168.980 80.445 169.200 ;
        RECT 72.525 168.300 81.805 168.980 ;
        RECT 81.815 168.300 83.185 169.080 ;
        RECT 83.430 168.300 88.245 168.980 ;
        RECT 88.255 168.300 89.625 169.080 ;
        RECT 89.645 168.385 90.075 169.170 ;
        RECT 90.095 168.980 91.025 169.210 ;
        RECT 94.235 168.980 95.165 169.210 ;
        RECT 101.575 168.980 102.505 169.210 ;
        RECT 106.635 168.980 107.565 169.210 ;
        RECT 110.230 168.980 111.150 169.210 ;
        RECT 90.095 168.300 93.995 168.980 ;
        RECT 94.235 168.300 98.135 168.980 ;
        RECT 98.605 168.300 102.505 168.980 ;
        RECT 103.665 168.300 107.565 168.980 ;
        RECT 107.685 168.300 111.150 168.980 ;
        RECT 111.255 168.300 113.085 168.980 ;
        RECT 113.095 168.300 114.465 169.080 ;
        RECT 114.475 168.300 115.845 169.110 ;
        RECT 14.795 168.090 14.965 168.300 ;
        RECT 16.175 168.250 16.345 168.280 ;
        RECT 16.175 168.140 16.350 168.250 ;
        RECT 16.175 168.090 16.345 168.140 ;
        RECT 17.555 168.110 17.725 168.300 ;
        RECT 18.935 168.110 19.105 168.300 ;
        RECT 19.395 168.110 19.565 168.300 ;
        RECT 26.110 168.090 26.280 168.280 ;
        RECT 30.895 168.090 31.065 168.280 ;
        RECT 31.410 168.140 31.530 168.250 ;
        RECT 31.815 168.110 31.985 168.300 ;
        RECT 32.735 168.145 32.895 168.255 ;
        RECT 33.195 168.110 33.365 168.300 ;
        RECT 34.575 168.110 34.745 168.300 ;
        RECT 38.770 168.140 38.890 168.250 ;
        RECT 40.555 168.090 40.725 168.280 ;
        RECT 41.015 168.090 41.185 168.280 ;
        RECT 41.475 168.110 41.645 168.300 ;
        RECT 50.675 168.110 50.845 168.300 ;
        RECT 52.055 168.110 52.225 168.300 ;
        RECT 52.515 168.110 52.685 168.300 ;
        RECT 56.190 168.110 56.360 168.300 ;
        RECT 58.035 168.110 58.205 168.300 ;
        RECT 60.335 168.090 60.505 168.280 ;
        RECT 63.095 168.090 63.265 168.280 ;
        RECT 63.555 168.110 63.725 168.300 ;
        RECT 65.855 168.090 66.025 168.300 ;
        RECT 66.315 168.090 66.485 168.300 ;
        RECT 69.130 168.140 69.250 168.250 ;
        RECT 70.915 168.090 71.085 168.280 ;
        RECT 71.835 168.110 72.005 168.300 ;
        RECT 72.295 168.090 72.465 168.280 ;
        RECT 76.160 168.090 76.330 168.280 ;
        RECT 78.275 168.090 78.445 168.280 ;
        RECT 78.790 168.140 78.910 168.250 ;
        RECT 79.195 168.090 79.365 168.280 ;
        RECT 81.495 168.110 81.665 168.300 ;
        RECT 81.955 168.110 82.125 168.300 ;
        RECT 87.935 168.110 88.105 168.300 ;
        RECT 88.855 168.135 89.015 168.245 ;
        RECT 89.315 168.090 89.485 168.300 ;
        RECT 90.510 168.110 90.680 168.300 ;
        RECT 90.695 168.090 90.865 168.280 ;
        RECT 94.650 168.110 94.820 168.300 ;
        RECT 101.920 168.110 102.090 168.300 ;
        RECT 102.195 168.090 102.365 168.280 ;
        RECT 103.115 168.250 103.275 168.255 ;
        RECT 103.115 168.145 103.290 168.250 ;
        RECT 103.170 168.140 103.290 168.145 ;
        RECT 103.575 168.090 103.745 168.280 ;
        RECT 106.980 168.110 107.150 168.300 ;
        RECT 107.715 168.110 107.885 168.300 ;
        RECT 112.775 168.110 112.945 168.300 ;
        RECT 113.695 168.090 113.865 168.280 ;
        RECT 114.155 168.250 114.325 168.300 ;
        RECT 114.155 168.140 114.330 168.250 ;
        RECT 114.155 168.110 114.325 168.140 ;
        RECT 115.535 168.090 115.705 168.300 ;
        RECT 14.655 167.280 16.025 168.090 ;
        RECT 16.035 167.410 25.225 168.090 ;
        RECT 20.545 167.190 21.475 167.410 ;
        RECT 24.305 167.180 25.225 167.410 ;
        RECT 25.245 167.220 25.675 168.005 ;
        RECT 25.695 167.410 29.595 168.090 ;
        RECT 25.695 167.180 26.625 167.410 ;
        RECT 29.835 167.310 31.205 168.090 ;
        RECT 31.675 167.410 40.865 168.090 ;
        RECT 40.875 167.410 49.980 168.090 ;
        RECT 31.675 167.180 32.595 167.410 ;
        RECT 35.425 167.190 36.355 167.410 ;
        RECT 51.005 167.220 51.435 168.005 ;
        RECT 51.455 167.410 60.645 168.090 ;
        RECT 60.665 167.410 63.405 168.090 ;
        RECT 63.425 167.410 66.165 168.090 ;
        RECT 51.455 167.180 52.375 167.410 ;
        RECT 55.205 167.190 56.135 167.410 ;
        RECT 66.175 167.180 68.895 168.090 ;
        RECT 69.395 167.280 71.225 168.090 ;
        RECT 71.245 167.180 72.595 168.090 ;
        RECT 72.845 167.410 76.745 168.090 ;
        RECT 75.815 167.180 76.745 167.410 ;
        RECT 76.765 167.220 77.195 168.005 ;
        RECT 77.225 167.180 78.575 168.090 ;
        RECT 79.055 167.410 88.160 168.090 ;
        RECT 89.185 167.180 90.535 168.090 ;
        RECT 90.555 167.410 99.660 168.090 ;
        RECT 100.415 167.280 102.505 168.090 ;
        RECT 102.525 167.220 102.955 168.005 ;
        RECT 103.445 167.180 104.795 168.090 ;
        RECT 104.815 167.410 114.005 168.090 ;
        RECT 104.815 167.180 105.735 167.410 ;
        RECT 108.565 167.190 109.495 167.410 ;
        RECT 114.475 167.280 115.845 168.090 ;
      LAYER nwell ;
        RECT 14.460 164.060 116.040 166.890 ;
      LAYER pwell ;
        RECT 14.655 162.860 16.025 163.670 ;
        RECT 17.395 163.540 18.315 163.760 ;
        RECT 24.395 163.660 25.315 163.770 ;
        RECT 22.980 163.540 25.315 163.660 ;
        RECT 16.035 162.860 25.315 163.540 ;
        RECT 26.700 162.860 35.805 163.540 ;
        RECT 35.815 162.860 37.180 163.540 ;
        RECT 38.125 162.945 38.555 163.730 ;
        RECT 39.035 162.860 40.405 163.640 ;
        RECT 40.415 163.540 41.345 163.770 ;
        RECT 40.415 162.860 44.315 163.540 ;
        RECT 44.555 162.860 46.385 163.670 ;
        RECT 49.595 163.540 50.525 163.770 ;
        RECT 53.735 163.540 54.665 163.770 ;
        RECT 46.625 162.860 50.525 163.540 ;
        RECT 50.765 162.860 54.665 163.540 ;
        RECT 54.675 162.860 56.045 163.640 ;
        RECT 56.055 162.860 57.425 163.640 ;
        RECT 57.905 162.860 59.255 163.770 ;
        RECT 60.335 162.860 62.945 163.770 ;
        RECT 63.885 162.945 64.315 163.730 ;
        RECT 65.255 163.540 66.600 163.770 ;
        RECT 67.580 163.540 68.925 163.770 ;
        RECT 65.255 162.860 67.085 163.540 ;
        RECT 67.095 162.860 68.925 163.540 ;
        RECT 69.855 162.860 73.525 163.670 ;
        RECT 76.735 163.540 77.665 163.770 ;
        RECT 73.765 162.860 77.665 163.540 ;
        RECT 77.675 162.860 79.045 163.640 ;
        RECT 79.975 162.860 85.485 163.670 ;
        RECT 88.695 163.540 89.625 163.770 ;
        RECT 85.725 162.860 89.625 163.540 ;
        RECT 89.645 162.945 90.075 163.730 ;
        RECT 90.465 163.660 91.385 163.770 ;
        RECT 90.465 163.540 92.800 163.660 ;
        RECT 97.465 163.540 98.385 163.760 ;
        RECT 99.755 163.540 100.675 163.770 ;
        RECT 103.505 163.540 104.435 163.760 ;
        RECT 109.050 163.540 109.970 163.770 ;
        RECT 90.465 162.860 99.745 163.540 ;
        RECT 99.755 162.860 108.945 163.540 ;
        RECT 109.050 162.860 112.515 163.540 ;
        RECT 112.635 162.860 114.465 163.670 ;
        RECT 114.475 162.860 115.845 163.670 ;
        RECT 14.795 162.650 14.965 162.860 ;
        RECT 16.175 162.670 16.345 162.860 ;
        RECT 17.555 162.650 17.725 162.840 ;
        RECT 18.935 162.650 19.105 162.840 ;
        RECT 19.670 162.650 19.840 162.840 ;
        RECT 24.915 162.650 25.085 162.840 ;
        RECT 26.295 162.705 26.455 162.815 ;
        RECT 27.215 162.650 27.385 162.840 ;
        RECT 31.080 162.650 31.250 162.840 ;
        RECT 32.275 162.695 32.435 162.805 ;
        RECT 32.735 162.650 32.905 162.840 ;
        RECT 34.390 162.650 34.560 162.840 ;
        RECT 35.495 162.670 35.665 162.860 ;
        RECT 40.095 162.840 40.265 162.860 ;
        RECT 37.335 162.670 37.505 162.840 ;
        RECT 37.850 162.700 37.970 162.810 ;
        RECT 38.770 162.700 38.890 162.810 ;
        RECT 39.635 162.650 39.805 162.840 ;
        RECT 40.095 162.670 40.270 162.840 ;
        RECT 40.830 162.670 41.000 162.860 ;
        RECT 40.100 162.650 40.270 162.670 ;
        RECT 43.775 162.650 43.945 162.840 ;
        RECT 46.075 162.670 46.245 162.860 ;
        RECT 49.940 162.670 50.110 162.860 ;
        RECT 50.675 162.650 50.845 162.840 ;
        RECT 51.650 162.700 51.770 162.810 ;
        RECT 52.055 162.650 52.225 162.840 ;
        RECT 54.080 162.670 54.250 162.860 ;
        RECT 55.735 162.670 55.905 162.860 ;
        RECT 56.195 162.670 56.365 162.860 ;
        RECT 58.035 162.840 58.205 162.860 ;
        RECT 62.630 162.840 62.800 162.860 ;
        RECT 57.630 162.700 57.750 162.810 ;
        RECT 58.030 162.670 58.205 162.840 ;
        RECT 58.955 162.695 59.115 162.805 ;
        RECT 59.875 162.705 60.035 162.815 ;
        RECT 58.030 162.650 58.200 162.670 ;
        RECT 60.795 162.650 60.965 162.840 ;
        RECT 62.630 162.670 62.805 162.840 ;
        RECT 62.635 162.650 62.805 162.670 ;
        RECT 63.095 162.650 63.265 162.840 ;
        RECT 63.555 162.705 63.715 162.815 ;
        RECT 64.935 162.810 65.095 162.815 ;
        RECT 64.935 162.705 65.110 162.810 ;
        RECT 64.990 162.700 65.110 162.705 ;
        RECT 66.775 162.650 66.945 162.860 ;
        RECT 67.235 162.650 67.405 162.860 ;
        RECT 69.080 162.650 69.250 162.840 ;
        RECT 69.535 162.705 69.695 162.815 ;
        RECT 73.215 162.670 73.385 162.860 ;
        RECT 76.160 162.650 76.330 162.840 ;
        RECT 77.080 162.670 77.250 162.860 ;
        RECT 77.815 162.670 77.985 162.860 ;
        RECT 78.735 162.650 78.905 162.840 ;
        RECT 79.655 162.705 79.815 162.815 ;
        RECT 80.115 162.650 80.285 162.840 ;
        RECT 80.575 162.650 80.745 162.840 ;
        RECT 82.415 162.695 82.575 162.805 ;
        RECT 85.175 162.670 85.345 162.860 ;
        RECT 89.040 162.670 89.210 162.860 ;
        RECT 92.075 162.650 92.245 162.840 ;
        RECT 93.455 162.650 93.625 162.840 ;
        RECT 94.375 162.695 94.535 162.805 ;
        RECT 98.055 162.650 98.225 162.840 ;
        RECT 99.435 162.670 99.605 162.860 ;
        RECT 101.730 162.650 101.900 162.840 ;
        RECT 102.250 162.700 102.370 162.810 ;
        RECT 103.575 162.695 103.735 162.805 ;
        RECT 107.440 162.650 107.610 162.840 ;
        RECT 108.635 162.670 108.805 162.860 ;
        RECT 111.390 162.650 111.560 162.840 ;
        RECT 111.855 162.650 112.025 162.840 ;
        RECT 112.315 162.670 112.485 162.860 ;
        RECT 114.155 162.650 114.325 162.860 ;
        RECT 115.535 162.650 115.705 162.860 ;
        RECT 14.655 161.840 16.025 162.650 ;
        RECT 16.035 161.840 17.865 162.650 ;
        RECT 17.885 161.740 19.235 162.650 ;
        RECT 19.255 161.970 23.155 162.650 ;
        RECT 19.255 161.740 20.185 161.970 ;
        RECT 23.395 161.840 25.225 162.650 ;
        RECT 25.245 161.780 25.675 162.565 ;
        RECT 25.695 161.840 27.525 162.650 ;
        RECT 27.765 161.970 31.665 162.650 ;
        RECT 30.735 161.740 31.665 161.970 ;
        RECT 32.595 161.870 33.965 162.650 ;
        RECT 33.975 161.970 37.875 162.650 ;
        RECT 33.975 161.740 34.905 161.970 ;
        RECT 38.115 161.840 39.945 162.650 ;
        RECT 39.955 161.740 43.430 162.650 ;
        RECT 43.745 161.970 47.210 162.650 ;
        RECT 46.290 161.740 47.210 161.970 ;
        RECT 47.410 161.970 50.875 162.650 ;
        RECT 47.410 161.740 48.330 161.970 ;
        RECT 51.005 161.780 51.435 162.565 ;
        RECT 52.025 161.970 55.490 162.650 ;
        RECT 54.570 161.740 55.490 161.970 ;
        RECT 55.735 161.740 58.345 162.650 ;
        RECT 59.275 161.970 61.105 162.650 ;
        RECT 61.115 161.970 62.945 162.650 ;
        RECT 62.955 161.970 64.785 162.650 ;
        RECT 59.275 161.740 60.620 161.970 ;
        RECT 61.115 161.740 62.460 161.970 ;
        RECT 63.440 161.740 64.785 161.970 ;
        RECT 65.255 161.970 67.085 162.650 ;
        RECT 67.095 161.970 68.925 162.650 ;
        RECT 65.255 161.740 66.600 161.970 ;
        RECT 67.580 161.740 68.925 161.970 ;
        RECT 68.935 161.740 72.410 162.650 ;
        RECT 72.845 161.970 76.745 162.650 ;
        RECT 75.815 161.740 76.745 161.970 ;
        RECT 76.765 161.780 77.195 162.565 ;
        RECT 77.215 161.840 79.045 162.650 ;
        RECT 79.065 161.740 80.415 162.650 ;
        RECT 80.435 161.870 81.805 162.650 ;
        RECT 83.105 161.970 92.385 162.650 ;
        RECT 83.105 161.850 85.440 161.970 ;
        RECT 83.105 161.740 84.025 161.850 ;
        RECT 90.105 161.750 91.025 161.970 ;
        RECT 92.395 161.870 93.765 162.650 ;
        RECT 94.790 161.970 98.255 162.650 ;
        RECT 94.790 161.740 95.710 161.970 ;
        RECT 98.570 161.740 102.045 162.650 ;
        RECT 102.525 161.780 102.955 162.565 ;
        RECT 104.125 161.970 108.025 162.650 ;
        RECT 107.095 161.740 108.025 161.970 ;
        RECT 109.095 161.740 111.705 162.650 ;
        RECT 111.715 161.870 113.085 162.650 ;
        RECT 113.095 161.840 114.465 162.650 ;
        RECT 114.475 161.840 115.845 162.650 ;
      LAYER nwell ;
        RECT 14.460 158.620 116.040 161.450 ;
      LAYER pwell ;
        RECT 14.655 157.420 16.025 158.230 ;
        RECT 16.865 158.220 17.785 158.330 ;
        RECT 16.865 158.100 19.200 158.220 ;
        RECT 23.865 158.100 24.785 158.320 ;
        RECT 16.865 157.420 26.145 158.100 ;
        RECT 27.085 157.420 28.435 158.330 ;
        RECT 28.825 158.220 29.745 158.330 ;
        RECT 28.825 158.100 31.160 158.220 ;
        RECT 35.825 158.100 36.745 158.320 ;
        RECT 28.825 157.420 38.105 158.100 ;
        RECT 38.125 157.505 38.555 158.290 ;
        RECT 39.035 157.420 41.785 158.230 ;
        RECT 41.795 157.420 45.270 158.330 ;
        RECT 45.475 157.420 48.950 158.330 ;
        RECT 49.155 157.420 52.630 158.330 ;
        RECT 52.835 157.420 54.665 158.230 ;
        RECT 54.760 157.420 63.865 158.100 ;
        RECT 63.885 157.505 64.315 158.290 ;
        RECT 65.740 158.100 67.085 158.330 ;
        RECT 65.255 157.420 67.085 158.100 ;
        RECT 67.290 157.420 70.765 158.330 ;
        RECT 70.775 157.420 74.250 158.330 ;
        RECT 75.285 158.220 76.205 158.330 ;
        RECT 75.285 158.100 77.620 158.220 ;
        RECT 82.285 158.100 83.205 158.320 ;
        RECT 75.285 157.420 84.565 158.100 ;
        RECT 84.575 157.420 85.945 158.230 ;
        RECT 85.965 157.420 87.315 158.330 ;
        RECT 88.255 157.420 89.625 158.200 ;
        RECT 89.645 157.505 90.075 158.290 ;
        RECT 91.015 158.130 91.960 158.330 ;
        RECT 91.015 157.450 93.765 158.130 ;
        RECT 91.015 157.420 91.960 157.450 ;
        RECT 14.795 157.210 14.965 157.420 ;
        RECT 16.230 157.260 16.350 157.370 ;
        RECT 18.475 157.210 18.645 157.400 ;
        RECT 19.855 157.210 20.025 157.400 ;
        RECT 23.720 157.210 23.890 157.400 ;
        RECT 24.915 157.255 25.075 157.365 ;
        RECT 25.835 157.230 26.005 157.420 ;
        RECT 26.295 157.255 26.455 157.365 ;
        RECT 26.755 157.265 26.915 157.375 ;
        RECT 27.215 157.230 27.385 157.420 ;
        RECT 29.975 157.210 30.145 157.400 ;
        RECT 30.440 157.210 30.610 157.400 ;
        RECT 35.495 157.210 35.665 157.400 ;
        RECT 37.795 157.230 37.965 157.420 ;
        RECT 38.770 157.260 38.890 157.370 ;
        RECT 39.170 157.210 39.340 157.400 ;
        RECT 41.475 157.230 41.645 157.420 ;
        RECT 41.940 157.230 42.110 157.420 ;
        RECT 45.620 157.400 45.790 157.420 ;
        RECT 42.850 157.210 43.020 157.400 ;
        RECT 45.615 157.230 45.790 157.400 ;
        RECT 45.615 157.210 45.785 157.230 ;
        RECT 46.075 157.210 46.245 157.400 ;
        RECT 49.300 157.230 49.470 157.420 ;
        RECT 49.755 157.210 49.925 157.400 ;
        RECT 50.675 157.255 50.835 157.365 ;
        RECT 51.650 157.260 51.770 157.370 ;
        RECT 53.435 157.210 53.605 157.400 ;
        RECT 53.895 157.210 54.065 157.400 ;
        RECT 54.355 157.230 54.525 157.420 ;
        RECT 63.555 157.230 63.725 157.420 ;
        RECT 64.475 157.210 64.645 157.400 ;
        RECT 64.935 157.265 65.095 157.375 ;
        RECT 65.395 157.230 65.565 157.420 ;
        RECT 65.855 157.210 66.025 157.400 ;
        RECT 66.315 157.210 66.485 157.400 ;
        RECT 68.155 157.210 68.325 157.400 ;
        RECT 70.450 157.230 70.620 157.420 ;
        RECT 70.920 157.230 71.090 157.420 ;
        RECT 71.375 157.255 71.535 157.365 ;
        RECT 74.650 157.260 74.770 157.370 ;
        RECT 75.050 157.210 75.220 157.400 ;
        RECT 76.435 157.210 76.605 157.400 ;
        RECT 77.815 157.255 77.975 157.365 ;
        RECT 83.335 157.210 83.505 157.400 ;
        RECT 84.255 157.230 84.425 157.420 ;
        RECT 85.635 157.230 85.805 157.420 ;
        RECT 86.095 157.230 86.265 157.420 ;
        RECT 87.935 157.265 88.095 157.375 ;
        RECT 88.395 157.230 88.565 157.420 ;
        RECT 88.855 157.210 89.025 157.400 ;
        RECT 89.320 157.210 89.490 157.400 ;
        RECT 90.695 157.265 90.855 157.375 ;
        RECT 93.450 157.230 93.620 157.450 ;
        RECT 94.695 157.420 98.170 158.330 ;
        RECT 99.030 157.420 102.505 158.330 ;
        RECT 102.515 157.420 105.125 158.330 ;
        RECT 107.930 158.100 108.850 158.330 ;
        RECT 105.385 157.420 108.850 158.100 ;
        RECT 108.955 157.420 114.465 158.230 ;
        RECT 114.475 157.420 115.845 158.230 ;
        RECT 93.920 157.210 94.090 157.400 ;
        RECT 94.375 157.265 94.535 157.375 ;
        RECT 94.840 157.230 95.010 157.420 ;
        RECT 98.570 157.260 98.690 157.370 ;
        RECT 100.810 157.210 100.980 157.400 ;
        RECT 101.275 157.210 101.445 157.400 ;
        RECT 102.190 157.230 102.360 157.420 ;
        RECT 102.660 157.230 102.830 157.420 ;
        RECT 104.035 157.210 104.205 157.400 ;
        RECT 105.415 157.230 105.585 157.420 ;
        RECT 107.715 157.210 107.885 157.400 ;
        RECT 109.095 157.210 109.265 157.400 ;
        RECT 110.015 157.255 110.175 157.365 ;
        RECT 110.475 157.210 110.645 157.400 ;
        RECT 114.155 157.210 114.325 157.420 ;
        RECT 115.535 157.210 115.705 157.420 ;
        RECT 14.655 156.400 16.025 157.210 ;
        RECT 16.035 156.400 18.785 157.210 ;
        RECT 18.795 156.430 20.165 157.210 ;
        RECT 20.405 156.530 24.305 157.210 ;
        RECT 23.375 156.300 24.305 156.530 ;
        RECT 25.245 156.340 25.675 157.125 ;
        RECT 26.615 156.400 30.285 157.210 ;
        RECT 30.295 156.300 33.770 157.210 ;
        RECT 33.975 156.400 35.805 157.210 ;
        RECT 36.010 156.300 39.485 157.210 ;
        RECT 39.690 156.300 43.165 157.210 ;
        RECT 43.175 156.400 45.925 157.210 ;
        RECT 45.945 156.300 47.295 157.210 ;
        RECT 47.975 156.400 50.065 157.210 ;
        RECT 51.005 156.340 51.435 157.125 ;
        RECT 51.915 156.400 53.745 157.210 ;
        RECT 53.755 156.430 55.125 157.210 ;
        RECT 55.505 156.530 64.785 157.210 ;
        RECT 55.505 156.410 57.840 156.530 ;
        RECT 55.505 156.300 56.425 156.410 ;
        RECT 62.505 156.310 63.425 156.530 ;
        RECT 64.795 156.400 66.165 157.210 ;
        RECT 66.175 156.530 68.005 157.210 ;
        RECT 66.660 156.300 68.005 156.530 ;
        RECT 68.015 156.300 70.735 157.210 ;
        RECT 71.890 156.300 75.365 157.210 ;
        RECT 75.375 156.400 76.745 157.210 ;
        RECT 76.765 156.340 77.195 157.125 ;
        RECT 78.135 156.400 83.645 157.210 ;
        RECT 83.655 156.400 89.165 157.210 ;
        RECT 89.175 156.300 92.650 157.210 ;
        RECT 93.775 156.300 97.250 157.210 ;
        RECT 97.650 156.300 101.125 157.210 ;
        RECT 101.135 156.430 102.505 157.210 ;
        RECT 102.525 156.340 102.955 157.125 ;
        RECT 102.975 156.400 104.345 157.210 ;
        RECT 104.355 156.400 108.025 157.210 ;
        RECT 108.045 156.300 109.395 157.210 ;
        RECT 110.335 156.430 111.705 157.210 ;
        RECT 111.715 156.400 114.465 157.210 ;
        RECT 114.475 156.400 115.845 157.210 ;
      LAYER nwell ;
        RECT 14.460 153.180 116.040 156.010 ;
      LAYER pwell ;
        RECT 14.655 151.980 16.025 152.790 ;
        RECT 16.405 152.780 17.325 152.890 ;
        RECT 16.405 152.660 18.740 152.780 ;
        RECT 23.405 152.660 24.325 152.880 ;
        RECT 16.405 151.980 25.685 152.660 ;
        RECT 25.695 151.980 27.065 152.760 ;
        RECT 27.995 152.690 28.940 152.890 ;
        RECT 27.995 152.010 30.745 152.690 ;
        RECT 27.995 151.980 28.940 152.010 ;
        RECT 14.795 151.770 14.965 151.980 ;
        RECT 19.395 151.770 19.565 151.960 ;
        RECT 19.855 151.770 20.025 151.960 ;
        RECT 21.510 151.770 21.680 151.960 ;
        RECT 25.375 151.790 25.545 151.980 ;
        RECT 26.755 151.770 26.925 151.980 ;
        RECT 27.215 151.770 27.385 151.960 ;
        RECT 27.675 151.825 27.835 151.935 ;
        RECT 29.055 151.815 29.215 151.925 ;
        RECT 30.430 151.790 30.600 152.010 ;
        RECT 30.755 151.980 34.230 152.890 ;
        RECT 34.630 151.980 38.105 152.890 ;
        RECT 38.125 152.065 38.555 152.850 ;
        RECT 40.380 152.690 41.325 152.890 ;
        RECT 38.575 152.010 41.325 152.690 ;
        RECT 30.900 151.790 31.070 151.980 ;
        RECT 32.920 151.770 33.090 151.960 ;
        RECT 33.660 151.770 33.830 151.960 ;
        RECT 37.790 151.790 37.960 151.980 ;
        RECT 38.720 151.960 38.890 152.010 ;
        RECT 40.380 151.980 41.325 152.010 ;
        RECT 41.795 152.690 42.740 152.890 ;
        RECT 41.795 152.010 44.545 152.690 ;
        RECT 47.210 152.660 48.130 152.890 ;
        RECT 41.795 151.980 42.740 152.010 ;
        RECT 38.715 151.790 38.890 151.960 ;
        RECT 38.715 151.770 38.885 151.790 ;
        RECT 14.655 150.960 16.025 151.770 ;
        RECT 16.035 150.960 19.705 151.770 ;
        RECT 19.725 150.860 21.075 151.770 ;
        RECT 21.095 151.090 24.995 151.770 ;
        RECT 21.095 150.860 22.025 151.090 ;
        RECT 25.245 150.900 25.675 151.685 ;
        RECT 25.695 150.960 27.065 151.770 ;
        RECT 27.085 150.860 28.435 151.770 ;
        RECT 29.605 151.090 33.505 151.770 ;
        RECT 32.575 150.860 33.505 151.090 ;
        RECT 33.515 150.860 36.990 151.770 ;
        RECT 37.195 150.960 39.025 151.770 ;
        RECT 39.180 151.740 39.350 151.960 ;
        RECT 41.530 151.820 41.650 151.930 ;
        RECT 41.940 151.770 42.110 151.960 ;
        RECT 44.230 151.790 44.400 152.010 ;
        RECT 44.665 151.980 48.130 152.660 ;
        RECT 48.235 152.660 49.155 152.890 ;
        RECT 51.985 152.660 52.915 152.880 ;
        RECT 48.235 151.980 57.425 152.660 ;
        RECT 57.435 151.980 60.910 152.890 ;
        RECT 61.125 151.980 63.865 152.660 ;
        RECT 63.885 152.065 64.315 152.850 ;
        RECT 66.990 152.660 67.910 152.890 ;
        RECT 64.445 151.980 67.910 152.660 ;
        RECT 68.015 151.980 71.225 152.890 ;
        RECT 74.480 152.660 75.825 152.890 ;
        RECT 71.235 151.980 73.975 152.660 ;
        RECT 73.995 151.980 75.825 152.660 ;
        RECT 76.305 151.980 77.655 152.890 ;
        RECT 80.875 152.660 81.805 152.890 ;
        RECT 77.905 151.980 81.805 152.660 ;
        RECT 82.275 151.980 83.645 152.760 ;
        RECT 87.775 152.660 88.705 152.890 ;
        RECT 84.805 151.980 88.705 152.660 ;
        RECT 89.645 152.065 90.075 152.850 ;
        RECT 90.555 151.980 92.385 152.790 ;
        RECT 92.395 151.980 95.870 152.890 ;
        RECT 96.075 151.980 99.550 152.890 ;
        RECT 99.755 151.980 101.125 152.790 ;
        RECT 104.335 152.660 105.265 152.890 ;
        RECT 101.365 151.980 105.265 152.660 ;
        RECT 105.275 152.660 106.195 152.890 ;
        RECT 109.025 152.660 109.955 152.880 ;
        RECT 105.275 151.980 114.465 152.660 ;
        RECT 114.475 151.980 115.845 152.790 ;
        RECT 44.695 151.790 44.865 151.980 ;
        RECT 49.020 151.770 49.190 151.960 ;
        RECT 50.675 151.770 50.845 151.960 ;
        RECT 52.055 151.815 52.215 151.925 ;
        RECT 52.790 151.770 52.960 151.960 ;
        RECT 57.115 151.790 57.285 151.980 ;
        RECT 57.580 151.790 57.750 151.980 ;
        RECT 58.955 151.770 59.125 151.960 ;
        RECT 63.555 151.790 63.725 151.980 ;
        RECT 64.475 151.790 64.645 151.980 ;
        RECT 68.615 151.770 68.785 151.960 ;
        RECT 69.535 151.815 69.695 151.925 ;
        RECT 70.915 151.790 71.085 151.980 ;
        RECT 71.375 151.790 71.545 151.980 ;
        RECT 40.840 151.740 41.785 151.770 ;
        RECT 39.035 151.060 41.785 151.740 ;
        RECT 40.840 150.860 41.785 151.060 ;
        RECT 41.795 150.860 45.270 151.770 ;
        RECT 45.705 151.090 49.605 151.770 ;
        RECT 48.675 150.860 49.605 151.090 ;
        RECT 49.615 150.960 50.985 151.770 ;
        RECT 51.005 150.900 51.435 151.685 ;
        RECT 52.375 151.090 56.275 151.770 ;
        RECT 52.375 150.860 53.305 151.090 ;
        RECT 56.515 150.960 59.265 151.770 ;
        RECT 59.645 151.090 68.925 151.770 ;
        RECT 69.855 151.740 70.800 151.770 ;
        RECT 72.290 151.740 72.460 151.960 ;
        RECT 72.760 151.770 72.930 151.960 ;
        RECT 74.135 151.790 74.305 151.980 ;
        RECT 76.030 151.820 76.150 151.930 ;
        RECT 76.490 151.820 76.610 151.930 ;
        RECT 77.355 151.790 77.525 151.980 ;
        RECT 81.220 151.790 81.390 151.980 ;
        RECT 82.010 151.820 82.130 151.930 ;
        RECT 82.415 151.790 82.585 151.980 ;
        RECT 84.255 151.825 84.415 151.935 ;
        RECT 86.555 151.770 86.725 151.960 ;
        RECT 87.015 151.770 87.185 151.960 ;
        RECT 88.120 151.790 88.290 151.980 ;
        RECT 89.315 151.825 89.475 151.935 ;
        RECT 90.290 151.820 90.410 151.930 ;
        RECT 92.075 151.790 92.245 151.980 ;
        RECT 92.540 151.790 92.710 151.980 ;
        RECT 96.220 151.960 96.390 151.980 ;
        RECT 96.215 151.790 96.390 151.960 ;
        RECT 96.215 151.770 96.385 151.790 ;
        RECT 59.645 150.970 61.980 151.090 ;
        RECT 59.645 150.860 60.565 150.970 ;
        RECT 66.645 150.870 67.565 151.090 ;
        RECT 69.855 151.060 72.605 151.740 ;
        RECT 69.855 150.860 70.800 151.060 ;
        RECT 72.615 150.860 76.090 151.770 ;
        RECT 76.765 150.900 77.195 151.685 ;
        RECT 77.585 151.090 86.865 151.770 ;
        RECT 86.875 151.090 96.065 151.770 ;
        RECT 96.185 151.090 99.650 151.770 ;
        RECT 99.900 151.740 100.070 151.960 ;
        RECT 100.815 151.790 100.985 151.980 ;
        RECT 103.170 151.820 103.290 151.930 ;
        RECT 104.680 151.790 104.850 151.980 ;
        RECT 104.955 151.770 105.125 151.960 ;
        RECT 108.820 151.770 108.990 151.960 ;
        RECT 112.775 151.770 112.945 151.960 ;
        RECT 114.155 151.770 114.325 151.980 ;
        RECT 115.535 151.770 115.705 151.980 ;
        RECT 101.560 151.740 102.505 151.770 ;
        RECT 77.585 150.970 79.920 151.090 ;
        RECT 77.585 150.860 78.505 150.970 ;
        RECT 84.585 150.870 85.505 151.090 ;
        RECT 91.385 150.870 92.315 151.090 ;
        RECT 95.145 150.860 96.065 151.090 ;
        RECT 98.730 150.860 99.650 151.090 ;
        RECT 99.755 151.060 102.505 151.740 ;
        RECT 101.560 150.860 102.505 151.060 ;
        RECT 102.525 150.900 102.955 151.685 ;
        RECT 103.435 150.960 105.265 151.770 ;
        RECT 105.505 151.090 109.405 151.770 ;
        RECT 108.475 150.860 109.405 151.090 ;
        RECT 109.510 151.090 112.975 151.770 ;
        RECT 109.510 150.860 110.430 151.090 ;
        RECT 113.095 150.990 114.465 151.770 ;
        RECT 114.475 150.960 115.845 151.770 ;
      LAYER nwell ;
        RECT 14.460 147.740 116.040 150.570 ;
      LAYER pwell ;
        RECT 14.655 146.540 16.025 147.350 ;
        RECT 16.035 146.540 19.705 147.350 ;
        RECT 19.725 146.540 21.075 147.450 ;
        RECT 21.095 146.540 22.465 147.350 ;
        RECT 24.225 147.340 25.145 147.450 ;
        RECT 22.475 146.540 23.845 147.320 ;
        RECT 24.225 147.220 26.560 147.340 ;
        RECT 31.225 147.220 32.145 147.440 ;
        RECT 24.225 146.540 33.505 147.220 ;
        RECT 33.515 146.540 34.885 147.320 ;
        RECT 34.895 146.540 36.725 147.350 ;
        RECT 36.745 146.540 38.095 147.450 ;
        RECT 38.125 146.625 38.555 147.410 ;
        RECT 38.945 147.340 39.865 147.450 ;
        RECT 38.945 147.220 41.280 147.340 ;
        RECT 45.945 147.220 46.865 147.440 ;
        RECT 38.945 146.540 48.225 147.220 ;
        RECT 48.235 146.540 51.710 147.450 ;
        RECT 51.915 146.540 53.285 147.320 ;
        RECT 54.215 146.540 57.885 147.350 ;
        RECT 58.090 146.540 61.565 147.450 ;
        RECT 62.505 146.540 63.855 147.450 ;
        RECT 63.885 146.625 64.315 147.410 ;
        RECT 64.335 146.540 65.705 147.320 ;
        RECT 66.200 147.220 67.545 147.450 ;
        RECT 68.040 147.220 69.385 147.450 ;
        RECT 65.715 146.540 67.545 147.220 ;
        RECT 67.555 146.540 69.385 147.220 ;
        RECT 69.855 147.250 70.800 147.450 ;
        RECT 69.855 146.570 72.605 147.250 ;
        RECT 69.855 146.540 70.800 146.570 ;
        RECT 14.795 146.330 14.965 146.540 ;
        RECT 19.395 146.330 19.565 146.540 ;
        RECT 20.775 146.350 20.945 146.540 ;
        RECT 22.155 146.350 22.325 146.540 ;
        RECT 22.615 146.350 22.785 146.540 ;
        RECT 24.915 146.330 25.085 146.520 ;
        RECT 29.055 146.330 29.225 146.520 ;
        RECT 33.195 146.350 33.365 146.540 ;
        RECT 34.575 146.330 34.745 146.540 ;
        RECT 35.035 146.330 35.205 146.520 ;
        RECT 36.415 146.350 36.585 146.540 ;
        RECT 36.875 146.350 37.045 146.540 ;
        RECT 14.655 145.520 16.025 146.330 ;
        RECT 16.035 145.520 19.705 146.330 ;
        RECT 19.715 145.520 25.225 146.330 ;
        RECT 25.245 145.460 25.675 146.245 ;
        RECT 25.695 145.520 29.365 146.330 ;
        RECT 29.375 145.520 34.885 146.330 ;
        RECT 34.895 145.650 44.175 146.330 ;
        RECT 36.255 145.430 37.175 145.650 ;
        RECT 41.840 145.530 44.175 145.650 ;
        RECT 43.255 145.420 44.175 145.530 ;
        RECT 44.555 146.300 45.500 146.330 ;
        RECT 46.990 146.300 47.160 146.520 ;
        RECT 47.460 146.330 47.630 146.520 ;
        RECT 47.915 146.350 48.085 146.540 ;
        RECT 48.380 146.350 48.550 146.540 ;
        RECT 52.515 146.330 52.685 146.520 ;
        RECT 52.975 146.350 53.145 146.540 ;
        RECT 53.895 146.385 54.055 146.495 ;
        RECT 56.195 146.330 56.365 146.520 ;
        RECT 57.575 146.350 57.745 146.540 ;
        RECT 60.060 146.330 60.230 146.520 ;
        RECT 61.250 146.350 61.420 146.540 ;
        RECT 62.175 146.385 62.335 146.495 ;
        RECT 62.635 146.350 62.805 146.540 ;
        RECT 64.475 146.350 64.645 146.540 ;
        RECT 65.855 146.350 66.025 146.540 ;
        RECT 67.695 146.350 67.865 146.540 ;
        RECT 69.590 146.380 69.710 146.490 ;
        RECT 69.995 146.330 70.165 146.520 ;
        RECT 70.915 146.375 71.075 146.485 ;
        RECT 72.290 146.350 72.460 146.570 ;
        RECT 72.615 146.540 76.090 147.450 ;
        RECT 76.755 146.540 79.505 147.350 ;
        RECT 79.525 146.540 80.875 147.450 ;
        RECT 80.895 146.540 82.265 147.320 ;
        RECT 83.195 146.540 86.865 147.350 ;
        RECT 86.885 146.540 88.235 147.450 ;
        RECT 88.255 146.540 89.625 147.320 ;
        RECT 89.645 146.625 90.075 147.410 ;
        RECT 90.095 146.540 92.845 147.350 ;
        RECT 92.855 147.250 93.800 147.450 ;
        RECT 92.855 146.570 95.605 147.250 ;
        RECT 92.855 146.540 93.800 146.570 ;
        RECT 72.760 146.350 72.930 146.540 ;
        RECT 76.435 146.490 76.605 146.520 ;
        RECT 76.435 146.380 76.610 146.490 ;
        RECT 76.435 146.330 76.605 146.380 ;
        RECT 79.195 146.350 79.365 146.540 ;
        RECT 79.655 146.350 79.825 146.540 ;
        RECT 81.035 146.350 81.205 146.540 ;
        RECT 82.875 146.385 83.035 146.495 ;
        RECT 86.555 146.330 86.725 146.540 ;
        RECT 87.015 146.350 87.185 146.540 ;
        RECT 87.475 146.375 87.635 146.485 ;
        RECT 89.315 146.350 89.485 146.540 ;
        RECT 92.535 146.350 92.705 146.540 ;
        RECT 92.995 146.330 93.165 146.520 ;
        RECT 95.290 146.350 95.460 146.570 ;
        RECT 95.615 146.540 99.090 147.450 ;
        RECT 99.490 146.540 102.965 147.450 ;
        RECT 102.975 146.540 104.805 147.350 ;
        RECT 105.185 147.340 106.105 147.450 ;
        RECT 105.185 147.220 107.520 147.340 ;
        RECT 112.185 147.220 113.105 147.440 ;
        RECT 105.185 146.540 114.465 147.220 ;
        RECT 114.475 146.540 115.845 147.350 ;
        RECT 95.760 146.520 95.930 146.540 ;
        RECT 95.750 146.350 95.930 146.520 ;
        RECT 44.555 145.620 47.305 146.300 ;
        RECT 44.555 145.420 45.500 145.620 ;
        RECT 47.315 145.420 50.790 146.330 ;
        RECT 51.005 145.460 51.435 146.245 ;
        RECT 51.455 145.520 52.825 146.330 ;
        RECT 52.835 145.520 56.505 146.330 ;
        RECT 56.745 145.650 60.645 146.330 ;
        RECT 59.715 145.420 60.645 145.650 ;
        RECT 61.025 145.650 70.305 146.330 ;
        RECT 61.025 145.530 63.360 145.650 ;
        RECT 61.025 145.420 61.945 145.530 ;
        RECT 68.025 145.430 68.945 145.650 ;
        RECT 71.235 145.520 76.745 146.330 ;
        RECT 76.765 145.460 77.195 146.245 ;
        RECT 77.585 145.650 86.865 146.330 ;
        RECT 77.585 145.530 79.920 145.650 ;
        RECT 77.585 145.420 78.505 145.530 ;
        RECT 84.585 145.430 85.505 145.650 ;
        RECT 87.795 145.520 93.305 146.330 ;
        RECT 93.315 146.300 94.260 146.330 ;
        RECT 95.750 146.300 95.920 146.350 ;
        RECT 96.220 146.330 96.390 146.520 ;
        RECT 102.195 146.330 102.365 146.520 ;
        RECT 102.650 146.350 102.820 146.540 ;
        RECT 104.495 146.350 104.665 146.540 ;
        RECT 105.415 146.330 105.585 146.520 ;
        RECT 105.875 146.330 106.045 146.520 ;
        RECT 107.255 146.330 107.425 146.520 ;
        RECT 109.555 146.330 109.725 146.520 ;
        RECT 110.475 146.375 110.635 146.485 ;
        RECT 114.155 146.330 114.325 146.540 ;
        RECT 115.535 146.330 115.705 146.540 ;
        RECT 93.315 145.620 96.065 146.300 ;
        RECT 93.315 145.420 94.260 145.620 ;
        RECT 96.075 145.420 99.550 146.330 ;
        RECT 99.755 145.520 102.505 146.330 ;
        RECT 102.525 145.460 102.955 146.245 ;
        RECT 102.975 145.520 105.725 146.330 ;
        RECT 105.745 145.420 107.095 146.330 ;
        RECT 107.125 145.420 108.475 146.330 ;
        RECT 108.505 145.420 109.855 146.330 ;
        RECT 110.795 145.520 114.465 146.330 ;
        RECT 114.475 145.520 115.845 146.330 ;
      LAYER nwell ;
        RECT 14.460 142.300 116.040 145.130 ;
      LAYER pwell ;
        RECT 14.655 141.100 16.025 141.910 ;
        RECT 16.405 141.900 17.325 142.010 ;
        RECT 16.405 141.780 18.740 141.900 ;
        RECT 23.405 141.780 24.325 142.000 ;
        RECT 16.405 141.100 25.685 141.780 ;
        RECT 26.155 141.100 29.825 141.910 ;
        RECT 29.835 141.810 30.780 142.010 ;
        RECT 32.595 141.810 33.540 142.010 ;
        RECT 29.835 141.130 32.585 141.810 ;
        RECT 32.595 141.130 35.345 141.810 ;
        RECT 29.835 141.100 30.780 141.130 ;
        RECT 14.795 140.890 14.965 141.100 ;
        RECT 17.095 140.890 17.265 141.080 ;
        RECT 20.775 140.890 20.945 141.080 ;
        RECT 21.235 140.890 21.405 141.080 ;
        RECT 22.615 140.890 22.785 141.080 ;
        RECT 24.915 140.890 25.085 141.080 ;
        RECT 25.375 140.910 25.545 141.100 ;
        RECT 25.890 140.940 26.010 141.050 ;
        RECT 26.755 140.890 26.925 141.080 ;
        RECT 28.135 140.890 28.305 141.080 ;
        RECT 29.515 140.890 29.685 141.100 ;
        RECT 29.975 140.910 30.145 141.080 ;
        RECT 32.270 140.910 32.440 141.130 ;
        RECT 32.595 141.100 33.540 141.130 ;
        RECT 35.030 140.910 35.200 141.130 ;
        RECT 35.355 141.100 36.725 141.910 ;
        RECT 36.745 141.100 38.095 142.010 ;
        RECT 38.125 141.185 38.555 141.970 ;
        RECT 38.575 141.100 39.945 141.910 ;
        RECT 39.955 141.100 41.325 141.880 ;
        RECT 41.335 141.780 42.265 142.010 ;
        RECT 41.335 141.100 45.235 141.780 ;
        RECT 45.935 141.100 47.765 141.910 ;
        RECT 48.145 141.900 49.065 142.010 ;
        RECT 48.145 141.780 50.480 141.900 ;
        RECT 55.145 141.780 56.065 142.000 ;
        RECT 48.145 141.100 57.425 141.780 ;
        RECT 57.435 141.100 60.910 142.010 ;
        RECT 61.115 141.100 63.865 141.910 ;
        RECT 63.885 141.185 64.315 141.970 ;
        RECT 64.345 141.100 65.695 142.010 ;
        RECT 65.715 141.100 67.085 141.880 ;
        RECT 67.095 141.100 70.765 141.910 ;
        RECT 70.775 141.100 76.285 141.910 ;
        RECT 79.495 141.780 80.425 142.010 ;
        RECT 76.525 141.100 80.425 141.780 ;
        RECT 81.355 141.100 86.865 141.910 ;
        RECT 86.875 141.810 87.820 142.010 ;
        RECT 86.875 141.130 89.625 141.810 ;
        RECT 89.645 141.185 90.075 141.970 ;
        RECT 86.875 141.100 87.820 141.130 ;
        RECT 29.995 140.890 30.145 140.910 ;
        RECT 35.495 140.890 35.665 141.080 ;
        RECT 36.415 140.910 36.585 141.100 ;
        RECT 36.875 140.910 37.045 141.100 ;
        RECT 39.635 140.910 39.805 141.100 ;
        RECT 41.015 140.890 41.185 141.100 ;
        RECT 41.750 140.910 41.920 141.100 ;
        RECT 45.670 140.940 45.790 141.050 ;
        RECT 46.535 140.890 46.705 141.080 ;
        RECT 47.455 140.910 47.625 141.100 ;
        RECT 50.400 140.890 50.570 141.080 ;
        RECT 52.515 140.890 52.685 141.080 ;
        RECT 53.030 140.940 53.150 141.050 ;
        RECT 53.435 140.890 53.605 141.080 ;
        RECT 56.195 140.890 56.365 141.080 ;
        RECT 56.660 140.890 56.830 141.080 ;
        RECT 57.115 140.910 57.285 141.100 ;
        RECT 57.580 140.910 57.750 141.100 ;
        RECT 60.390 140.940 60.510 141.050 ;
        RECT 63.555 140.910 63.725 141.100 ;
        RECT 64.200 140.890 64.370 141.080 ;
        RECT 65.395 140.910 65.565 141.100 ;
        RECT 65.855 140.910 66.025 141.100 ;
        RECT 67.235 140.890 67.405 141.080 ;
        RECT 70.455 140.910 70.625 141.100 ;
        RECT 72.755 140.890 72.925 141.080 ;
        RECT 75.975 140.910 76.145 141.100 ;
        RECT 76.430 140.890 76.600 141.080 ;
        RECT 77.355 140.890 77.525 141.080 ;
        RECT 79.655 140.890 79.825 141.080 ;
        RECT 79.840 140.910 80.010 141.100 ;
        RECT 81.035 140.945 81.195 141.055 ;
        RECT 86.555 140.910 86.725 141.100 ;
        RECT 89.310 141.080 89.480 141.130 ;
        RECT 90.095 141.100 93.570 142.010 ;
        RECT 93.775 141.780 94.705 142.010 ;
        RECT 93.775 141.100 97.675 141.780 ;
        RECT 97.915 141.100 100.665 141.910 ;
        RECT 103.875 141.780 104.805 142.010 ;
        RECT 100.905 141.100 104.805 141.780 ;
        RECT 105.185 141.900 106.105 142.010 ;
        RECT 105.185 141.780 107.520 141.900 ;
        RECT 112.185 141.780 113.105 142.000 ;
        RECT 105.185 141.100 114.465 141.780 ;
        RECT 114.475 141.100 115.845 141.910 ;
        RECT 89.310 140.910 89.485 141.080 ;
        RECT 90.240 140.910 90.410 141.100 ;
        RECT 94.190 140.910 94.360 141.100 ;
        RECT 89.315 140.890 89.485 140.910 ;
        RECT 98.975 140.890 99.145 141.080 ;
        RECT 100.355 140.910 100.525 141.100 ;
        RECT 14.655 140.080 16.025 140.890 ;
        RECT 16.035 140.080 17.405 140.890 ;
        RECT 17.415 140.080 21.085 140.890 ;
        RECT 21.105 139.980 22.455 140.890 ;
        RECT 22.475 140.110 23.845 140.890 ;
        RECT 23.855 140.080 25.225 140.890 ;
        RECT 25.245 140.020 25.675 140.805 ;
        RECT 25.695 140.080 27.065 140.890 ;
        RECT 27.075 140.110 28.445 140.890 ;
        RECT 28.455 140.080 29.825 140.890 ;
        RECT 29.995 140.070 31.925 140.890 ;
        RECT 32.135 140.080 35.805 140.890 ;
        RECT 35.815 140.080 41.325 140.890 ;
        RECT 41.335 140.080 46.845 140.890 ;
        RECT 47.085 140.210 50.985 140.890 ;
        RECT 30.975 139.980 31.925 140.070 ;
        RECT 50.055 139.980 50.985 140.210 ;
        RECT 51.005 140.020 51.435 140.805 ;
        RECT 51.465 139.980 52.815 140.890 ;
        RECT 53.295 140.110 54.665 140.890 ;
        RECT 54.675 140.080 56.505 140.890 ;
        RECT 56.515 139.980 59.990 140.890 ;
        RECT 60.885 140.210 64.785 140.890 ;
        RECT 63.855 139.980 64.785 140.210 ;
        RECT 64.795 140.080 67.545 140.890 ;
        RECT 67.555 140.080 73.065 140.890 ;
        RECT 73.270 139.980 76.745 140.890 ;
        RECT 76.765 140.020 77.195 140.805 ;
        RECT 77.215 140.110 78.585 140.890 ;
        RECT 78.605 139.980 79.955 140.890 ;
        RECT 80.345 140.210 89.625 140.890 ;
        RECT 90.005 140.210 99.285 140.890 ;
        RECT 99.295 140.860 100.240 140.890 ;
        RECT 101.730 140.860 101.900 141.080 ;
        RECT 102.250 140.940 102.370 141.050 ;
        RECT 104.220 140.910 104.390 141.100 ;
        RECT 112.315 140.890 112.485 141.080 ;
        RECT 113.695 140.890 113.865 141.080 ;
        RECT 114.155 141.050 114.325 141.100 ;
        RECT 114.155 140.940 114.330 141.050 ;
        RECT 114.155 140.910 114.325 140.940 ;
        RECT 115.535 140.890 115.705 141.100 ;
        RECT 80.345 140.090 82.680 140.210 ;
        RECT 80.345 139.980 81.265 140.090 ;
        RECT 87.345 139.990 88.265 140.210 ;
        RECT 90.005 140.090 92.340 140.210 ;
        RECT 90.005 139.980 90.925 140.090 ;
        RECT 97.005 139.990 97.925 140.210 ;
        RECT 99.295 140.180 102.045 140.860 ;
        RECT 99.295 139.980 100.240 140.180 ;
        RECT 102.525 140.020 102.955 140.805 ;
        RECT 103.345 140.210 112.625 140.890 ;
        RECT 103.345 140.090 105.680 140.210 ;
        RECT 103.345 139.980 104.265 140.090 ;
        RECT 110.345 139.990 111.265 140.210 ;
        RECT 112.635 140.110 114.005 140.890 ;
        RECT 114.475 140.080 115.845 140.890 ;
      LAYER nwell ;
        RECT 14.460 136.860 116.040 139.690 ;
      LAYER pwell ;
        RECT 14.655 135.660 16.025 136.470 ;
        RECT 16.035 135.660 17.405 136.470 ;
        RECT 17.425 135.660 18.775 136.570 ;
        RECT 19.165 136.460 20.085 136.570 ;
        RECT 19.165 136.340 21.500 136.460 ;
        RECT 26.165 136.340 27.085 136.560 ;
        RECT 29.595 136.480 30.545 136.570 ;
        RECT 31.895 136.480 32.845 136.570 ;
        RECT 34.195 136.480 35.145 136.570 ;
        RECT 36.955 136.480 37.905 136.570 ;
        RECT 19.165 135.660 28.445 136.340 ;
        RECT 28.615 135.660 30.545 136.480 ;
        RECT 30.915 135.660 32.845 136.480 ;
        RECT 33.215 135.660 35.145 136.480 ;
        RECT 35.975 135.660 37.905 136.480 ;
        RECT 38.125 135.745 38.555 136.530 ;
        RECT 38.575 136.370 39.520 136.570 ;
        RECT 38.575 135.690 41.325 136.370 ;
        RECT 38.575 135.660 39.520 135.690 ;
        RECT 14.795 135.450 14.965 135.660 ;
        RECT 16.230 135.500 16.350 135.610 ;
        RECT 17.095 135.470 17.265 135.660 ;
        RECT 17.555 135.470 17.725 135.660 ;
        RECT 19.855 135.450 20.025 135.640 ;
        RECT 23.720 135.450 23.890 135.640 ;
        RECT 24.915 135.495 25.075 135.605 ;
        RECT 25.890 135.500 26.010 135.610 ;
        RECT 26.570 135.450 26.740 135.640 ;
        RECT 28.135 135.470 28.305 135.660 ;
        RECT 28.615 135.640 28.765 135.660 ;
        RECT 30.915 135.640 31.065 135.660 ;
        RECT 33.215 135.640 33.365 135.660 ;
        RECT 35.975 135.640 36.125 135.660 ;
        RECT 28.595 135.470 28.765 135.640 ;
        RECT 30.435 135.450 30.605 135.640 ;
        RECT 30.895 135.470 31.065 135.640 ;
        RECT 33.195 135.470 33.365 135.640 ;
        RECT 35.220 135.450 35.390 135.640 ;
        RECT 35.550 135.500 35.670 135.610 ;
        RECT 35.955 135.470 36.125 135.640 ;
        RECT 37.335 135.450 37.505 135.640 ;
        RECT 14.655 134.640 16.025 135.450 ;
        RECT 16.495 134.640 20.165 135.450 ;
        RECT 20.405 134.770 24.305 135.450 ;
        RECT 23.375 134.540 24.305 134.770 ;
        RECT 25.245 134.580 25.675 135.365 ;
        RECT 26.155 134.770 30.055 135.450 ;
        RECT 26.155 134.540 27.085 134.770 ;
        RECT 30.305 134.540 31.655 135.450 ;
        RECT 31.905 134.770 35.805 135.450 ;
        RECT 34.875 134.540 35.805 134.770 ;
        RECT 35.815 134.640 37.645 135.450 ;
        RECT 37.655 135.420 38.600 135.450 ;
        RECT 40.090 135.420 40.260 135.640 ;
        RECT 41.010 135.470 41.180 135.690 ;
        RECT 41.335 135.660 46.845 136.470 ;
        RECT 46.855 135.660 50.330 136.570 ;
        RECT 51.465 135.660 52.815 136.570 ;
        RECT 53.295 135.660 56.965 136.470 ;
        RECT 56.975 135.660 62.485 136.470 ;
        RECT 62.505 135.660 63.855 136.570 ;
        RECT 63.885 135.745 64.315 136.530 ;
        RECT 64.335 135.660 65.705 136.470 ;
        RECT 68.475 136.370 69.420 136.570 ;
        RECT 65.715 135.660 67.545 136.340 ;
        RECT 68.475 135.690 71.225 136.370 ;
        RECT 68.475 135.660 69.420 135.690 ;
        RECT 40.415 135.420 41.360 135.450 ;
        RECT 42.850 135.420 43.020 135.640 ;
        RECT 43.320 135.450 43.490 135.640 ;
        RECT 46.535 135.470 46.705 135.660 ;
        RECT 47.000 135.470 47.170 135.660 ;
        RECT 50.400 135.450 50.570 135.640 ;
        RECT 51.135 135.505 51.295 135.615 ;
        RECT 51.595 135.610 51.765 135.660 ;
        RECT 51.595 135.500 51.770 135.610 ;
        RECT 51.595 135.470 51.765 135.500 ;
        RECT 52.055 135.450 52.225 135.640 ;
        RECT 53.030 135.500 53.150 135.610 ;
        RECT 56.655 135.470 56.825 135.660 ;
        RECT 56.840 135.450 57.010 135.640 ;
        RECT 58.495 135.450 58.665 135.640 ;
        RECT 62.175 135.470 62.345 135.660 ;
        RECT 63.555 135.470 63.725 135.660 ;
        RECT 65.395 135.470 65.565 135.660 ;
        RECT 67.235 135.470 67.405 135.660 ;
        RECT 68.155 135.450 68.325 135.640 ;
        RECT 70.910 135.470 71.080 135.690 ;
        RECT 71.235 135.660 74.710 136.570 ;
        RECT 75.285 136.460 76.205 136.570 ;
        RECT 75.285 136.340 77.620 136.460 ;
        RECT 82.285 136.340 83.205 136.560 ;
        RECT 87.775 136.340 88.705 136.570 ;
        RECT 75.285 135.660 84.565 136.340 ;
        RECT 84.805 135.660 88.705 136.340 ;
        RECT 89.645 135.745 90.075 136.530 ;
        RECT 90.095 135.660 91.465 136.470 ;
        RECT 91.485 135.660 92.835 136.570 ;
        RECT 95.815 136.480 96.765 136.570 ;
        RECT 92.855 135.660 94.225 136.470 ;
        RECT 94.235 135.660 95.605 136.440 ;
        RECT 95.815 135.660 97.745 136.480 ;
        RECT 97.915 135.660 99.285 136.470 ;
        RECT 99.295 135.660 102.965 136.470 ;
        RECT 106.175 136.340 107.105 136.570 ;
        RECT 103.205 135.660 107.105 136.340 ;
        RECT 107.575 135.660 108.945 136.440 ;
        RECT 108.955 135.660 114.465 136.470 ;
        RECT 114.475 135.660 115.845 136.470 ;
        RECT 71.380 135.470 71.550 135.660 ;
        RECT 71.835 135.450 72.005 135.640 ;
        RECT 37.655 134.740 40.405 135.420 ;
        RECT 40.415 134.740 43.165 135.420 ;
        RECT 37.655 134.540 38.600 134.740 ;
        RECT 40.415 134.540 41.360 134.740 ;
        RECT 43.175 134.540 46.650 135.450 ;
        RECT 47.085 134.770 50.985 135.450 ;
        RECT 50.055 134.540 50.985 134.770 ;
        RECT 51.005 134.580 51.435 135.365 ;
        RECT 51.915 134.670 53.285 135.450 ;
        RECT 53.525 134.770 57.425 135.450 ;
        RECT 56.495 134.540 57.425 134.770 ;
        RECT 57.435 134.640 58.805 135.450 ;
        RECT 59.185 134.770 68.465 135.450 ;
        RECT 59.185 134.650 61.520 134.770 ;
        RECT 59.185 134.540 60.105 134.650 ;
        RECT 66.185 134.550 67.105 134.770 ;
        RECT 68.475 134.640 72.145 135.450 ;
        RECT 72.155 135.420 73.100 135.450 ;
        RECT 74.590 135.420 74.760 135.640 ;
        RECT 76.435 135.450 76.605 135.640 ;
        RECT 77.630 135.450 77.800 135.640 ;
        RECT 81.550 135.500 81.670 135.610 ;
        RECT 83.335 135.450 83.505 135.640 ;
        RECT 84.255 135.470 84.425 135.660 ;
        RECT 84.715 135.450 84.885 135.640 ;
        RECT 85.635 135.495 85.795 135.605 ;
        RECT 87.015 135.450 87.185 135.640 ;
        RECT 88.120 135.470 88.290 135.660 ;
        RECT 88.395 135.450 88.565 135.640 ;
        RECT 89.315 135.505 89.475 135.615 ;
        RECT 89.775 135.450 89.945 135.640 ;
        RECT 91.155 135.470 91.325 135.660 ;
        RECT 91.615 135.470 91.785 135.660 ;
        RECT 92.075 135.470 92.245 135.640 ;
        RECT 93.915 135.470 94.085 135.660 ;
        RECT 94.375 135.470 94.545 135.660 ;
        RECT 97.595 135.640 97.745 135.660 ;
        RECT 95.295 135.495 95.455 135.605 ;
        RECT 97.595 135.470 97.765 135.640 ;
        RECT 92.075 135.450 92.225 135.470 ;
        RECT 94.375 135.450 94.525 135.470 ;
        RECT 98.055 135.450 98.225 135.640 ;
        RECT 98.515 135.470 98.685 135.640 ;
        RECT 98.975 135.470 99.145 135.660 ;
        RECT 98.535 135.450 98.685 135.470 ;
        RECT 102.195 135.450 102.365 135.640 ;
        RECT 102.655 135.470 102.825 135.660 ;
        RECT 103.170 135.500 103.290 135.610 ;
        RECT 106.520 135.470 106.690 135.660 ;
        RECT 107.310 135.500 107.430 135.610 ;
        RECT 107.715 135.470 107.885 135.660 ;
        RECT 108.635 135.450 108.805 135.640 ;
        RECT 114.155 135.450 114.325 135.660 ;
        RECT 115.535 135.450 115.705 135.660 ;
        RECT 72.155 134.740 74.905 135.420 ;
        RECT 72.155 134.540 73.100 134.740 ;
        RECT 74.915 134.640 76.745 135.450 ;
        RECT 76.765 134.580 77.195 135.365 ;
        RECT 77.215 134.770 81.115 135.450 ;
        RECT 77.215 134.540 78.145 134.770 ;
        RECT 81.815 134.640 83.645 135.450 ;
        RECT 83.665 134.540 85.015 135.450 ;
        RECT 85.955 134.670 87.325 135.450 ;
        RECT 87.335 134.670 88.705 135.450 ;
        RECT 88.715 134.640 90.085 135.450 ;
        RECT 90.295 134.630 92.225 135.450 ;
        RECT 92.595 134.630 94.525 135.450 ;
        RECT 95.625 134.770 98.365 135.450 ;
        RECT 98.535 134.630 100.465 135.450 ;
        RECT 100.675 134.640 102.505 135.450 ;
        RECT 90.295 134.540 91.245 134.630 ;
        RECT 92.595 134.540 93.545 134.630 ;
        RECT 99.515 134.540 100.465 134.630 ;
        RECT 102.525 134.580 102.955 135.365 ;
        RECT 103.435 134.640 108.945 135.450 ;
        RECT 108.955 134.640 114.465 135.450 ;
        RECT 114.475 134.640 115.845 135.450 ;
      LAYER nwell ;
        RECT 14.460 131.420 116.040 134.250 ;
      LAYER pwell ;
        RECT 14.655 130.220 16.025 131.030 ;
        RECT 16.865 131.020 17.785 131.130 ;
        RECT 16.865 130.900 19.200 131.020 ;
        RECT 23.865 130.900 24.785 131.120 ;
        RECT 16.865 130.220 26.145 130.900 ;
        RECT 26.165 130.220 27.515 131.130 ;
        RECT 27.905 131.020 28.825 131.130 ;
        RECT 27.905 130.900 30.240 131.020 ;
        RECT 34.905 130.900 35.825 131.120 ;
        RECT 27.905 130.220 37.185 130.900 ;
        RECT 38.125 130.305 38.555 131.090 ;
        RECT 39.715 131.040 40.665 131.130 ;
        RECT 38.735 130.220 40.665 131.040 ;
        RECT 42.455 131.040 43.405 131.130 ;
        RECT 40.875 130.220 42.245 131.030 ;
        RECT 42.455 130.220 44.385 131.040 ;
        RECT 44.555 130.220 48.030 131.130 ;
        RECT 48.605 131.020 49.525 131.130 ;
        RECT 48.605 130.900 50.940 131.020 ;
        RECT 55.605 130.900 56.525 131.120 ;
        RECT 62.015 130.900 62.945 131.130 ;
        RECT 48.605 130.220 57.885 130.900 ;
        RECT 59.045 130.220 62.945 130.900 ;
        RECT 63.885 130.305 64.315 131.090 ;
        RECT 65.455 131.040 66.405 131.130 ;
        RECT 72.355 131.040 73.305 131.130 ;
        RECT 65.455 130.220 67.385 131.040 ;
        RECT 67.555 130.220 69.385 130.900 ;
        RECT 69.395 130.220 70.765 131.000 ;
        RECT 70.775 130.220 72.145 131.030 ;
        RECT 72.355 130.220 74.285 131.040 ;
        RECT 74.455 130.220 75.825 131.030 ;
        RECT 85.035 130.900 85.965 131.130 ;
        RECT 75.920 130.220 85.025 130.900 ;
        RECT 85.035 130.220 88.935 130.900 ;
        RECT 89.645 130.305 90.075 131.090 ;
        RECT 100.435 131.040 101.385 131.130 ;
        RECT 90.180 130.220 99.285 130.900 ;
        RECT 99.455 130.220 101.385 131.040 ;
        RECT 104.795 130.900 105.725 131.130 ;
        RECT 101.825 130.220 105.725 130.900 ;
        RECT 105.735 130.220 107.565 131.030 ;
        RECT 107.585 130.220 108.935 131.130 ;
        RECT 109.415 130.220 110.785 131.000 ;
        RECT 110.795 130.220 114.465 131.030 ;
        RECT 114.475 130.220 115.845 131.030 ;
        RECT 14.795 130.010 14.965 130.220 ;
        RECT 16.230 130.060 16.350 130.170 ;
        RECT 18.475 130.010 18.645 130.200 ;
        RECT 18.935 130.010 19.105 130.200 ;
        RECT 20.590 130.010 20.760 130.200 ;
        RECT 24.915 130.055 25.075 130.165 ;
        RECT 25.835 130.030 26.005 130.220 ;
        RECT 26.295 130.030 26.465 130.220 ;
        RECT 35.495 130.010 35.665 130.200 ;
        RECT 36.875 130.010 37.045 130.220 ;
        RECT 38.735 130.200 38.885 130.220 ;
        RECT 37.795 130.065 37.955 130.175 ;
        RECT 38.715 130.030 38.885 130.200 ;
        RECT 40.740 130.010 40.910 130.200 ;
        RECT 41.475 130.010 41.645 130.200 ;
        RECT 41.935 130.030 42.105 130.220 ;
        RECT 44.235 130.200 44.385 130.220 ;
        RECT 44.235 130.030 44.405 130.200 ;
        RECT 44.700 130.030 44.870 130.220 ;
        RECT 50.730 130.060 50.850 130.170 ;
        RECT 52.975 130.010 53.145 130.200 ;
        RECT 57.575 130.030 57.745 130.220 ;
        RECT 58.495 130.065 58.655 130.175 ;
        RECT 62.360 130.030 62.530 130.220 ;
        RECT 67.235 130.200 67.385 130.220 ;
        RECT 62.635 130.010 62.805 130.200 ;
        RECT 63.555 130.065 63.715 130.175 ;
        RECT 64.935 130.065 65.095 130.175 ;
        RECT 65.395 130.010 65.565 130.200 ;
        RECT 65.855 130.010 66.025 130.200 ;
        RECT 67.235 130.030 67.405 130.200 ;
        RECT 67.695 130.030 67.865 130.220 ;
        RECT 69.995 130.010 70.165 130.200 ;
        RECT 70.455 130.030 70.625 130.220 ;
        RECT 71.835 130.030 72.005 130.220 ;
        RECT 74.135 130.200 74.285 130.220 ;
        RECT 72.295 130.030 72.465 130.200 ;
        RECT 74.135 130.030 74.305 130.200 ;
        RECT 75.515 130.030 75.685 130.220 ;
        RECT 72.295 130.010 72.445 130.030 ;
        RECT 76.160 130.010 76.330 130.200 ;
        RECT 79.195 130.030 79.365 130.200 ;
        RECT 79.195 130.010 79.345 130.030 ;
        RECT 82.875 130.010 83.045 130.200 ;
        RECT 83.335 130.010 83.505 130.200 ;
        RECT 84.715 130.030 84.885 130.220 ;
        RECT 85.450 130.030 85.620 130.220 ;
        RECT 89.370 130.060 89.490 130.170 ;
        RECT 94.375 130.010 94.545 130.200 ;
        RECT 96.675 130.030 96.845 130.200 ;
        RECT 96.675 130.010 96.825 130.030 ;
        RECT 98.055 130.010 98.225 130.200 ;
        RECT 98.975 130.030 99.145 130.220 ;
        RECT 99.455 130.200 99.605 130.220 ;
        RECT 99.435 130.030 99.605 130.200 ;
        RECT 101.920 130.010 102.090 130.200 ;
        RECT 103.170 130.060 103.290 130.170 ;
        RECT 104.495 130.010 104.665 130.200 ;
        RECT 105.140 130.030 105.310 130.220 ;
        RECT 107.255 130.030 107.425 130.220 ;
        RECT 107.715 130.030 107.885 130.220 ;
        RECT 109.150 130.060 109.270 130.170 ;
        RECT 109.555 130.030 109.725 130.220 ;
        RECT 114.155 130.010 114.325 130.220 ;
        RECT 115.535 130.010 115.705 130.220 ;
        RECT 14.655 129.200 16.025 130.010 ;
        RECT 16.035 129.200 18.785 130.010 ;
        RECT 18.795 129.230 20.165 130.010 ;
        RECT 20.175 129.330 24.075 130.010 ;
        RECT 20.175 129.100 21.105 129.330 ;
        RECT 25.245 129.140 25.675 129.925 ;
        RECT 26.700 129.330 35.805 130.010 ;
        RECT 35.815 129.230 37.185 130.010 ;
        RECT 37.425 129.330 41.325 130.010 ;
        RECT 41.335 129.330 50.440 130.010 ;
        RECT 40.395 129.100 41.325 129.330 ;
        RECT 51.005 129.140 51.435 129.925 ;
        RECT 51.455 129.200 53.285 130.010 ;
        RECT 53.665 129.330 62.945 130.010 ;
        RECT 62.965 129.330 65.705 130.010 ;
        RECT 65.715 129.330 68.455 130.010 ;
        RECT 53.665 129.210 56.000 129.330 ;
        RECT 53.665 129.100 54.585 129.210 ;
        RECT 60.665 129.110 61.585 129.330 ;
        RECT 68.475 129.200 70.305 130.010 ;
        RECT 70.515 129.190 72.445 130.010 ;
        RECT 72.845 129.330 76.745 130.010 ;
        RECT 70.515 129.100 71.465 129.190 ;
        RECT 75.815 129.100 76.745 129.330 ;
        RECT 76.765 129.140 77.195 129.925 ;
        RECT 77.415 129.190 79.345 130.010 ;
        RECT 79.515 129.200 83.185 130.010 ;
        RECT 83.195 129.330 92.475 130.010 ;
        RECT 77.415 129.100 78.365 129.190 ;
        RECT 84.555 129.110 85.475 129.330 ;
        RECT 90.140 129.210 92.475 129.330 ;
        RECT 91.555 129.100 92.475 129.210 ;
        RECT 92.855 129.200 94.685 130.010 ;
        RECT 94.895 129.190 96.825 130.010 ;
        RECT 96.995 129.200 98.365 130.010 ;
        RECT 98.605 129.330 102.505 130.010 ;
        RECT 94.895 129.100 95.845 129.190 ;
        RECT 101.575 129.100 102.505 129.330 ;
        RECT 102.525 129.140 102.955 129.925 ;
        RECT 103.445 129.100 104.795 130.010 ;
        RECT 105.185 129.330 114.465 130.010 ;
        RECT 105.185 129.210 107.520 129.330 ;
        RECT 105.185 129.100 106.105 129.210 ;
        RECT 112.185 129.110 113.105 129.330 ;
        RECT 114.475 129.200 115.845 130.010 ;
      LAYER nwell ;
        RECT 14.460 125.980 116.040 128.810 ;
      LAYER pwell ;
        RECT 14.655 124.780 16.025 125.590 ;
        RECT 16.865 125.580 17.785 125.690 ;
        RECT 16.865 125.460 19.200 125.580 ;
        RECT 23.865 125.460 24.785 125.680 ;
        RECT 16.865 124.780 26.145 125.460 ;
        RECT 27.075 124.780 28.445 125.560 ;
        RECT 29.815 125.460 30.735 125.680 ;
        RECT 36.815 125.580 37.735 125.690 ;
        RECT 35.400 125.460 37.735 125.580 ;
        RECT 28.455 124.780 37.735 125.460 ;
        RECT 38.125 124.865 38.555 125.650 ;
        RECT 39.515 124.780 50.525 125.690 ;
        RECT 50.735 125.600 51.685 125.690 ;
        RECT 50.735 124.780 52.665 125.600 ;
        RECT 53.295 124.780 56.965 125.590 ;
        RECT 56.985 124.780 58.335 125.690 ;
        RECT 58.355 124.780 59.725 125.560 ;
        RECT 60.195 124.780 63.865 125.590 ;
        RECT 63.885 124.865 64.315 125.650 ;
        RECT 64.335 124.780 67.085 125.590 ;
        RECT 67.095 125.460 68.025 125.690 ;
        RECT 71.435 125.600 72.385 125.690 ;
        RECT 67.095 124.780 70.995 125.460 ;
        RECT 71.435 124.780 73.365 125.600 ;
        RECT 73.905 125.580 74.825 125.690 ;
        RECT 73.905 125.460 76.240 125.580 ;
        RECT 80.905 125.460 81.825 125.680 ;
        RECT 73.905 124.780 83.185 125.460 ;
        RECT 83.195 124.780 84.565 125.560 ;
        RECT 85.035 124.780 86.865 125.590 ;
        RECT 86.885 124.780 88.235 125.690 ;
        RECT 88.255 124.780 89.625 125.590 ;
        RECT 89.645 124.865 90.075 125.650 ;
        RECT 90.095 125.460 91.025 125.690 ;
        RECT 90.095 124.780 93.995 125.460 ;
        RECT 94.235 124.780 95.605 125.590 ;
        RECT 98.815 125.460 99.745 125.690 ;
        RECT 95.845 124.780 99.745 125.460 ;
        RECT 100.125 125.580 101.045 125.690 ;
        RECT 100.125 125.460 102.460 125.580 ;
        RECT 107.125 125.460 108.045 125.680 ;
        RECT 100.125 124.780 109.405 125.460 ;
        RECT 109.415 124.780 110.785 125.560 ;
        RECT 110.795 124.780 114.465 125.590 ;
        RECT 114.475 124.780 115.845 125.590 ;
        RECT 14.795 124.570 14.965 124.780 ;
        RECT 16.230 124.620 16.350 124.730 ;
        RECT 17.555 124.570 17.725 124.760 ;
        RECT 18.015 124.570 18.185 124.760 ;
        RECT 19.395 124.570 19.565 124.760 ;
        RECT 21.050 124.570 21.220 124.760 ;
        RECT 24.970 124.620 25.090 124.730 ;
        RECT 25.835 124.590 26.005 124.780 ;
        RECT 26.295 124.615 26.455 124.725 ;
        RECT 26.755 124.625 26.915 124.735 ;
        RECT 27.030 124.570 27.200 124.760 ;
        RECT 28.135 124.590 28.305 124.780 ;
        RECT 28.595 124.590 28.765 124.780 ;
        RECT 31.355 124.615 31.515 124.725 ;
        RECT 32.735 124.570 32.905 124.760 ;
        RECT 34.575 124.590 34.745 124.760 ;
        RECT 39.175 124.625 39.335 124.735 ;
        RECT 44.235 124.570 44.405 124.760 ;
        RECT 46.535 124.590 46.705 124.760 ;
        RECT 50.210 124.590 50.380 124.780 ;
        RECT 52.515 124.760 52.665 124.780 ;
        RECT 46.535 124.570 46.685 124.590 ;
        RECT 50.400 124.570 50.570 124.760 ;
        RECT 51.650 124.620 51.770 124.730 ;
        RECT 52.515 124.590 52.685 124.760 ;
        RECT 53.030 124.620 53.150 124.730 ;
        RECT 53.435 124.570 53.605 124.760 ;
        RECT 53.895 124.570 54.065 124.760 ;
        RECT 56.655 124.590 56.825 124.780 ;
        RECT 57.570 124.570 57.740 124.760 ;
        RECT 58.035 124.590 58.205 124.780 ;
        RECT 58.495 124.590 58.665 124.780 ;
        RECT 59.930 124.620 60.050 124.730 ;
        RECT 61.255 124.570 61.425 124.760 ;
        RECT 61.715 124.570 61.885 124.760 ;
        RECT 63.555 124.590 63.725 124.780 ;
        RECT 66.775 124.590 66.945 124.780 ;
        RECT 67.510 124.590 67.680 124.780 ;
        RECT 73.215 124.760 73.365 124.780 ;
        RECT 73.215 124.590 73.385 124.760 ;
        RECT 74.780 124.570 74.950 124.760 ;
        RECT 76.435 124.570 76.605 124.760 ;
        RECT 78.275 124.570 78.445 124.760 ;
        RECT 79.195 124.615 79.355 124.725 ;
        RECT 82.875 124.590 83.045 124.780 ;
        RECT 83.060 124.570 83.230 124.760 ;
        RECT 84.255 124.590 84.425 124.780 ;
        RECT 84.770 124.620 84.890 124.730 ;
        RECT 86.555 124.590 86.725 124.780 ;
        RECT 87.015 124.590 87.185 124.780 ;
        RECT 89.315 124.590 89.485 124.780 ;
        RECT 90.510 124.590 90.680 124.780 ;
        RECT 92.995 124.570 93.165 124.760 ;
        RECT 94.375 124.570 94.545 124.760 ;
        RECT 94.835 124.570 95.005 124.760 ;
        RECT 95.295 124.590 95.465 124.780 ;
        RECT 99.160 124.590 99.330 124.780 ;
        RECT 99.620 124.570 99.790 124.760 ;
        RECT 100.815 124.615 100.975 124.725 ;
        RECT 101.275 124.570 101.445 124.760 ;
        RECT 109.095 124.590 109.265 124.780 ;
        RECT 109.555 124.590 109.725 124.780 ;
        RECT 112.315 124.570 112.485 124.760 ;
        RECT 114.155 124.570 114.325 124.780 ;
        RECT 115.535 124.570 115.705 124.780 ;
        RECT 14.655 123.760 16.025 124.570 ;
        RECT 16.505 123.660 17.855 124.570 ;
        RECT 17.885 123.660 19.235 124.570 ;
        RECT 19.255 123.790 20.625 124.570 ;
        RECT 20.635 123.890 24.535 124.570 ;
        RECT 20.635 123.660 21.565 123.890 ;
        RECT 25.245 123.700 25.675 124.485 ;
        RECT 26.615 123.890 30.515 124.570 ;
        RECT 26.615 123.660 27.545 123.890 ;
        RECT 31.675 123.790 33.045 124.570 ;
        RECT 33.055 123.890 34.420 124.570 ;
        RECT 35.265 123.890 44.545 124.570 ;
        RECT 35.265 123.770 37.600 123.890 ;
        RECT 35.265 123.660 36.185 123.770 ;
        RECT 42.265 123.670 43.185 123.890 ;
        RECT 44.755 123.750 46.685 124.570 ;
        RECT 47.085 123.890 50.985 124.570 ;
        RECT 44.755 123.660 45.705 123.750 ;
        RECT 50.055 123.660 50.985 123.890 ;
        RECT 51.005 123.700 51.435 124.485 ;
        RECT 51.915 123.760 53.745 124.570 ;
        RECT 53.765 123.660 55.115 124.570 ;
        RECT 55.275 123.660 57.885 124.570 ;
        RECT 57.895 123.760 61.565 124.570 ;
        RECT 61.575 123.890 70.855 124.570 ;
        RECT 71.465 123.890 75.365 124.570 ;
        RECT 62.935 123.670 63.855 123.890 ;
        RECT 68.520 123.770 70.855 123.890 ;
        RECT 69.935 123.660 70.855 123.770 ;
        RECT 74.435 123.660 75.365 123.890 ;
        RECT 75.375 123.760 76.745 124.570 ;
        RECT 76.765 123.700 77.195 124.485 ;
        RECT 77.225 123.660 78.575 124.570 ;
        RECT 79.745 123.890 83.645 124.570 ;
        RECT 82.715 123.660 83.645 123.890 ;
        RECT 84.025 123.890 93.305 124.570 ;
        RECT 84.025 123.770 86.360 123.890 ;
        RECT 84.025 123.660 84.945 123.770 ;
        RECT 91.025 123.670 91.945 123.890 ;
        RECT 93.315 123.760 94.685 124.570 ;
        RECT 94.705 123.660 96.055 124.570 ;
        RECT 96.305 123.890 100.205 124.570 ;
        RECT 99.275 123.660 100.205 123.890 ;
        RECT 101.135 123.790 102.505 124.570 ;
        RECT 102.525 123.700 102.955 124.485 ;
        RECT 103.345 123.890 112.625 124.570 ;
        RECT 103.345 123.770 105.680 123.890 ;
        RECT 103.345 123.660 104.265 123.770 ;
        RECT 110.345 123.670 111.265 123.890 ;
        RECT 112.635 123.760 114.465 124.570 ;
        RECT 114.475 123.760 115.845 124.570 ;
      LAYER nwell ;
        RECT 14.460 120.540 116.040 123.370 ;
      LAYER pwell ;
        RECT 14.655 119.340 16.025 120.150 ;
        RECT 16.035 119.340 17.865 120.150 ;
        RECT 17.875 119.340 23.385 120.150 ;
        RECT 24.755 120.020 25.675 120.240 ;
        RECT 31.755 120.140 32.675 120.250 ;
        RECT 30.340 120.020 32.675 120.140 ;
        RECT 23.395 119.340 32.675 120.020 ;
        RECT 33.975 120.020 34.905 120.250 ;
        RECT 33.975 119.340 37.875 120.020 ;
        RECT 38.125 119.425 38.555 120.210 ;
        RECT 39.715 120.160 40.665 120.250 ;
        RECT 38.735 119.340 40.665 120.160 ;
        RECT 41.245 120.140 42.165 120.250 ;
        RECT 41.245 120.020 43.580 120.140 ;
        RECT 48.245 120.020 49.165 120.240 ;
        RECT 50.905 120.140 51.825 120.250 ;
        RECT 50.905 120.020 53.240 120.140 ;
        RECT 57.905 120.020 58.825 120.240 ;
        RECT 41.245 119.340 50.525 120.020 ;
        RECT 50.905 119.340 60.185 120.020 ;
        RECT 60.195 119.340 63.865 120.150 ;
        RECT 63.885 119.425 64.315 120.210 ;
        RECT 64.345 119.340 65.695 120.250 ;
        RECT 66.085 120.140 67.005 120.250 ;
        RECT 66.085 120.020 68.420 120.140 ;
        RECT 73.085 120.020 74.005 120.240 ;
        RECT 77.125 120.140 78.045 120.250 ;
        RECT 66.085 119.340 75.365 120.020 ;
        RECT 75.375 119.340 76.745 120.120 ;
        RECT 77.125 120.020 79.460 120.140 ;
        RECT 84.125 120.020 85.045 120.240 ;
        RECT 77.125 119.340 86.405 120.020 ;
        RECT 86.415 119.340 87.785 120.120 ;
        RECT 87.795 119.340 89.625 120.150 ;
        RECT 89.645 119.425 90.075 120.210 ;
        RECT 92.305 120.140 93.225 120.250 ;
        RECT 90.555 119.340 91.925 120.120 ;
        RECT 92.305 120.020 94.640 120.140 ;
        RECT 99.305 120.020 100.225 120.240 ;
        RECT 92.305 119.340 101.585 120.020 ;
        RECT 102.055 119.340 105.725 120.150 ;
        RECT 105.745 119.340 107.095 120.250 ;
        RECT 107.115 119.340 108.945 120.150 ;
        RECT 108.955 119.340 114.465 120.150 ;
        RECT 114.475 119.340 115.845 120.150 ;
        RECT 14.795 119.130 14.965 119.340 ;
        RECT 17.555 119.150 17.725 119.340 ;
        RECT 19.395 119.130 19.565 119.320 ;
        RECT 23.075 119.150 23.245 119.340 ;
        RECT 23.535 119.150 23.705 119.340 ;
        RECT 24.915 119.130 25.085 119.320 ;
        RECT 26.295 119.175 26.455 119.285 ;
        RECT 31.815 119.130 31.985 119.320 ;
        RECT 33.195 119.130 33.365 119.320 ;
        RECT 33.655 119.185 33.815 119.295 ;
        RECT 34.115 119.175 34.275 119.285 ;
        RECT 34.390 119.150 34.560 119.340 ;
        RECT 38.735 119.320 38.885 119.340 ;
        RECT 37.795 119.130 37.965 119.320 ;
        RECT 38.255 119.130 38.425 119.320 ;
        RECT 38.715 119.150 38.885 119.320 ;
        RECT 39.635 119.130 39.805 119.320 ;
        RECT 41.070 119.180 41.190 119.290 ;
        RECT 43.775 119.130 43.945 119.320 ;
        RECT 44.235 119.130 44.405 119.320 ;
        RECT 45.615 119.130 45.785 119.320 ;
        RECT 47.270 119.130 47.440 119.320 ;
        RECT 50.215 119.150 50.385 119.340 ;
        RECT 51.650 119.180 51.770 119.290 ;
        RECT 55.275 119.130 55.445 119.320 ;
        RECT 55.735 119.130 55.905 119.320 ;
        RECT 58.035 119.130 58.205 119.320 ;
        RECT 59.875 119.150 60.045 119.340 ;
        RECT 61.715 119.130 61.885 119.320 ;
        RECT 63.555 119.150 63.725 119.340 ;
        RECT 64.475 119.150 64.645 119.340 ;
        RECT 67.235 119.130 67.405 119.320 ;
        RECT 68.615 119.130 68.785 119.320 ;
        RECT 69.075 119.130 69.245 119.320 ;
        RECT 70.915 119.175 71.075 119.285 ;
        RECT 75.055 119.150 75.225 119.340 ;
        RECT 76.435 119.130 76.605 119.340 ;
        RECT 77.410 119.180 77.530 119.290 ;
        RECT 80.115 119.130 80.285 119.320 ;
        RECT 81.495 119.130 81.665 119.320 ;
        RECT 83.335 119.130 83.505 119.320 ;
        RECT 83.795 119.130 83.965 119.320 ;
        RECT 86.095 119.150 86.265 119.340 ;
        RECT 87.475 119.130 87.645 119.340 ;
        RECT 89.315 119.150 89.485 119.340 ;
        RECT 90.290 119.180 90.410 119.290 ;
        RECT 90.695 119.150 90.865 119.340 ;
        RECT 92.995 119.130 93.165 119.320 ;
        RECT 98.515 119.130 98.685 119.320 ;
        RECT 99.895 119.130 100.065 119.320 ;
        RECT 100.410 119.180 100.530 119.290 ;
        RECT 101.275 119.150 101.445 119.340 ;
        RECT 101.790 119.180 101.910 119.290 ;
        RECT 102.195 119.130 102.365 119.320 ;
        RECT 104.035 119.130 104.205 119.320 ;
        RECT 105.415 119.150 105.585 119.340 ;
        RECT 105.875 119.150 106.045 119.340 ;
        RECT 107.715 119.130 107.885 119.320 ;
        RECT 108.175 119.130 108.345 119.320 ;
        RECT 108.635 119.150 108.805 119.340 ;
        RECT 114.155 119.320 114.325 119.340 ;
        RECT 110.475 119.130 110.645 119.320 ;
        RECT 111.855 119.130 112.025 119.320 ;
        RECT 112.775 119.175 112.935 119.285 ;
        RECT 114.145 119.150 114.325 119.320 ;
        RECT 114.145 119.130 114.315 119.150 ;
        RECT 115.535 119.130 115.705 119.340 ;
        RECT 14.655 118.320 16.025 119.130 ;
        RECT 16.035 118.320 19.705 119.130 ;
        RECT 19.715 118.320 25.225 119.130 ;
        RECT 25.245 118.260 25.675 119.045 ;
        RECT 26.615 118.320 32.125 119.130 ;
        RECT 32.145 118.220 33.495 119.130 ;
        RECT 34.435 118.320 38.105 119.130 ;
        RECT 38.125 118.220 39.475 119.130 ;
        RECT 39.495 118.350 40.865 119.130 ;
        RECT 41.335 118.320 44.085 119.130 ;
        RECT 44.105 118.220 45.455 119.130 ;
        RECT 45.475 118.350 46.845 119.130 ;
        RECT 46.855 118.450 50.755 119.130 ;
        RECT 46.855 118.220 47.785 118.450 ;
        RECT 51.005 118.260 51.435 119.045 ;
        RECT 51.915 118.320 55.585 119.130 ;
        RECT 55.595 118.350 56.965 119.130 ;
        RECT 56.975 118.320 58.345 119.130 ;
        RECT 58.355 118.320 62.025 119.130 ;
        RECT 62.035 118.320 67.545 119.130 ;
        RECT 67.555 118.350 68.925 119.130 ;
        RECT 68.945 118.220 70.295 119.130 ;
        RECT 71.235 118.320 76.745 119.130 ;
        RECT 76.765 118.260 77.195 119.045 ;
        RECT 77.675 118.320 80.425 119.130 ;
        RECT 80.445 118.220 81.795 119.130 ;
        RECT 81.815 118.320 83.645 119.130 ;
        RECT 83.665 118.220 85.015 119.130 ;
        RECT 85.035 118.320 87.785 119.130 ;
        RECT 87.795 118.320 93.305 119.130 ;
        RECT 93.315 118.320 98.825 119.130 ;
        RECT 98.835 118.350 100.205 119.130 ;
        RECT 100.675 118.320 102.505 119.130 ;
        RECT 102.525 118.260 102.955 119.045 ;
        RECT 102.975 118.320 104.345 119.130 ;
        RECT 104.355 118.320 108.025 119.130 ;
        RECT 108.045 118.220 109.395 119.130 ;
        RECT 109.415 118.350 110.785 119.130 ;
        RECT 110.795 118.350 112.165 119.130 ;
        RECT 113.095 118.350 114.465 119.130 ;
        RECT 114.475 118.320 115.845 119.130 ;
      LAYER nwell ;
        RECT 14.460 115.100 116.040 117.930 ;
      LAYER pwell ;
        RECT 14.655 113.900 16.025 114.710 ;
        RECT 17.155 114.580 19.365 114.810 ;
        RECT 22.085 114.580 23.015 114.800 ;
        RECT 17.155 113.900 27.525 114.580 ;
        RECT 28.005 113.900 29.355 114.810 ;
        RECT 29.375 113.900 30.745 114.680 ;
        RECT 31.215 113.900 32.585 114.680 ;
        RECT 33.055 113.900 34.425 114.680 ;
        RECT 34.435 113.900 38.105 114.710 ;
        RECT 38.125 113.985 38.555 114.770 ;
        RECT 39.035 113.900 41.785 114.710 ;
        RECT 41.795 113.900 47.305 114.710 ;
        RECT 47.315 113.900 48.685 114.680 ;
        RECT 49.155 113.900 51.905 114.710 ;
        RECT 51.915 113.900 57.425 114.710 ;
        RECT 57.435 113.900 60.045 114.810 ;
        RECT 60.195 113.900 63.865 114.710 ;
        RECT 63.885 113.985 64.315 114.770 ;
        RECT 64.795 113.900 68.465 114.710 ;
        RECT 68.485 113.900 69.835 114.810 ;
        RECT 69.855 113.900 71.225 114.680 ;
        RECT 71.245 113.900 72.595 114.810 ;
        RECT 73.535 113.900 76.145 114.810 ;
        RECT 77.215 113.900 80.885 114.710 ;
        RECT 80.895 113.900 86.405 114.710 ;
        RECT 86.415 113.900 87.785 114.680 ;
        RECT 87.795 113.900 89.625 114.710 ;
        RECT 89.645 113.985 90.075 114.770 ;
        RECT 90.095 113.900 91.925 114.710 ;
        RECT 91.935 113.900 93.305 114.680 ;
        RECT 93.315 113.900 96.985 114.710 ;
        RECT 96.995 113.900 98.365 114.680 ;
        RECT 98.835 113.900 100.205 114.680 ;
        RECT 100.215 113.900 101.585 114.680 ;
        RECT 102.055 113.900 103.885 114.710 ;
        RECT 108.405 114.580 109.335 114.800 ;
        RECT 112.055 114.580 114.265 114.810 ;
        RECT 103.895 113.900 114.265 114.580 ;
        RECT 114.475 113.900 115.845 114.710 ;
        RECT 14.795 113.690 14.965 113.900 ;
        RECT 16.635 113.745 16.795 113.855 ;
        RECT 19.395 113.690 19.565 113.880 ;
        RECT 20.775 113.690 20.945 113.880 ;
        RECT 22.155 113.690 22.325 113.880 ;
        RECT 23.535 113.690 23.705 113.880 ;
        RECT 23.995 113.690 24.165 113.880 ;
        RECT 25.890 113.740 26.010 113.850 ;
        RECT 27.215 113.710 27.385 113.900 ;
        RECT 27.730 113.740 27.850 113.850 ;
        RECT 28.135 113.710 28.305 113.900 ;
        RECT 30.435 113.710 30.605 113.900 ;
        RECT 30.950 113.740 31.070 113.850 ;
        RECT 32.275 113.710 32.445 113.900 ;
        RECT 32.790 113.740 32.910 113.850 ;
        RECT 33.195 113.710 33.365 113.900 ;
        RECT 36.415 113.690 36.585 113.880 ;
        RECT 37.335 113.735 37.495 113.845 ;
        RECT 37.795 113.710 37.965 113.900 ;
        RECT 38.715 113.850 38.885 113.880 ;
        RECT 38.715 113.740 38.890 113.850 ;
        RECT 38.715 113.690 38.885 113.740 ;
        RECT 39.175 113.690 39.345 113.880 ;
        RECT 41.475 113.710 41.645 113.900 ;
        RECT 46.995 113.710 47.165 113.900 ;
        RECT 47.455 113.710 47.625 113.900 ;
        RECT 48.890 113.740 49.010 113.850 ;
        RECT 50.675 113.690 50.845 113.880 ;
        RECT 51.595 113.710 51.765 113.900 ;
        RECT 52.055 113.735 52.215 113.845 ;
        RECT 52.515 113.690 52.685 113.880 ;
        RECT 57.115 113.710 57.285 113.900 ;
        RECT 57.580 113.710 57.750 113.900 ;
        RECT 63.555 113.710 63.725 113.900 ;
        RECT 64.015 113.690 64.185 113.880 ;
        RECT 64.475 113.850 64.645 113.880 ;
        RECT 64.475 113.740 64.650 113.850 ;
        RECT 64.475 113.690 64.645 113.740 ;
        RECT 68.155 113.710 68.325 113.900 ;
        RECT 69.535 113.710 69.705 113.900 ;
        RECT 69.995 113.710 70.165 113.900 ;
        RECT 72.295 113.710 72.465 113.900 ;
        RECT 73.215 113.745 73.375 113.855 ;
        RECT 73.680 113.710 73.850 113.900 ;
        RECT 75.975 113.690 76.145 113.880 ;
        RECT 76.490 113.740 76.610 113.850 ;
        RECT 76.895 113.745 77.055 113.855 ;
        RECT 78.275 113.690 78.445 113.880 ;
        RECT 79.195 113.735 79.355 113.845 ;
        RECT 79.655 113.690 79.825 113.880 ;
        RECT 80.575 113.710 80.745 113.900 ;
        RECT 86.095 113.710 86.265 113.900 ;
        RECT 86.555 113.710 86.725 113.900 ;
        RECT 89.315 113.710 89.485 113.900 ;
        RECT 91.155 113.690 91.325 113.880 ;
        RECT 91.615 113.710 91.785 113.900 ;
        RECT 92.075 113.710 92.245 113.900 ;
        RECT 96.675 113.710 96.845 113.900 ;
        RECT 97.135 113.710 97.305 113.900 ;
        RECT 98.570 113.740 98.690 113.850 ;
        RECT 98.975 113.710 99.145 113.900 ;
        RECT 100.355 113.710 100.525 113.900 ;
        RECT 101.735 113.850 101.905 113.880 ;
        RECT 101.735 113.740 101.910 113.850 ;
        RECT 102.250 113.740 102.370 113.850 ;
        RECT 101.735 113.690 101.905 113.740 ;
        RECT 103.115 113.690 103.285 113.880 ;
        RECT 103.575 113.710 103.745 113.900 ;
        RECT 104.035 113.710 104.205 113.900 ;
        RECT 114.155 113.735 114.315 113.845 ;
        RECT 115.535 113.690 115.705 113.900 ;
        RECT 14.655 112.880 16.025 113.690 ;
        RECT 16.035 112.880 19.705 113.690 ;
        RECT 19.725 112.780 21.075 113.690 ;
        RECT 21.105 112.780 22.455 113.690 ;
        RECT 22.485 112.780 23.835 113.690 ;
        RECT 23.855 112.910 25.225 113.690 ;
        RECT 25.245 112.820 25.675 113.605 ;
        RECT 26.355 113.010 36.725 113.690 ;
        RECT 26.355 112.780 28.565 113.010 ;
        RECT 31.285 112.790 32.215 113.010 ;
        RECT 37.655 112.910 39.025 113.690 ;
        RECT 39.035 112.910 40.405 113.690 ;
        RECT 40.615 113.010 50.985 113.690 ;
        RECT 40.615 112.780 42.825 113.010 ;
        RECT 45.545 112.790 46.475 113.010 ;
        RECT 51.005 112.820 51.435 113.605 ;
        RECT 52.375 112.910 53.745 113.690 ;
        RECT 53.955 113.010 64.325 113.690 ;
        RECT 53.955 112.780 56.165 113.010 ;
        RECT 58.885 112.790 59.815 113.010 ;
        RECT 64.335 112.910 65.705 113.690 ;
        RECT 65.915 113.010 76.285 113.690 ;
        RECT 65.915 112.780 68.125 113.010 ;
        RECT 70.845 112.790 71.775 113.010 ;
        RECT 76.765 112.820 77.195 113.605 ;
        RECT 77.215 112.910 78.585 113.690 ;
        RECT 79.515 112.910 80.885 113.690 ;
        RECT 81.095 113.010 91.465 113.690 ;
        RECT 91.675 113.010 102.045 113.690 ;
        RECT 81.095 112.780 83.305 113.010 ;
        RECT 86.025 112.790 86.955 113.010 ;
        RECT 91.675 112.780 93.885 113.010 ;
        RECT 96.605 112.790 97.535 113.010 ;
        RECT 102.525 112.820 102.955 113.605 ;
        RECT 102.975 113.010 113.345 113.690 ;
        RECT 107.485 112.790 108.415 113.010 ;
        RECT 111.135 112.780 113.345 113.010 ;
        RECT 114.475 112.880 115.845 113.690 ;
      LAYER nwell ;
        RECT 14.460 109.660 116.040 112.490 ;
      LAYER pwell ;
        RECT 14.655 108.460 16.025 109.270 ;
        RECT 17.155 109.140 19.365 109.370 ;
        RECT 22.085 109.140 23.015 109.360 ;
        RECT 27.735 109.140 29.945 109.370 ;
        RECT 32.665 109.140 33.595 109.360 ;
        RECT 17.155 108.460 27.525 109.140 ;
        RECT 27.735 108.460 38.105 109.140 ;
        RECT 38.125 108.545 38.555 109.330 ;
        RECT 38.585 108.460 39.935 109.370 ;
        RECT 40.885 108.460 42.235 109.370 ;
        RECT 43.175 108.460 46.845 109.270 ;
        RECT 46.865 108.460 48.215 109.370 ;
        RECT 48.435 109.140 50.645 109.370 ;
        RECT 53.365 109.140 54.295 109.360 ;
        RECT 48.435 108.460 58.805 109.140 ;
        RECT 59.735 108.460 61.105 109.240 ;
        RECT 61.125 108.460 62.475 109.370 ;
        RECT 62.495 108.460 63.865 109.270 ;
        RECT 63.885 108.545 64.315 109.330 ;
        RECT 64.535 109.140 66.745 109.370 ;
        RECT 69.465 109.140 70.395 109.360 ;
        RECT 76.035 109.140 78.245 109.370 ;
        RECT 80.965 109.140 81.895 109.360 ;
        RECT 64.535 108.460 74.905 109.140 ;
        RECT 76.035 108.460 86.405 109.140 ;
        RECT 86.425 108.460 87.775 109.370 ;
        RECT 88.265 108.460 89.615 109.370 ;
        RECT 89.645 108.545 90.075 109.330 ;
        RECT 90.295 109.140 92.505 109.370 ;
        RECT 95.225 109.140 96.155 109.360 ;
        RECT 100.875 109.140 103.085 109.370 ;
        RECT 105.805 109.140 106.735 109.360 ;
        RECT 90.295 108.460 100.665 109.140 ;
        RECT 100.875 108.460 111.245 109.140 ;
        RECT 111.265 108.460 112.615 109.370 ;
        RECT 112.645 108.460 113.995 109.370 ;
        RECT 114.475 108.460 115.845 109.270 ;
        RECT 14.795 108.250 14.965 108.460 ;
        RECT 16.635 108.305 16.795 108.415 ;
        RECT 19.395 108.250 19.565 108.440 ;
        RECT 24.915 108.250 25.085 108.440 ;
        RECT 27.215 108.270 27.385 108.460 ;
        RECT 35.955 108.250 36.125 108.440 ;
        RECT 37.795 108.250 37.965 108.460 ;
        RECT 39.635 108.270 39.805 108.460 ;
        RECT 40.555 108.305 40.715 108.415 ;
        RECT 41.015 108.270 41.185 108.460 ;
        RECT 42.855 108.305 43.015 108.415 ;
        RECT 46.535 108.270 46.705 108.460 ;
        RECT 47.915 108.270 48.085 108.460 ;
        RECT 48.835 108.250 49.005 108.440 ;
        RECT 50.675 108.250 50.845 108.440 ;
        RECT 52.515 108.250 52.685 108.440 ;
        RECT 53.895 108.250 54.065 108.440 ;
        RECT 57.575 108.250 57.745 108.440 ;
        RECT 58.495 108.270 58.665 108.460 ;
        RECT 58.955 108.250 59.125 108.440 ;
        RECT 59.415 108.305 59.575 108.415 ;
        RECT 59.875 108.270 60.045 108.460 ;
        RECT 61.255 108.270 61.425 108.460 ;
        RECT 63.555 108.250 63.725 108.460 ;
        RECT 65.855 108.250 66.025 108.440 ;
        RECT 74.595 108.270 74.765 108.460 ;
        RECT 75.515 108.305 75.675 108.415 ;
        RECT 76.435 108.250 76.605 108.440 ;
        RECT 78.275 108.250 78.445 108.440 ;
        RECT 79.655 108.250 79.825 108.440 ;
        RECT 81.035 108.250 81.205 108.440 ;
        RECT 83.795 108.250 83.965 108.440 ;
        RECT 86.095 108.270 86.265 108.460 ;
        RECT 87.475 108.270 87.645 108.460 ;
        RECT 87.990 108.300 88.110 108.410 ;
        RECT 88.395 108.270 88.565 108.460 ;
        RECT 89.315 108.250 89.485 108.440 ;
        RECT 95.295 108.250 95.465 108.440 ;
        RECT 96.675 108.250 96.845 108.440 ;
        RECT 97.190 108.300 97.310 108.410 ;
        RECT 99.895 108.250 100.065 108.440 ;
        RECT 100.355 108.250 100.525 108.460 ;
        RECT 102.195 108.295 102.355 108.405 ;
        RECT 103.575 108.295 103.735 108.405 ;
        RECT 104.035 108.250 104.205 108.440 ;
        RECT 110.935 108.270 111.105 108.460 ;
        RECT 112.315 108.270 112.485 108.460 ;
        RECT 112.775 108.270 112.945 108.460 ;
        RECT 114.210 108.300 114.330 108.410 ;
        RECT 115.535 108.250 115.705 108.460 ;
        RECT 14.655 107.440 16.025 108.250 ;
        RECT 16.035 107.440 19.705 108.250 ;
        RECT 19.715 107.440 25.225 108.250 ;
        RECT 25.245 107.380 25.675 108.165 ;
        RECT 25.895 107.570 36.265 108.250 ;
        RECT 25.895 107.340 28.105 107.570 ;
        RECT 30.825 107.350 31.755 107.570 ;
        RECT 36.275 107.440 38.105 108.250 ;
        RECT 38.125 107.380 38.555 108.165 ;
        RECT 38.775 107.570 49.145 108.250 ;
        RECT 38.775 107.340 40.985 107.570 ;
        RECT 43.705 107.350 44.635 107.570 ;
        RECT 49.155 107.440 50.985 108.250 ;
        RECT 51.005 107.380 51.435 108.165 ;
        RECT 51.455 107.440 52.825 108.250 ;
        RECT 52.845 107.340 54.195 108.250 ;
        RECT 54.215 107.440 57.885 108.250 ;
        RECT 57.905 107.340 59.255 108.250 ;
        RECT 60.195 107.440 63.865 108.250 ;
        RECT 63.885 107.380 64.315 108.165 ;
        RECT 64.335 107.440 66.165 108.250 ;
        RECT 66.375 107.570 76.745 108.250 ;
        RECT 66.375 107.340 68.585 107.570 ;
        RECT 71.305 107.350 72.235 107.570 ;
        RECT 76.765 107.380 77.195 108.165 ;
        RECT 77.225 107.340 78.575 108.250 ;
        RECT 78.595 107.440 79.965 108.250 ;
        RECT 79.985 107.340 81.335 108.250 ;
        RECT 81.355 107.440 84.105 108.250 ;
        RECT 84.115 107.440 89.625 108.250 ;
        RECT 89.645 107.380 90.075 108.165 ;
        RECT 90.095 107.440 95.605 108.250 ;
        RECT 95.625 107.340 96.975 108.250 ;
        RECT 97.455 107.440 100.205 108.250 ;
        RECT 100.225 107.340 101.575 108.250 ;
        RECT 102.525 107.380 102.955 108.165 ;
        RECT 103.895 107.570 114.265 108.250 ;
        RECT 108.405 107.350 109.335 107.570 ;
        RECT 112.055 107.340 114.265 107.570 ;
        RECT 114.475 107.440 115.845 108.250 ;
      LAYER nwell ;
        RECT 14.460 105.445 116.040 107.050 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 14.650 206.190 115.850 206.360 ;
        RECT 14.735 205.440 15.945 206.190 ;
        RECT 14.735 204.900 15.255 205.440 ;
        RECT 16.115 205.420 19.625 206.190 ;
        RECT 19.800 205.645 25.145 206.190 ;
        RECT 15.425 204.730 15.945 205.270 ;
        RECT 14.735 203.640 15.945 204.730 ;
        RECT 16.115 204.730 17.805 205.250 ;
        RECT 17.975 204.900 19.625 205.420 ;
        RECT 16.115 203.640 19.625 204.730 ;
        RECT 21.390 204.075 21.740 205.325 ;
        RECT 23.220 204.815 23.560 205.645 ;
        RECT 25.315 205.465 25.605 206.190 ;
        RECT 25.775 205.440 26.985 206.190 ;
        RECT 27.160 205.645 32.505 206.190 ;
        RECT 32.680 205.645 38.025 206.190 ;
        RECT 19.800 203.640 25.145 204.075 ;
        RECT 25.315 203.640 25.605 204.805 ;
        RECT 25.775 204.730 26.295 205.270 ;
        RECT 26.465 204.900 26.985 205.440 ;
        RECT 25.775 203.640 26.985 204.730 ;
        RECT 28.750 204.075 29.100 205.325 ;
        RECT 30.580 204.815 30.920 205.645 ;
        RECT 34.270 204.075 34.620 205.325 ;
        RECT 36.100 204.815 36.440 205.645 ;
        RECT 38.195 205.465 38.485 206.190 ;
        RECT 38.655 205.440 39.865 206.190 ;
        RECT 40.040 205.645 45.385 206.190 ;
        RECT 45.560 205.645 50.905 206.190 ;
        RECT 27.160 203.640 32.505 204.075 ;
        RECT 32.680 203.640 38.025 204.075 ;
        RECT 38.195 203.640 38.485 204.805 ;
        RECT 38.655 204.730 39.175 205.270 ;
        RECT 39.345 204.900 39.865 205.440 ;
        RECT 38.655 203.640 39.865 204.730 ;
        RECT 41.630 204.075 41.980 205.325 ;
        RECT 43.460 204.815 43.800 205.645 ;
        RECT 47.150 204.075 47.500 205.325 ;
        RECT 48.980 204.815 49.320 205.645 ;
        RECT 51.075 205.465 51.365 206.190 ;
        RECT 51.535 205.440 52.745 206.190 ;
        RECT 52.920 205.645 58.265 206.190 ;
        RECT 58.440 205.645 63.785 206.190 ;
        RECT 40.040 203.640 45.385 204.075 ;
        RECT 45.560 203.640 50.905 204.075 ;
        RECT 51.075 203.640 51.365 204.805 ;
        RECT 51.535 204.730 52.055 205.270 ;
        RECT 52.225 204.900 52.745 205.440 ;
        RECT 51.535 203.640 52.745 204.730 ;
        RECT 54.510 204.075 54.860 205.325 ;
        RECT 56.340 204.815 56.680 205.645 ;
        RECT 60.030 204.075 60.380 205.325 ;
        RECT 61.860 204.815 62.200 205.645 ;
        RECT 63.955 205.465 64.245 206.190 ;
        RECT 64.415 205.440 65.625 206.190 ;
        RECT 65.800 205.645 71.145 206.190 ;
        RECT 71.320 205.645 76.665 206.190 ;
        RECT 52.920 203.640 58.265 204.075 ;
        RECT 58.440 203.640 63.785 204.075 ;
        RECT 63.955 203.640 64.245 204.805 ;
        RECT 64.415 204.730 64.935 205.270 ;
        RECT 65.105 204.900 65.625 205.440 ;
        RECT 64.415 203.640 65.625 204.730 ;
        RECT 67.390 204.075 67.740 205.325 ;
        RECT 69.220 204.815 69.560 205.645 ;
        RECT 72.910 204.075 73.260 205.325 ;
        RECT 74.740 204.815 75.080 205.645 ;
        RECT 76.835 205.465 77.125 206.190 ;
        RECT 77.295 205.440 78.505 206.190 ;
        RECT 78.680 205.645 84.025 206.190 ;
        RECT 84.200 205.645 89.545 206.190 ;
        RECT 65.800 203.640 71.145 204.075 ;
        RECT 71.320 203.640 76.665 204.075 ;
        RECT 76.835 203.640 77.125 204.805 ;
        RECT 77.295 204.730 77.815 205.270 ;
        RECT 77.985 204.900 78.505 205.440 ;
        RECT 77.295 203.640 78.505 204.730 ;
        RECT 80.270 204.075 80.620 205.325 ;
        RECT 82.100 204.815 82.440 205.645 ;
        RECT 85.790 204.075 86.140 205.325 ;
        RECT 87.620 204.815 87.960 205.645 ;
        RECT 89.715 205.465 90.005 206.190 ;
        RECT 90.175 205.440 91.385 206.190 ;
        RECT 91.560 205.645 96.905 206.190 ;
        RECT 97.080 205.645 102.425 206.190 ;
        RECT 78.680 203.640 84.025 204.075 ;
        RECT 84.200 203.640 89.545 204.075 ;
        RECT 89.715 203.640 90.005 204.805 ;
        RECT 90.175 204.730 90.695 205.270 ;
        RECT 90.865 204.900 91.385 205.440 ;
        RECT 90.175 203.640 91.385 204.730 ;
        RECT 93.150 204.075 93.500 205.325 ;
        RECT 94.980 204.815 95.320 205.645 ;
        RECT 98.670 204.075 99.020 205.325 ;
        RECT 100.500 204.815 100.840 205.645 ;
        RECT 102.595 205.465 102.885 206.190 ;
        RECT 103.520 205.645 108.865 206.190 ;
        RECT 109.040 205.645 114.385 206.190 ;
        RECT 91.560 203.640 96.905 204.075 ;
        RECT 97.080 203.640 102.425 204.075 ;
        RECT 102.595 203.640 102.885 204.805 ;
        RECT 105.110 204.075 105.460 205.325 ;
        RECT 106.940 204.815 107.280 205.645 ;
        RECT 110.630 204.075 110.980 205.325 ;
        RECT 112.460 204.815 112.800 205.645 ;
        RECT 114.555 205.440 115.765 206.190 ;
        RECT 114.555 204.730 115.075 205.270 ;
        RECT 115.245 204.900 115.765 205.440 ;
        RECT 103.520 203.640 108.865 204.075 ;
        RECT 109.040 203.640 114.385 204.075 ;
        RECT 114.555 203.640 115.765 204.730 ;
        RECT 14.650 203.470 115.850 203.640 ;
        RECT 14.735 202.380 15.945 203.470 ;
        RECT 16.120 203.035 21.465 203.470 ;
        RECT 21.640 203.035 26.985 203.470 ;
        RECT 27.160 203.035 32.505 203.470 ;
        RECT 32.680 203.035 38.025 203.470 ;
        RECT 14.735 201.670 15.255 202.210 ;
        RECT 15.425 201.840 15.945 202.380 ;
        RECT 17.710 201.785 18.060 203.035 ;
        RECT 14.735 200.920 15.945 201.670 ;
        RECT 19.540 201.465 19.880 202.295 ;
        RECT 23.230 201.785 23.580 203.035 ;
        RECT 25.060 201.465 25.400 202.295 ;
        RECT 28.750 201.785 29.100 203.035 ;
        RECT 30.580 201.465 30.920 202.295 ;
        RECT 34.270 201.785 34.620 203.035 ;
        RECT 38.195 202.305 38.485 203.470 ;
        RECT 38.660 203.035 44.005 203.470 ;
        RECT 44.180 203.035 49.525 203.470 ;
        RECT 49.700 203.035 55.045 203.470 ;
        RECT 55.220 203.035 60.565 203.470 ;
        RECT 36.100 201.465 36.440 202.295 ;
        RECT 40.250 201.785 40.600 203.035 ;
        RECT 16.120 200.920 21.465 201.465 ;
        RECT 21.640 200.920 26.985 201.465 ;
        RECT 27.160 200.920 32.505 201.465 ;
        RECT 32.680 200.920 38.025 201.465 ;
        RECT 38.195 200.920 38.485 201.645 ;
        RECT 42.080 201.465 42.420 202.295 ;
        RECT 45.770 201.785 46.120 203.035 ;
        RECT 47.600 201.465 47.940 202.295 ;
        RECT 51.290 201.785 51.640 203.035 ;
        RECT 53.120 201.465 53.460 202.295 ;
        RECT 56.810 201.785 57.160 203.035 ;
        RECT 60.775 202.330 61.005 203.470 ;
        RECT 61.175 202.320 61.505 203.300 ;
        RECT 61.675 202.330 61.885 203.470 ;
        RECT 62.205 202.540 62.375 203.300 ;
        RECT 62.590 202.710 62.920 203.470 ;
        RECT 62.205 202.370 62.920 202.540 ;
        RECT 63.090 202.395 63.345 203.300 ;
        RECT 58.640 201.465 58.980 202.295 ;
        RECT 60.755 201.910 61.085 202.160 ;
        RECT 38.660 200.920 44.005 201.465 ;
        RECT 44.180 200.920 49.525 201.465 ;
        RECT 49.700 200.920 55.045 201.465 ;
        RECT 55.220 200.920 60.565 201.465 ;
        RECT 60.775 200.920 61.005 201.740 ;
        RECT 61.255 201.720 61.505 202.320 ;
        RECT 62.115 201.820 62.470 202.190 ;
        RECT 62.750 202.160 62.920 202.370 ;
        RECT 62.750 201.830 63.005 202.160 ;
        RECT 61.175 201.090 61.505 201.720 ;
        RECT 61.675 200.920 61.885 201.740 ;
        RECT 62.750 201.640 62.920 201.830 ;
        RECT 63.175 201.665 63.345 202.395 ;
        RECT 63.520 202.320 63.780 203.470 ;
        RECT 63.955 202.305 64.245 203.470 ;
        RECT 64.415 202.395 64.685 203.300 ;
        RECT 64.855 202.710 65.185 203.470 ;
        RECT 65.365 202.540 65.535 203.300 ;
        RECT 66.260 203.045 66.595 203.470 ;
        RECT 66.765 202.865 66.950 203.270 ;
        RECT 62.205 201.470 62.920 201.640 ;
        RECT 62.205 201.090 62.375 201.470 ;
        RECT 62.590 200.920 62.920 201.300 ;
        RECT 63.090 201.090 63.345 201.665 ;
        RECT 63.520 200.920 63.780 201.760 ;
        RECT 63.955 200.920 64.245 201.645 ;
        RECT 64.415 201.595 64.585 202.395 ;
        RECT 64.870 202.370 65.535 202.540 ;
        RECT 66.285 202.690 66.950 202.865 ;
        RECT 67.155 202.690 67.485 203.470 ;
        RECT 64.870 202.225 65.040 202.370 ;
        RECT 64.755 201.895 65.040 202.225 ;
        RECT 64.870 201.640 65.040 201.895 ;
        RECT 65.275 201.820 65.605 202.190 ;
        RECT 66.285 201.660 66.625 202.690 ;
        RECT 67.655 202.500 67.925 203.270 ;
        RECT 66.795 202.330 67.925 202.500 ;
        RECT 66.795 201.830 67.045 202.330 ;
        RECT 64.415 201.090 64.675 201.595 ;
        RECT 64.870 201.470 65.535 201.640 ;
        RECT 66.285 201.490 66.970 201.660 ;
        RECT 67.225 201.580 67.585 202.160 ;
        RECT 64.855 200.920 65.185 201.300 ;
        RECT 65.365 201.090 65.535 201.470 ;
        RECT 66.260 200.920 66.595 201.320 ;
        RECT 66.765 201.090 66.970 201.490 ;
        RECT 67.755 201.420 67.925 202.330 ;
        RECT 68.555 202.380 70.225 203.470 ;
        RECT 68.555 201.860 69.305 202.380 ;
        RECT 70.400 202.280 70.655 203.160 ;
        RECT 70.825 202.330 71.130 203.470 ;
        RECT 71.470 203.090 71.800 203.470 ;
        RECT 71.980 202.920 72.150 203.210 ;
        RECT 72.320 203.010 72.570 203.470 ;
        RECT 71.350 202.750 72.150 202.920 ;
        RECT 72.740 202.960 73.610 203.300 ;
        RECT 69.475 201.690 70.225 202.210 ;
        RECT 67.180 200.920 67.455 201.400 ;
        RECT 67.665 201.090 67.925 201.420 ;
        RECT 68.555 200.920 70.225 201.690 ;
        RECT 70.400 201.630 70.610 202.280 ;
        RECT 71.350 202.160 71.520 202.750 ;
        RECT 72.740 202.580 72.910 202.960 ;
        RECT 73.845 202.840 74.015 203.300 ;
        RECT 74.185 203.010 74.555 203.470 ;
        RECT 74.850 202.870 75.020 203.210 ;
        RECT 75.190 203.040 75.520 203.470 ;
        RECT 75.755 202.870 75.925 203.210 ;
        RECT 71.690 202.410 72.910 202.580 ;
        RECT 73.080 202.500 73.540 202.790 ;
        RECT 73.845 202.670 74.405 202.840 ;
        RECT 74.850 202.700 75.925 202.870 ;
        RECT 76.095 202.970 76.775 203.300 ;
        RECT 76.990 202.970 77.240 203.300 ;
        RECT 77.410 203.010 77.660 203.470 ;
        RECT 74.235 202.530 74.405 202.670 ;
        RECT 73.080 202.490 74.045 202.500 ;
        RECT 72.740 202.320 72.910 202.410 ;
        RECT 73.370 202.330 74.045 202.490 ;
        RECT 70.780 202.130 71.520 202.160 ;
        RECT 70.780 201.830 71.695 202.130 ;
        RECT 71.370 201.655 71.695 201.830 ;
        RECT 70.400 201.100 70.655 201.630 ;
        RECT 70.825 200.920 71.130 201.380 ;
        RECT 71.375 201.300 71.695 201.655 ;
        RECT 71.865 201.870 72.405 202.240 ;
        RECT 72.740 202.150 73.145 202.320 ;
        RECT 71.865 201.470 72.105 201.870 ;
        RECT 72.585 201.700 72.805 201.980 ;
        RECT 72.275 201.530 72.805 201.700 ;
        RECT 72.275 201.300 72.445 201.530 ;
        RECT 72.975 201.370 73.145 202.150 ;
        RECT 73.315 201.540 73.665 202.160 ;
        RECT 73.835 201.540 74.045 202.330 ;
        RECT 74.235 202.360 75.735 202.530 ;
        RECT 74.235 201.670 74.405 202.360 ;
        RECT 76.095 202.190 76.265 202.970 ;
        RECT 77.070 202.840 77.240 202.970 ;
        RECT 74.575 202.020 76.265 202.190 ;
        RECT 76.435 202.410 76.900 202.800 ;
        RECT 77.070 202.670 77.465 202.840 ;
        RECT 74.575 201.840 74.745 202.020 ;
        RECT 71.375 201.130 72.445 201.300 ;
        RECT 72.615 200.920 72.805 201.360 ;
        RECT 72.975 201.090 73.925 201.370 ;
        RECT 74.235 201.280 74.495 201.670 ;
        RECT 74.915 201.600 75.705 201.850 ;
        RECT 74.145 201.110 74.495 201.280 ;
        RECT 74.705 200.920 75.035 201.380 ;
        RECT 75.910 201.310 76.080 202.020 ;
        RECT 76.435 201.820 76.605 202.410 ;
        RECT 76.250 201.600 76.605 201.820 ;
        RECT 76.775 201.600 77.125 202.220 ;
        RECT 77.295 201.310 77.465 202.670 ;
        RECT 77.830 202.500 78.155 203.285 ;
        RECT 77.635 201.450 78.095 202.500 ;
        RECT 75.910 201.140 76.765 201.310 ;
        RECT 76.970 201.140 77.465 201.310 ;
        RECT 77.635 200.920 77.965 201.280 ;
        RECT 78.325 201.180 78.495 203.300 ;
        RECT 78.665 202.970 78.995 203.470 ;
        RECT 79.165 202.800 79.420 203.300 ;
        RECT 78.670 202.630 79.420 202.800 ;
        RECT 78.670 201.640 78.900 202.630 ;
        RECT 79.070 201.810 79.420 202.460 ;
        RECT 80.515 202.380 84.025 203.470 ;
        RECT 84.200 203.035 89.545 203.470 ;
        RECT 80.515 201.860 82.205 202.380 ;
        RECT 82.375 201.690 84.025 202.210 ;
        RECT 85.790 201.785 86.140 203.035 ;
        RECT 89.715 202.305 90.005 203.470 ;
        RECT 90.635 202.380 92.305 203.470 ;
        RECT 92.480 203.035 97.825 203.470 ;
        RECT 98.000 203.035 103.345 203.470 ;
        RECT 103.520 203.035 108.865 203.470 ;
        RECT 109.040 203.035 114.385 203.470 ;
        RECT 78.670 201.470 79.420 201.640 ;
        RECT 78.665 200.920 78.995 201.300 ;
        RECT 79.165 201.180 79.420 201.470 ;
        RECT 80.515 200.920 84.025 201.690 ;
        RECT 87.620 201.465 87.960 202.295 ;
        RECT 90.635 201.860 91.385 202.380 ;
        RECT 91.555 201.690 92.305 202.210 ;
        RECT 94.070 201.785 94.420 203.035 ;
        RECT 84.200 200.920 89.545 201.465 ;
        RECT 89.715 200.920 90.005 201.645 ;
        RECT 90.635 200.920 92.305 201.690 ;
        RECT 95.900 201.465 96.240 202.295 ;
        RECT 99.590 201.785 99.940 203.035 ;
        RECT 101.420 201.465 101.760 202.295 ;
        RECT 105.110 201.785 105.460 203.035 ;
        RECT 106.940 201.465 107.280 202.295 ;
        RECT 110.630 201.785 110.980 203.035 ;
        RECT 114.555 202.380 115.765 203.470 ;
        RECT 112.460 201.465 112.800 202.295 ;
        RECT 114.555 201.840 115.075 202.380 ;
        RECT 115.245 201.670 115.765 202.210 ;
        RECT 92.480 200.920 97.825 201.465 ;
        RECT 98.000 200.920 103.345 201.465 ;
        RECT 103.520 200.920 108.865 201.465 ;
        RECT 109.040 200.920 114.385 201.465 ;
        RECT 114.555 200.920 115.765 201.670 ;
        RECT 14.650 200.750 115.850 200.920 ;
        RECT 14.735 200.000 15.945 200.750 ;
        RECT 14.735 199.460 15.255 200.000 ;
        RECT 16.115 199.980 19.625 200.750 ;
        RECT 19.800 200.205 25.145 200.750 ;
        RECT 15.425 199.290 15.945 199.830 ;
        RECT 14.735 198.200 15.945 199.290 ;
        RECT 16.115 199.290 17.805 199.810 ;
        RECT 17.975 199.460 19.625 199.980 ;
        RECT 16.115 198.200 19.625 199.290 ;
        RECT 21.390 198.635 21.740 199.885 ;
        RECT 23.220 199.375 23.560 200.205 ;
        RECT 25.315 200.025 25.605 200.750 ;
        RECT 26.235 199.980 28.825 200.750 ;
        RECT 29.000 200.205 34.345 200.750 ;
        RECT 34.520 200.205 39.865 200.750 ;
        RECT 40.040 200.205 45.385 200.750 ;
        RECT 45.560 200.205 50.905 200.750 ;
        RECT 19.800 198.200 25.145 198.635 ;
        RECT 25.315 198.200 25.605 199.365 ;
        RECT 26.235 199.290 27.445 199.810 ;
        RECT 27.615 199.460 28.825 199.980 ;
        RECT 26.235 198.200 28.825 199.290 ;
        RECT 30.590 198.635 30.940 199.885 ;
        RECT 32.420 199.375 32.760 200.205 ;
        RECT 36.110 198.635 36.460 199.885 ;
        RECT 37.940 199.375 38.280 200.205 ;
        RECT 41.630 198.635 41.980 199.885 ;
        RECT 43.460 199.375 43.800 200.205 ;
        RECT 47.150 198.635 47.500 199.885 ;
        RECT 48.980 199.375 49.320 200.205 ;
        RECT 51.075 200.025 51.365 200.750 ;
        RECT 52.460 200.205 57.805 200.750 ;
        RECT 29.000 198.200 34.345 198.635 ;
        RECT 34.520 198.200 39.865 198.635 ;
        RECT 40.040 198.200 45.385 198.635 ;
        RECT 45.560 198.200 50.905 198.635 ;
        RECT 51.075 198.200 51.365 199.365 ;
        RECT 54.050 198.635 54.400 199.885 ;
        RECT 55.880 199.375 56.220 200.205 ;
        RECT 58.035 199.930 58.245 200.750 ;
        RECT 58.415 199.950 58.745 200.580 ;
        RECT 58.415 199.350 58.665 199.950 ;
        RECT 58.915 199.930 59.145 200.750 ;
        RECT 59.360 200.040 59.615 200.570 ;
        RECT 59.785 200.290 60.090 200.750 ;
        RECT 60.335 200.370 61.405 200.540 ;
        RECT 58.835 199.510 59.165 199.760 ;
        RECT 59.360 199.390 59.570 200.040 ;
        RECT 60.335 200.015 60.655 200.370 ;
        RECT 60.330 199.840 60.655 200.015 ;
        RECT 59.740 199.540 60.655 199.840 ;
        RECT 60.825 199.800 61.065 200.200 ;
        RECT 61.235 200.140 61.405 200.370 ;
        RECT 61.575 200.310 61.765 200.750 ;
        RECT 61.935 200.300 62.885 200.580 ;
        RECT 63.105 200.390 63.455 200.560 ;
        RECT 61.235 199.970 61.765 200.140 ;
        RECT 59.740 199.510 60.480 199.540 ;
        RECT 52.460 198.200 57.805 198.635 ;
        RECT 58.035 198.200 58.245 199.340 ;
        RECT 58.415 198.370 58.745 199.350 ;
        RECT 58.915 198.200 59.145 199.340 ;
        RECT 59.360 198.510 59.615 199.390 ;
        RECT 59.785 198.200 60.090 199.340 ;
        RECT 60.310 198.920 60.480 199.510 ;
        RECT 60.825 199.430 61.365 199.800 ;
        RECT 61.545 199.690 61.765 199.970 ;
        RECT 61.935 199.520 62.105 200.300 ;
        RECT 61.700 199.350 62.105 199.520 ;
        RECT 62.275 199.510 62.625 200.130 ;
        RECT 61.700 199.260 61.870 199.350 ;
        RECT 62.795 199.340 63.005 200.130 ;
        RECT 60.650 199.090 61.870 199.260 ;
        RECT 62.330 199.180 63.005 199.340 ;
        RECT 60.310 198.750 61.110 198.920 ;
        RECT 60.430 198.200 60.760 198.580 ;
        RECT 60.940 198.460 61.110 198.750 ;
        RECT 61.700 198.710 61.870 199.090 ;
        RECT 62.040 199.170 63.005 199.180 ;
        RECT 63.195 200.000 63.455 200.390 ;
        RECT 63.665 200.290 63.995 200.750 ;
        RECT 64.870 200.360 65.725 200.530 ;
        RECT 65.930 200.360 66.425 200.530 ;
        RECT 66.595 200.390 66.925 200.750 ;
        RECT 63.195 199.310 63.365 200.000 ;
        RECT 63.535 199.650 63.705 199.830 ;
        RECT 63.875 199.820 64.665 200.070 ;
        RECT 64.870 199.650 65.040 200.360 ;
        RECT 65.210 199.850 65.565 200.070 ;
        RECT 63.535 199.480 65.225 199.650 ;
        RECT 62.040 198.880 62.500 199.170 ;
        RECT 63.195 199.140 64.695 199.310 ;
        RECT 63.195 199.000 63.365 199.140 ;
        RECT 62.805 198.830 63.365 199.000 ;
        RECT 61.280 198.200 61.530 198.660 ;
        RECT 61.700 198.370 62.570 198.710 ;
        RECT 62.805 198.370 62.975 198.830 ;
        RECT 63.810 198.800 64.885 198.970 ;
        RECT 63.145 198.200 63.515 198.660 ;
        RECT 63.810 198.460 63.980 198.800 ;
        RECT 64.150 198.200 64.480 198.630 ;
        RECT 64.715 198.460 64.885 198.800 ;
        RECT 65.055 198.700 65.225 199.480 ;
        RECT 65.395 199.260 65.565 199.850 ;
        RECT 65.735 199.450 66.085 200.070 ;
        RECT 65.395 198.870 65.860 199.260 ;
        RECT 66.255 199.000 66.425 200.360 ;
        RECT 66.595 199.170 67.055 200.220 ;
        RECT 66.030 198.830 66.425 199.000 ;
        RECT 66.030 198.700 66.200 198.830 ;
        RECT 65.055 198.370 65.735 198.700 ;
        RECT 65.950 198.370 66.200 198.700 ;
        RECT 66.370 198.200 66.620 198.660 ;
        RECT 66.790 198.385 67.115 199.170 ;
        RECT 67.285 198.370 67.455 200.490 ;
        RECT 67.625 200.370 67.955 200.750 ;
        RECT 68.125 200.200 68.380 200.490 ;
        RECT 67.630 200.030 68.380 200.200 ;
        RECT 67.630 199.040 67.860 200.030 ;
        RECT 69.475 200.010 69.795 200.490 ;
        RECT 69.965 200.180 70.195 200.580 ;
        RECT 70.365 200.360 70.715 200.750 ;
        RECT 69.965 200.100 70.475 200.180 ;
        RECT 70.885 200.100 71.215 200.580 ;
        RECT 69.965 200.010 71.215 200.100 ;
        RECT 68.030 199.210 68.380 199.860 ;
        RECT 69.475 199.080 69.645 200.010 ;
        RECT 70.305 199.930 71.215 200.010 ;
        RECT 71.385 199.930 71.555 200.750 ;
        RECT 72.060 200.010 72.525 200.555 ;
        RECT 72.860 200.240 73.100 200.750 ;
        RECT 73.280 200.240 73.560 200.570 ;
        RECT 73.790 200.240 74.005 200.750 ;
        RECT 69.815 199.420 69.985 199.840 ;
        RECT 70.215 199.590 70.815 199.760 ;
        RECT 69.815 199.250 70.475 199.420 ;
        RECT 67.630 198.870 68.380 199.040 ;
        RECT 69.475 198.880 70.135 199.080 ;
        RECT 70.305 199.050 70.475 199.250 ;
        RECT 70.645 199.390 70.815 199.590 ;
        RECT 70.985 199.560 71.680 199.760 ;
        RECT 71.940 199.390 72.185 199.840 ;
        RECT 70.645 199.220 72.185 199.390 ;
        RECT 72.355 199.050 72.525 200.010 ;
        RECT 72.755 199.510 73.110 200.070 ;
        RECT 73.280 199.340 73.450 200.240 ;
        RECT 73.620 199.510 73.885 200.070 ;
        RECT 74.175 200.010 74.790 200.580 ;
        RECT 75.085 200.200 75.255 200.580 ;
        RECT 75.435 200.370 75.765 200.750 ;
        RECT 75.085 200.030 75.750 200.200 ;
        RECT 75.945 200.075 76.205 200.580 ;
        RECT 74.135 199.340 74.305 199.840 ;
        RECT 70.305 198.880 72.525 199.050 ;
        RECT 72.880 199.170 74.305 199.340 ;
        RECT 72.880 198.995 73.270 199.170 ;
        RECT 67.625 198.200 67.955 198.700 ;
        RECT 68.125 198.370 68.380 198.870 ;
        RECT 69.965 198.710 70.135 198.880 ;
        RECT 69.495 198.200 69.795 198.710 ;
        RECT 69.965 198.540 70.345 198.710 ;
        RECT 70.925 198.200 71.555 198.710 ;
        RECT 71.725 198.370 72.055 198.880 ;
        RECT 72.225 198.200 72.525 198.710 ;
        RECT 73.755 198.200 74.085 199.000 ;
        RECT 74.475 198.990 74.790 200.010 ;
        RECT 75.015 199.480 75.345 199.850 ;
        RECT 75.580 199.775 75.750 200.030 ;
        RECT 75.580 199.445 75.865 199.775 ;
        RECT 75.580 199.300 75.750 199.445 ;
        RECT 74.255 198.370 74.790 198.990 ;
        RECT 75.085 199.130 75.750 199.300 ;
        RECT 76.035 199.275 76.205 200.075 ;
        RECT 76.835 200.025 77.125 200.750 ;
        RECT 77.295 200.100 77.555 200.580 ;
        RECT 77.725 200.210 77.975 200.750 ;
        RECT 75.085 198.370 75.255 199.130 ;
        RECT 75.435 198.200 75.765 198.960 ;
        RECT 75.935 198.370 76.205 199.275 ;
        RECT 76.835 198.200 77.125 199.365 ;
        RECT 77.295 199.070 77.465 200.100 ;
        RECT 78.145 200.045 78.365 200.530 ;
        RECT 77.635 199.450 77.865 199.845 ;
        RECT 78.035 199.620 78.365 200.045 ;
        RECT 78.535 200.370 79.425 200.540 ;
        RECT 78.535 199.645 78.705 200.370 ;
        RECT 78.875 199.815 79.425 200.200 ;
        RECT 79.655 199.930 79.865 200.750 ;
        RECT 80.035 199.950 80.365 200.580 ;
        RECT 78.535 199.575 79.425 199.645 ;
        RECT 78.530 199.550 79.425 199.575 ;
        RECT 78.520 199.535 79.425 199.550 ;
        RECT 78.515 199.520 79.425 199.535 ;
        RECT 78.505 199.515 79.425 199.520 ;
        RECT 78.500 199.505 79.425 199.515 ;
        RECT 78.495 199.495 79.425 199.505 ;
        RECT 78.485 199.490 79.425 199.495 ;
        RECT 78.475 199.480 79.425 199.490 ;
        RECT 78.465 199.475 79.425 199.480 ;
        RECT 78.465 199.470 78.800 199.475 ;
        RECT 78.450 199.465 78.800 199.470 ;
        RECT 78.435 199.455 78.800 199.465 ;
        RECT 78.410 199.450 78.800 199.455 ;
        RECT 77.635 199.445 78.800 199.450 ;
        RECT 77.635 199.410 78.770 199.445 ;
        RECT 77.635 199.385 78.735 199.410 ;
        RECT 77.635 199.355 78.705 199.385 ;
        RECT 77.635 199.325 78.685 199.355 ;
        RECT 77.635 199.295 78.665 199.325 ;
        RECT 77.635 199.285 78.595 199.295 ;
        RECT 77.635 199.275 78.570 199.285 ;
        RECT 77.635 199.260 78.550 199.275 ;
        RECT 77.635 199.245 78.530 199.260 ;
        RECT 77.740 199.235 78.525 199.245 ;
        RECT 77.740 199.200 78.510 199.235 ;
        RECT 77.295 198.370 77.570 199.070 ;
        RECT 77.740 198.950 78.495 199.200 ;
        RECT 78.665 198.880 78.995 199.125 ;
        RECT 79.165 199.025 79.425 199.475 ;
        RECT 80.035 199.350 80.285 199.950 ;
        RECT 80.535 199.930 80.765 200.750 ;
        RECT 81.015 199.930 81.245 200.750 ;
        RECT 81.415 199.950 81.745 200.580 ;
        RECT 80.455 199.510 80.785 199.760 ;
        RECT 80.995 199.510 81.325 199.760 ;
        RECT 81.495 199.350 81.745 199.950 ;
        RECT 81.915 199.930 82.125 200.750 ;
        RECT 82.415 199.930 82.625 200.750 ;
        RECT 82.795 199.950 83.125 200.580 ;
        RECT 78.810 198.855 78.995 198.880 ;
        RECT 78.810 198.755 79.425 198.855 ;
        RECT 77.740 198.200 77.995 198.745 ;
        RECT 78.165 198.370 78.645 198.710 ;
        RECT 78.820 198.200 79.425 198.755 ;
        RECT 79.655 198.200 79.865 199.340 ;
        RECT 80.035 198.370 80.365 199.350 ;
        RECT 80.535 198.200 80.765 199.340 ;
        RECT 81.015 198.200 81.245 199.340 ;
        RECT 81.415 198.370 81.745 199.350 ;
        RECT 82.795 199.350 83.045 199.950 ;
        RECT 83.295 199.930 83.525 200.750 ;
        RECT 84.195 199.980 85.865 200.750 ;
        RECT 86.040 200.205 91.385 200.750 ;
        RECT 91.560 200.205 96.905 200.750 ;
        RECT 97.080 200.205 102.425 200.750 ;
        RECT 83.215 199.510 83.545 199.760 ;
        RECT 81.915 198.200 82.125 199.340 ;
        RECT 82.415 198.200 82.625 199.340 ;
        RECT 82.795 198.370 83.125 199.350 ;
        RECT 83.295 198.200 83.525 199.340 ;
        RECT 84.195 199.290 84.945 199.810 ;
        RECT 85.115 199.460 85.865 199.980 ;
        RECT 84.195 198.200 85.865 199.290 ;
        RECT 87.630 198.635 87.980 199.885 ;
        RECT 89.460 199.375 89.800 200.205 ;
        RECT 93.150 198.635 93.500 199.885 ;
        RECT 94.980 199.375 95.320 200.205 ;
        RECT 98.670 198.635 99.020 199.885 ;
        RECT 100.500 199.375 100.840 200.205 ;
        RECT 102.595 200.025 102.885 200.750 ;
        RECT 103.520 200.205 108.865 200.750 ;
        RECT 109.040 200.205 114.385 200.750 ;
        RECT 86.040 198.200 91.385 198.635 ;
        RECT 91.560 198.200 96.905 198.635 ;
        RECT 97.080 198.200 102.425 198.635 ;
        RECT 102.595 198.200 102.885 199.365 ;
        RECT 105.110 198.635 105.460 199.885 ;
        RECT 106.940 199.375 107.280 200.205 ;
        RECT 110.630 198.635 110.980 199.885 ;
        RECT 112.460 199.375 112.800 200.205 ;
        RECT 114.555 200.000 115.765 200.750 ;
        RECT 114.555 199.290 115.075 199.830 ;
        RECT 115.245 199.460 115.765 200.000 ;
        RECT 103.520 198.200 108.865 198.635 ;
        RECT 109.040 198.200 114.385 198.635 ;
        RECT 114.555 198.200 115.765 199.290 ;
        RECT 14.650 198.030 115.850 198.200 ;
        RECT 14.735 196.940 15.945 198.030 ;
        RECT 16.120 197.595 21.465 198.030 ;
        RECT 21.640 197.595 26.985 198.030 ;
        RECT 27.160 197.595 32.505 198.030 ;
        RECT 32.680 197.595 38.025 198.030 ;
        RECT 14.735 196.230 15.255 196.770 ;
        RECT 15.425 196.400 15.945 196.940 ;
        RECT 17.710 196.345 18.060 197.595 ;
        RECT 14.735 195.480 15.945 196.230 ;
        RECT 19.540 196.025 19.880 196.855 ;
        RECT 23.230 196.345 23.580 197.595 ;
        RECT 25.060 196.025 25.400 196.855 ;
        RECT 28.750 196.345 29.100 197.595 ;
        RECT 30.580 196.025 30.920 196.855 ;
        RECT 34.270 196.345 34.620 197.595 ;
        RECT 38.195 196.865 38.485 198.030 ;
        RECT 38.655 196.940 42.165 198.030 ;
        RECT 42.340 197.595 47.685 198.030 ;
        RECT 47.860 197.595 53.205 198.030 ;
        RECT 36.100 196.025 36.440 196.855 ;
        RECT 38.655 196.420 40.345 196.940 ;
        RECT 40.515 196.250 42.165 196.770 ;
        RECT 43.930 196.345 44.280 197.595 ;
        RECT 16.120 195.480 21.465 196.025 ;
        RECT 21.640 195.480 26.985 196.025 ;
        RECT 27.160 195.480 32.505 196.025 ;
        RECT 32.680 195.480 38.025 196.025 ;
        RECT 38.195 195.480 38.485 196.205 ;
        RECT 38.655 195.480 42.165 196.250 ;
        RECT 45.760 196.025 46.100 196.855 ;
        RECT 49.450 196.345 49.800 197.595 ;
        RECT 53.380 197.360 53.635 197.860 ;
        RECT 53.805 197.530 54.135 198.030 ;
        RECT 53.380 197.190 54.130 197.360 ;
        RECT 51.280 196.025 51.620 196.855 ;
        RECT 53.380 196.370 53.730 197.020 ;
        RECT 53.900 196.200 54.130 197.190 ;
        RECT 53.380 196.030 54.130 196.200 ;
        RECT 42.340 195.480 47.685 196.025 ;
        RECT 47.860 195.480 53.205 196.025 ;
        RECT 53.380 195.740 53.635 196.030 ;
        RECT 53.805 195.480 54.135 195.860 ;
        RECT 54.305 195.740 54.475 197.860 ;
        RECT 54.645 197.060 54.970 197.845 ;
        RECT 55.140 197.570 55.390 198.030 ;
        RECT 55.560 197.530 55.810 197.860 ;
        RECT 56.025 197.530 56.705 197.860 ;
        RECT 55.560 197.400 55.730 197.530 ;
        RECT 55.335 197.230 55.730 197.400 ;
        RECT 54.705 196.010 55.165 197.060 ;
        RECT 55.335 195.870 55.505 197.230 ;
        RECT 55.900 196.970 56.365 197.360 ;
        RECT 55.675 196.160 56.025 196.780 ;
        RECT 56.195 196.380 56.365 196.970 ;
        RECT 56.535 196.750 56.705 197.530 ;
        RECT 56.875 197.430 57.045 197.770 ;
        RECT 57.280 197.600 57.610 198.030 ;
        RECT 57.780 197.430 57.950 197.770 ;
        RECT 58.245 197.570 58.615 198.030 ;
        RECT 56.875 197.260 57.950 197.430 ;
        RECT 58.785 197.400 58.955 197.860 ;
        RECT 59.190 197.520 60.060 197.860 ;
        RECT 60.230 197.570 60.480 198.030 ;
        RECT 58.395 197.230 58.955 197.400 ;
        RECT 58.395 197.090 58.565 197.230 ;
        RECT 57.065 196.920 58.565 197.090 ;
        RECT 59.260 197.060 59.720 197.350 ;
        RECT 56.535 196.580 58.225 196.750 ;
        RECT 56.195 196.160 56.550 196.380 ;
        RECT 56.720 195.870 56.890 196.580 ;
        RECT 57.095 196.160 57.885 196.410 ;
        RECT 58.055 196.400 58.225 196.580 ;
        RECT 58.395 196.230 58.565 196.920 ;
        RECT 54.835 195.480 55.165 195.840 ;
        RECT 55.335 195.700 55.830 195.870 ;
        RECT 56.035 195.700 56.890 195.870 ;
        RECT 57.765 195.480 58.095 195.940 ;
        RECT 58.305 195.840 58.565 196.230 ;
        RECT 58.755 197.050 59.720 197.060 ;
        RECT 59.890 197.140 60.060 197.520 ;
        RECT 60.650 197.480 60.820 197.770 ;
        RECT 61.000 197.650 61.330 198.030 ;
        RECT 60.650 197.310 61.450 197.480 ;
        RECT 58.755 196.890 59.430 197.050 ;
        RECT 59.890 196.970 61.110 197.140 ;
        RECT 58.755 196.100 58.965 196.890 ;
        RECT 59.890 196.880 60.060 196.970 ;
        RECT 59.135 196.100 59.485 196.720 ;
        RECT 59.655 196.710 60.060 196.880 ;
        RECT 59.655 195.930 59.825 196.710 ;
        RECT 59.995 196.260 60.215 196.540 ;
        RECT 60.395 196.430 60.935 196.800 ;
        RECT 61.280 196.690 61.450 197.310 ;
        RECT 61.625 196.970 61.795 198.030 ;
        RECT 62.005 197.020 62.295 197.860 ;
        RECT 62.465 197.190 62.635 198.030 ;
        RECT 62.845 197.020 63.095 197.860 ;
        RECT 63.305 197.190 63.475 198.030 ;
        RECT 62.005 196.850 63.730 197.020 ;
        RECT 63.955 196.865 64.245 198.030 ;
        RECT 59.995 196.090 60.525 196.260 ;
        RECT 58.305 195.670 58.655 195.840 ;
        RECT 58.875 195.650 59.825 195.930 ;
        RECT 59.995 195.480 60.185 195.920 ;
        RECT 60.355 195.860 60.525 196.090 ;
        RECT 60.695 196.030 60.935 196.430 ;
        RECT 61.105 196.680 61.450 196.690 ;
        RECT 61.105 196.470 63.135 196.680 ;
        RECT 61.105 196.215 61.430 196.470 ;
        RECT 63.320 196.300 63.730 196.850 ;
        RECT 61.105 195.860 61.425 196.215 ;
        RECT 60.355 195.690 61.425 195.860 ;
        RECT 61.625 195.480 61.795 196.290 ;
        RECT 61.965 196.130 63.730 196.300 ;
        RECT 61.965 195.650 62.295 196.130 ;
        RECT 62.465 195.480 62.635 195.950 ;
        RECT 62.805 195.650 63.135 196.130 ;
        RECT 63.305 195.480 63.475 195.950 ;
        RECT 63.955 195.480 64.245 196.205 ;
        RECT 65.335 195.650 65.595 197.860 ;
        RECT 65.765 197.650 66.095 198.030 ;
        RECT 66.520 197.480 66.690 197.860 ;
        RECT 66.950 197.650 67.280 198.030 ;
        RECT 67.475 197.480 67.645 197.860 ;
        RECT 67.855 197.650 68.185 198.030 ;
        RECT 68.435 197.480 68.625 197.860 ;
        RECT 68.865 197.650 69.195 198.030 ;
        RECT 69.505 197.530 69.765 197.860 ;
        RECT 65.765 197.310 67.715 197.480 ;
        RECT 65.765 196.390 65.935 197.310 ;
        RECT 66.305 196.720 66.500 197.030 ;
        RECT 66.770 196.720 66.955 197.030 ;
        RECT 66.245 196.390 66.500 196.720 ;
        RECT 66.725 196.390 66.955 196.720 ;
        RECT 65.765 195.480 66.095 195.860 ;
        RECT 66.305 195.815 66.500 196.390 ;
        RECT 66.770 195.810 66.955 196.390 ;
        RECT 67.205 195.820 67.375 196.720 ;
        RECT 67.545 196.320 67.715 197.310 ;
        RECT 67.885 197.310 68.625 197.480 ;
        RECT 67.885 196.800 68.055 197.310 ;
        RECT 68.225 196.970 68.805 197.140 ;
        RECT 69.075 197.020 69.425 197.350 ;
        RECT 68.635 196.850 68.805 196.970 ;
        RECT 69.595 196.850 69.765 197.530 ;
        RECT 69.935 196.890 70.195 198.030 ;
        RECT 70.365 197.060 70.695 197.860 ;
        RECT 70.865 197.230 71.035 198.030 ;
        RECT 71.235 197.060 71.565 197.860 ;
        RECT 71.765 197.230 72.045 198.030 ;
        RECT 70.365 196.890 71.645 197.060 ;
        RECT 67.885 196.630 68.455 196.800 ;
        RECT 68.635 196.680 69.765 196.850 ;
        RECT 67.545 195.990 68.095 196.320 ;
        RECT 68.285 196.150 68.455 196.630 ;
        RECT 68.625 196.340 69.245 196.510 ;
        RECT 69.035 196.160 69.245 196.340 ;
        RECT 68.285 195.820 68.685 196.150 ;
        RECT 69.595 195.980 69.765 196.680 ;
        RECT 69.960 196.390 70.245 196.720 ;
        RECT 70.445 196.390 70.825 196.720 ;
        RECT 70.995 196.390 71.305 196.720 ;
        RECT 67.205 195.650 68.685 195.820 ;
        RECT 68.865 195.480 69.195 195.860 ;
        RECT 69.505 195.650 69.765 195.980 ;
        RECT 69.940 195.480 70.275 196.220 ;
        RECT 70.445 195.695 70.660 196.390 ;
        RECT 70.995 196.220 71.200 196.390 ;
        RECT 71.475 196.220 71.645 196.890 ;
        RECT 71.825 196.390 72.065 197.060 ;
        RECT 73.160 196.840 73.415 197.720 ;
        RECT 73.585 196.890 73.890 198.030 ;
        RECT 74.230 197.650 74.560 198.030 ;
        RECT 74.740 197.480 74.910 197.770 ;
        RECT 75.080 197.570 75.330 198.030 ;
        RECT 74.110 197.310 74.910 197.480 ;
        RECT 75.500 197.520 76.370 197.860 ;
        RECT 70.850 195.695 71.200 196.220 ;
        RECT 71.370 195.650 72.065 196.220 ;
        RECT 73.160 196.190 73.370 196.840 ;
        RECT 74.110 196.720 74.280 197.310 ;
        RECT 75.500 197.140 75.670 197.520 ;
        RECT 76.605 197.400 76.775 197.860 ;
        RECT 76.945 197.570 77.315 198.030 ;
        RECT 77.610 197.430 77.780 197.770 ;
        RECT 77.950 197.600 78.280 198.030 ;
        RECT 78.515 197.430 78.685 197.770 ;
        RECT 74.450 196.970 75.670 197.140 ;
        RECT 75.840 197.060 76.300 197.350 ;
        RECT 76.605 197.230 77.165 197.400 ;
        RECT 77.610 197.260 78.685 197.430 ;
        RECT 78.855 197.530 79.535 197.860 ;
        RECT 79.750 197.530 80.000 197.860 ;
        RECT 80.170 197.570 80.420 198.030 ;
        RECT 76.995 197.090 77.165 197.230 ;
        RECT 75.840 197.050 76.805 197.060 ;
        RECT 75.500 196.880 75.670 196.970 ;
        RECT 76.130 196.890 76.805 197.050 ;
        RECT 73.540 196.690 74.280 196.720 ;
        RECT 73.540 196.390 74.455 196.690 ;
        RECT 74.130 196.215 74.455 196.390 ;
        RECT 73.160 195.660 73.415 196.190 ;
        RECT 73.585 195.480 73.890 195.940 ;
        RECT 74.135 195.860 74.455 196.215 ;
        RECT 74.625 196.430 75.165 196.800 ;
        RECT 75.500 196.710 75.905 196.880 ;
        RECT 74.625 196.030 74.865 196.430 ;
        RECT 75.345 196.260 75.565 196.540 ;
        RECT 75.035 196.090 75.565 196.260 ;
        RECT 75.035 195.860 75.205 196.090 ;
        RECT 75.735 195.930 75.905 196.710 ;
        RECT 76.075 196.100 76.425 196.720 ;
        RECT 76.595 196.100 76.805 196.890 ;
        RECT 76.995 196.920 78.495 197.090 ;
        RECT 76.995 196.230 77.165 196.920 ;
        RECT 78.855 196.750 79.025 197.530 ;
        RECT 79.830 197.400 80.000 197.530 ;
        RECT 77.335 196.580 79.025 196.750 ;
        RECT 79.195 196.970 79.660 197.360 ;
        RECT 79.830 197.230 80.225 197.400 ;
        RECT 77.335 196.400 77.505 196.580 ;
        RECT 74.135 195.690 75.205 195.860 ;
        RECT 75.375 195.480 75.565 195.920 ;
        RECT 75.735 195.650 76.685 195.930 ;
        RECT 76.995 195.840 77.255 196.230 ;
        RECT 77.675 196.160 78.465 196.410 ;
        RECT 76.905 195.670 77.255 195.840 ;
        RECT 77.465 195.480 77.795 195.940 ;
        RECT 78.670 195.870 78.840 196.580 ;
        RECT 79.195 196.380 79.365 196.970 ;
        RECT 79.010 196.160 79.365 196.380 ;
        RECT 79.535 196.160 79.885 196.780 ;
        RECT 80.055 195.870 80.225 197.230 ;
        RECT 80.590 197.060 80.915 197.845 ;
        RECT 80.395 196.010 80.855 197.060 ;
        RECT 78.670 195.700 79.525 195.870 ;
        RECT 79.730 195.700 80.225 195.870 ;
        RECT 80.395 195.480 80.725 195.840 ;
        RECT 81.085 195.740 81.255 197.860 ;
        RECT 81.425 197.530 81.755 198.030 ;
        RECT 81.925 197.360 82.180 197.860 ;
        RECT 81.430 197.190 82.180 197.360 ;
        RECT 81.430 196.200 81.660 197.190 ;
        RECT 81.830 196.370 82.180 197.020 ;
        RECT 82.355 196.940 84.025 198.030 ;
        RECT 84.200 197.595 89.545 198.030 ;
        RECT 82.355 196.420 83.105 196.940 ;
        RECT 83.275 196.250 84.025 196.770 ;
        RECT 85.790 196.345 86.140 197.595 ;
        RECT 89.715 196.865 90.005 198.030 ;
        RECT 90.175 196.940 93.685 198.030 ;
        RECT 93.970 197.400 94.255 197.860 ;
        RECT 94.425 197.570 94.695 198.030 ;
        RECT 93.970 197.180 94.925 197.400 ;
        RECT 81.430 196.030 82.180 196.200 ;
        RECT 81.425 195.480 81.755 195.860 ;
        RECT 81.925 195.740 82.180 196.030 ;
        RECT 82.355 195.480 84.025 196.250 ;
        RECT 87.620 196.025 87.960 196.855 ;
        RECT 90.175 196.420 91.865 196.940 ;
        RECT 92.035 196.250 93.685 196.770 ;
        RECT 93.855 196.450 94.545 197.010 ;
        RECT 94.715 196.280 94.925 197.180 ;
        RECT 84.200 195.480 89.545 196.025 ;
        RECT 89.715 195.480 90.005 196.205 ;
        RECT 90.175 195.480 93.685 196.250 ;
        RECT 93.970 196.110 94.925 196.280 ;
        RECT 95.095 197.010 95.495 197.860 ;
        RECT 95.685 197.400 95.965 197.860 ;
        RECT 96.485 197.570 96.810 198.030 ;
        RECT 95.685 197.180 96.810 197.400 ;
        RECT 95.095 196.450 96.190 197.010 ;
        RECT 96.360 196.720 96.810 197.180 ;
        RECT 96.980 196.890 97.365 197.860 ;
        RECT 93.970 195.650 94.255 196.110 ;
        RECT 94.425 195.480 94.695 195.940 ;
        RECT 95.095 195.650 95.495 196.450 ;
        RECT 96.360 196.390 96.915 196.720 ;
        RECT 96.360 196.280 96.810 196.390 ;
        RECT 95.685 196.110 96.810 196.280 ;
        RECT 97.085 196.220 97.365 196.890 ;
        RECT 95.685 195.650 95.965 196.110 ;
        RECT 96.485 195.480 96.810 195.940 ;
        RECT 96.980 195.650 97.365 196.220 ;
        RECT 97.540 196.840 97.795 197.720 ;
        RECT 97.965 196.890 98.270 198.030 ;
        RECT 98.610 197.650 98.940 198.030 ;
        RECT 99.120 197.480 99.290 197.770 ;
        RECT 99.460 197.570 99.710 198.030 ;
        RECT 98.490 197.310 99.290 197.480 ;
        RECT 99.880 197.520 100.750 197.860 ;
        RECT 97.540 196.190 97.750 196.840 ;
        RECT 98.490 196.720 98.660 197.310 ;
        RECT 99.880 197.140 100.050 197.520 ;
        RECT 100.985 197.400 101.155 197.860 ;
        RECT 101.325 197.570 101.695 198.030 ;
        RECT 101.990 197.430 102.160 197.770 ;
        RECT 102.330 197.600 102.660 198.030 ;
        RECT 102.895 197.430 103.065 197.770 ;
        RECT 98.830 196.970 100.050 197.140 ;
        RECT 100.220 197.060 100.680 197.350 ;
        RECT 100.985 197.230 101.545 197.400 ;
        RECT 101.990 197.260 103.065 197.430 ;
        RECT 103.235 197.530 103.915 197.860 ;
        RECT 104.130 197.530 104.380 197.860 ;
        RECT 104.550 197.570 104.800 198.030 ;
        RECT 101.375 197.090 101.545 197.230 ;
        RECT 100.220 197.050 101.185 197.060 ;
        RECT 99.880 196.880 100.050 196.970 ;
        RECT 100.510 196.890 101.185 197.050 ;
        RECT 97.920 196.690 98.660 196.720 ;
        RECT 97.920 196.390 98.835 196.690 ;
        RECT 98.510 196.215 98.835 196.390 ;
        RECT 97.540 195.660 97.795 196.190 ;
        RECT 97.965 195.480 98.270 195.940 ;
        RECT 98.515 195.860 98.835 196.215 ;
        RECT 99.005 196.430 99.545 196.800 ;
        RECT 99.880 196.710 100.285 196.880 ;
        RECT 99.005 196.030 99.245 196.430 ;
        RECT 99.725 196.260 99.945 196.540 ;
        RECT 99.415 196.090 99.945 196.260 ;
        RECT 99.415 195.860 99.585 196.090 ;
        RECT 100.115 195.930 100.285 196.710 ;
        RECT 100.455 196.100 100.805 196.720 ;
        RECT 100.975 196.100 101.185 196.890 ;
        RECT 101.375 196.920 102.875 197.090 ;
        RECT 101.375 196.230 101.545 196.920 ;
        RECT 103.235 196.750 103.405 197.530 ;
        RECT 104.210 197.400 104.380 197.530 ;
        RECT 101.715 196.580 103.405 196.750 ;
        RECT 103.575 196.970 104.040 197.360 ;
        RECT 104.210 197.230 104.605 197.400 ;
        RECT 101.715 196.400 101.885 196.580 ;
        RECT 98.515 195.690 99.585 195.860 ;
        RECT 99.755 195.480 99.945 195.920 ;
        RECT 100.115 195.650 101.065 195.930 ;
        RECT 101.375 195.840 101.635 196.230 ;
        RECT 102.055 196.160 102.845 196.410 ;
        RECT 101.285 195.670 101.635 195.840 ;
        RECT 101.845 195.480 102.175 195.940 ;
        RECT 103.050 195.870 103.220 196.580 ;
        RECT 103.575 196.380 103.745 196.970 ;
        RECT 103.390 196.160 103.745 196.380 ;
        RECT 103.915 196.160 104.265 196.780 ;
        RECT 104.435 195.870 104.605 197.230 ;
        RECT 104.970 197.060 105.295 197.845 ;
        RECT 104.775 196.010 105.235 197.060 ;
        RECT 103.050 195.700 103.905 195.870 ;
        RECT 104.110 195.700 104.605 195.870 ;
        RECT 104.775 195.480 105.105 195.840 ;
        RECT 105.465 195.740 105.635 197.860 ;
        RECT 105.805 197.530 106.135 198.030 ;
        RECT 106.305 197.360 106.560 197.860 ;
        RECT 105.810 197.190 106.560 197.360 ;
        RECT 105.810 196.200 106.040 197.190 ;
        RECT 106.210 196.370 106.560 197.020 ;
        RECT 107.195 196.940 108.865 198.030 ;
        RECT 109.040 197.595 114.385 198.030 ;
        RECT 107.195 196.420 107.945 196.940 ;
        RECT 108.115 196.250 108.865 196.770 ;
        RECT 110.630 196.345 110.980 197.595 ;
        RECT 114.555 196.940 115.765 198.030 ;
        RECT 105.810 196.030 106.560 196.200 ;
        RECT 105.805 195.480 106.135 195.860 ;
        RECT 106.305 195.740 106.560 196.030 ;
        RECT 107.195 195.480 108.865 196.250 ;
        RECT 112.460 196.025 112.800 196.855 ;
        RECT 114.555 196.400 115.075 196.940 ;
        RECT 115.245 196.230 115.765 196.770 ;
        RECT 109.040 195.480 114.385 196.025 ;
        RECT 114.555 195.480 115.765 196.230 ;
        RECT 14.650 195.310 115.850 195.480 ;
        RECT 14.735 194.560 15.945 195.310 ;
        RECT 14.735 194.020 15.255 194.560 ;
        RECT 16.115 194.540 19.625 195.310 ;
        RECT 19.800 194.765 25.145 195.310 ;
        RECT 15.425 193.850 15.945 194.390 ;
        RECT 14.735 192.760 15.945 193.850 ;
        RECT 16.115 193.850 17.805 194.370 ;
        RECT 17.975 194.020 19.625 194.540 ;
        RECT 16.115 192.760 19.625 193.850 ;
        RECT 21.390 193.195 21.740 194.445 ;
        RECT 23.220 193.935 23.560 194.765 ;
        RECT 25.315 194.585 25.605 195.310 ;
        RECT 26.235 194.540 29.745 195.310 ;
        RECT 29.920 194.765 35.265 195.310 ;
        RECT 35.440 194.765 40.785 195.310 ;
        RECT 19.800 192.760 25.145 193.195 ;
        RECT 25.315 192.760 25.605 193.925 ;
        RECT 26.235 193.850 27.925 194.370 ;
        RECT 28.095 194.020 29.745 194.540 ;
        RECT 26.235 192.760 29.745 193.850 ;
        RECT 31.510 193.195 31.860 194.445 ;
        RECT 33.340 193.935 33.680 194.765 ;
        RECT 37.030 193.195 37.380 194.445 ;
        RECT 38.860 193.935 39.200 194.765 ;
        RECT 41.070 194.680 41.355 195.140 ;
        RECT 41.525 194.850 41.795 195.310 ;
        RECT 41.070 194.510 42.025 194.680 ;
        RECT 40.955 193.780 41.645 194.340 ;
        RECT 41.815 193.610 42.025 194.510 ;
        RECT 41.070 193.390 42.025 193.610 ;
        RECT 42.195 194.340 42.595 195.140 ;
        RECT 42.785 194.680 43.065 195.140 ;
        RECT 43.585 194.850 43.910 195.310 ;
        RECT 42.785 194.510 43.910 194.680 ;
        RECT 44.080 194.570 44.465 195.140 ;
        RECT 43.460 194.400 43.910 194.510 ;
        RECT 42.195 193.780 43.290 194.340 ;
        RECT 43.460 194.070 44.015 194.400 ;
        RECT 29.920 192.760 35.265 193.195 ;
        RECT 35.440 192.760 40.785 193.195 ;
        RECT 41.070 192.930 41.355 193.390 ;
        RECT 41.525 192.760 41.795 193.220 ;
        RECT 42.195 192.930 42.595 193.780 ;
        RECT 43.460 193.610 43.910 194.070 ;
        RECT 44.185 193.900 44.465 194.570 ;
        RECT 45.095 194.540 47.685 195.310 ;
        RECT 42.785 193.390 43.910 193.610 ;
        RECT 42.785 192.930 43.065 193.390 ;
        RECT 43.585 192.760 43.910 193.220 ;
        RECT 44.080 192.930 44.465 193.900 ;
        RECT 45.095 193.850 46.305 194.370 ;
        RECT 46.475 194.020 47.685 194.540 ;
        RECT 47.915 194.490 48.125 195.310 ;
        RECT 48.295 194.510 48.625 195.140 ;
        RECT 48.295 193.910 48.545 194.510 ;
        RECT 48.795 194.490 49.025 195.310 ;
        RECT 49.235 194.635 49.495 195.140 ;
        RECT 49.675 194.930 50.005 195.310 ;
        RECT 50.185 194.760 50.355 195.140 ;
        RECT 48.715 194.070 49.045 194.320 ;
        RECT 45.095 192.760 47.685 193.850 ;
        RECT 47.915 192.760 48.125 193.900 ;
        RECT 48.295 192.930 48.625 193.910 ;
        RECT 48.795 192.760 49.025 193.900 ;
        RECT 49.235 193.835 49.405 194.635 ;
        RECT 49.690 194.590 50.355 194.760 ;
        RECT 49.690 194.335 49.860 194.590 ;
        RECT 51.075 194.585 51.365 195.310 ;
        RECT 51.995 194.540 55.505 195.310 ;
        RECT 55.680 194.765 61.025 195.310 ;
        RECT 61.525 194.910 61.855 195.310 ;
        RECT 49.575 194.005 49.860 194.335 ;
        RECT 50.095 194.040 50.425 194.410 ;
        RECT 49.690 193.860 49.860 194.005 ;
        RECT 49.235 192.930 49.505 193.835 ;
        RECT 49.690 193.690 50.355 193.860 ;
        RECT 49.675 192.760 50.005 193.520 ;
        RECT 50.185 192.930 50.355 193.690 ;
        RECT 51.075 192.760 51.365 193.925 ;
        RECT 51.995 193.850 53.685 194.370 ;
        RECT 53.855 194.020 55.505 194.540 ;
        RECT 51.995 192.760 55.505 193.850 ;
        RECT 57.270 193.195 57.620 194.445 ;
        RECT 59.100 193.935 59.440 194.765 ;
        RECT 62.025 194.740 62.355 195.080 ;
        RECT 63.405 194.910 63.735 195.310 ;
        RECT 61.370 194.570 63.735 194.740 ;
        RECT 63.905 194.585 64.235 195.095 ;
        RECT 61.370 193.570 61.540 194.570 ;
        RECT 63.565 194.400 63.735 194.570 ;
        RECT 61.710 193.740 61.955 194.400 ;
        RECT 62.170 193.740 62.435 194.400 ;
        RECT 62.630 193.740 62.915 194.400 ;
        RECT 63.090 194.070 63.395 194.400 ;
        RECT 63.565 194.070 63.875 194.400 ;
        RECT 63.090 193.740 63.305 194.070 ;
        RECT 61.370 193.400 61.825 193.570 ;
        RECT 55.680 192.760 61.025 193.195 ;
        RECT 61.495 192.970 61.825 193.400 ;
        RECT 62.005 193.400 63.295 193.570 ;
        RECT 62.005 192.980 62.255 193.400 ;
        RECT 62.485 192.760 62.815 193.230 ;
        RECT 63.045 192.980 63.295 193.400 ;
        RECT 63.485 192.760 63.735 193.900 ;
        RECT 64.045 193.820 64.235 194.585 ;
        RECT 64.500 194.740 64.675 195.140 ;
        RECT 64.845 194.930 65.175 195.310 ;
        RECT 65.420 194.810 65.650 195.140 ;
        RECT 64.500 194.570 65.130 194.740 ;
        RECT 64.960 194.400 65.130 194.570 ;
        RECT 63.905 192.970 64.235 193.820 ;
        RECT 64.415 193.720 64.780 194.400 ;
        RECT 64.960 194.070 65.310 194.400 ;
        RECT 64.960 193.550 65.130 194.070 ;
        RECT 64.500 193.380 65.130 193.550 ;
        RECT 65.480 193.520 65.650 194.810 ;
        RECT 65.850 193.700 66.130 194.975 ;
        RECT 66.355 194.630 66.625 194.975 ;
        RECT 67.085 194.930 67.415 195.310 ;
        RECT 67.585 195.055 67.920 195.100 ;
        RECT 66.315 194.460 66.625 194.630 ;
        RECT 66.355 193.700 66.625 194.460 ;
        RECT 66.815 193.700 67.155 194.730 ;
        RECT 67.585 194.590 67.925 195.055 ;
        RECT 67.325 194.070 67.585 194.400 ;
        RECT 67.325 193.520 67.495 194.070 ;
        RECT 67.755 193.900 67.925 194.590 ;
        RECT 68.095 194.560 69.305 195.310 ;
        RECT 64.500 192.930 64.675 193.380 ;
        RECT 65.480 193.350 67.495 193.520 ;
        RECT 64.845 192.760 65.175 193.200 ;
        RECT 65.480 192.930 65.650 193.350 ;
        RECT 65.885 192.760 66.555 193.170 ;
        RECT 66.770 192.930 66.940 193.350 ;
        RECT 67.140 192.760 67.470 193.170 ;
        RECT 67.665 192.930 67.925 193.900 ;
        RECT 68.095 193.850 68.615 194.390 ;
        RECT 68.785 194.020 69.305 194.560 ;
        RECT 69.590 194.680 69.875 195.140 ;
        RECT 70.045 194.850 70.315 195.310 ;
        RECT 69.590 194.510 70.545 194.680 ;
        RECT 68.095 192.760 69.305 193.850 ;
        RECT 69.475 193.780 70.165 194.340 ;
        RECT 70.335 193.610 70.545 194.510 ;
        RECT 69.590 193.390 70.545 193.610 ;
        RECT 70.715 194.340 71.115 195.140 ;
        RECT 71.305 194.680 71.585 195.140 ;
        RECT 72.105 194.850 72.430 195.310 ;
        RECT 71.305 194.510 72.430 194.680 ;
        RECT 72.600 194.570 72.985 195.140 ;
        RECT 71.980 194.400 72.430 194.510 ;
        RECT 70.715 193.780 71.810 194.340 ;
        RECT 71.980 194.070 72.535 194.400 ;
        RECT 69.590 192.930 69.875 193.390 ;
        RECT 70.045 192.760 70.315 193.220 ;
        RECT 70.715 192.930 71.115 193.780 ;
        RECT 71.980 193.610 72.430 194.070 ;
        RECT 72.705 193.900 72.985 194.570 ;
        RECT 71.305 193.390 72.430 193.610 ;
        RECT 71.305 192.930 71.585 193.390 ;
        RECT 72.105 192.760 72.430 193.220 ;
        RECT 72.600 192.930 72.985 193.900 ;
        RECT 73.155 194.660 73.415 195.140 ;
        RECT 73.585 194.770 73.835 195.310 ;
        RECT 73.155 193.630 73.325 194.660 ;
        RECT 74.005 194.630 74.225 195.090 ;
        RECT 73.975 194.605 74.225 194.630 ;
        RECT 73.495 194.010 73.725 194.405 ;
        RECT 73.895 194.180 74.225 194.605 ;
        RECT 74.395 194.930 75.285 195.100 ;
        RECT 74.395 194.205 74.565 194.930 ;
        RECT 74.735 194.375 75.285 194.760 ;
        RECT 75.455 194.510 76.150 195.140 ;
        RECT 76.355 194.510 76.665 195.310 ;
        RECT 76.835 194.585 77.125 195.310 ;
        RECT 77.760 194.765 83.105 195.310 ;
        RECT 74.395 194.135 75.285 194.205 ;
        RECT 74.390 194.110 75.285 194.135 ;
        RECT 74.380 194.095 75.285 194.110 ;
        RECT 74.375 194.080 75.285 194.095 ;
        RECT 74.365 194.075 75.285 194.080 ;
        RECT 74.360 194.065 75.285 194.075 ;
        RECT 75.475 194.070 75.810 194.320 ;
        RECT 74.355 194.055 75.285 194.065 ;
        RECT 74.345 194.050 75.285 194.055 ;
        RECT 74.335 194.040 75.285 194.050 ;
        RECT 74.325 194.035 75.285 194.040 ;
        RECT 74.325 194.030 74.660 194.035 ;
        RECT 74.310 194.025 74.660 194.030 ;
        RECT 74.295 194.015 74.660 194.025 ;
        RECT 74.270 194.010 74.660 194.015 ;
        RECT 73.495 194.005 74.660 194.010 ;
        RECT 73.495 193.970 74.630 194.005 ;
        RECT 73.495 193.945 74.595 193.970 ;
        RECT 73.495 193.915 74.565 193.945 ;
        RECT 73.495 193.885 74.545 193.915 ;
        RECT 73.495 193.855 74.525 193.885 ;
        RECT 73.495 193.845 74.455 193.855 ;
        RECT 73.495 193.835 74.430 193.845 ;
        RECT 73.495 193.820 74.410 193.835 ;
        RECT 73.495 193.805 74.390 193.820 ;
        RECT 73.600 193.795 74.385 193.805 ;
        RECT 73.600 193.760 74.370 193.795 ;
        RECT 73.155 192.930 73.430 193.630 ;
        RECT 73.600 193.510 74.355 193.760 ;
        RECT 74.525 193.440 74.855 193.685 ;
        RECT 75.025 193.585 75.285 194.035 ;
        RECT 75.980 193.910 76.150 194.510 ;
        RECT 76.320 194.070 76.655 194.340 ;
        RECT 74.670 193.415 74.855 193.440 ;
        RECT 74.670 193.315 75.285 193.415 ;
        RECT 73.600 192.760 73.855 193.305 ;
        RECT 74.025 192.930 74.505 193.270 ;
        RECT 74.680 192.760 75.285 193.315 ;
        RECT 75.455 192.760 75.715 193.900 ;
        RECT 75.885 192.930 76.215 193.910 ;
        RECT 76.385 192.760 76.665 193.900 ;
        RECT 76.835 192.760 77.125 193.925 ;
        RECT 79.350 193.195 79.700 194.445 ;
        RECT 81.180 193.935 81.520 194.765 ;
        RECT 83.365 194.760 83.535 195.140 ;
        RECT 83.715 194.930 84.045 195.310 ;
        RECT 83.365 194.590 84.030 194.760 ;
        RECT 84.225 194.635 84.485 195.140 ;
        RECT 83.295 194.040 83.625 194.410 ;
        RECT 83.860 194.335 84.030 194.590 ;
        RECT 83.860 194.005 84.145 194.335 ;
        RECT 83.860 193.860 84.030 194.005 ;
        RECT 83.365 193.690 84.030 193.860 ;
        RECT 84.315 193.835 84.485 194.635 ;
        RECT 84.655 194.560 85.865 195.310 ;
        RECT 77.760 192.760 83.105 193.195 ;
        RECT 83.365 192.930 83.535 193.690 ;
        RECT 83.715 192.760 84.045 193.520 ;
        RECT 84.215 192.930 84.485 193.835 ;
        RECT 84.655 193.850 85.175 194.390 ;
        RECT 85.345 194.020 85.865 194.560 ;
        RECT 86.075 194.490 86.305 195.310 ;
        RECT 86.475 194.510 86.805 195.140 ;
        RECT 86.055 194.070 86.385 194.320 ;
        RECT 86.555 193.910 86.805 194.510 ;
        RECT 86.975 194.490 87.185 195.310 ;
        RECT 87.420 194.760 87.675 195.050 ;
        RECT 87.845 194.930 88.175 195.310 ;
        RECT 87.420 194.590 88.170 194.760 ;
        RECT 84.655 192.760 85.865 193.850 ;
        RECT 86.075 192.760 86.305 193.900 ;
        RECT 86.475 192.930 86.805 193.910 ;
        RECT 86.975 192.760 87.185 193.900 ;
        RECT 87.420 193.770 87.770 194.420 ;
        RECT 87.940 193.600 88.170 194.590 ;
        RECT 87.420 193.430 88.170 193.600 ;
        RECT 87.420 192.930 87.675 193.430 ;
        RECT 87.845 192.760 88.175 193.260 ;
        RECT 88.345 192.930 88.515 195.050 ;
        RECT 88.875 194.950 89.205 195.310 ;
        RECT 89.375 194.920 89.870 195.090 ;
        RECT 90.075 194.920 90.930 195.090 ;
        RECT 88.745 193.730 89.205 194.780 ;
        RECT 88.685 192.945 89.010 193.730 ;
        RECT 89.375 193.560 89.545 194.920 ;
        RECT 89.715 194.010 90.065 194.630 ;
        RECT 90.235 194.410 90.590 194.630 ;
        RECT 90.235 193.820 90.405 194.410 ;
        RECT 90.760 194.210 90.930 194.920 ;
        RECT 91.805 194.850 92.135 195.310 ;
        RECT 92.345 194.950 92.695 195.120 ;
        RECT 91.135 194.380 91.925 194.630 ;
        RECT 92.345 194.560 92.605 194.950 ;
        RECT 92.915 194.860 93.865 195.140 ;
        RECT 94.035 194.870 94.225 195.310 ;
        RECT 94.395 194.930 95.465 195.100 ;
        RECT 92.095 194.210 92.265 194.390 ;
        RECT 89.375 193.390 89.770 193.560 ;
        RECT 89.940 193.430 90.405 193.820 ;
        RECT 90.575 194.040 92.265 194.210 ;
        RECT 89.600 193.260 89.770 193.390 ;
        RECT 90.575 193.260 90.745 194.040 ;
        RECT 92.435 193.870 92.605 194.560 ;
        RECT 91.105 193.700 92.605 193.870 ;
        RECT 92.795 193.900 93.005 194.690 ;
        RECT 93.175 194.070 93.525 194.690 ;
        RECT 93.695 194.080 93.865 194.860 ;
        RECT 94.395 194.700 94.565 194.930 ;
        RECT 94.035 194.530 94.565 194.700 ;
        RECT 94.035 194.250 94.255 194.530 ;
        RECT 94.735 194.360 94.975 194.760 ;
        RECT 93.695 193.910 94.100 194.080 ;
        RECT 94.435 193.990 94.975 194.360 ;
        RECT 95.145 194.575 95.465 194.930 ;
        RECT 95.710 194.850 96.015 195.310 ;
        RECT 96.185 194.600 96.440 195.130 ;
        RECT 95.145 194.400 95.470 194.575 ;
        RECT 95.145 194.100 96.060 194.400 ;
        RECT 95.320 194.070 96.060 194.100 ;
        RECT 92.795 193.740 93.470 193.900 ;
        RECT 93.930 193.820 94.100 193.910 ;
        RECT 92.795 193.730 93.760 193.740 ;
        RECT 92.435 193.560 92.605 193.700 ;
        RECT 89.180 192.760 89.430 193.220 ;
        RECT 89.600 192.930 89.850 193.260 ;
        RECT 90.065 192.930 90.745 193.260 ;
        RECT 90.915 193.360 91.990 193.530 ;
        RECT 92.435 193.390 92.995 193.560 ;
        RECT 93.300 193.440 93.760 193.730 ;
        RECT 93.930 193.650 95.150 193.820 ;
        RECT 90.915 193.020 91.085 193.360 ;
        RECT 91.320 192.760 91.650 193.190 ;
        RECT 91.820 193.020 91.990 193.360 ;
        RECT 92.285 192.760 92.655 193.220 ;
        RECT 92.825 192.930 92.995 193.390 ;
        RECT 93.930 193.270 94.100 193.650 ;
        RECT 95.320 193.480 95.490 194.070 ;
        RECT 96.230 193.950 96.440 194.600 ;
        RECT 97.115 194.490 97.345 195.310 ;
        RECT 97.515 194.510 97.845 195.140 ;
        RECT 97.095 194.070 97.425 194.320 ;
        RECT 93.230 192.930 94.100 193.270 ;
        RECT 94.690 193.310 95.490 193.480 ;
        RECT 94.270 192.760 94.520 193.220 ;
        RECT 94.690 193.020 94.860 193.310 ;
        RECT 95.040 192.760 95.370 193.140 ;
        RECT 95.710 192.760 96.015 193.900 ;
        RECT 96.185 193.070 96.440 193.950 ;
        RECT 97.595 193.910 97.845 194.510 ;
        RECT 98.015 194.490 98.225 195.310 ;
        RECT 98.730 194.500 98.975 195.105 ;
        RECT 99.195 194.775 99.705 195.310 ;
        RECT 97.115 192.760 97.345 193.900 ;
        RECT 97.515 192.930 97.845 193.910 ;
        RECT 98.455 194.330 99.685 194.500 ;
        RECT 98.015 192.760 98.225 193.900 ;
        RECT 98.455 193.520 98.795 194.330 ;
        RECT 98.965 193.765 99.715 193.955 ;
        RECT 98.455 193.110 98.970 193.520 ;
        RECT 99.205 192.760 99.375 193.520 ;
        RECT 99.545 193.100 99.715 193.765 ;
        RECT 99.885 193.780 100.075 195.140 ;
        RECT 100.245 194.970 100.520 195.140 ;
        RECT 100.245 194.800 100.525 194.970 ;
        RECT 100.245 193.980 100.520 194.800 ;
        RECT 100.710 194.775 101.240 195.140 ;
        RECT 101.665 194.910 101.995 195.310 ;
        RECT 101.065 194.740 101.240 194.775 ;
        RECT 100.725 193.780 100.895 194.580 ;
        RECT 99.885 193.610 100.895 193.780 ;
        RECT 101.065 194.570 101.995 194.740 ;
        RECT 102.165 194.570 102.420 195.140 ;
        RECT 102.595 194.585 102.885 195.310 ;
        RECT 103.170 194.680 103.455 195.140 ;
        RECT 103.625 194.850 103.895 195.310 ;
        RECT 101.065 193.440 101.235 194.570 ;
        RECT 101.825 194.400 101.995 194.570 ;
        RECT 100.110 193.270 101.235 193.440 ;
        RECT 101.405 194.070 101.600 194.400 ;
        RECT 101.825 194.070 102.080 194.400 ;
        RECT 101.405 193.100 101.575 194.070 ;
        RECT 102.250 193.900 102.420 194.570 ;
        RECT 103.170 194.510 104.125 194.680 ;
        RECT 99.545 192.930 101.575 193.100 ;
        RECT 101.745 192.760 101.915 193.900 ;
        RECT 102.085 192.930 102.420 193.900 ;
        RECT 102.595 192.760 102.885 193.925 ;
        RECT 103.055 193.780 103.745 194.340 ;
        RECT 103.915 193.610 104.125 194.510 ;
        RECT 103.170 193.390 104.125 193.610 ;
        RECT 104.295 194.340 104.695 195.140 ;
        RECT 104.885 194.680 105.165 195.140 ;
        RECT 105.685 194.850 106.010 195.310 ;
        RECT 104.885 194.510 106.010 194.680 ;
        RECT 106.180 194.570 106.565 195.140 ;
        RECT 105.560 194.400 106.010 194.510 ;
        RECT 104.295 193.780 105.390 194.340 ;
        RECT 105.560 194.070 106.115 194.400 ;
        RECT 103.170 192.930 103.455 193.390 ;
        RECT 103.625 192.760 103.895 193.220 ;
        RECT 104.295 192.930 104.695 193.780 ;
        RECT 105.560 193.610 106.010 194.070 ;
        RECT 106.285 193.900 106.565 194.570 ;
        RECT 106.775 194.490 107.005 195.310 ;
        RECT 107.175 194.510 107.505 195.140 ;
        RECT 106.755 194.070 107.085 194.320 ;
        RECT 107.255 193.910 107.505 194.510 ;
        RECT 107.675 194.490 107.885 195.310 ;
        RECT 108.205 194.760 108.375 195.140 ;
        RECT 108.555 194.930 108.885 195.310 ;
        RECT 108.205 194.590 108.870 194.760 ;
        RECT 109.065 194.635 109.325 195.140 ;
        RECT 108.135 194.040 108.465 194.410 ;
        RECT 108.700 194.335 108.870 194.590 ;
        RECT 104.885 193.390 106.010 193.610 ;
        RECT 104.885 192.930 105.165 193.390 ;
        RECT 105.685 192.760 106.010 193.220 ;
        RECT 106.180 192.930 106.565 193.900 ;
        RECT 106.775 192.760 107.005 193.900 ;
        RECT 107.175 192.930 107.505 193.910 ;
        RECT 108.700 194.005 108.985 194.335 ;
        RECT 107.675 192.760 107.885 193.900 ;
        RECT 108.700 193.860 108.870 194.005 ;
        RECT 108.205 193.690 108.870 193.860 ;
        RECT 109.155 193.835 109.325 194.635 ;
        RECT 109.495 194.560 110.705 195.310 ;
        RECT 108.205 192.930 108.375 193.690 ;
        RECT 108.555 192.760 108.885 193.520 ;
        RECT 109.055 192.930 109.325 193.835 ;
        RECT 109.495 193.850 110.015 194.390 ;
        RECT 110.185 194.020 110.705 194.560 ;
        RECT 110.875 194.540 114.385 195.310 ;
        RECT 114.555 194.560 115.765 195.310 ;
        RECT 110.875 193.850 112.565 194.370 ;
        RECT 112.735 194.020 114.385 194.540 ;
        RECT 114.555 193.850 115.075 194.390 ;
        RECT 115.245 194.020 115.765 194.560 ;
        RECT 109.495 192.760 110.705 193.850 ;
        RECT 110.875 192.760 114.385 193.850 ;
        RECT 114.555 192.760 115.765 193.850 ;
        RECT 14.650 192.590 115.850 192.760 ;
        RECT 14.735 191.500 15.945 192.590 ;
        RECT 14.735 190.790 15.255 191.330 ;
        RECT 15.425 190.960 15.945 191.500 ;
        RECT 16.115 191.500 17.325 192.590 ;
        RECT 17.495 191.500 21.005 192.590 ;
        RECT 21.180 192.155 26.525 192.590 ;
        RECT 16.115 190.960 16.635 191.500 ;
        RECT 16.805 190.790 17.325 191.330 ;
        RECT 17.495 190.980 19.185 191.500 ;
        RECT 19.355 190.810 21.005 191.330 ;
        RECT 22.770 190.905 23.120 192.155 ;
        RECT 26.810 191.960 27.095 192.420 ;
        RECT 27.265 192.130 27.535 192.590 ;
        RECT 26.810 191.740 27.765 191.960 ;
        RECT 14.735 190.040 15.945 190.790 ;
        RECT 16.115 190.040 17.325 190.790 ;
        RECT 17.495 190.040 21.005 190.810 ;
        RECT 24.600 190.585 24.940 191.415 ;
        RECT 26.695 191.010 27.385 191.570 ;
        RECT 27.555 190.840 27.765 191.740 ;
        RECT 26.810 190.670 27.765 190.840 ;
        RECT 27.935 191.570 28.335 192.420 ;
        RECT 28.525 191.960 28.805 192.420 ;
        RECT 29.325 192.130 29.650 192.590 ;
        RECT 28.525 191.740 29.650 191.960 ;
        RECT 27.935 191.010 29.030 191.570 ;
        RECT 29.200 191.280 29.650 191.740 ;
        RECT 29.820 191.450 30.205 192.420 ;
        RECT 21.180 190.040 26.525 190.585 ;
        RECT 26.810 190.210 27.095 190.670 ;
        RECT 27.265 190.040 27.535 190.500 ;
        RECT 27.935 190.210 28.335 191.010 ;
        RECT 29.200 190.950 29.755 191.280 ;
        RECT 29.200 190.840 29.650 190.950 ;
        RECT 28.525 190.670 29.650 190.840 ;
        RECT 29.925 190.780 30.205 191.450 ;
        RECT 30.835 191.500 32.505 192.590 ;
        RECT 30.835 190.980 31.585 191.500 ;
        RECT 32.715 191.450 32.945 192.590 ;
        RECT 33.115 191.440 33.445 192.420 ;
        RECT 33.615 191.450 33.825 192.590 ;
        RECT 34.055 191.830 34.570 192.240 ;
        RECT 34.805 191.830 34.975 192.590 ;
        RECT 35.145 192.250 37.175 192.420 ;
        RECT 31.755 190.810 32.505 191.330 ;
        RECT 32.695 191.030 33.025 191.280 ;
        RECT 28.525 190.210 28.805 190.670 ;
        RECT 29.325 190.040 29.650 190.500 ;
        RECT 29.820 190.210 30.205 190.780 ;
        RECT 30.835 190.040 32.505 190.810 ;
        RECT 32.715 190.040 32.945 190.860 ;
        RECT 33.195 190.840 33.445 191.440 ;
        RECT 34.055 191.020 34.395 191.830 ;
        RECT 35.145 191.585 35.315 192.250 ;
        RECT 35.710 191.910 36.835 192.080 ;
        RECT 34.565 191.395 35.315 191.585 ;
        RECT 35.485 191.570 36.495 191.740 ;
        RECT 33.115 190.210 33.445 190.840 ;
        RECT 33.615 190.040 33.825 190.860 ;
        RECT 34.055 190.850 35.285 191.020 ;
        RECT 34.330 190.245 34.575 190.850 ;
        RECT 34.795 190.040 35.305 190.575 ;
        RECT 35.485 190.210 35.675 191.570 ;
        RECT 35.845 190.890 36.120 191.370 ;
        RECT 35.845 190.720 36.125 190.890 ;
        RECT 36.325 190.770 36.495 191.570 ;
        RECT 36.665 190.780 36.835 191.910 ;
        RECT 37.005 191.280 37.175 192.250 ;
        RECT 37.345 191.450 37.515 192.590 ;
        RECT 37.685 191.450 38.020 192.420 ;
        RECT 37.005 190.950 37.200 191.280 ;
        RECT 37.425 190.950 37.680 191.280 ;
        RECT 37.425 190.780 37.595 190.950 ;
        RECT 37.850 190.780 38.020 191.450 ;
        RECT 38.195 191.425 38.485 192.590 ;
        RECT 38.745 191.660 38.915 192.420 ;
        RECT 39.095 191.830 39.425 192.590 ;
        RECT 38.745 191.490 39.410 191.660 ;
        RECT 39.595 191.515 39.865 192.420 ;
        RECT 39.240 191.345 39.410 191.490 ;
        RECT 38.675 190.940 39.005 191.310 ;
        RECT 39.240 191.015 39.525 191.345 ;
        RECT 35.845 190.210 36.120 190.720 ;
        RECT 36.665 190.610 37.595 190.780 ;
        RECT 36.665 190.575 36.840 190.610 ;
        RECT 36.310 190.210 36.840 190.575 ;
        RECT 37.265 190.040 37.595 190.440 ;
        RECT 37.765 190.210 38.020 190.780 ;
        RECT 38.195 190.040 38.485 190.765 ;
        RECT 39.240 190.760 39.410 191.015 ;
        RECT 38.745 190.590 39.410 190.760 ;
        RECT 39.695 190.715 39.865 191.515 ;
        RECT 38.745 190.210 38.915 190.590 ;
        RECT 39.095 190.040 39.425 190.420 ;
        RECT 39.605 190.210 39.865 190.715 ;
        RECT 40.500 191.400 40.755 192.280 ;
        RECT 40.925 191.450 41.230 192.590 ;
        RECT 41.570 192.210 41.900 192.590 ;
        RECT 42.080 192.040 42.250 192.330 ;
        RECT 42.420 192.130 42.670 192.590 ;
        RECT 41.450 191.870 42.250 192.040 ;
        RECT 42.840 192.080 43.710 192.420 ;
        RECT 40.500 190.750 40.710 191.400 ;
        RECT 41.450 191.280 41.620 191.870 ;
        RECT 42.840 191.700 43.010 192.080 ;
        RECT 43.945 191.960 44.115 192.420 ;
        RECT 44.285 192.130 44.655 192.590 ;
        RECT 44.950 191.990 45.120 192.330 ;
        RECT 45.290 192.160 45.620 192.590 ;
        RECT 45.855 191.990 46.025 192.330 ;
        RECT 41.790 191.530 43.010 191.700 ;
        RECT 43.180 191.620 43.640 191.910 ;
        RECT 43.945 191.790 44.505 191.960 ;
        RECT 44.950 191.820 46.025 191.990 ;
        RECT 46.195 192.090 46.875 192.420 ;
        RECT 47.090 192.090 47.340 192.420 ;
        RECT 47.510 192.130 47.760 192.590 ;
        RECT 44.335 191.650 44.505 191.790 ;
        RECT 43.180 191.610 44.145 191.620 ;
        RECT 42.840 191.440 43.010 191.530 ;
        RECT 43.470 191.450 44.145 191.610 ;
        RECT 40.880 191.250 41.620 191.280 ;
        RECT 40.880 190.950 41.795 191.250 ;
        RECT 41.470 190.775 41.795 190.950 ;
        RECT 40.500 190.220 40.755 190.750 ;
        RECT 40.925 190.040 41.230 190.500 ;
        RECT 41.475 190.420 41.795 190.775 ;
        RECT 41.965 190.990 42.505 191.360 ;
        RECT 42.840 191.270 43.245 191.440 ;
        RECT 41.965 190.590 42.205 190.990 ;
        RECT 42.685 190.820 42.905 191.100 ;
        RECT 42.375 190.650 42.905 190.820 ;
        RECT 42.375 190.420 42.545 190.650 ;
        RECT 43.075 190.490 43.245 191.270 ;
        RECT 43.415 190.660 43.765 191.280 ;
        RECT 43.935 190.660 44.145 191.450 ;
        RECT 44.335 191.480 45.835 191.650 ;
        RECT 44.335 190.790 44.505 191.480 ;
        RECT 46.195 191.310 46.365 192.090 ;
        RECT 47.170 191.960 47.340 192.090 ;
        RECT 44.675 191.140 46.365 191.310 ;
        RECT 46.535 191.530 47.000 191.920 ;
        RECT 47.170 191.790 47.565 191.960 ;
        RECT 44.675 190.960 44.845 191.140 ;
        RECT 41.475 190.250 42.545 190.420 ;
        RECT 42.715 190.040 42.905 190.480 ;
        RECT 43.075 190.210 44.025 190.490 ;
        RECT 44.335 190.400 44.595 190.790 ;
        RECT 45.015 190.720 45.805 190.970 ;
        RECT 44.245 190.230 44.595 190.400 ;
        RECT 44.805 190.040 45.135 190.500 ;
        RECT 46.010 190.430 46.180 191.140 ;
        RECT 46.535 190.940 46.705 191.530 ;
        RECT 46.350 190.720 46.705 190.940 ;
        RECT 46.875 190.720 47.225 191.340 ;
        RECT 47.395 190.430 47.565 191.790 ;
        RECT 47.930 191.620 48.255 192.405 ;
        RECT 47.735 190.570 48.195 191.620 ;
        RECT 46.010 190.260 46.865 190.430 ;
        RECT 47.070 190.260 47.565 190.430 ;
        RECT 47.735 190.040 48.065 190.400 ;
        RECT 48.425 190.300 48.595 192.420 ;
        RECT 48.765 192.090 49.095 192.590 ;
        RECT 49.265 191.920 49.520 192.420 ;
        RECT 48.770 191.750 49.520 191.920 ;
        RECT 48.770 190.760 49.000 191.750 ;
        RECT 49.170 190.930 49.520 191.580 ;
        RECT 49.700 191.400 49.955 192.280 ;
        RECT 50.125 191.450 50.430 192.590 ;
        RECT 50.770 192.210 51.100 192.590 ;
        RECT 51.280 192.040 51.450 192.330 ;
        RECT 51.620 192.130 51.870 192.590 ;
        RECT 50.650 191.870 51.450 192.040 ;
        RECT 52.040 192.080 52.910 192.420 ;
        RECT 48.770 190.590 49.520 190.760 ;
        RECT 48.765 190.040 49.095 190.420 ;
        RECT 49.265 190.300 49.520 190.590 ;
        RECT 49.700 190.750 49.910 191.400 ;
        RECT 50.650 191.280 50.820 191.870 ;
        RECT 52.040 191.700 52.210 192.080 ;
        RECT 53.145 191.960 53.315 192.420 ;
        RECT 53.485 192.130 53.855 192.590 ;
        RECT 54.150 191.990 54.320 192.330 ;
        RECT 54.490 192.160 54.820 192.590 ;
        RECT 55.055 191.990 55.225 192.330 ;
        RECT 50.990 191.530 52.210 191.700 ;
        RECT 52.380 191.620 52.840 191.910 ;
        RECT 53.145 191.790 53.705 191.960 ;
        RECT 54.150 191.820 55.225 191.990 ;
        RECT 55.395 192.090 56.075 192.420 ;
        RECT 56.290 192.090 56.540 192.420 ;
        RECT 56.710 192.130 56.960 192.590 ;
        RECT 53.535 191.650 53.705 191.790 ;
        RECT 52.380 191.610 53.345 191.620 ;
        RECT 52.040 191.440 52.210 191.530 ;
        RECT 52.670 191.450 53.345 191.610 ;
        RECT 50.080 191.250 50.820 191.280 ;
        RECT 50.080 190.950 50.995 191.250 ;
        RECT 50.670 190.775 50.995 190.950 ;
        RECT 49.700 190.220 49.955 190.750 ;
        RECT 50.125 190.040 50.430 190.500 ;
        RECT 50.675 190.420 50.995 190.775 ;
        RECT 51.165 190.990 51.705 191.360 ;
        RECT 52.040 191.270 52.445 191.440 ;
        RECT 51.165 190.590 51.405 190.990 ;
        RECT 51.885 190.820 52.105 191.100 ;
        RECT 51.575 190.650 52.105 190.820 ;
        RECT 51.575 190.420 51.745 190.650 ;
        RECT 52.275 190.490 52.445 191.270 ;
        RECT 52.615 190.660 52.965 191.280 ;
        RECT 53.135 190.660 53.345 191.450 ;
        RECT 53.535 191.480 55.035 191.650 ;
        RECT 53.535 190.790 53.705 191.480 ;
        RECT 55.395 191.310 55.565 192.090 ;
        RECT 56.370 191.960 56.540 192.090 ;
        RECT 53.875 191.140 55.565 191.310 ;
        RECT 55.735 191.530 56.200 191.920 ;
        RECT 56.370 191.790 56.765 191.960 ;
        RECT 53.875 190.960 54.045 191.140 ;
        RECT 50.675 190.250 51.745 190.420 ;
        RECT 51.915 190.040 52.105 190.480 ;
        RECT 52.275 190.210 53.225 190.490 ;
        RECT 53.535 190.400 53.795 190.790 ;
        RECT 54.215 190.720 55.005 190.970 ;
        RECT 53.445 190.230 53.795 190.400 ;
        RECT 54.005 190.040 54.335 190.500 ;
        RECT 55.210 190.430 55.380 191.140 ;
        RECT 55.735 190.940 55.905 191.530 ;
        RECT 55.550 190.720 55.905 190.940 ;
        RECT 56.075 190.720 56.425 191.340 ;
        RECT 56.595 190.430 56.765 191.790 ;
        RECT 57.130 191.620 57.455 192.405 ;
        RECT 56.935 190.570 57.395 191.620 ;
        RECT 55.210 190.260 56.065 190.430 ;
        RECT 56.270 190.260 56.765 190.430 ;
        RECT 56.935 190.040 57.265 190.400 ;
        RECT 57.625 190.300 57.795 192.420 ;
        RECT 57.965 192.090 58.295 192.590 ;
        RECT 58.465 191.920 58.720 192.420 ;
        RECT 57.970 191.750 58.720 191.920 ;
        RECT 57.970 190.760 58.200 191.750 ;
        RECT 58.370 190.930 58.720 191.580 ;
        RECT 58.935 191.450 59.165 192.590 ;
        RECT 59.335 191.440 59.665 192.420 ;
        RECT 59.835 191.450 60.045 192.590 ;
        RECT 60.390 191.960 60.675 192.420 ;
        RECT 60.845 192.130 61.115 192.590 ;
        RECT 60.390 191.740 61.345 191.960 ;
        RECT 58.915 191.030 59.245 191.280 ;
        RECT 57.970 190.590 58.720 190.760 ;
        RECT 57.965 190.040 58.295 190.420 ;
        RECT 58.465 190.300 58.720 190.590 ;
        RECT 58.935 190.040 59.165 190.860 ;
        RECT 59.415 190.840 59.665 191.440 ;
        RECT 60.275 191.010 60.965 191.570 ;
        RECT 59.335 190.210 59.665 190.840 ;
        RECT 59.835 190.040 60.045 190.860 ;
        RECT 61.135 190.840 61.345 191.740 ;
        RECT 60.390 190.670 61.345 190.840 ;
        RECT 61.515 191.570 61.915 192.420 ;
        RECT 62.105 191.960 62.385 192.420 ;
        RECT 62.905 192.130 63.230 192.590 ;
        RECT 62.105 191.740 63.230 191.960 ;
        RECT 61.515 191.010 62.610 191.570 ;
        RECT 62.780 191.280 63.230 191.740 ;
        RECT 63.400 191.450 63.785 192.420 ;
        RECT 60.390 190.210 60.675 190.670 ;
        RECT 60.845 190.040 61.115 190.500 ;
        RECT 61.515 190.210 61.915 191.010 ;
        RECT 62.780 190.950 63.335 191.280 ;
        RECT 62.780 190.840 63.230 190.950 ;
        RECT 62.105 190.670 63.230 190.840 ;
        RECT 63.505 190.780 63.785 191.450 ;
        RECT 63.955 191.425 64.245 192.590 ;
        RECT 64.415 191.500 66.085 192.590 ;
        RECT 64.415 190.980 65.165 191.500 ;
        RECT 66.255 191.450 66.515 192.590 ;
        RECT 66.755 192.080 68.370 192.410 ;
        RECT 65.335 190.810 66.085 191.330 ;
        RECT 66.765 191.280 66.935 191.840 ;
        RECT 67.195 191.740 68.370 191.910 ;
        RECT 68.540 191.790 68.820 192.590 ;
        RECT 67.195 191.450 67.525 191.740 ;
        RECT 68.200 191.620 68.370 191.740 ;
        RECT 67.695 191.280 67.940 191.570 ;
        RECT 68.200 191.450 68.860 191.620 ;
        RECT 69.030 191.450 69.305 192.420 ;
        RECT 69.475 191.450 69.735 192.590 ;
        RECT 69.975 192.080 71.590 192.410 ;
        RECT 68.690 191.280 68.860 191.450 ;
        RECT 66.260 191.030 66.595 191.280 ;
        RECT 66.765 190.950 67.480 191.280 ;
        RECT 67.695 190.950 68.520 191.280 ;
        RECT 68.690 190.950 68.965 191.280 ;
        RECT 66.765 190.860 67.015 190.950 ;
        RECT 62.105 190.210 62.385 190.670 ;
        RECT 62.905 190.040 63.230 190.500 ;
        RECT 63.400 190.210 63.785 190.780 ;
        RECT 63.955 190.040 64.245 190.765 ;
        RECT 64.415 190.040 66.085 190.810 ;
        RECT 66.255 190.040 66.515 190.860 ;
        RECT 66.685 190.440 67.015 190.860 ;
        RECT 68.690 190.780 68.860 190.950 ;
        RECT 67.195 190.610 68.860 190.780 ;
        RECT 69.135 190.715 69.305 191.450 ;
        RECT 69.985 191.280 70.155 191.840 ;
        RECT 70.415 191.740 71.590 191.910 ;
        RECT 71.760 191.790 72.040 192.590 ;
        RECT 70.415 191.450 70.745 191.740 ;
        RECT 71.420 191.620 71.590 191.740 ;
        RECT 70.915 191.280 71.160 191.570 ;
        RECT 71.420 191.450 72.080 191.620 ;
        RECT 72.250 191.450 72.525 192.420 ;
        RECT 71.910 191.280 72.080 191.450 ;
        RECT 69.480 191.030 69.815 191.280 ;
        RECT 69.985 190.950 70.700 191.280 ;
        RECT 70.915 190.950 71.740 191.280 ;
        RECT 71.910 190.950 72.185 191.280 ;
        RECT 69.985 190.860 70.235 190.950 ;
        RECT 67.195 190.210 67.455 190.610 ;
        RECT 67.625 190.040 67.955 190.440 ;
        RECT 68.125 190.260 68.295 190.610 ;
        RECT 68.465 190.040 68.840 190.440 ;
        RECT 69.030 190.370 69.305 190.715 ;
        RECT 69.475 190.040 69.735 190.860 ;
        RECT 69.905 190.440 70.235 190.860 ;
        RECT 71.910 190.780 72.080 190.950 ;
        RECT 70.415 190.610 72.080 190.780 ;
        RECT 72.355 190.715 72.525 191.450 ;
        RECT 70.415 190.210 70.675 190.610 ;
        RECT 70.845 190.040 71.175 190.440 ;
        RECT 71.345 190.260 71.515 190.610 ;
        RECT 71.685 190.040 72.060 190.440 ;
        RECT 72.250 190.370 72.525 190.715 ;
        RECT 72.695 191.620 72.965 192.390 ;
        RECT 73.135 191.810 73.465 192.590 ;
        RECT 73.670 191.985 73.855 192.390 ;
        RECT 74.025 192.165 74.360 192.590 ;
        RECT 73.670 191.810 74.335 191.985 ;
        RECT 72.695 191.450 73.825 191.620 ;
        RECT 72.695 190.540 72.865 191.450 ;
        RECT 73.035 190.700 73.395 191.280 ;
        RECT 73.575 190.950 73.825 191.450 ;
        RECT 73.995 190.780 74.335 191.810 ;
        RECT 74.995 191.500 77.585 192.590 ;
        RECT 78.130 191.610 78.385 192.280 ;
        RECT 78.565 191.790 78.850 192.590 ;
        RECT 79.030 191.870 79.360 192.380 ;
        RECT 74.995 190.980 76.205 191.500 ;
        RECT 76.375 190.810 77.585 191.330 ;
        RECT 73.650 190.610 74.335 190.780 ;
        RECT 72.695 190.210 72.955 190.540 ;
        RECT 73.165 190.040 73.440 190.520 ;
        RECT 73.650 190.210 73.855 190.610 ;
        RECT 74.025 190.040 74.360 190.440 ;
        RECT 74.995 190.040 77.585 190.810 ;
        RECT 78.130 190.750 78.310 191.610 ;
        RECT 79.030 191.280 79.280 191.870 ;
        RECT 79.630 191.720 79.800 192.330 ;
        RECT 79.970 191.900 80.300 192.590 ;
        RECT 80.530 192.040 80.770 192.330 ;
        RECT 80.970 192.210 81.390 192.590 ;
        RECT 81.570 192.120 82.200 192.370 ;
        RECT 82.670 192.210 83.000 192.590 ;
        RECT 81.570 192.040 81.740 192.120 ;
        RECT 83.170 192.040 83.340 192.330 ;
        RECT 83.520 192.210 83.900 192.590 ;
        RECT 84.140 192.205 84.970 192.375 ;
        RECT 80.530 191.870 81.740 192.040 ;
        RECT 78.480 190.950 79.280 191.280 ;
        RECT 78.130 190.550 78.385 190.750 ;
        RECT 78.045 190.380 78.385 190.550 ;
        RECT 78.130 190.220 78.385 190.380 ;
        RECT 78.565 190.040 78.850 190.500 ;
        RECT 79.030 190.300 79.280 190.950 ;
        RECT 79.480 191.700 79.800 191.720 ;
        RECT 79.480 191.530 81.400 191.700 ;
        RECT 79.480 190.635 79.670 191.530 ;
        RECT 81.570 191.360 81.740 191.870 ;
        RECT 81.910 191.610 82.430 191.920 ;
        RECT 79.840 191.190 81.740 191.360 ;
        RECT 79.840 191.130 80.170 191.190 ;
        RECT 80.320 190.960 80.650 191.020 ;
        RECT 79.990 190.690 80.650 190.960 ;
        RECT 79.480 190.305 79.800 190.635 ;
        RECT 79.980 190.040 80.640 190.520 ;
        RECT 80.840 190.430 81.010 191.190 ;
        RECT 81.910 191.020 82.090 191.430 ;
        RECT 81.180 190.850 81.510 190.970 ;
        RECT 82.260 190.850 82.430 191.610 ;
        RECT 81.180 190.680 82.430 190.850 ;
        RECT 82.600 191.790 83.970 192.040 ;
        RECT 82.600 191.020 82.790 191.790 ;
        RECT 83.720 191.530 83.970 191.790 ;
        RECT 82.960 191.360 83.210 191.520 ;
        RECT 84.140 191.360 84.310 192.205 ;
        RECT 85.205 191.920 85.375 192.420 ;
        RECT 85.545 192.090 85.875 192.590 ;
        RECT 84.480 191.530 84.980 191.910 ;
        RECT 85.205 191.750 85.900 191.920 ;
        RECT 82.960 191.190 84.310 191.360 ;
        RECT 83.890 191.150 84.310 191.190 ;
        RECT 82.600 190.680 83.020 191.020 ;
        RECT 83.310 190.690 83.720 191.020 ;
        RECT 80.840 190.260 81.690 190.430 ;
        RECT 82.250 190.040 82.570 190.500 ;
        RECT 82.770 190.250 83.020 190.680 ;
        RECT 83.310 190.040 83.720 190.480 ;
        RECT 83.890 190.420 84.060 191.150 ;
        RECT 84.230 190.600 84.580 190.970 ;
        RECT 84.760 190.660 84.980 191.530 ;
        RECT 85.150 190.960 85.560 191.580 ;
        RECT 85.730 190.780 85.900 191.750 ;
        RECT 85.205 190.590 85.900 190.780 ;
        RECT 83.890 190.220 84.905 190.420 ;
        RECT 85.205 190.260 85.375 190.590 ;
        RECT 85.545 190.040 85.875 190.420 ;
        RECT 86.090 190.300 86.315 192.420 ;
        RECT 86.485 192.090 86.815 192.590 ;
        RECT 86.985 191.920 87.155 192.420 ;
        RECT 86.490 191.750 87.155 191.920 ;
        RECT 86.490 190.760 86.720 191.750 ;
        RECT 86.890 190.930 87.240 191.580 ;
        RECT 88.335 191.515 88.605 192.420 ;
        RECT 88.775 191.830 89.105 192.590 ;
        RECT 89.285 191.660 89.455 192.420 ;
        RECT 86.490 190.590 87.155 190.760 ;
        RECT 86.485 190.040 86.815 190.420 ;
        RECT 86.985 190.300 87.155 190.590 ;
        RECT 88.335 190.715 88.505 191.515 ;
        RECT 88.790 191.490 89.455 191.660 ;
        RECT 88.790 191.345 88.960 191.490 ;
        RECT 89.715 191.425 90.005 192.590 ;
        RECT 90.180 191.450 90.515 192.420 ;
        RECT 90.685 191.450 90.855 192.590 ;
        RECT 91.025 192.250 93.055 192.420 ;
        RECT 88.675 191.015 88.960 191.345 ;
        RECT 88.790 190.760 88.960 191.015 ;
        RECT 89.195 190.940 89.525 191.310 ;
        RECT 90.180 190.780 90.350 191.450 ;
        RECT 91.025 191.280 91.195 192.250 ;
        RECT 90.520 190.950 90.775 191.280 ;
        RECT 91.000 190.950 91.195 191.280 ;
        RECT 91.365 191.910 92.490 192.080 ;
        RECT 90.605 190.780 90.775 190.950 ;
        RECT 91.365 190.780 91.535 191.910 ;
        RECT 88.335 190.210 88.595 190.715 ;
        RECT 88.790 190.590 89.455 190.760 ;
        RECT 88.775 190.040 89.105 190.420 ;
        RECT 89.285 190.210 89.455 190.590 ;
        RECT 89.715 190.040 90.005 190.765 ;
        RECT 90.180 190.210 90.435 190.780 ;
        RECT 90.605 190.610 91.535 190.780 ;
        RECT 91.705 191.570 92.715 191.740 ;
        RECT 91.705 190.770 91.875 191.570 ;
        RECT 91.360 190.575 91.535 190.610 ;
        RECT 90.605 190.040 90.935 190.440 ;
        RECT 91.360 190.210 91.890 190.575 ;
        RECT 92.080 190.550 92.355 191.370 ;
        RECT 92.075 190.380 92.355 190.550 ;
        RECT 92.080 190.210 92.355 190.380 ;
        RECT 92.525 190.210 92.715 191.570 ;
        RECT 92.885 191.585 93.055 192.250 ;
        RECT 93.225 191.830 93.395 192.590 ;
        RECT 93.630 191.830 94.145 192.240 ;
        RECT 92.885 191.395 93.635 191.585 ;
        RECT 93.805 191.020 94.145 191.830 ;
        RECT 92.915 190.850 94.145 191.020 ;
        RECT 94.315 191.500 96.905 192.590 ;
        RECT 94.315 190.980 95.525 191.500 ;
        RECT 97.080 191.450 97.415 192.420 ;
        RECT 97.585 191.450 97.755 192.590 ;
        RECT 97.925 192.250 99.955 192.420 ;
        RECT 92.895 190.040 93.405 190.575 ;
        RECT 93.625 190.245 93.870 190.850 ;
        RECT 95.695 190.810 96.905 191.330 ;
        RECT 94.315 190.040 96.905 190.810 ;
        RECT 97.080 190.780 97.250 191.450 ;
        RECT 97.925 191.280 98.095 192.250 ;
        RECT 97.420 190.950 97.675 191.280 ;
        RECT 97.900 190.950 98.095 191.280 ;
        RECT 98.265 191.910 99.390 192.080 ;
        RECT 97.505 190.780 97.675 190.950 ;
        RECT 98.265 190.780 98.435 191.910 ;
        RECT 97.080 190.210 97.335 190.780 ;
        RECT 97.505 190.610 98.435 190.780 ;
        RECT 98.605 191.570 99.615 191.740 ;
        RECT 98.605 190.770 98.775 191.570 ;
        RECT 98.980 190.890 99.255 191.370 ;
        RECT 98.975 190.720 99.255 190.890 ;
        RECT 98.260 190.575 98.435 190.610 ;
        RECT 97.505 190.040 97.835 190.440 ;
        RECT 98.260 190.210 98.790 190.575 ;
        RECT 98.980 190.210 99.255 190.720 ;
        RECT 99.425 190.210 99.615 191.570 ;
        RECT 99.785 191.585 99.955 192.250 ;
        RECT 100.125 191.830 100.295 192.590 ;
        RECT 100.530 191.830 101.045 192.240 ;
        RECT 99.785 191.395 100.535 191.585 ;
        RECT 100.705 191.020 101.045 191.830 ;
        RECT 99.815 190.850 101.045 191.020 ;
        RECT 101.220 191.400 101.475 192.280 ;
        RECT 101.645 191.450 101.950 192.590 ;
        RECT 102.290 192.210 102.620 192.590 ;
        RECT 102.800 192.040 102.970 192.330 ;
        RECT 103.140 192.130 103.390 192.590 ;
        RECT 102.170 191.870 102.970 192.040 ;
        RECT 103.560 192.080 104.430 192.420 ;
        RECT 99.795 190.040 100.305 190.575 ;
        RECT 100.525 190.245 100.770 190.850 ;
        RECT 101.220 190.750 101.430 191.400 ;
        RECT 102.170 191.280 102.340 191.870 ;
        RECT 103.560 191.700 103.730 192.080 ;
        RECT 104.665 191.960 104.835 192.420 ;
        RECT 105.005 192.130 105.375 192.590 ;
        RECT 105.670 191.990 105.840 192.330 ;
        RECT 106.010 192.160 106.340 192.590 ;
        RECT 106.575 191.990 106.745 192.330 ;
        RECT 102.510 191.530 103.730 191.700 ;
        RECT 103.900 191.620 104.360 191.910 ;
        RECT 104.665 191.790 105.225 191.960 ;
        RECT 105.670 191.820 106.745 191.990 ;
        RECT 106.915 192.090 107.595 192.420 ;
        RECT 107.810 192.090 108.060 192.420 ;
        RECT 108.230 192.130 108.480 192.590 ;
        RECT 105.055 191.650 105.225 191.790 ;
        RECT 103.900 191.610 104.865 191.620 ;
        RECT 103.560 191.440 103.730 191.530 ;
        RECT 104.190 191.450 104.865 191.610 ;
        RECT 101.600 191.250 102.340 191.280 ;
        RECT 101.600 190.950 102.515 191.250 ;
        RECT 102.190 190.775 102.515 190.950 ;
        RECT 101.220 190.220 101.475 190.750 ;
        RECT 101.645 190.040 101.950 190.500 ;
        RECT 102.195 190.420 102.515 190.775 ;
        RECT 102.685 190.990 103.225 191.360 ;
        RECT 103.560 191.270 103.965 191.440 ;
        RECT 102.685 190.590 102.925 190.990 ;
        RECT 103.405 190.820 103.625 191.100 ;
        RECT 103.095 190.650 103.625 190.820 ;
        RECT 103.095 190.420 103.265 190.650 ;
        RECT 103.795 190.490 103.965 191.270 ;
        RECT 104.135 190.660 104.485 191.280 ;
        RECT 104.655 190.660 104.865 191.450 ;
        RECT 105.055 191.480 106.555 191.650 ;
        RECT 105.055 190.790 105.225 191.480 ;
        RECT 106.915 191.310 107.085 192.090 ;
        RECT 107.890 191.960 108.060 192.090 ;
        RECT 105.395 191.140 107.085 191.310 ;
        RECT 107.255 191.530 107.720 191.920 ;
        RECT 107.890 191.790 108.285 191.960 ;
        RECT 105.395 190.960 105.565 191.140 ;
        RECT 102.195 190.250 103.265 190.420 ;
        RECT 103.435 190.040 103.625 190.480 ;
        RECT 103.795 190.210 104.745 190.490 ;
        RECT 105.055 190.400 105.315 190.790 ;
        RECT 105.735 190.720 106.525 190.970 ;
        RECT 104.965 190.230 105.315 190.400 ;
        RECT 105.525 190.040 105.855 190.500 ;
        RECT 106.730 190.430 106.900 191.140 ;
        RECT 107.255 190.940 107.425 191.530 ;
        RECT 107.070 190.720 107.425 190.940 ;
        RECT 107.595 190.720 107.945 191.340 ;
        RECT 108.115 190.430 108.285 191.790 ;
        RECT 108.650 191.620 108.975 192.405 ;
        RECT 108.455 190.570 108.915 191.620 ;
        RECT 106.730 190.260 107.585 190.430 ;
        RECT 107.790 190.260 108.285 190.430 ;
        RECT 108.455 190.040 108.785 190.400 ;
        RECT 109.145 190.300 109.315 192.420 ;
        RECT 109.485 192.090 109.815 192.590 ;
        RECT 109.985 191.920 110.240 192.420 ;
        RECT 109.490 191.750 110.240 191.920 ;
        RECT 109.490 190.760 109.720 191.750 ;
        RECT 109.890 190.930 110.240 191.580 ;
        RECT 110.875 191.500 114.385 192.590 ;
        RECT 114.555 191.500 115.765 192.590 ;
        RECT 110.875 190.980 112.565 191.500 ;
        RECT 112.735 190.810 114.385 191.330 ;
        RECT 114.555 190.960 115.075 191.500 ;
        RECT 109.490 190.590 110.240 190.760 ;
        RECT 109.485 190.040 109.815 190.420 ;
        RECT 109.985 190.300 110.240 190.590 ;
        RECT 110.875 190.040 114.385 190.810 ;
        RECT 115.245 190.790 115.765 191.330 ;
        RECT 114.555 190.040 115.765 190.790 ;
        RECT 14.650 189.870 115.850 190.040 ;
        RECT 14.735 189.120 15.945 189.870 ;
        RECT 14.735 188.580 15.255 189.120 ;
        RECT 16.115 189.100 19.625 189.870 ;
        RECT 19.800 189.325 25.145 189.870 ;
        RECT 15.425 188.410 15.945 188.950 ;
        RECT 14.735 187.320 15.945 188.410 ;
        RECT 16.115 188.410 17.805 188.930 ;
        RECT 17.975 188.580 19.625 189.100 ;
        RECT 16.115 187.320 19.625 188.410 ;
        RECT 21.390 187.755 21.740 189.005 ;
        RECT 23.220 188.495 23.560 189.325 ;
        RECT 25.315 189.145 25.605 189.870 ;
        RECT 26.695 189.195 26.955 189.700 ;
        RECT 27.135 189.490 27.465 189.870 ;
        RECT 27.645 189.320 27.815 189.700 ;
        RECT 19.800 187.320 25.145 187.755 ;
        RECT 25.315 187.320 25.605 188.485 ;
        RECT 26.695 188.395 26.865 189.195 ;
        RECT 27.150 189.150 27.815 189.320 ;
        RECT 28.190 189.240 28.475 189.700 ;
        RECT 28.645 189.410 28.915 189.870 ;
        RECT 27.150 188.895 27.320 189.150 ;
        RECT 28.190 189.070 29.145 189.240 ;
        RECT 27.035 188.565 27.320 188.895 ;
        RECT 27.555 188.600 27.885 188.970 ;
        RECT 27.150 188.420 27.320 188.565 ;
        RECT 26.695 187.490 26.965 188.395 ;
        RECT 27.150 188.250 27.815 188.420 ;
        RECT 28.075 188.340 28.765 188.900 ;
        RECT 27.135 187.320 27.465 188.080 ;
        RECT 27.645 187.490 27.815 188.250 ;
        RECT 28.935 188.170 29.145 189.070 ;
        RECT 28.190 187.950 29.145 188.170 ;
        RECT 29.315 188.900 29.715 189.700 ;
        RECT 29.905 189.240 30.185 189.700 ;
        RECT 30.705 189.410 31.030 189.870 ;
        RECT 29.905 189.070 31.030 189.240 ;
        RECT 31.200 189.130 31.585 189.700 ;
        RECT 30.580 188.960 31.030 189.070 ;
        RECT 29.315 188.340 30.410 188.900 ;
        RECT 30.580 188.630 31.135 188.960 ;
        RECT 28.190 187.490 28.475 187.950 ;
        RECT 28.645 187.320 28.915 187.780 ;
        RECT 29.315 187.490 29.715 188.340 ;
        RECT 30.580 188.170 31.030 188.630 ;
        RECT 31.305 188.460 31.585 189.130 ;
        RECT 29.905 187.950 31.030 188.170 ;
        RECT 29.905 187.490 30.185 187.950 ;
        RECT 30.705 187.320 31.030 187.780 ;
        RECT 31.200 187.490 31.585 188.460 ;
        RECT 32.130 189.160 32.385 189.690 ;
        RECT 32.565 189.410 32.850 189.870 ;
        RECT 32.130 188.300 32.310 189.160 ;
        RECT 33.030 188.960 33.280 189.610 ;
        RECT 32.480 188.630 33.280 188.960 ;
        RECT 32.130 187.830 32.385 188.300 ;
        RECT 32.045 187.660 32.385 187.830 ;
        RECT 32.130 187.630 32.385 187.660 ;
        RECT 32.565 187.320 32.850 188.120 ;
        RECT 33.030 188.040 33.280 188.630 ;
        RECT 33.480 189.275 33.800 189.605 ;
        RECT 33.980 189.390 34.640 189.870 ;
        RECT 34.840 189.480 35.690 189.650 ;
        RECT 33.480 188.380 33.670 189.275 ;
        RECT 33.990 188.950 34.650 189.220 ;
        RECT 34.320 188.890 34.650 188.950 ;
        RECT 33.840 188.720 34.170 188.780 ;
        RECT 34.840 188.720 35.010 189.480 ;
        RECT 36.250 189.410 36.570 189.870 ;
        RECT 36.770 189.230 37.020 189.660 ;
        RECT 37.310 189.430 37.720 189.870 ;
        RECT 37.890 189.490 38.905 189.690 ;
        RECT 35.180 189.060 36.430 189.230 ;
        RECT 35.180 188.940 35.510 189.060 ;
        RECT 33.840 188.550 35.740 188.720 ;
        RECT 33.480 188.210 35.400 188.380 ;
        RECT 33.480 188.190 33.800 188.210 ;
        RECT 33.030 187.530 33.360 188.040 ;
        RECT 33.630 187.580 33.800 188.190 ;
        RECT 35.570 188.040 35.740 188.550 ;
        RECT 35.910 188.480 36.090 188.890 ;
        RECT 36.260 188.300 36.430 189.060 ;
        RECT 33.970 187.320 34.300 188.010 ;
        RECT 34.530 187.870 35.740 188.040 ;
        RECT 35.910 187.990 36.430 188.300 ;
        RECT 36.600 188.890 37.020 189.230 ;
        RECT 37.310 188.890 37.720 189.220 ;
        RECT 36.600 188.120 36.790 188.890 ;
        RECT 37.890 188.760 38.060 189.490 ;
        RECT 39.205 189.320 39.375 189.650 ;
        RECT 39.545 189.490 39.875 189.870 ;
        RECT 38.230 188.940 38.580 189.310 ;
        RECT 37.890 188.720 38.310 188.760 ;
        RECT 36.960 188.550 38.310 188.720 ;
        RECT 36.960 188.390 37.210 188.550 ;
        RECT 37.720 188.120 37.970 188.380 ;
        RECT 36.600 187.870 37.970 188.120 ;
        RECT 34.530 187.580 34.770 187.870 ;
        RECT 35.570 187.790 35.740 187.870 ;
        RECT 34.970 187.320 35.390 187.700 ;
        RECT 35.570 187.540 36.200 187.790 ;
        RECT 36.670 187.320 37.000 187.700 ;
        RECT 37.170 187.580 37.340 187.870 ;
        RECT 38.140 187.705 38.310 188.550 ;
        RECT 38.760 188.380 38.980 189.250 ;
        RECT 39.205 189.130 39.900 189.320 ;
        RECT 38.480 188.000 38.980 188.380 ;
        RECT 39.150 188.330 39.560 188.950 ;
        RECT 39.730 188.160 39.900 189.130 ;
        RECT 39.205 187.990 39.900 188.160 ;
        RECT 37.520 187.320 37.900 187.700 ;
        RECT 38.140 187.535 38.970 187.705 ;
        RECT 39.205 187.490 39.375 187.990 ;
        RECT 39.545 187.320 39.875 187.820 ;
        RECT 40.090 187.490 40.315 189.610 ;
        RECT 40.485 189.490 40.815 189.870 ;
        RECT 40.985 189.320 41.155 189.610 ;
        RECT 40.490 189.150 41.155 189.320 ;
        RECT 41.415 189.195 41.675 189.700 ;
        RECT 41.855 189.490 42.185 189.870 ;
        RECT 42.365 189.320 42.535 189.700 ;
        RECT 40.490 188.160 40.720 189.150 ;
        RECT 40.890 188.330 41.240 188.980 ;
        RECT 41.415 188.395 41.585 189.195 ;
        RECT 41.870 189.150 42.535 189.320 ;
        RECT 41.870 188.895 42.040 189.150 ;
        RECT 43.070 189.060 43.315 189.665 ;
        RECT 43.535 189.335 44.045 189.870 ;
        RECT 41.755 188.565 42.040 188.895 ;
        RECT 42.275 188.600 42.605 188.970 ;
        RECT 42.795 188.890 44.025 189.060 ;
        RECT 41.870 188.420 42.040 188.565 ;
        RECT 40.490 187.990 41.155 188.160 ;
        RECT 40.485 187.320 40.815 187.820 ;
        RECT 40.985 187.490 41.155 187.990 ;
        RECT 41.415 187.490 41.685 188.395 ;
        RECT 41.870 188.250 42.535 188.420 ;
        RECT 41.855 187.320 42.185 188.080 ;
        RECT 42.365 187.490 42.535 188.250 ;
        RECT 42.795 188.080 43.135 188.890 ;
        RECT 43.305 188.325 44.055 188.515 ;
        RECT 42.795 187.670 43.310 188.080 ;
        RECT 43.545 187.320 43.715 188.080 ;
        RECT 43.885 187.660 44.055 188.325 ;
        RECT 44.225 188.340 44.415 189.700 ;
        RECT 44.585 188.850 44.860 189.700 ;
        RECT 45.050 189.335 45.580 189.700 ;
        RECT 46.005 189.470 46.335 189.870 ;
        RECT 45.405 189.300 45.580 189.335 ;
        RECT 44.585 188.680 44.865 188.850 ;
        RECT 44.585 188.540 44.860 188.680 ;
        RECT 45.065 188.340 45.235 189.140 ;
        RECT 44.225 188.170 45.235 188.340 ;
        RECT 45.405 189.130 46.335 189.300 ;
        RECT 46.505 189.130 46.760 189.700 ;
        RECT 45.405 188.000 45.575 189.130 ;
        RECT 46.165 188.960 46.335 189.130 ;
        RECT 44.450 187.830 45.575 188.000 ;
        RECT 45.745 188.630 45.940 188.960 ;
        RECT 46.165 188.630 46.420 188.960 ;
        RECT 45.745 187.660 45.915 188.630 ;
        RECT 46.590 188.460 46.760 189.130 ;
        RECT 47.210 189.060 47.455 189.665 ;
        RECT 47.675 189.335 48.185 189.870 ;
        RECT 43.885 187.490 45.915 187.660 ;
        RECT 46.085 187.320 46.255 188.460 ;
        RECT 46.425 187.490 46.760 188.460 ;
        RECT 46.935 188.890 48.165 189.060 ;
        RECT 46.935 188.080 47.275 188.890 ;
        RECT 47.445 188.325 48.195 188.515 ;
        RECT 46.935 187.670 47.450 188.080 ;
        RECT 47.685 187.320 47.855 188.080 ;
        RECT 48.025 187.660 48.195 188.325 ;
        RECT 48.365 188.340 48.555 189.700 ;
        RECT 48.725 189.190 49.000 189.700 ;
        RECT 49.190 189.335 49.720 189.700 ;
        RECT 50.145 189.470 50.475 189.870 ;
        RECT 49.545 189.300 49.720 189.335 ;
        RECT 48.725 189.020 49.005 189.190 ;
        RECT 48.725 188.540 49.000 189.020 ;
        RECT 49.205 188.340 49.375 189.140 ;
        RECT 48.365 188.170 49.375 188.340 ;
        RECT 49.545 189.130 50.475 189.300 ;
        RECT 50.645 189.130 50.900 189.700 ;
        RECT 51.075 189.145 51.365 189.870 ;
        RECT 49.545 188.000 49.715 189.130 ;
        RECT 50.305 188.960 50.475 189.130 ;
        RECT 48.590 187.830 49.715 188.000 ;
        RECT 49.885 188.630 50.080 188.960 ;
        RECT 50.305 188.630 50.560 188.960 ;
        RECT 49.885 187.660 50.055 188.630 ;
        RECT 50.730 188.460 50.900 189.130 ;
        RECT 51.535 189.120 52.745 189.870 ;
        RECT 48.025 187.490 50.055 187.660 ;
        RECT 50.225 187.320 50.395 188.460 ;
        RECT 50.565 187.490 50.900 188.460 ;
        RECT 51.075 187.320 51.365 188.485 ;
        RECT 51.535 188.410 52.055 188.950 ;
        RECT 52.225 188.580 52.745 189.120 ;
        RECT 52.975 189.050 53.185 189.870 ;
        RECT 53.355 189.070 53.685 189.700 ;
        RECT 53.355 188.470 53.605 189.070 ;
        RECT 53.855 189.050 54.085 189.870 ;
        RECT 54.845 189.320 55.015 189.700 ;
        RECT 55.195 189.490 55.525 189.870 ;
        RECT 54.845 189.150 55.510 189.320 ;
        RECT 55.705 189.195 55.965 189.700 ;
        RECT 53.775 188.630 54.105 188.880 ;
        RECT 54.775 188.600 55.105 188.970 ;
        RECT 55.340 188.895 55.510 189.150 ;
        RECT 55.340 188.565 55.625 188.895 ;
        RECT 51.535 187.320 52.745 188.410 ;
        RECT 52.975 187.320 53.185 188.460 ;
        RECT 53.355 187.490 53.685 188.470 ;
        RECT 53.855 187.320 54.085 188.460 ;
        RECT 55.340 188.420 55.510 188.565 ;
        RECT 54.845 188.250 55.510 188.420 ;
        RECT 55.795 188.395 55.965 189.195 ;
        RECT 56.595 189.100 58.265 189.870 ;
        RECT 54.845 187.490 55.015 188.250 ;
        RECT 55.195 187.320 55.525 188.080 ;
        RECT 55.695 187.490 55.965 188.395 ;
        RECT 56.595 188.410 57.345 188.930 ;
        RECT 57.515 188.580 58.265 189.100 ;
        RECT 58.440 189.160 58.695 189.690 ;
        RECT 58.865 189.410 59.170 189.870 ;
        RECT 59.415 189.490 60.485 189.660 ;
        RECT 58.440 188.510 58.650 189.160 ;
        RECT 59.415 189.135 59.735 189.490 ;
        RECT 59.410 188.960 59.735 189.135 ;
        RECT 58.820 188.660 59.735 188.960 ;
        RECT 59.905 188.920 60.145 189.320 ;
        RECT 60.315 189.260 60.485 189.490 ;
        RECT 60.655 189.430 60.845 189.870 ;
        RECT 61.015 189.420 61.965 189.700 ;
        RECT 62.185 189.510 62.535 189.680 ;
        RECT 60.315 189.090 60.845 189.260 ;
        RECT 58.820 188.630 59.560 188.660 ;
        RECT 56.595 187.320 58.265 188.410 ;
        RECT 58.440 187.630 58.695 188.510 ;
        RECT 58.865 187.320 59.170 188.460 ;
        RECT 59.390 188.040 59.560 188.630 ;
        RECT 59.905 188.550 60.445 188.920 ;
        RECT 60.625 188.810 60.845 189.090 ;
        RECT 61.015 188.640 61.185 189.420 ;
        RECT 60.780 188.470 61.185 188.640 ;
        RECT 61.355 188.630 61.705 189.250 ;
        RECT 60.780 188.380 60.950 188.470 ;
        RECT 61.875 188.460 62.085 189.250 ;
        RECT 59.730 188.210 60.950 188.380 ;
        RECT 61.410 188.300 62.085 188.460 ;
        RECT 59.390 187.870 60.190 188.040 ;
        RECT 59.510 187.320 59.840 187.700 ;
        RECT 60.020 187.580 60.190 187.870 ;
        RECT 60.780 187.830 60.950 188.210 ;
        RECT 61.120 188.290 62.085 188.300 ;
        RECT 62.275 189.120 62.535 189.510 ;
        RECT 62.745 189.410 63.075 189.870 ;
        RECT 63.950 189.480 64.805 189.650 ;
        RECT 65.010 189.480 65.505 189.650 ;
        RECT 65.675 189.510 66.005 189.870 ;
        RECT 62.275 188.430 62.445 189.120 ;
        RECT 62.615 188.770 62.785 188.950 ;
        RECT 62.955 188.940 63.745 189.190 ;
        RECT 63.950 188.770 64.120 189.480 ;
        RECT 64.290 188.970 64.645 189.190 ;
        RECT 62.615 188.600 64.305 188.770 ;
        RECT 61.120 188.000 61.580 188.290 ;
        RECT 62.275 188.260 63.775 188.430 ;
        RECT 62.275 188.120 62.445 188.260 ;
        RECT 61.885 187.950 62.445 188.120 ;
        RECT 60.360 187.320 60.610 187.780 ;
        RECT 60.780 187.490 61.650 187.830 ;
        RECT 61.885 187.490 62.055 187.950 ;
        RECT 62.890 187.920 63.965 188.090 ;
        RECT 62.225 187.320 62.595 187.780 ;
        RECT 62.890 187.580 63.060 187.920 ;
        RECT 63.230 187.320 63.560 187.750 ;
        RECT 63.795 187.580 63.965 187.920 ;
        RECT 64.135 187.820 64.305 188.600 ;
        RECT 64.475 188.380 64.645 188.970 ;
        RECT 64.815 188.570 65.165 189.190 ;
        RECT 64.475 187.990 64.940 188.380 ;
        RECT 65.335 188.120 65.505 189.480 ;
        RECT 65.675 188.290 66.135 189.340 ;
        RECT 65.110 187.950 65.505 188.120 ;
        RECT 65.110 187.820 65.280 187.950 ;
        RECT 64.135 187.490 64.815 187.820 ;
        RECT 65.030 187.490 65.280 187.820 ;
        RECT 65.450 187.320 65.700 187.780 ;
        RECT 65.870 187.505 66.195 188.290 ;
        RECT 66.365 187.490 66.535 189.610 ;
        RECT 66.705 189.490 67.035 189.870 ;
        RECT 67.205 189.320 67.460 189.610 ;
        RECT 66.710 189.150 67.460 189.320 ;
        RECT 66.710 188.160 66.940 189.150 ;
        RECT 67.635 189.130 67.955 189.610 ;
        RECT 68.125 189.300 68.355 189.700 ;
        RECT 68.525 189.480 68.875 189.870 ;
        RECT 68.125 189.220 68.635 189.300 ;
        RECT 69.045 189.220 69.375 189.700 ;
        RECT 68.125 189.130 69.375 189.220 ;
        RECT 67.110 188.330 67.460 188.980 ;
        RECT 67.635 188.200 67.805 189.130 ;
        RECT 68.465 189.050 69.375 189.130 ;
        RECT 69.545 189.050 69.715 189.870 ;
        RECT 70.220 189.130 70.685 189.675 ;
        RECT 71.320 189.325 76.665 189.870 ;
        RECT 67.975 188.540 68.145 188.960 ;
        RECT 68.375 188.710 68.975 188.880 ;
        RECT 67.975 188.370 68.635 188.540 ;
        RECT 66.710 187.990 67.460 188.160 ;
        RECT 67.635 188.000 68.295 188.200 ;
        RECT 68.465 188.170 68.635 188.370 ;
        RECT 68.805 188.510 68.975 188.710 ;
        RECT 69.145 188.680 69.840 188.880 ;
        RECT 70.100 188.510 70.345 188.960 ;
        RECT 68.805 188.340 70.345 188.510 ;
        RECT 70.515 188.170 70.685 189.130 ;
        RECT 68.465 188.000 70.685 188.170 ;
        RECT 66.705 187.320 67.035 187.820 ;
        RECT 67.205 187.490 67.460 187.990 ;
        RECT 68.125 187.830 68.295 188.000 ;
        RECT 67.655 187.320 67.955 187.830 ;
        RECT 68.125 187.660 68.505 187.830 ;
        RECT 69.085 187.320 69.715 187.830 ;
        RECT 69.885 187.490 70.215 188.000 ;
        RECT 70.385 187.320 70.685 187.830 ;
        RECT 72.910 187.755 73.260 189.005 ;
        RECT 74.740 188.495 75.080 189.325 ;
        RECT 76.835 189.145 77.125 189.870 ;
        RECT 77.355 189.050 77.565 189.870 ;
        RECT 77.735 189.070 78.065 189.700 ;
        RECT 71.320 187.320 76.665 187.755 ;
        RECT 76.835 187.320 77.125 188.485 ;
        RECT 77.735 188.470 77.985 189.070 ;
        RECT 78.235 189.050 78.465 189.870 ;
        RECT 78.950 189.060 79.195 189.665 ;
        RECT 79.415 189.335 79.925 189.870 ;
        RECT 78.675 188.890 79.905 189.060 ;
        RECT 78.155 188.630 78.485 188.880 ;
        RECT 77.355 187.320 77.565 188.460 ;
        RECT 77.735 187.490 78.065 188.470 ;
        RECT 78.235 187.320 78.465 188.460 ;
        RECT 78.675 188.080 79.015 188.890 ;
        RECT 79.185 188.325 79.935 188.515 ;
        RECT 78.675 187.670 79.190 188.080 ;
        RECT 79.425 187.320 79.595 188.080 ;
        RECT 79.765 187.660 79.935 188.325 ;
        RECT 80.105 188.340 80.295 189.700 ;
        RECT 80.465 189.190 80.740 189.700 ;
        RECT 80.930 189.335 81.460 189.700 ;
        RECT 81.885 189.470 82.215 189.870 ;
        RECT 81.285 189.300 81.460 189.335 ;
        RECT 80.465 189.020 80.745 189.190 ;
        RECT 80.465 188.540 80.740 189.020 ;
        RECT 80.945 188.340 81.115 189.140 ;
        RECT 80.105 188.170 81.115 188.340 ;
        RECT 81.285 189.130 82.215 189.300 ;
        RECT 82.385 189.130 82.640 189.700 ;
        RECT 81.285 188.000 81.455 189.130 ;
        RECT 82.045 188.960 82.215 189.130 ;
        RECT 80.330 187.830 81.455 188.000 ;
        RECT 81.625 188.630 81.820 188.960 ;
        RECT 82.045 188.630 82.300 188.960 ;
        RECT 81.625 187.660 81.795 188.630 ;
        RECT 82.470 188.460 82.640 189.130 ;
        RECT 82.875 189.050 83.085 189.870 ;
        RECT 83.255 189.070 83.585 189.700 ;
        RECT 83.255 188.470 83.505 189.070 ;
        RECT 83.755 189.050 83.985 189.870 ;
        RECT 84.195 189.120 85.405 189.870 ;
        RECT 83.675 188.630 84.005 188.880 ;
        RECT 79.765 187.490 81.795 187.660 ;
        RECT 81.965 187.320 82.135 188.460 ;
        RECT 82.305 187.490 82.640 188.460 ;
        RECT 82.875 187.320 83.085 188.460 ;
        RECT 83.255 187.490 83.585 188.470 ;
        RECT 83.755 187.320 83.985 188.460 ;
        RECT 84.195 188.410 84.715 188.950 ;
        RECT 84.885 188.580 85.405 189.120 ;
        RECT 85.575 189.100 89.085 189.870 ;
        RECT 85.575 188.410 87.265 188.930 ;
        RECT 87.435 188.580 89.085 189.100 ;
        RECT 89.295 189.050 89.525 189.870 ;
        RECT 89.695 189.070 90.025 189.700 ;
        RECT 89.275 188.630 89.605 188.880 ;
        RECT 89.775 188.470 90.025 189.070 ;
        RECT 90.195 189.050 90.405 189.870 ;
        RECT 90.635 189.130 91.020 189.700 ;
        RECT 91.190 189.410 91.515 189.870 ;
        RECT 92.035 189.240 92.315 189.700 ;
        RECT 84.195 187.320 85.405 188.410 ;
        RECT 85.575 187.320 89.085 188.410 ;
        RECT 89.295 187.320 89.525 188.460 ;
        RECT 89.695 187.490 90.025 188.470 ;
        RECT 90.635 188.460 90.915 189.130 ;
        RECT 91.190 189.070 92.315 189.240 ;
        RECT 91.190 188.960 91.640 189.070 ;
        RECT 91.085 188.630 91.640 188.960 ;
        RECT 92.505 188.900 92.905 189.700 ;
        RECT 93.305 189.410 93.575 189.870 ;
        RECT 93.745 189.240 94.030 189.700 ;
        RECT 90.195 187.320 90.405 188.460 ;
        RECT 90.635 187.490 91.020 188.460 ;
        RECT 91.190 188.170 91.640 188.630 ;
        RECT 91.810 188.340 92.905 188.900 ;
        RECT 91.190 187.950 92.315 188.170 ;
        RECT 91.190 187.320 91.515 187.780 ;
        RECT 92.035 187.490 92.315 187.950 ;
        RECT 92.505 187.490 92.905 188.340 ;
        RECT 93.075 189.070 94.030 189.240 ;
        RECT 94.865 189.320 95.035 189.700 ;
        RECT 95.215 189.490 95.545 189.870 ;
        RECT 94.865 189.150 95.530 189.320 ;
        RECT 95.725 189.195 95.985 189.700 ;
        RECT 93.075 188.170 93.285 189.070 ;
        RECT 93.455 188.340 94.145 188.900 ;
        RECT 94.795 188.600 95.125 188.970 ;
        RECT 95.360 188.895 95.530 189.150 ;
        RECT 95.360 188.565 95.645 188.895 ;
        RECT 95.360 188.420 95.530 188.565 ;
        RECT 94.865 188.250 95.530 188.420 ;
        RECT 95.815 188.395 95.985 189.195 ;
        RECT 93.075 187.950 94.030 188.170 ;
        RECT 93.305 187.320 93.575 187.780 ;
        RECT 93.745 187.490 94.030 187.950 ;
        RECT 94.865 187.490 95.035 188.250 ;
        RECT 95.215 187.320 95.545 188.080 ;
        RECT 95.715 187.490 95.985 188.395 ;
        RECT 96.155 189.130 96.540 189.700 ;
        RECT 96.710 189.410 97.035 189.870 ;
        RECT 97.555 189.240 97.835 189.700 ;
        RECT 96.155 188.460 96.435 189.130 ;
        RECT 96.710 189.070 97.835 189.240 ;
        RECT 96.710 188.960 97.160 189.070 ;
        RECT 96.605 188.630 97.160 188.960 ;
        RECT 98.025 188.900 98.425 189.700 ;
        RECT 98.825 189.410 99.095 189.870 ;
        RECT 99.265 189.240 99.550 189.700 ;
        RECT 96.155 187.490 96.540 188.460 ;
        RECT 96.710 188.170 97.160 188.630 ;
        RECT 97.330 188.340 98.425 188.900 ;
        RECT 96.710 187.950 97.835 188.170 ;
        RECT 96.710 187.320 97.035 187.780 ;
        RECT 97.555 187.490 97.835 187.950 ;
        RECT 98.025 187.490 98.425 188.340 ;
        RECT 98.595 189.070 99.550 189.240 ;
        RECT 98.595 188.170 98.805 189.070 ;
        RECT 99.875 189.050 100.105 189.870 ;
        RECT 100.275 189.070 100.605 189.700 ;
        RECT 98.975 188.340 99.665 188.900 ;
        RECT 99.855 188.630 100.185 188.880 ;
        RECT 100.355 188.470 100.605 189.070 ;
        RECT 100.775 189.050 100.985 189.870 ;
        RECT 101.255 189.050 101.485 189.870 ;
        RECT 101.655 189.070 101.985 189.700 ;
        RECT 101.235 188.630 101.565 188.880 ;
        RECT 101.735 188.470 101.985 189.070 ;
        RECT 102.155 189.050 102.365 189.870 ;
        RECT 102.595 189.145 102.885 189.870 ;
        RECT 103.055 189.130 103.440 189.700 ;
        RECT 103.610 189.410 103.935 189.870 ;
        RECT 104.455 189.240 104.735 189.700 ;
        RECT 98.595 187.950 99.550 188.170 ;
        RECT 98.825 187.320 99.095 187.780 ;
        RECT 99.265 187.490 99.550 187.950 ;
        RECT 99.875 187.320 100.105 188.460 ;
        RECT 100.275 187.490 100.605 188.470 ;
        RECT 100.775 187.320 100.985 188.460 ;
        RECT 101.255 187.320 101.485 188.460 ;
        RECT 101.655 187.490 101.985 188.470 ;
        RECT 102.155 187.320 102.365 188.460 ;
        RECT 102.595 187.320 102.885 188.485 ;
        RECT 103.055 188.460 103.335 189.130 ;
        RECT 103.610 189.070 104.735 189.240 ;
        RECT 103.610 188.960 104.060 189.070 ;
        RECT 103.505 188.630 104.060 188.960 ;
        RECT 104.925 188.900 105.325 189.700 ;
        RECT 105.725 189.410 105.995 189.870 ;
        RECT 106.165 189.240 106.450 189.700 ;
        RECT 103.055 187.490 103.440 188.460 ;
        RECT 103.610 188.170 104.060 188.630 ;
        RECT 104.230 188.340 105.325 188.900 ;
        RECT 103.610 187.950 104.735 188.170 ;
        RECT 103.610 187.320 103.935 187.780 ;
        RECT 104.455 187.490 104.735 187.950 ;
        RECT 104.925 187.490 105.325 188.340 ;
        RECT 105.495 189.070 106.450 189.240 ;
        RECT 107.195 189.100 108.865 189.870 ;
        RECT 109.040 189.325 114.385 189.870 ;
        RECT 105.495 188.170 105.705 189.070 ;
        RECT 105.875 188.340 106.565 188.900 ;
        RECT 107.195 188.410 107.945 188.930 ;
        RECT 108.115 188.580 108.865 189.100 ;
        RECT 105.495 187.950 106.450 188.170 ;
        RECT 105.725 187.320 105.995 187.780 ;
        RECT 106.165 187.490 106.450 187.950 ;
        RECT 107.195 187.320 108.865 188.410 ;
        RECT 110.630 187.755 110.980 189.005 ;
        RECT 112.460 188.495 112.800 189.325 ;
        RECT 114.555 189.120 115.765 189.870 ;
        RECT 114.555 188.410 115.075 188.950 ;
        RECT 115.245 188.580 115.765 189.120 ;
        RECT 109.040 187.320 114.385 187.755 ;
        RECT 114.555 187.320 115.765 188.410 ;
        RECT 14.650 187.150 115.850 187.320 ;
        RECT 14.735 186.060 15.945 187.150 ;
        RECT 14.735 185.350 15.255 185.890 ;
        RECT 15.425 185.520 15.945 186.060 ;
        RECT 16.575 186.060 19.165 187.150 ;
        RECT 16.575 185.540 17.785 186.060 ;
        RECT 19.375 186.010 19.605 187.150 ;
        RECT 19.775 186.000 20.105 186.980 ;
        RECT 20.275 186.010 20.485 187.150 ;
        RECT 20.830 186.520 21.115 186.980 ;
        RECT 21.285 186.690 21.555 187.150 ;
        RECT 20.830 186.300 21.785 186.520 ;
        RECT 17.955 185.370 19.165 185.890 ;
        RECT 19.355 185.590 19.685 185.840 ;
        RECT 14.735 184.600 15.945 185.350 ;
        RECT 16.575 184.600 19.165 185.370 ;
        RECT 19.375 184.600 19.605 185.420 ;
        RECT 19.855 185.400 20.105 186.000 ;
        RECT 20.715 185.570 21.405 186.130 ;
        RECT 19.775 184.770 20.105 185.400 ;
        RECT 20.275 184.600 20.485 185.420 ;
        RECT 21.575 185.400 21.785 186.300 ;
        RECT 20.830 185.230 21.785 185.400 ;
        RECT 21.955 186.130 22.355 186.980 ;
        RECT 22.545 186.520 22.825 186.980 ;
        RECT 23.345 186.690 23.670 187.150 ;
        RECT 22.545 186.300 23.670 186.520 ;
        RECT 21.955 185.570 23.050 186.130 ;
        RECT 23.220 185.840 23.670 186.300 ;
        RECT 23.840 186.010 24.225 186.980 ;
        RECT 24.400 186.480 24.655 186.980 ;
        RECT 24.825 186.650 25.155 187.150 ;
        RECT 24.400 186.310 25.150 186.480 ;
        RECT 20.830 184.770 21.115 185.230 ;
        RECT 21.285 184.600 21.555 185.060 ;
        RECT 21.955 184.770 22.355 185.570 ;
        RECT 23.220 185.510 23.775 185.840 ;
        RECT 23.220 185.400 23.670 185.510 ;
        RECT 22.545 185.230 23.670 185.400 ;
        RECT 23.945 185.340 24.225 186.010 ;
        RECT 24.400 185.490 24.750 186.140 ;
        RECT 22.545 184.770 22.825 185.230 ;
        RECT 23.345 184.600 23.670 185.060 ;
        RECT 23.840 184.770 24.225 185.340 ;
        RECT 24.920 185.320 25.150 186.310 ;
        RECT 24.400 185.150 25.150 185.320 ;
        RECT 24.400 184.860 24.655 185.150 ;
        RECT 24.825 184.600 25.155 184.980 ;
        RECT 25.325 184.860 25.495 186.980 ;
        RECT 25.665 186.180 25.990 186.965 ;
        RECT 26.160 186.690 26.410 187.150 ;
        RECT 26.580 186.650 26.830 186.980 ;
        RECT 27.045 186.650 27.725 186.980 ;
        RECT 26.580 186.520 26.750 186.650 ;
        RECT 26.355 186.350 26.750 186.520 ;
        RECT 25.725 185.130 26.185 186.180 ;
        RECT 26.355 184.990 26.525 186.350 ;
        RECT 26.920 186.090 27.385 186.480 ;
        RECT 26.695 185.280 27.045 185.900 ;
        RECT 27.215 185.500 27.385 186.090 ;
        RECT 27.555 185.870 27.725 186.650 ;
        RECT 27.895 186.550 28.065 186.890 ;
        RECT 28.300 186.720 28.630 187.150 ;
        RECT 28.800 186.550 28.970 186.890 ;
        RECT 29.265 186.690 29.635 187.150 ;
        RECT 27.895 186.380 28.970 186.550 ;
        RECT 29.805 186.520 29.975 186.980 ;
        RECT 30.210 186.640 31.080 186.980 ;
        RECT 31.250 186.690 31.500 187.150 ;
        RECT 29.415 186.350 29.975 186.520 ;
        RECT 29.415 186.210 29.585 186.350 ;
        RECT 28.085 186.040 29.585 186.210 ;
        RECT 30.280 186.180 30.740 186.470 ;
        RECT 27.555 185.700 29.245 185.870 ;
        RECT 27.215 185.280 27.570 185.500 ;
        RECT 27.740 184.990 27.910 185.700 ;
        RECT 28.115 185.280 28.905 185.530 ;
        RECT 29.075 185.520 29.245 185.700 ;
        RECT 29.415 185.350 29.585 186.040 ;
        RECT 25.855 184.600 26.185 184.960 ;
        RECT 26.355 184.820 26.850 184.990 ;
        RECT 27.055 184.820 27.910 184.990 ;
        RECT 28.785 184.600 29.115 185.060 ;
        RECT 29.325 184.960 29.585 185.350 ;
        RECT 29.775 186.170 30.740 186.180 ;
        RECT 30.910 186.260 31.080 186.640 ;
        RECT 31.670 186.600 31.840 186.890 ;
        RECT 32.020 186.770 32.350 187.150 ;
        RECT 31.670 186.430 32.470 186.600 ;
        RECT 29.775 186.010 30.450 186.170 ;
        RECT 30.910 186.090 32.130 186.260 ;
        RECT 29.775 185.220 29.985 186.010 ;
        RECT 30.910 186.000 31.080 186.090 ;
        RECT 30.155 185.220 30.505 185.840 ;
        RECT 30.675 185.830 31.080 186.000 ;
        RECT 30.675 185.050 30.845 185.830 ;
        RECT 31.015 185.380 31.235 185.660 ;
        RECT 31.415 185.550 31.955 185.920 ;
        RECT 32.300 185.840 32.470 186.430 ;
        RECT 32.690 186.010 32.995 187.150 ;
        RECT 33.165 185.960 33.420 186.840 ;
        RECT 34.720 186.180 35.050 186.980 ;
        RECT 35.220 186.350 35.550 187.150 ;
        RECT 35.850 186.180 36.180 186.980 ;
        RECT 36.825 186.350 37.075 187.150 ;
        RECT 34.720 186.010 37.155 186.180 ;
        RECT 37.345 186.010 37.515 187.150 ;
        RECT 37.685 186.010 38.025 186.980 ;
        RECT 32.300 185.810 33.040 185.840 ;
        RECT 31.015 185.210 31.545 185.380 ;
        RECT 29.325 184.790 29.675 184.960 ;
        RECT 29.895 184.770 30.845 185.050 ;
        RECT 31.015 184.600 31.205 185.040 ;
        RECT 31.375 184.980 31.545 185.210 ;
        RECT 31.715 185.150 31.955 185.550 ;
        RECT 32.125 185.510 33.040 185.810 ;
        RECT 32.125 185.335 32.450 185.510 ;
        RECT 32.125 184.980 32.445 185.335 ;
        RECT 33.210 185.310 33.420 185.960 ;
        RECT 34.515 185.590 34.865 185.840 ;
        RECT 35.050 185.380 35.220 186.010 ;
        RECT 35.390 185.590 35.720 185.790 ;
        RECT 35.890 185.590 36.220 185.790 ;
        RECT 36.390 185.590 36.810 185.790 ;
        RECT 36.985 185.760 37.155 186.010 ;
        RECT 36.985 185.590 37.680 185.760 ;
        RECT 31.375 184.810 32.445 184.980 ;
        RECT 32.690 184.600 32.995 185.060 ;
        RECT 33.165 184.780 33.420 185.310 ;
        RECT 34.720 184.770 35.220 185.380 ;
        RECT 35.850 185.250 37.075 185.420 ;
        RECT 37.850 185.400 38.025 186.010 ;
        RECT 38.195 185.985 38.485 187.150 ;
        RECT 39.120 186.010 39.455 186.980 ;
        RECT 39.625 186.010 39.795 187.150 ;
        RECT 39.965 186.810 41.995 186.980 ;
        RECT 35.850 184.770 36.180 185.250 ;
        RECT 36.350 184.600 36.575 185.060 ;
        RECT 36.745 184.770 37.075 185.250 ;
        RECT 37.265 184.600 37.515 185.400 ;
        RECT 37.685 184.770 38.025 185.400 ;
        RECT 39.120 185.340 39.290 186.010 ;
        RECT 39.965 185.840 40.135 186.810 ;
        RECT 39.460 185.510 39.715 185.840 ;
        RECT 39.940 185.510 40.135 185.840 ;
        RECT 40.305 186.470 41.430 186.640 ;
        RECT 39.545 185.340 39.715 185.510 ;
        RECT 40.305 185.340 40.475 186.470 ;
        RECT 38.195 184.600 38.485 185.325 ;
        RECT 39.120 184.770 39.375 185.340 ;
        RECT 39.545 185.170 40.475 185.340 ;
        RECT 40.645 186.130 41.655 186.300 ;
        RECT 40.645 185.330 40.815 186.130 ;
        RECT 41.020 185.790 41.295 185.930 ;
        RECT 41.015 185.620 41.295 185.790 ;
        RECT 40.300 185.135 40.475 185.170 ;
        RECT 39.545 184.600 39.875 185.000 ;
        RECT 40.300 184.770 40.830 185.135 ;
        RECT 41.020 184.770 41.295 185.620 ;
        RECT 41.465 184.770 41.655 186.130 ;
        RECT 41.825 186.145 41.995 186.810 ;
        RECT 42.165 186.390 42.335 187.150 ;
        RECT 42.570 186.390 43.085 186.800 ;
        RECT 41.825 185.955 42.575 186.145 ;
        RECT 42.745 185.580 43.085 186.390 ;
        RECT 41.855 185.410 43.085 185.580 ;
        RECT 43.260 185.960 43.515 186.840 ;
        RECT 43.685 186.010 43.990 187.150 ;
        RECT 44.330 186.770 44.660 187.150 ;
        RECT 44.840 186.600 45.010 186.890 ;
        RECT 45.180 186.690 45.430 187.150 ;
        RECT 44.210 186.430 45.010 186.600 ;
        RECT 45.600 186.640 46.470 186.980 ;
        RECT 41.835 184.600 42.345 185.135 ;
        RECT 42.565 184.805 42.810 185.410 ;
        RECT 43.260 185.310 43.470 185.960 ;
        RECT 44.210 185.840 44.380 186.430 ;
        RECT 45.600 186.260 45.770 186.640 ;
        RECT 46.705 186.520 46.875 186.980 ;
        RECT 47.045 186.690 47.415 187.150 ;
        RECT 47.710 186.550 47.880 186.890 ;
        RECT 48.050 186.720 48.380 187.150 ;
        RECT 48.615 186.550 48.785 186.890 ;
        RECT 44.550 186.090 45.770 186.260 ;
        RECT 45.940 186.180 46.400 186.470 ;
        RECT 46.705 186.350 47.265 186.520 ;
        RECT 47.710 186.380 48.785 186.550 ;
        RECT 48.955 186.650 49.635 186.980 ;
        RECT 49.850 186.650 50.100 186.980 ;
        RECT 50.270 186.690 50.520 187.150 ;
        RECT 47.095 186.210 47.265 186.350 ;
        RECT 45.940 186.170 46.905 186.180 ;
        RECT 45.600 186.000 45.770 186.090 ;
        RECT 46.230 186.010 46.905 186.170 ;
        RECT 43.640 185.810 44.380 185.840 ;
        RECT 43.640 185.510 44.555 185.810 ;
        RECT 44.230 185.335 44.555 185.510 ;
        RECT 43.260 184.780 43.515 185.310 ;
        RECT 43.685 184.600 43.990 185.060 ;
        RECT 44.235 184.980 44.555 185.335 ;
        RECT 44.725 185.550 45.265 185.920 ;
        RECT 45.600 185.830 46.005 186.000 ;
        RECT 44.725 185.150 44.965 185.550 ;
        RECT 45.445 185.380 45.665 185.660 ;
        RECT 45.135 185.210 45.665 185.380 ;
        RECT 45.135 184.980 45.305 185.210 ;
        RECT 45.835 185.050 46.005 185.830 ;
        RECT 46.175 185.220 46.525 185.840 ;
        RECT 46.695 185.220 46.905 186.010 ;
        RECT 47.095 186.040 48.595 186.210 ;
        RECT 47.095 185.350 47.265 186.040 ;
        RECT 48.955 185.870 49.125 186.650 ;
        RECT 49.930 186.520 50.100 186.650 ;
        RECT 47.435 185.700 49.125 185.870 ;
        RECT 49.295 186.090 49.760 186.480 ;
        RECT 49.930 186.350 50.325 186.520 ;
        RECT 47.435 185.520 47.605 185.700 ;
        RECT 44.235 184.810 45.305 184.980 ;
        RECT 45.475 184.600 45.665 185.040 ;
        RECT 45.835 184.770 46.785 185.050 ;
        RECT 47.095 184.960 47.355 185.350 ;
        RECT 47.775 185.280 48.565 185.530 ;
        RECT 47.005 184.790 47.355 184.960 ;
        RECT 47.565 184.600 47.895 185.060 ;
        RECT 48.770 184.990 48.940 185.700 ;
        RECT 49.295 185.500 49.465 186.090 ;
        RECT 49.110 185.280 49.465 185.500 ;
        RECT 49.635 185.280 49.985 185.900 ;
        RECT 50.155 184.990 50.325 186.350 ;
        RECT 50.690 186.180 51.015 186.965 ;
        RECT 50.495 185.130 50.955 186.180 ;
        RECT 48.770 184.820 49.625 184.990 ;
        RECT 49.830 184.820 50.325 184.990 ;
        RECT 50.495 184.600 50.825 184.960 ;
        RECT 51.185 184.860 51.355 186.980 ;
        RECT 51.525 186.650 51.855 187.150 ;
        RECT 52.025 186.480 52.280 186.980 ;
        RECT 52.920 186.715 58.265 187.150 ;
        RECT 58.440 186.715 63.785 187.150 ;
        RECT 51.530 186.310 52.280 186.480 ;
        RECT 51.530 185.320 51.760 186.310 ;
        RECT 51.930 185.490 52.280 186.140 ;
        RECT 54.510 185.465 54.860 186.715 ;
        RECT 51.530 185.150 52.280 185.320 ;
        RECT 51.525 184.600 51.855 184.980 ;
        RECT 52.025 184.860 52.280 185.150 ;
        RECT 56.340 185.145 56.680 185.975 ;
        RECT 60.030 185.465 60.380 186.715 ;
        RECT 63.955 185.985 64.245 187.150 ;
        RECT 64.420 186.715 69.765 187.150 ;
        RECT 69.940 186.715 75.285 187.150 ;
        RECT 61.860 185.145 62.200 185.975 ;
        RECT 66.010 185.465 66.360 186.715 ;
        RECT 52.920 184.600 58.265 185.145 ;
        RECT 58.440 184.600 63.785 185.145 ;
        RECT 63.955 184.600 64.245 185.325 ;
        RECT 67.840 185.145 68.180 185.975 ;
        RECT 71.530 185.465 71.880 186.715 ;
        RECT 75.830 186.170 76.085 186.840 ;
        RECT 76.265 186.350 76.550 187.150 ;
        RECT 76.730 186.430 77.060 186.940 ;
        RECT 73.360 185.145 73.700 185.975 ;
        RECT 75.830 185.310 76.010 186.170 ;
        RECT 76.730 185.840 76.980 186.430 ;
        RECT 77.330 186.280 77.500 186.890 ;
        RECT 77.670 186.460 78.000 187.150 ;
        RECT 78.230 186.600 78.470 186.890 ;
        RECT 78.670 186.770 79.090 187.150 ;
        RECT 79.270 186.680 79.900 186.930 ;
        RECT 80.370 186.770 80.700 187.150 ;
        RECT 79.270 186.600 79.440 186.680 ;
        RECT 80.870 186.600 81.040 186.890 ;
        RECT 81.220 186.770 81.600 187.150 ;
        RECT 81.840 186.765 82.670 186.935 ;
        RECT 78.230 186.430 79.440 186.600 ;
        RECT 76.180 185.510 76.980 185.840 ;
        RECT 64.420 184.600 69.765 185.145 ;
        RECT 69.940 184.600 75.285 185.145 ;
        RECT 75.830 185.110 76.085 185.310 ;
        RECT 75.745 184.940 76.085 185.110 ;
        RECT 75.830 184.780 76.085 184.940 ;
        RECT 76.265 184.600 76.550 185.060 ;
        RECT 76.730 184.860 76.980 185.510 ;
        RECT 77.180 186.260 77.500 186.280 ;
        RECT 77.180 186.090 79.100 186.260 ;
        RECT 77.180 185.195 77.370 186.090 ;
        RECT 79.270 185.920 79.440 186.430 ;
        RECT 79.610 186.170 80.130 186.480 ;
        RECT 77.540 185.750 79.440 185.920 ;
        RECT 77.540 185.690 77.870 185.750 ;
        RECT 78.020 185.520 78.350 185.580 ;
        RECT 77.690 185.250 78.350 185.520 ;
        RECT 77.180 184.865 77.500 185.195 ;
        RECT 77.680 184.600 78.340 185.080 ;
        RECT 78.540 184.990 78.710 185.750 ;
        RECT 79.610 185.580 79.790 185.990 ;
        RECT 78.880 185.410 79.210 185.530 ;
        RECT 79.960 185.410 80.130 186.170 ;
        RECT 78.880 185.240 80.130 185.410 ;
        RECT 80.300 186.350 81.670 186.600 ;
        RECT 80.300 185.580 80.490 186.350 ;
        RECT 81.420 186.090 81.670 186.350 ;
        RECT 80.660 185.920 80.910 186.080 ;
        RECT 81.840 185.920 82.010 186.765 ;
        RECT 82.905 186.480 83.075 186.980 ;
        RECT 83.245 186.650 83.575 187.150 ;
        RECT 82.180 186.090 82.680 186.470 ;
        RECT 82.905 186.310 83.600 186.480 ;
        RECT 80.660 185.750 82.010 185.920 ;
        RECT 81.590 185.710 82.010 185.750 ;
        RECT 80.300 185.240 80.720 185.580 ;
        RECT 81.010 185.250 81.420 185.580 ;
        RECT 78.540 184.820 79.390 184.990 ;
        RECT 79.950 184.600 80.270 185.060 ;
        RECT 80.470 184.810 80.720 185.240 ;
        RECT 81.010 184.600 81.420 185.040 ;
        RECT 81.590 184.980 81.760 185.710 ;
        RECT 81.930 185.160 82.280 185.530 ;
        RECT 82.460 185.220 82.680 186.090 ;
        RECT 82.850 185.520 83.260 186.140 ;
        RECT 83.430 185.340 83.600 186.310 ;
        RECT 82.905 185.150 83.600 185.340 ;
        RECT 81.590 184.780 82.605 184.980 ;
        RECT 82.905 184.820 83.075 185.150 ;
        RECT 83.245 184.600 83.575 184.980 ;
        RECT 83.790 184.860 84.015 186.980 ;
        RECT 84.185 186.650 84.515 187.150 ;
        RECT 84.685 186.480 84.855 186.980 ;
        RECT 84.190 186.310 84.855 186.480 ;
        RECT 84.190 185.320 84.420 186.310 ;
        RECT 84.590 185.490 84.940 186.140 ;
        RECT 85.115 186.075 85.385 186.980 ;
        RECT 85.555 186.390 85.885 187.150 ;
        RECT 86.065 186.220 86.235 186.980 ;
        RECT 84.190 185.150 84.855 185.320 ;
        RECT 84.185 184.600 84.515 184.980 ;
        RECT 84.685 184.860 84.855 185.150 ;
        RECT 85.115 185.275 85.285 186.075 ;
        RECT 85.570 186.050 86.235 186.220 ;
        RECT 86.495 186.060 87.705 187.150 ;
        RECT 85.570 185.905 85.740 186.050 ;
        RECT 85.455 185.575 85.740 185.905 ;
        RECT 85.570 185.320 85.740 185.575 ;
        RECT 85.975 185.500 86.305 185.870 ;
        RECT 86.495 185.520 87.015 186.060 ;
        RECT 87.915 186.010 88.145 187.150 ;
        RECT 88.315 186.000 88.645 186.980 ;
        RECT 88.815 186.010 89.025 187.150 ;
        RECT 87.185 185.350 87.705 185.890 ;
        RECT 87.895 185.590 88.225 185.840 ;
        RECT 85.115 184.770 85.375 185.275 ;
        RECT 85.570 185.150 86.235 185.320 ;
        RECT 85.555 184.600 85.885 184.980 ;
        RECT 86.065 184.770 86.235 185.150 ;
        RECT 86.495 184.600 87.705 185.350 ;
        RECT 87.915 184.600 88.145 185.420 ;
        RECT 88.395 185.400 88.645 186.000 ;
        RECT 89.715 185.985 90.005 187.150 ;
        RECT 90.180 185.960 90.435 186.840 ;
        RECT 90.605 186.010 90.910 187.150 ;
        RECT 91.250 186.770 91.580 187.150 ;
        RECT 91.760 186.600 91.930 186.890 ;
        RECT 92.100 186.690 92.350 187.150 ;
        RECT 91.130 186.430 91.930 186.600 ;
        RECT 92.520 186.640 93.390 186.980 ;
        RECT 88.315 184.770 88.645 185.400 ;
        RECT 88.815 184.600 89.025 185.420 ;
        RECT 89.715 184.600 90.005 185.325 ;
        RECT 90.180 185.310 90.390 185.960 ;
        RECT 91.130 185.840 91.300 186.430 ;
        RECT 92.520 186.260 92.690 186.640 ;
        RECT 93.625 186.520 93.795 186.980 ;
        RECT 93.965 186.690 94.335 187.150 ;
        RECT 94.630 186.550 94.800 186.890 ;
        RECT 94.970 186.720 95.300 187.150 ;
        RECT 95.535 186.550 95.705 186.890 ;
        RECT 91.470 186.090 92.690 186.260 ;
        RECT 92.860 186.180 93.320 186.470 ;
        RECT 93.625 186.350 94.185 186.520 ;
        RECT 94.630 186.380 95.705 186.550 ;
        RECT 95.875 186.650 96.555 186.980 ;
        RECT 96.770 186.650 97.020 186.980 ;
        RECT 97.190 186.690 97.440 187.150 ;
        RECT 94.015 186.210 94.185 186.350 ;
        RECT 92.860 186.170 93.825 186.180 ;
        RECT 92.520 186.000 92.690 186.090 ;
        RECT 93.150 186.010 93.825 186.170 ;
        RECT 90.560 185.810 91.300 185.840 ;
        RECT 90.560 185.510 91.475 185.810 ;
        RECT 91.150 185.335 91.475 185.510 ;
        RECT 90.180 184.780 90.435 185.310 ;
        RECT 90.605 184.600 90.910 185.060 ;
        RECT 91.155 184.980 91.475 185.335 ;
        RECT 91.645 185.550 92.185 185.920 ;
        RECT 92.520 185.830 92.925 186.000 ;
        RECT 91.645 185.150 91.885 185.550 ;
        RECT 92.365 185.380 92.585 185.660 ;
        RECT 92.055 185.210 92.585 185.380 ;
        RECT 92.055 184.980 92.225 185.210 ;
        RECT 92.755 185.050 92.925 185.830 ;
        RECT 93.095 185.220 93.445 185.840 ;
        RECT 93.615 185.220 93.825 186.010 ;
        RECT 94.015 186.040 95.515 186.210 ;
        RECT 94.015 185.350 94.185 186.040 ;
        RECT 95.875 185.870 96.045 186.650 ;
        RECT 96.850 186.520 97.020 186.650 ;
        RECT 94.355 185.700 96.045 185.870 ;
        RECT 96.215 186.090 96.680 186.480 ;
        RECT 96.850 186.350 97.245 186.520 ;
        RECT 94.355 185.520 94.525 185.700 ;
        RECT 91.155 184.810 92.225 184.980 ;
        RECT 92.395 184.600 92.585 185.040 ;
        RECT 92.755 184.770 93.705 185.050 ;
        RECT 94.015 184.960 94.275 185.350 ;
        RECT 94.695 185.280 95.485 185.530 ;
        RECT 93.925 184.790 94.275 184.960 ;
        RECT 94.485 184.600 94.815 185.060 ;
        RECT 95.690 184.990 95.860 185.700 ;
        RECT 96.215 185.500 96.385 186.090 ;
        RECT 96.030 185.280 96.385 185.500 ;
        RECT 96.555 185.280 96.905 185.900 ;
        RECT 97.075 184.990 97.245 186.350 ;
        RECT 97.610 186.180 97.935 186.965 ;
        RECT 97.415 185.130 97.875 186.180 ;
        RECT 95.690 184.820 96.545 184.990 ;
        RECT 96.750 184.820 97.245 184.990 ;
        RECT 97.415 184.600 97.745 184.960 ;
        RECT 98.105 184.860 98.275 186.980 ;
        RECT 98.445 186.650 98.775 187.150 ;
        RECT 98.945 186.480 99.200 186.980 ;
        RECT 98.450 186.310 99.200 186.480 ;
        RECT 98.450 185.320 98.680 186.310 ;
        RECT 98.850 185.490 99.200 186.140 ;
        RECT 99.375 186.010 99.760 186.980 ;
        RECT 99.930 186.690 100.255 187.150 ;
        RECT 100.775 186.520 101.055 186.980 ;
        RECT 99.930 186.300 101.055 186.520 ;
        RECT 99.375 185.340 99.655 186.010 ;
        RECT 99.930 185.840 100.380 186.300 ;
        RECT 101.245 186.130 101.645 186.980 ;
        RECT 102.045 186.690 102.315 187.150 ;
        RECT 102.485 186.520 102.770 186.980 ;
        RECT 99.825 185.510 100.380 185.840 ;
        RECT 100.550 185.570 101.645 186.130 ;
        RECT 99.930 185.400 100.380 185.510 ;
        RECT 98.450 185.150 99.200 185.320 ;
        RECT 98.445 184.600 98.775 184.980 ;
        RECT 98.945 184.860 99.200 185.150 ;
        RECT 99.375 184.770 99.760 185.340 ;
        RECT 99.930 185.230 101.055 185.400 ;
        RECT 99.930 184.600 100.255 185.060 ;
        RECT 100.775 184.770 101.055 185.230 ;
        RECT 101.245 184.770 101.645 185.570 ;
        RECT 101.815 186.300 102.770 186.520 ;
        RECT 101.815 185.400 102.025 186.300 ;
        RECT 102.195 185.570 102.885 186.130 ;
        RECT 103.980 185.960 104.235 186.840 ;
        RECT 104.405 186.010 104.710 187.150 ;
        RECT 105.050 186.770 105.380 187.150 ;
        RECT 105.560 186.600 105.730 186.890 ;
        RECT 105.900 186.690 106.150 187.150 ;
        RECT 104.930 186.430 105.730 186.600 ;
        RECT 106.320 186.640 107.190 186.980 ;
        RECT 101.815 185.230 102.770 185.400 ;
        RECT 102.045 184.600 102.315 185.060 ;
        RECT 102.485 184.770 102.770 185.230 ;
        RECT 103.980 185.310 104.190 185.960 ;
        RECT 104.930 185.840 105.100 186.430 ;
        RECT 106.320 186.260 106.490 186.640 ;
        RECT 107.425 186.520 107.595 186.980 ;
        RECT 107.765 186.690 108.135 187.150 ;
        RECT 108.430 186.550 108.600 186.890 ;
        RECT 108.770 186.720 109.100 187.150 ;
        RECT 109.335 186.550 109.505 186.890 ;
        RECT 105.270 186.090 106.490 186.260 ;
        RECT 106.660 186.180 107.120 186.470 ;
        RECT 107.425 186.350 107.985 186.520 ;
        RECT 108.430 186.380 109.505 186.550 ;
        RECT 109.675 186.650 110.355 186.980 ;
        RECT 110.570 186.650 110.820 186.980 ;
        RECT 110.990 186.690 111.240 187.150 ;
        RECT 107.815 186.210 107.985 186.350 ;
        RECT 106.660 186.170 107.625 186.180 ;
        RECT 106.320 186.000 106.490 186.090 ;
        RECT 106.950 186.010 107.625 186.170 ;
        RECT 104.360 185.810 105.100 185.840 ;
        RECT 104.360 185.510 105.275 185.810 ;
        RECT 104.950 185.335 105.275 185.510 ;
        RECT 103.980 184.780 104.235 185.310 ;
        RECT 104.405 184.600 104.710 185.060 ;
        RECT 104.955 184.980 105.275 185.335 ;
        RECT 105.445 185.550 105.985 185.920 ;
        RECT 106.320 185.830 106.725 186.000 ;
        RECT 105.445 185.150 105.685 185.550 ;
        RECT 106.165 185.380 106.385 185.660 ;
        RECT 105.855 185.210 106.385 185.380 ;
        RECT 105.855 184.980 106.025 185.210 ;
        RECT 106.555 185.050 106.725 185.830 ;
        RECT 106.895 185.220 107.245 185.840 ;
        RECT 107.415 185.220 107.625 186.010 ;
        RECT 107.815 186.040 109.315 186.210 ;
        RECT 107.815 185.350 107.985 186.040 ;
        RECT 109.675 185.870 109.845 186.650 ;
        RECT 110.650 186.520 110.820 186.650 ;
        RECT 108.155 185.700 109.845 185.870 ;
        RECT 110.015 186.090 110.480 186.480 ;
        RECT 110.650 186.350 111.045 186.520 ;
        RECT 108.155 185.520 108.325 185.700 ;
        RECT 104.955 184.810 106.025 184.980 ;
        RECT 106.195 184.600 106.385 185.040 ;
        RECT 106.555 184.770 107.505 185.050 ;
        RECT 107.815 184.960 108.075 185.350 ;
        RECT 108.495 185.280 109.285 185.530 ;
        RECT 107.725 184.790 108.075 184.960 ;
        RECT 108.285 184.600 108.615 185.060 ;
        RECT 109.490 184.990 109.660 185.700 ;
        RECT 110.015 185.500 110.185 186.090 ;
        RECT 109.830 185.280 110.185 185.500 ;
        RECT 110.355 185.280 110.705 185.900 ;
        RECT 110.875 184.990 111.045 186.350 ;
        RECT 111.410 186.180 111.735 186.965 ;
        RECT 111.215 185.130 111.675 186.180 ;
        RECT 109.490 184.820 110.345 184.990 ;
        RECT 110.550 184.820 111.045 184.990 ;
        RECT 111.215 184.600 111.545 184.960 ;
        RECT 111.905 184.860 112.075 186.980 ;
        RECT 112.245 186.650 112.575 187.150 ;
        RECT 112.745 186.480 113.000 186.980 ;
        RECT 112.250 186.310 113.000 186.480 ;
        RECT 112.250 185.320 112.480 186.310 ;
        RECT 112.650 185.490 113.000 186.140 ;
        RECT 113.175 186.060 114.385 187.150 ;
        RECT 114.555 186.060 115.765 187.150 ;
        RECT 113.175 185.520 113.695 186.060 ;
        RECT 113.865 185.350 114.385 185.890 ;
        RECT 114.555 185.520 115.075 186.060 ;
        RECT 115.245 185.350 115.765 185.890 ;
        RECT 112.250 185.150 113.000 185.320 ;
        RECT 112.245 184.600 112.575 184.980 ;
        RECT 112.745 184.860 113.000 185.150 ;
        RECT 113.175 184.600 114.385 185.350 ;
        RECT 114.555 184.600 115.765 185.350 ;
        RECT 14.650 184.430 115.850 184.600 ;
        RECT 14.735 183.680 15.945 184.430 ;
        RECT 14.735 183.140 15.255 183.680 ;
        RECT 16.115 183.660 17.785 184.430 ;
        RECT 15.425 182.970 15.945 183.510 ;
        RECT 14.735 181.880 15.945 182.970 ;
        RECT 16.115 182.970 16.865 183.490 ;
        RECT 17.035 183.140 17.785 183.660 ;
        RECT 18.070 183.800 18.355 184.260 ;
        RECT 18.525 183.970 18.795 184.430 ;
        RECT 18.070 183.630 19.025 183.800 ;
        RECT 16.115 181.880 17.785 182.970 ;
        RECT 17.955 182.900 18.645 183.460 ;
        RECT 18.815 182.730 19.025 183.630 ;
        RECT 18.070 182.510 19.025 182.730 ;
        RECT 19.195 183.460 19.595 184.260 ;
        RECT 19.785 183.800 20.065 184.260 ;
        RECT 20.585 183.970 20.910 184.430 ;
        RECT 19.785 183.630 20.910 183.800 ;
        RECT 21.080 183.690 21.465 184.260 ;
        RECT 20.460 183.520 20.910 183.630 ;
        RECT 19.195 182.900 20.290 183.460 ;
        RECT 20.460 183.190 21.015 183.520 ;
        RECT 18.070 182.050 18.355 182.510 ;
        RECT 18.525 181.880 18.795 182.340 ;
        RECT 19.195 182.050 19.595 182.900 ;
        RECT 20.460 182.730 20.910 183.190 ;
        RECT 21.185 183.020 21.465 183.690 ;
        RECT 21.750 183.800 22.035 184.260 ;
        RECT 22.205 183.970 22.475 184.430 ;
        RECT 21.750 183.630 22.705 183.800 ;
        RECT 19.785 182.510 20.910 182.730 ;
        RECT 19.785 182.050 20.065 182.510 ;
        RECT 20.585 181.880 20.910 182.340 ;
        RECT 21.080 182.050 21.465 183.020 ;
        RECT 21.635 182.900 22.325 183.460 ;
        RECT 22.495 182.730 22.705 183.630 ;
        RECT 21.750 182.510 22.705 182.730 ;
        RECT 22.875 183.460 23.275 184.260 ;
        RECT 23.465 183.800 23.745 184.260 ;
        RECT 24.265 183.970 24.590 184.430 ;
        RECT 23.465 183.630 24.590 183.800 ;
        RECT 24.760 183.690 25.145 184.260 ;
        RECT 25.315 183.705 25.605 184.430 ;
        RECT 24.140 183.520 24.590 183.630 ;
        RECT 22.875 182.900 23.970 183.460 ;
        RECT 24.140 183.190 24.695 183.520 ;
        RECT 21.750 182.050 22.035 182.510 ;
        RECT 22.205 181.880 22.475 182.340 ;
        RECT 22.875 182.050 23.275 182.900 ;
        RECT 24.140 182.730 24.590 183.190 ;
        RECT 24.865 183.020 25.145 183.690 ;
        RECT 25.835 183.610 26.045 184.430 ;
        RECT 26.215 183.630 26.545 184.260 ;
        RECT 23.465 182.510 24.590 182.730 ;
        RECT 23.465 182.050 23.745 182.510 ;
        RECT 24.265 181.880 24.590 182.340 ;
        RECT 24.760 182.050 25.145 183.020 ;
        RECT 25.315 181.880 25.605 183.045 ;
        RECT 26.215 183.030 26.465 183.630 ;
        RECT 26.715 183.610 26.945 184.430 ;
        RECT 27.155 183.680 28.365 184.430 ;
        RECT 26.635 183.190 26.965 183.440 ;
        RECT 25.835 181.880 26.045 183.020 ;
        RECT 26.215 182.050 26.545 183.030 ;
        RECT 26.715 181.880 26.945 183.020 ;
        RECT 27.155 182.970 27.675 183.510 ;
        RECT 27.845 183.140 28.365 183.680 ;
        RECT 28.540 183.690 28.795 184.260 ;
        RECT 28.965 184.030 29.295 184.430 ;
        RECT 29.720 183.895 30.250 184.260 ;
        RECT 29.720 183.860 29.895 183.895 ;
        RECT 28.965 183.690 29.895 183.860 ;
        RECT 30.440 183.750 30.715 184.260 ;
        RECT 28.540 183.020 28.710 183.690 ;
        RECT 28.965 183.520 29.135 183.690 ;
        RECT 28.880 183.190 29.135 183.520 ;
        RECT 29.360 183.190 29.555 183.520 ;
        RECT 27.155 181.880 28.365 182.970 ;
        RECT 28.540 182.050 28.875 183.020 ;
        RECT 29.045 181.880 29.215 183.020 ;
        RECT 29.385 182.220 29.555 183.190 ;
        RECT 29.725 182.560 29.895 183.690 ;
        RECT 30.065 182.900 30.235 183.700 ;
        RECT 30.435 183.580 30.715 183.750 ;
        RECT 30.440 183.100 30.715 183.580 ;
        RECT 30.885 182.900 31.075 184.260 ;
        RECT 31.255 183.895 31.765 184.430 ;
        RECT 31.985 183.620 32.230 184.225 ;
        RECT 33.600 183.720 33.855 184.250 ;
        RECT 34.025 183.970 34.330 184.430 ;
        RECT 34.575 184.050 35.645 184.220 ;
        RECT 31.275 183.450 32.505 183.620 ;
        RECT 30.065 182.730 31.075 182.900 ;
        RECT 31.245 182.885 31.995 183.075 ;
        RECT 29.725 182.390 30.850 182.560 ;
        RECT 31.245 182.220 31.415 182.885 ;
        RECT 32.165 182.640 32.505 183.450 ;
        RECT 29.385 182.050 31.415 182.220 ;
        RECT 31.585 181.880 31.755 182.640 ;
        RECT 31.990 182.230 32.505 182.640 ;
        RECT 33.600 183.070 33.810 183.720 ;
        RECT 34.575 183.695 34.895 184.050 ;
        RECT 34.570 183.520 34.895 183.695 ;
        RECT 33.980 183.220 34.895 183.520 ;
        RECT 35.065 183.480 35.305 183.880 ;
        RECT 35.475 183.820 35.645 184.050 ;
        RECT 35.815 183.990 36.005 184.430 ;
        RECT 36.175 183.980 37.125 184.260 ;
        RECT 37.345 184.070 37.695 184.240 ;
        RECT 35.475 183.650 36.005 183.820 ;
        RECT 33.980 183.190 34.720 183.220 ;
        RECT 33.600 182.190 33.855 183.070 ;
        RECT 34.025 181.880 34.330 183.020 ;
        RECT 34.550 182.600 34.720 183.190 ;
        RECT 35.065 183.110 35.605 183.480 ;
        RECT 35.785 183.370 36.005 183.650 ;
        RECT 36.175 183.200 36.345 183.980 ;
        RECT 35.940 183.030 36.345 183.200 ;
        RECT 36.515 183.190 36.865 183.810 ;
        RECT 35.940 182.940 36.110 183.030 ;
        RECT 37.035 183.020 37.245 183.810 ;
        RECT 34.890 182.770 36.110 182.940 ;
        RECT 36.570 182.860 37.245 183.020 ;
        RECT 34.550 182.430 35.350 182.600 ;
        RECT 34.670 181.880 35.000 182.260 ;
        RECT 35.180 182.140 35.350 182.430 ;
        RECT 35.940 182.390 36.110 182.770 ;
        RECT 36.280 182.850 37.245 182.860 ;
        RECT 37.435 183.680 37.695 184.070 ;
        RECT 37.905 183.970 38.235 184.430 ;
        RECT 39.110 184.040 39.965 184.210 ;
        RECT 40.170 184.040 40.665 184.210 ;
        RECT 40.835 184.070 41.165 184.430 ;
        RECT 37.435 182.990 37.605 183.680 ;
        RECT 37.775 183.330 37.945 183.510 ;
        RECT 38.115 183.500 38.905 183.750 ;
        RECT 39.110 183.330 39.280 184.040 ;
        RECT 39.450 183.530 39.805 183.750 ;
        RECT 37.775 183.160 39.465 183.330 ;
        RECT 36.280 182.560 36.740 182.850 ;
        RECT 37.435 182.820 38.935 182.990 ;
        RECT 37.435 182.680 37.605 182.820 ;
        RECT 37.045 182.510 37.605 182.680 ;
        RECT 35.520 181.880 35.770 182.340 ;
        RECT 35.940 182.050 36.810 182.390 ;
        RECT 37.045 182.050 37.215 182.510 ;
        RECT 38.050 182.480 39.125 182.650 ;
        RECT 37.385 181.880 37.755 182.340 ;
        RECT 38.050 182.140 38.220 182.480 ;
        RECT 38.390 181.880 38.720 182.310 ;
        RECT 38.955 182.140 39.125 182.480 ;
        RECT 39.295 182.380 39.465 183.160 ;
        RECT 39.635 182.940 39.805 183.530 ;
        RECT 39.975 183.130 40.325 183.750 ;
        RECT 39.635 182.550 40.100 182.940 ;
        RECT 40.495 182.680 40.665 184.040 ;
        RECT 40.835 182.850 41.295 183.900 ;
        RECT 40.270 182.510 40.665 182.680 ;
        RECT 40.270 182.380 40.440 182.510 ;
        RECT 39.295 182.050 39.975 182.380 ;
        RECT 40.190 182.050 40.440 182.380 ;
        RECT 40.610 181.880 40.860 182.340 ;
        RECT 41.030 182.065 41.355 182.850 ;
        RECT 41.525 182.050 41.695 184.170 ;
        RECT 41.865 184.050 42.195 184.430 ;
        RECT 42.365 183.880 42.620 184.170 ;
        RECT 41.870 183.710 42.620 183.880 ;
        RECT 41.870 182.720 42.100 183.710 ;
        RECT 43.315 183.610 43.525 184.430 ;
        RECT 43.695 183.630 44.025 184.260 ;
        RECT 42.270 182.890 42.620 183.540 ;
        RECT 43.695 183.030 43.945 183.630 ;
        RECT 44.195 183.610 44.425 184.430 ;
        RECT 44.725 183.880 44.895 184.260 ;
        RECT 45.075 184.050 45.405 184.430 ;
        RECT 44.725 183.710 45.390 183.880 ;
        RECT 45.585 183.755 45.845 184.260 ;
        RECT 44.115 183.190 44.445 183.440 ;
        RECT 44.655 183.160 44.985 183.530 ;
        RECT 45.220 183.455 45.390 183.710 ;
        RECT 45.220 183.125 45.505 183.455 ;
        RECT 41.870 182.550 42.620 182.720 ;
        RECT 41.865 181.880 42.195 182.380 ;
        RECT 42.365 182.050 42.620 182.550 ;
        RECT 43.315 181.880 43.525 183.020 ;
        RECT 43.695 182.050 44.025 183.030 ;
        RECT 44.195 181.880 44.425 183.020 ;
        RECT 45.220 182.980 45.390 183.125 ;
        RECT 44.725 182.810 45.390 182.980 ;
        RECT 45.675 182.955 45.845 183.755 ;
        RECT 46.130 183.800 46.415 184.260 ;
        RECT 46.585 183.970 46.855 184.430 ;
        RECT 46.130 183.630 47.085 183.800 ;
        RECT 44.725 182.050 44.895 182.810 ;
        RECT 45.075 181.880 45.405 182.640 ;
        RECT 45.575 182.050 45.845 182.955 ;
        RECT 46.015 182.900 46.705 183.460 ;
        RECT 46.875 182.730 47.085 183.630 ;
        RECT 46.130 182.510 47.085 182.730 ;
        RECT 47.255 183.460 47.655 184.260 ;
        RECT 47.845 183.800 48.125 184.260 ;
        RECT 48.645 183.970 48.970 184.430 ;
        RECT 47.845 183.630 48.970 183.800 ;
        RECT 49.140 183.690 49.525 184.260 ;
        RECT 48.520 183.520 48.970 183.630 ;
        RECT 47.255 182.900 48.350 183.460 ;
        RECT 48.520 183.190 49.075 183.520 ;
        RECT 46.130 182.050 46.415 182.510 ;
        RECT 46.585 181.880 46.855 182.340 ;
        RECT 47.255 182.050 47.655 182.900 ;
        RECT 48.520 182.730 48.970 183.190 ;
        RECT 49.245 183.020 49.525 183.690 ;
        RECT 49.735 183.610 49.965 184.430 ;
        RECT 50.135 183.630 50.465 184.260 ;
        RECT 49.715 183.190 50.045 183.440 ;
        RECT 50.215 183.030 50.465 183.630 ;
        RECT 50.635 183.610 50.845 184.430 ;
        RECT 51.075 183.705 51.365 184.430 ;
        RECT 51.535 183.690 51.920 184.260 ;
        RECT 52.090 183.970 52.415 184.430 ;
        RECT 52.935 183.800 53.215 184.260 ;
        RECT 47.845 182.510 48.970 182.730 ;
        RECT 47.845 182.050 48.125 182.510 ;
        RECT 48.645 181.880 48.970 182.340 ;
        RECT 49.140 182.050 49.525 183.020 ;
        RECT 49.735 181.880 49.965 183.020 ;
        RECT 50.135 182.050 50.465 183.030 ;
        RECT 50.635 181.880 50.845 183.020 ;
        RECT 51.075 181.880 51.365 183.045 ;
        RECT 51.535 183.020 51.815 183.690 ;
        RECT 52.090 183.630 53.215 183.800 ;
        RECT 52.090 183.520 52.540 183.630 ;
        RECT 51.985 183.190 52.540 183.520 ;
        RECT 53.405 183.460 53.805 184.260 ;
        RECT 54.205 183.970 54.475 184.430 ;
        RECT 54.645 183.800 54.930 184.260 ;
        RECT 55.220 183.885 60.565 184.430 ;
        RECT 60.740 183.885 66.085 184.430 ;
        RECT 66.525 184.035 66.855 184.430 ;
        RECT 51.535 182.050 51.920 183.020 ;
        RECT 52.090 182.730 52.540 183.190 ;
        RECT 52.710 182.900 53.805 183.460 ;
        RECT 52.090 182.510 53.215 182.730 ;
        RECT 52.090 181.880 52.415 182.340 ;
        RECT 52.935 182.050 53.215 182.510 ;
        RECT 53.405 182.050 53.805 182.900 ;
        RECT 53.975 183.630 54.930 183.800 ;
        RECT 53.975 182.730 54.185 183.630 ;
        RECT 54.355 182.900 55.045 183.460 ;
        RECT 53.975 182.510 54.930 182.730 ;
        RECT 54.205 181.880 54.475 182.340 ;
        RECT 54.645 182.050 54.930 182.510 ;
        RECT 56.810 182.315 57.160 183.565 ;
        RECT 58.640 183.055 58.980 183.885 ;
        RECT 62.330 182.315 62.680 183.565 ;
        RECT 64.160 183.055 64.500 183.885 ;
        RECT 67.025 183.860 67.225 184.215 ;
        RECT 67.395 184.030 67.725 184.430 ;
        RECT 67.895 183.860 68.095 184.205 ;
        RECT 66.255 183.690 68.095 183.860 ;
        RECT 68.265 183.690 68.595 184.430 ;
        RECT 68.830 183.860 69.000 184.110 ;
        RECT 68.830 183.690 69.305 183.860 ;
        RECT 55.220 181.880 60.565 182.315 ;
        RECT 60.740 181.880 66.085 182.315 ;
        RECT 66.255 182.065 66.515 183.690 ;
        RECT 66.695 182.720 66.915 183.520 ;
        RECT 67.155 182.900 67.455 183.520 ;
        RECT 67.625 182.900 67.955 183.520 ;
        RECT 68.125 182.900 68.445 183.520 ;
        RECT 68.615 182.900 68.965 183.520 ;
        RECT 69.135 182.720 69.305 183.690 ;
        RECT 69.935 183.660 72.525 184.430 ;
        RECT 66.695 182.510 69.305 182.720 ;
        RECT 69.935 182.970 71.145 183.490 ;
        RECT 71.315 183.140 72.525 183.660 ;
        RECT 72.970 183.620 73.215 184.225 ;
        RECT 73.435 183.895 73.945 184.430 ;
        RECT 72.695 183.450 73.925 183.620 ;
        RECT 68.265 181.880 68.595 182.330 ;
        RECT 69.935 181.880 72.525 182.970 ;
        RECT 72.695 182.640 73.035 183.450 ;
        RECT 73.205 182.885 73.955 183.075 ;
        RECT 72.695 182.230 73.210 182.640 ;
        RECT 73.445 181.880 73.615 182.640 ;
        RECT 73.785 182.220 73.955 182.885 ;
        RECT 74.125 182.900 74.315 184.260 ;
        RECT 74.485 183.410 74.760 184.260 ;
        RECT 74.950 183.895 75.480 184.260 ;
        RECT 75.905 184.030 76.235 184.430 ;
        RECT 75.305 183.860 75.480 183.895 ;
        RECT 74.485 183.240 74.765 183.410 ;
        RECT 74.485 183.100 74.760 183.240 ;
        RECT 74.965 182.900 75.135 183.700 ;
        RECT 74.125 182.730 75.135 182.900 ;
        RECT 75.305 183.690 76.235 183.860 ;
        RECT 76.405 183.690 76.660 184.260 ;
        RECT 76.835 183.705 77.125 184.430 ;
        RECT 75.305 182.560 75.475 183.690 ;
        RECT 76.065 183.520 76.235 183.690 ;
        RECT 74.350 182.390 75.475 182.560 ;
        RECT 75.645 183.190 75.840 183.520 ;
        RECT 76.065 183.190 76.320 183.520 ;
        RECT 75.645 182.220 75.815 183.190 ;
        RECT 76.490 183.020 76.660 183.690 ;
        RECT 77.355 183.610 77.565 184.430 ;
        RECT 77.735 183.630 78.065 184.260 ;
        RECT 73.785 182.050 75.815 182.220 ;
        RECT 75.985 181.880 76.155 183.020 ;
        RECT 76.325 182.050 76.660 183.020 ;
        RECT 76.835 181.880 77.125 183.045 ;
        RECT 77.735 183.030 77.985 183.630 ;
        RECT 78.235 183.610 78.465 184.430 ;
        RECT 78.950 183.620 79.195 184.225 ;
        RECT 79.415 183.895 79.925 184.430 ;
        RECT 78.675 183.450 79.905 183.620 ;
        RECT 78.155 183.190 78.485 183.440 ;
        RECT 77.355 181.880 77.565 183.020 ;
        RECT 77.735 182.050 78.065 183.030 ;
        RECT 78.235 181.880 78.465 183.020 ;
        RECT 78.675 182.640 79.015 183.450 ;
        RECT 79.185 182.885 79.935 183.075 ;
        RECT 78.675 182.230 79.190 182.640 ;
        RECT 79.425 181.880 79.595 182.640 ;
        RECT 79.765 182.220 79.935 182.885 ;
        RECT 80.105 182.900 80.295 184.260 ;
        RECT 80.465 183.410 80.740 184.260 ;
        RECT 80.930 183.895 81.460 184.260 ;
        RECT 81.885 184.030 82.215 184.430 ;
        RECT 81.285 183.860 81.460 183.895 ;
        RECT 80.465 183.240 80.745 183.410 ;
        RECT 80.465 183.100 80.740 183.240 ;
        RECT 80.945 182.900 81.115 183.700 ;
        RECT 80.105 182.730 81.115 182.900 ;
        RECT 81.285 183.690 82.215 183.860 ;
        RECT 82.385 183.690 82.640 184.260 ;
        RECT 82.905 183.880 83.075 184.260 ;
        RECT 83.255 184.050 83.585 184.430 ;
        RECT 82.905 183.710 83.570 183.880 ;
        RECT 83.765 183.755 84.025 184.260 ;
        RECT 81.285 182.560 81.455 183.690 ;
        RECT 82.045 183.520 82.215 183.690 ;
        RECT 80.330 182.390 81.455 182.560 ;
        RECT 81.625 183.190 81.820 183.520 ;
        RECT 82.045 183.190 82.300 183.520 ;
        RECT 81.625 182.220 81.795 183.190 ;
        RECT 82.470 183.020 82.640 183.690 ;
        RECT 82.835 183.160 83.165 183.530 ;
        RECT 83.400 183.455 83.570 183.710 ;
        RECT 79.765 182.050 81.795 182.220 ;
        RECT 81.965 181.880 82.135 183.020 ;
        RECT 82.305 182.050 82.640 183.020 ;
        RECT 83.400 183.125 83.685 183.455 ;
        RECT 83.400 182.980 83.570 183.125 ;
        RECT 82.905 182.810 83.570 182.980 ;
        RECT 83.855 182.955 84.025 183.755 ;
        RECT 85.120 183.880 85.375 184.170 ;
        RECT 85.545 184.050 85.875 184.430 ;
        RECT 85.120 183.710 85.870 183.880 ;
        RECT 82.905 182.050 83.075 182.810 ;
        RECT 83.255 181.880 83.585 182.640 ;
        RECT 83.755 182.050 84.025 182.955 ;
        RECT 85.120 182.890 85.470 183.540 ;
        RECT 85.640 182.720 85.870 183.710 ;
        RECT 85.120 182.550 85.870 182.720 ;
        RECT 85.120 182.050 85.375 182.550 ;
        RECT 85.545 181.880 85.875 182.380 ;
        RECT 86.045 182.050 86.215 184.170 ;
        RECT 86.575 184.070 86.905 184.430 ;
        RECT 87.075 184.040 87.570 184.210 ;
        RECT 87.775 184.040 88.630 184.210 ;
        RECT 86.445 182.850 86.905 183.900 ;
        RECT 86.385 182.065 86.710 182.850 ;
        RECT 87.075 182.680 87.245 184.040 ;
        RECT 87.415 183.130 87.765 183.750 ;
        RECT 87.935 183.530 88.290 183.750 ;
        RECT 87.935 182.940 88.105 183.530 ;
        RECT 88.460 183.330 88.630 184.040 ;
        RECT 89.505 183.970 89.835 184.430 ;
        RECT 90.045 184.070 90.395 184.240 ;
        RECT 88.835 183.500 89.625 183.750 ;
        RECT 90.045 183.680 90.305 184.070 ;
        RECT 90.615 183.980 91.565 184.260 ;
        RECT 91.735 183.990 91.925 184.430 ;
        RECT 92.095 184.050 93.165 184.220 ;
        RECT 89.795 183.330 89.965 183.510 ;
        RECT 87.075 182.510 87.470 182.680 ;
        RECT 87.640 182.550 88.105 182.940 ;
        RECT 88.275 183.160 89.965 183.330 ;
        RECT 87.300 182.380 87.470 182.510 ;
        RECT 88.275 182.380 88.445 183.160 ;
        RECT 90.135 182.990 90.305 183.680 ;
        RECT 88.805 182.820 90.305 182.990 ;
        RECT 90.495 183.020 90.705 183.810 ;
        RECT 90.875 183.190 91.225 183.810 ;
        RECT 91.395 183.200 91.565 183.980 ;
        RECT 92.095 183.820 92.265 184.050 ;
        RECT 91.735 183.650 92.265 183.820 ;
        RECT 91.735 183.370 91.955 183.650 ;
        RECT 92.435 183.480 92.675 183.880 ;
        RECT 91.395 183.030 91.800 183.200 ;
        RECT 92.135 183.110 92.675 183.480 ;
        RECT 92.845 183.695 93.165 184.050 ;
        RECT 93.410 183.970 93.715 184.430 ;
        RECT 93.885 183.720 94.140 184.250 ;
        RECT 92.845 183.520 93.170 183.695 ;
        RECT 92.845 183.220 93.760 183.520 ;
        RECT 93.020 183.190 93.760 183.220 ;
        RECT 90.495 182.860 91.170 183.020 ;
        RECT 91.630 182.940 91.800 183.030 ;
        RECT 90.495 182.850 91.460 182.860 ;
        RECT 90.135 182.680 90.305 182.820 ;
        RECT 86.880 181.880 87.130 182.340 ;
        RECT 87.300 182.050 87.550 182.380 ;
        RECT 87.765 182.050 88.445 182.380 ;
        RECT 88.615 182.480 89.690 182.650 ;
        RECT 90.135 182.510 90.695 182.680 ;
        RECT 91.000 182.560 91.460 182.850 ;
        RECT 91.630 182.770 92.850 182.940 ;
        RECT 88.615 182.140 88.785 182.480 ;
        RECT 89.020 181.880 89.350 182.310 ;
        RECT 89.520 182.140 89.690 182.480 ;
        RECT 89.985 181.880 90.355 182.340 ;
        RECT 90.525 182.050 90.695 182.510 ;
        RECT 91.630 182.390 91.800 182.770 ;
        RECT 93.020 182.600 93.190 183.190 ;
        RECT 93.930 183.070 94.140 183.720 ;
        RECT 94.590 183.620 94.835 184.225 ;
        RECT 95.055 183.895 95.565 184.430 ;
        RECT 90.930 182.050 91.800 182.390 ;
        RECT 92.390 182.430 93.190 182.600 ;
        RECT 91.970 181.880 92.220 182.340 ;
        RECT 92.390 182.140 92.560 182.430 ;
        RECT 92.740 181.880 93.070 182.260 ;
        RECT 93.410 181.880 93.715 183.020 ;
        RECT 93.885 182.190 94.140 183.070 ;
        RECT 94.315 183.450 95.545 183.620 ;
        RECT 94.315 182.640 94.655 183.450 ;
        RECT 94.825 182.885 95.575 183.075 ;
        RECT 94.315 182.230 94.830 182.640 ;
        RECT 95.065 181.880 95.235 182.640 ;
        RECT 95.405 182.220 95.575 182.885 ;
        RECT 95.745 182.900 95.935 184.260 ;
        RECT 96.105 184.090 96.380 184.260 ;
        RECT 96.105 183.920 96.385 184.090 ;
        RECT 96.105 183.100 96.380 183.920 ;
        RECT 96.570 183.895 97.100 184.260 ;
        RECT 97.525 184.030 97.855 184.430 ;
        RECT 96.925 183.860 97.100 183.895 ;
        RECT 96.585 182.900 96.755 183.700 ;
        RECT 95.745 182.730 96.755 182.900 ;
        RECT 96.925 183.690 97.855 183.860 ;
        RECT 98.025 183.690 98.280 184.260 ;
        RECT 96.925 182.560 97.095 183.690 ;
        RECT 97.685 183.520 97.855 183.690 ;
        RECT 95.970 182.390 97.095 182.560 ;
        RECT 97.265 183.190 97.460 183.520 ;
        RECT 97.685 183.190 97.940 183.520 ;
        RECT 97.265 182.220 97.435 183.190 ;
        RECT 98.110 183.020 98.280 183.690 ;
        RECT 98.730 183.620 98.975 184.225 ;
        RECT 99.195 183.895 99.705 184.430 ;
        RECT 95.405 182.050 97.435 182.220 ;
        RECT 97.605 181.880 97.775 183.020 ;
        RECT 97.945 182.050 98.280 183.020 ;
        RECT 98.455 183.450 99.685 183.620 ;
        RECT 98.455 182.640 98.795 183.450 ;
        RECT 98.965 182.885 99.715 183.075 ;
        RECT 98.455 182.230 98.970 182.640 ;
        RECT 99.205 181.880 99.375 182.640 ;
        RECT 99.545 182.220 99.715 182.885 ;
        RECT 99.885 182.900 100.075 184.260 ;
        RECT 100.245 184.090 100.520 184.260 ;
        RECT 100.245 183.920 100.525 184.090 ;
        RECT 100.245 183.100 100.520 183.920 ;
        RECT 100.710 183.895 101.240 184.260 ;
        RECT 101.665 184.030 101.995 184.430 ;
        RECT 101.065 183.860 101.240 183.895 ;
        RECT 100.725 182.900 100.895 183.700 ;
        RECT 99.885 182.730 100.895 182.900 ;
        RECT 101.065 183.690 101.995 183.860 ;
        RECT 102.165 183.690 102.420 184.260 ;
        RECT 102.595 183.705 102.885 184.430 ;
        RECT 103.060 183.720 103.315 184.250 ;
        RECT 103.485 183.970 103.790 184.430 ;
        RECT 104.035 184.050 105.105 184.220 ;
        RECT 101.065 182.560 101.235 183.690 ;
        RECT 101.825 183.520 101.995 183.690 ;
        RECT 100.110 182.390 101.235 182.560 ;
        RECT 101.405 183.190 101.600 183.520 ;
        RECT 101.825 183.190 102.080 183.520 ;
        RECT 101.405 182.220 101.575 183.190 ;
        RECT 102.250 183.020 102.420 183.690 ;
        RECT 103.060 183.070 103.270 183.720 ;
        RECT 104.035 183.695 104.355 184.050 ;
        RECT 104.030 183.520 104.355 183.695 ;
        RECT 103.440 183.220 104.355 183.520 ;
        RECT 104.525 183.480 104.765 183.880 ;
        RECT 104.935 183.820 105.105 184.050 ;
        RECT 105.275 183.990 105.465 184.430 ;
        RECT 105.635 183.980 106.585 184.260 ;
        RECT 106.805 184.070 107.155 184.240 ;
        RECT 104.935 183.650 105.465 183.820 ;
        RECT 103.440 183.190 104.180 183.220 ;
        RECT 99.545 182.050 101.575 182.220 ;
        RECT 101.745 181.880 101.915 183.020 ;
        RECT 102.085 182.050 102.420 183.020 ;
        RECT 102.595 181.880 102.885 183.045 ;
        RECT 103.060 182.190 103.315 183.070 ;
        RECT 103.485 181.880 103.790 183.020 ;
        RECT 104.010 182.600 104.180 183.190 ;
        RECT 104.525 183.110 105.065 183.480 ;
        RECT 105.245 183.370 105.465 183.650 ;
        RECT 105.635 183.200 105.805 183.980 ;
        RECT 105.400 183.030 105.805 183.200 ;
        RECT 105.975 183.190 106.325 183.810 ;
        RECT 105.400 182.940 105.570 183.030 ;
        RECT 106.495 183.020 106.705 183.810 ;
        RECT 104.350 182.770 105.570 182.940 ;
        RECT 106.030 182.860 106.705 183.020 ;
        RECT 104.010 182.430 104.810 182.600 ;
        RECT 104.130 181.880 104.460 182.260 ;
        RECT 104.640 182.140 104.810 182.430 ;
        RECT 105.400 182.390 105.570 182.770 ;
        RECT 105.740 182.850 106.705 182.860 ;
        RECT 106.895 183.680 107.155 184.070 ;
        RECT 107.365 183.970 107.695 184.430 ;
        RECT 108.570 184.040 109.425 184.210 ;
        RECT 109.630 184.040 110.125 184.210 ;
        RECT 110.295 184.070 110.625 184.430 ;
        RECT 106.895 182.990 107.065 183.680 ;
        RECT 107.235 183.330 107.405 183.510 ;
        RECT 107.575 183.500 108.365 183.750 ;
        RECT 108.570 183.330 108.740 184.040 ;
        RECT 108.910 183.530 109.265 183.750 ;
        RECT 107.235 183.160 108.925 183.330 ;
        RECT 105.740 182.560 106.200 182.850 ;
        RECT 106.895 182.820 108.395 182.990 ;
        RECT 106.895 182.680 107.065 182.820 ;
        RECT 106.505 182.510 107.065 182.680 ;
        RECT 104.980 181.880 105.230 182.340 ;
        RECT 105.400 182.050 106.270 182.390 ;
        RECT 106.505 182.050 106.675 182.510 ;
        RECT 107.510 182.480 108.585 182.650 ;
        RECT 106.845 181.880 107.215 182.340 ;
        RECT 107.510 182.140 107.680 182.480 ;
        RECT 107.850 181.880 108.180 182.310 ;
        RECT 108.415 182.140 108.585 182.480 ;
        RECT 108.755 182.380 108.925 183.160 ;
        RECT 109.095 182.940 109.265 183.530 ;
        RECT 109.435 183.130 109.785 183.750 ;
        RECT 109.095 182.550 109.560 182.940 ;
        RECT 109.955 182.680 110.125 184.040 ;
        RECT 110.295 182.850 110.755 183.900 ;
        RECT 109.730 182.510 110.125 182.680 ;
        RECT 109.730 182.380 109.900 182.510 ;
        RECT 108.755 182.050 109.435 182.380 ;
        RECT 109.650 182.050 109.900 182.380 ;
        RECT 110.070 181.880 110.320 182.340 ;
        RECT 110.490 182.065 110.815 182.850 ;
        RECT 110.985 182.050 111.155 184.170 ;
        RECT 111.325 184.050 111.655 184.430 ;
        RECT 111.825 183.880 112.080 184.170 ;
        RECT 111.330 183.710 112.080 183.880 ;
        RECT 111.330 182.720 111.560 183.710 ;
        RECT 112.715 183.660 114.385 184.430 ;
        RECT 114.555 183.680 115.765 184.430 ;
        RECT 111.730 182.890 112.080 183.540 ;
        RECT 112.715 182.970 113.465 183.490 ;
        RECT 113.635 183.140 114.385 183.660 ;
        RECT 114.555 182.970 115.075 183.510 ;
        RECT 115.245 183.140 115.765 183.680 ;
        RECT 111.330 182.550 112.080 182.720 ;
        RECT 111.325 181.880 111.655 182.380 ;
        RECT 111.825 182.050 112.080 182.550 ;
        RECT 112.715 181.880 114.385 182.970 ;
        RECT 114.555 181.880 115.765 182.970 ;
        RECT 14.650 181.710 115.850 181.880 ;
        RECT 14.735 180.620 15.945 181.710 ;
        RECT 14.735 179.910 15.255 180.450 ;
        RECT 15.425 180.080 15.945 180.620 ;
        RECT 16.575 180.620 18.245 181.710 ;
        RECT 18.530 181.080 18.815 181.540 ;
        RECT 18.985 181.250 19.255 181.710 ;
        RECT 18.530 180.860 19.485 181.080 ;
        RECT 16.575 180.100 17.325 180.620 ;
        RECT 17.495 179.930 18.245 180.450 ;
        RECT 18.415 180.130 19.105 180.690 ;
        RECT 19.275 179.960 19.485 180.860 ;
        RECT 14.735 179.160 15.945 179.910 ;
        RECT 16.575 179.160 18.245 179.930 ;
        RECT 18.530 179.790 19.485 179.960 ;
        RECT 19.655 180.690 20.055 181.540 ;
        RECT 20.245 181.080 20.525 181.540 ;
        RECT 21.045 181.250 21.370 181.710 ;
        RECT 20.245 180.860 21.370 181.080 ;
        RECT 19.655 180.130 20.750 180.690 ;
        RECT 20.920 180.400 21.370 180.860 ;
        RECT 21.540 180.570 21.925 181.540 ;
        RECT 18.530 179.330 18.815 179.790 ;
        RECT 18.985 179.160 19.255 179.620 ;
        RECT 19.655 179.330 20.055 180.130 ;
        RECT 20.920 180.070 21.475 180.400 ;
        RECT 20.920 179.960 21.370 180.070 ;
        RECT 20.245 179.790 21.370 179.960 ;
        RECT 21.645 179.900 21.925 180.570 ;
        RECT 20.245 179.330 20.525 179.790 ;
        RECT 21.045 179.160 21.370 179.620 ;
        RECT 21.540 179.330 21.925 179.900 ;
        RECT 22.100 180.520 22.355 181.400 ;
        RECT 22.525 180.570 22.830 181.710 ;
        RECT 23.170 181.330 23.500 181.710 ;
        RECT 23.680 181.160 23.850 181.450 ;
        RECT 24.020 181.250 24.270 181.710 ;
        RECT 23.050 180.990 23.850 181.160 ;
        RECT 24.440 181.200 25.310 181.540 ;
        RECT 22.100 179.870 22.310 180.520 ;
        RECT 23.050 180.400 23.220 180.990 ;
        RECT 24.440 180.820 24.610 181.200 ;
        RECT 25.545 181.080 25.715 181.540 ;
        RECT 25.885 181.250 26.255 181.710 ;
        RECT 26.550 181.110 26.720 181.450 ;
        RECT 26.890 181.280 27.220 181.710 ;
        RECT 27.455 181.110 27.625 181.450 ;
        RECT 23.390 180.650 24.610 180.820 ;
        RECT 24.780 180.740 25.240 181.030 ;
        RECT 25.545 180.910 26.105 181.080 ;
        RECT 26.550 180.940 27.625 181.110 ;
        RECT 27.795 181.210 28.475 181.540 ;
        RECT 28.690 181.210 28.940 181.540 ;
        RECT 29.110 181.250 29.360 181.710 ;
        RECT 25.935 180.770 26.105 180.910 ;
        RECT 24.780 180.730 25.745 180.740 ;
        RECT 24.440 180.560 24.610 180.650 ;
        RECT 25.070 180.570 25.745 180.730 ;
        RECT 22.480 180.370 23.220 180.400 ;
        RECT 22.480 180.070 23.395 180.370 ;
        RECT 23.070 179.895 23.395 180.070 ;
        RECT 22.100 179.340 22.355 179.870 ;
        RECT 22.525 179.160 22.830 179.620 ;
        RECT 23.075 179.540 23.395 179.895 ;
        RECT 23.565 180.110 24.105 180.480 ;
        RECT 24.440 180.390 24.845 180.560 ;
        RECT 23.565 179.710 23.805 180.110 ;
        RECT 24.285 179.940 24.505 180.220 ;
        RECT 23.975 179.770 24.505 179.940 ;
        RECT 23.975 179.540 24.145 179.770 ;
        RECT 24.675 179.610 24.845 180.390 ;
        RECT 25.015 179.780 25.365 180.400 ;
        RECT 25.535 179.780 25.745 180.570 ;
        RECT 25.935 180.600 27.435 180.770 ;
        RECT 25.935 179.910 26.105 180.600 ;
        RECT 27.795 180.430 27.965 181.210 ;
        RECT 28.770 181.080 28.940 181.210 ;
        RECT 26.275 180.260 27.965 180.430 ;
        RECT 28.135 180.650 28.600 181.040 ;
        RECT 28.770 180.910 29.165 181.080 ;
        RECT 26.275 180.080 26.445 180.260 ;
        RECT 23.075 179.370 24.145 179.540 ;
        RECT 24.315 179.160 24.505 179.600 ;
        RECT 24.675 179.330 25.625 179.610 ;
        RECT 25.935 179.520 26.195 179.910 ;
        RECT 26.615 179.840 27.405 180.090 ;
        RECT 25.845 179.350 26.195 179.520 ;
        RECT 26.405 179.160 26.735 179.620 ;
        RECT 27.610 179.550 27.780 180.260 ;
        RECT 28.135 180.060 28.305 180.650 ;
        RECT 27.950 179.840 28.305 180.060 ;
        RECT 28.475 179.840 28.825 180.460 ;
        RECT 28.995 179.550 29.165 180.910 ;
        RECT 29.530 180.740 29.855 181.525 ;
        RECT 29.335 179.690 29.795 180.740 ;
        RECT 27.610 179.380 28.465 179.550 ;
        RECT 28.670 179.380 29.165 179.550 ;
        RECT 29.335 179.160 29.665 179.520 ;
        RECT 30.025 179.420 30.195 181.540 ;
        RECT 30.365 181.210 30.695 181.710 ;
        RECT 30.865 181.040 31.120 181.540 ;
        RECT 30.370 180.870 31.120 181.040 ;
        RECT 30.370 179.880 30.600 180.870 ;
        RECT 30.770 180.050 31.120 180.700 ;
        RECT 31.295 180.620 32.965 181.710 ;
        RECT 31.295 180.100 32.045 180.620 ;
        RECT 33.175 180.570 33.405 181.710 ;
        RECT 33.575 180.560 33.905 181.540 ;
        RECT 34.075 180.570 34.285 181.710 ;
        RECT 34.630 181.080 34.915 181.540 ;
        RECT 35.085 181.250 35.355 181.710 ;
        RECT 34.630 180.860 35.585 181.080 ;
        RECT 32.215 179.930 32.965 180.450 ;
        RECT 33.155 180.150 33.485 180.400 ;
        RECT 30.370 179.710 31.120 179.880 ;
        RECT 30.365 179.160 30.695 179.540 ;
        RECT 30.865 179.420 31.120 179.710 ;
        RECT 31.295 179.160 32.965 179.930 ;
        RECT 33.175 179.160 33.405 179.980 ;
        RECT 33.655 179.960 33.905 180.560 ;
        RECT 34.515 180.130 35.205 180.690 ;
        RECT 33.575 179.330 33.905 179.960 ;
        RECT 34.075 179.160 34.285 179.980 ;
        RECT 35.375 179.960 35.585 180.860 ;
        RECT 34.630 179.790 35.585 179.960 ;
        RECT 35.755 180.690 36.155 181.540 ;
        RECT 36.345 181.080 36.625 181.540 ;
        RECT 37.145 181.250 37.470 181.710 ;
        RECT 36.345 180.860 37.470 181.080 ;
        RECT 35.755 180.130 36.850 180.690 ;
        RECT 37.020 180.400 37.470 180.860 ;
        RECT 37.640 180.570 38.025 181.540 ;
        RECT 34.630 179.330 34.915 179.790 ;
        RECT 35.085 179.160 35.355 179.620 ;
        RECT 35.755 179.330 36.155 180.130 ;
        RECT 37.020 180.070 37.575 180.400 ;
        RECT 37.020 179.960 37.470 180.070 ;
        RECT 36.345 179.790 37.470 179.960 ;
        RECT 37.745 179.900 38.025 180.570 ;
        RECT 38.195 180.545 38.485 181.710 ;
        RECT 39.575 180.570 39.915 181.540 ;
        RECT 40.085 180.570 40.255 181.710 ;
        RECT 40.525 180.910 40.775 181.710 ;
        RECT 41.420 180.740 41.750 181.540 ;
        RECT 42.050 180.910 42.380 181.710 ;
        RECT 42.550 180.740 42.880 181.540 ;
        RECT 40.445 180.570 42.880 180.740 ;
        RECT 43.255 180.950 43.770 181.360 ;
        RECT 44.005 180.950 44.175 181.710 ;
        RECT 44.345 181.370 46.375 181.540 ;
        RECT 36.345 179.330 36.625 179.790 ;
        RECT 37.145 179.160 37.470 179.620 ;
        RECT 37.640 179.330 38.025 179.900 ;
        RECT 39.575 179.960 39.750 180.570 ;
        RECT 40.445 180.320 40.615 180.570 ;
        RECT 39.920 180.150 40.615 180.320 ;
        RECT 40.790 180.150 41.210 180.350 ;
        RECT 41.380 180.150 41.710 180.350 ;
        RECT 41.880 180.150 42.210 180.350 ;
        RECT 38.195 179.160 38.485 179.885 ;
        RECT 39.575 179.330 39.915 179.960 ;
        RECT 40.085 179.160 40.335 179.960 ;
        RECT 40.525 179.810 41.750 179.980 ;
        RECT 40.525 179.330 40.855 179.810 ;
        RECT 41.025 179.160 41.250 179.620 ;
        RECT 41.420 179.330 41.750 179.810 ;
        RECT 42.380 179.940 42.550 180.570 ;
        RECT 42.735 180.150 43.085 180.400 ;
        RECT 43.255 180.140 43.595 180.950 ;
        RECT 44.345 180.705 44.515 181.370 ;
        RECT 44.910 181.030 46.035 181.200 ;
        RECT 43.765 180.515 44.515 180.705 ;
        RECT 44.685 180.690 45.695 180.860 ;
        RECT 43.255 179.970 44.485 180.140 ;
        RECT 42.380 179.330 42.880 179.940 ;
        RECT 43.530 179.365 43.775 179.970 ;
        RECT 43.995 179.160 44.505 179.695 ;
        RECT 44.685 179.330 44.875 180.690 ;
        RECT 45.045 180.350 45.320 180.490 ;
        RECT 45.045 180.180 45.325 180.350 ;
        RECT 45.045 179.330 45.320 180.180 ;
        RECT 45.525 179.890 45.695 180.690 ;
        RECT 45.865 179.900 46.035 181.030 ;
        RECT 46.205 180.400 46.375 181.370 ;
        RECT 46.545 180.570 46.715 181.710 ;
        RECT 46.885 180.570 47.220 181.540 ;
        RECT 46.205 180.070 46.400 180.400 ;
        RECT 46.625 180.070 46.880 180.400 ;
        RECT 46.625 179.900 46.795 180.070 ;
        RECT 47.050 179.900 47.220 180.570 ;
        RECT 45.865 179.730 46.795 179.900 ;
        RECT 45.865 179.695 46.040 179.730 ;
        RECT 45.510 179.330 46.040 179.695 ;
        RECT 46.465 179.160 46.795 179.560 ;
        RECT 46.965 179.330 47.220 179.900 ;
        RECT 47.400 180.520 47.655 181.400 ;
        RECT 47.825 180.570 48.130 181.710 ;
        RECT 48.470 181.330 48.800 181.710 ;
        RECT 48.980 181.160 49.150 181.450 ;
        RECT 49.320 181.250 49.570 181.710 ;
        RECT 48.350 180.990 49.150 181.160 ;
        RECT 49.740 181.200 50.610 181.540 ;
        RECT 47.400 179.870 47.610 180.520 ;
        RECT 48.350 180.400 48.520 180.990 ;
        RECT 49.740 180.820 49.910 181.200 ;
        RECT 50.845 181.080 51.015 181.540 ;
        RECT 51.185 181.250 51.555 181.710 ;
        RECT 51.850 181.110 52.020 181.450 ;
        RECT 52.190 181.280 52.520 181.710 ;
        RECT 52.755 181.110 52.925 181.450 ;
        RECT 48.690 180.650 49.910 180.820 ;
        RECT 50.080 180.740 50.540 181.030 ;
        RECT 50.845 180.910 51.405 181.080 ;
        RECT 51.850 180.940 52.925 181.110 ;
        RECT 53.095 181.210 53.775 181.540 ;
        RECT 53.990 181.210 54.240 181.540 ;
        RECT 54.410 181.250 54.660 181.710 ;
        RECT 51.235 180.770 51.405 180.910 ;
        RECT 50.080 180.730 51.045 180.740 ;
        RECT 49.740 180.560 49.910 180.650 ;
        RECT 50.370 180.570 51.045 180.730 ;
        RECT 47.780 180.370 48.520 180.400 ;
        RECT 47.780 180.070 48.695 180.370 ;
        RECT 48.370 179.895 48.695 180.070 ;
        RECT 47.400 179.340 47.655 179.870 ;
        RECT 47.825 179.160 48.130 179.620 ;
        RECT 48.375 179.540 48.695 179.895 ;
        RECT 48.865 180.110 49.405 180.480 ;
        RECT 49.740 180.390 50.145 180.560 ;
        RECT 48.865 179.710 49.105 180.110 ;
        RECT 49.585 179.940 49.805 180.220 ;
        RECT 49.275 179.770 49.805 179.940 ;
        RECT 49.275 179.540 49.445 179.770 ;
        RECT 49.975 179.610 50.145 180.390 ;
        RECT 50.315 179.780 50.665 180.400 ;
        RECT 50.835 179.780 51.045 180.570 ;
        RECT 51.235 180.600 52.735 180.770 ;
        RECT 51.235 179.910 51.405 180.600 ;
        RECT 53.095 180.430 53.265 181.210 ;
        RECT 54.070 181.080 54.240 181.210 ;
        RECT 51.575 180.260 53.265 180.430 ;
        RECT 53.435 180.650 53.900 181.040 ;
        RECT 54.070 180.910 54.465 181.080 ;
        RECT 51.575 180.080 51.745 180.260 ;
        RECT 48.375 179.370 49.445 179.540 ;
        RECT 49.615 179.160 49.805 179.600 ;
        RECT 49.975 179.330 50.925 179.610 ;
        RECT 51.235 179.520 51.495 179.910 ;
        RECT 51.915 179.840 52.705 180.090 ;
        RECT 51.145 179.350 51.495 179.520 ;
        RECT 51.705 179.160 52.035 179.620 ;
        RECT 52.910 179.550 53.080 180.260 ;
        RECT 53.435 180.060 53.605 180.650 ;
        RECT 53.250 179.840 53.605 180.060 ;
        RECT 53.775 179.840 54.125 180.460 ;
        RECT 54.295 179.550 54.465 180.910 ;
        RECT 54.830 180.740 55.155 181.525 ;
        RECT 54.635 179.690 55.095 180.740 ;
        RECT 52.910 179.380 53.765 179.550 ;
        RECT 53.970 179.380 54.465 179.550 ;
        RECT 54.635 179.160 54.965 179.520 ;
        RECT 55.325 179.420 55.495 181.540 ;
        RECT 55.665 181.210 55.995 181.710 ;
        RECT 56.165 181.040 56.420 181.540 ;
        RECT 55.670 180.870 56.420 181.040 ;
        RECT 55.670 179.880 55.900 180.870 ;
        RECT 56.070 180.050 56.420 180.700 ;
        RECT 56.595 180.620 57.805 181.710 ;
        RECT 57.985 180.730 58.315 181.540 ;
        RECT 58.485 180.910 58.725 181.710 ;
        RECT 56.595 180.080 57.115 180.620 ;
        RECT 57.985 180.560 58.700 180.730 ;
        RECT 57.285 179.910 57.805 180.450 ;
        RECT 57.980 180.150 58.360 180.390 ;
        RECT 58.530 180.320 58.700 180.560 ;
        RECT 58.905 180.690 59.075 181.540 ;
        RECT 59.245 180.910 59.575 181.710 ;
        RECT 59.745 180.690 59.915 181.540 ;
        RECT 58.905 180.520 59.915 180.690 ;
        RECT 60.085 180.560 60.415 181.710 ;
        RECT 58.530 180.150 59.030 180.320 ;
        RECT 58.530 179.980 58.700 180.150 ;
        RECT 59.420 179.980 59.915 180.520 ;
        RECT 55.670 179.710 56.420 179.880 ;
        RECT 55.665 179.160 55.995 179.540 ;
        RECT 56.165 179.420 56.420 179.710 ;
        RECT 56.595 179.160 57.805 179.910 ;
        RECT 58.065 179.810 58.700 179.980 ;
        RECT 58.905 179.810 59.915 179.980 ;
        RECT 58.065 179.330 58.235 179.810 ;
        RECT 58.415 179.160 58.655 179.640 ;
        RECT 58.905 179.330 59.075 179.810 ;
        RECT 59.245 179.160 59.575 179.640 ;
        RECT 59.745 179.330 59.915 179.810 ;
        RECT 60.085 179.160 60.415 179.960 ;
        RECT 60.735 179.900 60.995 181.525 ;
        RECT 62.745 181.260 63.075 181.710 ;
        RECT 61.175 180.870 63.785 181.080 ;
        RECT 61.175 180.070 61.395 180.870 ;
        RECT 61.635 180.070 61.935 180.690 ;
        RECT 62.105 180.070 62.435 180.690 ;
        RECT 62.605 180.070 62.925 180.690 ;
        RECT 63.095 180.070 63.445 180.690 ;
        RECT 63.615 179.900 63.785 180.870 ;
        RECT 63.955 180.545 64.245 181.710 ;
        RECT 64.415 180.620 65.625 181.710 ;
        RECT 65.795 181.210 66.055 181.540 ;
        RECT 66.365 181.330 66.695 181.710 ;
        RECT 64.415 180.080 64.935 180.620 ;
        RECT 65.795 180.530 65.965 181.210 ;
        RECT 66.935 181.160 67.125 181.540 ;
        RECT 67.375 181.330 67.705 181.710 ;
        RECT 67.915 181.160 68.085 181.540 ;
        RECT 68.280 181.330 68.610 181.710 ;
        RECT 68.870 181.160 69.040 181.540 ;
        RECT 69.465 181.330 69.795 181.710 ;
        RECT 66.135 180.700 66.485 181.030 ;
        RECT 66.935 180.990 67.675 181.160 ;
        RECT 66.755 180.650 67.335 180.820 ;
        RECT 66.755 180.530 66.925 180.650 ;
        RECT 65.105 179.910 65.625 180.450 ;
        RECT 60.735 179.730 62.575 179.900 ;
        RECT 61.005 179.160 61.335 179.555 ;
        RECT 61.505 179.375 61.705 179.730 ;
        RECT 61.875 179.160 62.205 179.560 ;
        RECT 62.375 179.385 62.575 179.730 ;
        RECT 62.745 179.160 63.075 179.900 ;
        RECT 63.310 179.730 63.785 179.900 ;
        RECT 63.310 179.480 63.480 179.730 ;
        RECT 63.955 179.160 64.245 179.885 ;
        RECT 64.415 179.160 65.625 179.910 ;
        RECT 65.795 180.360 66.925 180.530 ;
        RECT 67.505 180.480 67.675 180.990 ;
        RECT 65.795 179.660 65.965 180.360 ;
        RECT 67.105 180.310 67.675 180.480 ;
        RECT 67.845 180.990 69.795 181.160 ;
        RECT 66.315 180.020 66.935 180.190 ;
        RECT 66.315 179.840 66.525 180.020 ;
        RECT 67.105 179.830 67.275 180.310 ;
        RECT 67.845 180.000 68.015 180.990 ;
        RECT 68.605 180.400 68.790 180.710 ;
        RECT 69.060 180.400 69.255 180.710 ;
        RECT 65.795 179.330 66.055 179.660 ;
        RECT 66.365 179.160 66.695 179.540 ;
        RECT 66.875 179.500 67.275 179.830 ;
        RECT 67.465 179.670 68.015 180.000 ;
        RECT 68.185 179.500 68.355 180.400 ;
        RECT 66.875 179.330 68.355 179.500 ;
        RECT 68.605 180.070 68.835 180.400 ;
        RECT 69.060 180.070 69.315 180.400 ;
        RECT 69.625 180.070 69.795 180.990 ;
        RECT 68.605 179.490 68.790 180.070 ;
        RECT 69.060 179.495 69.255 180.070 ;
        RECT 69.465 179.160 69.795 179.540 ;
        RECT 69.965 179.330 70.225 181.540 ;
        RECT 70.395 180.740 70.705 181.540 ;
        RECT 70.875 180.910 71.185 181.710 ;
        RECT 71.355 181.080 71.615 181.540 ;
        RECT 71.785 181.250 72.040 181.710 ;
        RECT 72.215 181.080 72.475 181.540 ;
        RECT 71.355 180.910 72.475 181.080 ;
        RECT 70.395 180.570 71.425 180.740 ;
        RECT 70.395 179.660 70.565 180.570 ;
        RECT 70.735 179.830 71.085 180.400 ;
        RECT 71.255 180.320 71.425 180.570 ;
        RECT 72.215 180.660 72.475 180.910 ;
        RECT 72.645 180.840 72.930 181.710 ;
        RECT 72.215 180.490 72.970 180.660 ;
        RECT 71.255 180.150 72.395 180.320 ;
        RECT 72.565 179.980 72.970 180.490 ;
        RECT 71.320 179.810 72.970 179.980 ;
        RECT 73.155 180.570 73.540 181.540 ;
        RECT 73.710 181.250 74.035 181.710 ;
        RECT 74.555 181.080 74.835 181.540 ;
        RECT 73.710 180.860 74.835 181.080 ;
        RECT 73.155 179.900 73.435 180.570 ;
        RECT 73.710 180.400 74.160 180.860 ;
        RECT 75.025 180.690 75.425 181.540 ;
        RECT 75.825 181.250 76.095 181.710 ;
        RECT 76.265 181.080 76.550 181.540 ;
        RECT 73.605 180.070 74.160 180.400 ;
        RECT 74.330 180.130 75.425 180.690 ;
        RECT 73.710 179.960 74.160 180.070 ;
        RECT 70.395 179.330 70.695 179.660 ;
        RECT 70.865 179.160 71.140 179.640 ;
        RECT 71.320 179.420 71.615 179.810 ;
        RECT 71.785 179.160 72.040 179.640 ;
        RECT 72.215 179.420 72.475 179.810 ;
        RECT 72.645 179.160 72.925 179.640 ;
        RECT 73.155 179.330 73.540 179.900 ;
        RECT 73.710 179.790 74.835 179.960 ;
        RECT 73.710 179.160 74.035 179.620 ;
        RECT 74.555 179.330 74.835 179.790 ;
        RECT 75.025 179.330 75.425 180.130 ;
        RECT 75.595 180.860 76.550 181.080 ;
        RECT 75.595 179.960 75.805 180.860 ;
        RECT 75.975 180.130 76.665 180.690 ;
        RECT 76.840 180.520 77.095 181.400 ;
        RECT 77.265 180.570 77.570 181.710 ;
        RECT 77.910 181.330 78.240 181.710 ;
        RECT 78.420 181.160 78.590 181.450 ;
        RECT 78.760 181.250 79.010 181.710 ;
        RECT 77.790 180.990 78.590 181.160 ;
        RECT 79.180 181.200 80.050 181.540 ;
        RECT 75.595 179.790 76.550 179.960 ;
        RECT 75.825 179.160 76.095 179.620 ;
        RECT 76.265 179.330 76.550 179.790 ;
        RECT 76.840 179.870 77.050 180.520 ;
        RECT 77.790 180.400 77.960 180.990 ;
        RECT 79.180 180.820 79.350 181.200 ;
        RECT 80.285 181.080 80.455 181.540 ;
        RECT 80.625 181.250 80.995 181.710 ;
        RECT 81.290 181.110 81.460 181.450 ;
        RECT 81.630 181.280 81.960 181.710 ;
        RECT 82.195 181.110 82.365 181.450 ;
        RECT 78.130 180.650 79.350 180.820 ;
        RECT 79.520 180.740 79.980 181.030 ;
        RECT 80.285 180.910 80.845 181.080 ;
        RECT 81.290 180.940 82.365 181.110 ;
        RECT 82.535 181.210 83.215 181.540 ;
        RECT 83.430 181.210 83.680 181.540 ;
        RECT 83.850 181.250 84.100 181.710 ;
        RECT 80.675 180.770 80.845 180.910 ;
        RECT 79.520 180.730 80.485 180.740 ;
        RECT 79.180 180.560 79.350 180.650 ;
        RECT 79.810 180.570 80.485 180.730 ;
        RECT 77.220 180.370 77.960 180.400 ;
        RECT 77.220 180.070 78.135 180.370 ;
        RECT 77.810 179.895 78.135 180.070 ;
        RECT 76.840 179.340 77.095 179.870 ;
        RECT 77.265 179.160 77.570 179.620 ;
        RECT 77.815 179.540 78.135 179.895 ;
        RECT 78.305 180.110 78.845 180.480 ;
        RECT 79.180 180.390 79.585 180.560 ;
        RECT 78.305 179.710 78.545 180.110 ;
        RECT 79.025 179.940 79.245 180.220 ;
        RECT 78.715 179.770 79.245 179.940 ;
        RECT 78.715 179.540 78.885 179.770 ;
        RECT 79.415 179.610 79.585 180.390 ;
        RECT 79.755 179.780 80.105 180.400 ;
        RECT 80.275 179.780 80.485 180.570 ;
        RECT 80.675 180.600 82.175 180.770 ;
        RECT 80.675 179.910 80.845 180.600 ;
        RECT 82.535 180.430 82.705 181.210 ;
        RECT 83.510 181.080 83.680 181.210 ;
        RECT 81.015 180.260 82.705 180.430 ;
        RECT 82.875 180.650 83.340 181.040 ;
        RECT 83.510 180.910 83.905 181.080 ;
        RECT 81.015 180.080 81.185 180.260 ;
        RECT 77.815 179.370 78.885 179.540 ;
        RECT 79.055 179.160 79.245 179.600 ;
        RECT 79.415 179.330 80.365 179.610 ;
        RECT 80.675 179.520 80.935 179.910 ;
        RECT 81.355 179.840 82.145 180.090 ;
        RECT 80.585 179.350 80.935 179.520 ;
        RECT 81.145 179.160 81.475 179.620 ;
        RECT 82.350 179.550 82.520 180.260 ;
        RECT 82.875 180.060 83.045 180.650 ;
        RECT 82.690 179.840 83.045 180.060 ;
        RECT 83.215 179.840 83.565 180.460 ;
        RECT 83.735 179.550 83.905 180.910 ;
        RECT 84.270 180.740 84.595 181.525 ;
        RECT 84.075 179.690 84.535 180.740 ;
        RECT 82.350 179.380 83.205 179.550 ;
        RECT 83.410 179.380 83.905 179.550 ;
        RECT 84.075 179.160 84.405 179.520 ;
        RECT 84.765 179.420 84.935 181.540 ;
        RECT 85.105 181.210 85.435 181.710 ;
        RECT 85.605 181.040 85.860 181.540 ;
        RECT 85.110 180.870 85.860 181.040 ;
        RECT 86.150 181.080 86.435 181.540 ;
        RECT 86.605 181.250 86.875 181.710 ;
        RECT 85.110 179.880 85.340 180.870 ;
        RECT 86.150 180.860 87.105 181.080 ;
        RECT 85.510 180.050 85.860 180.700 ;
        RECT 86.035 180.130 86.725 180.690 ;
        RECT 86.895 179.960 87.105 180.860 ;
        RECT 85.110 179.710 85.860 179.880 ;
        RECT 85.105 179.160 85.435 179.540 ;
        RECT 85.605 179.420 85.860 179.710 ;
        RECT 86.150 179.790 87.105 179.960 ;
        RECT 87.275 180.690 87.675 181.540 ;
        RECT 87.865 181.080 88.145 181.540 ;
        RECT 88.665 181.250 88.990 181.710 ;
        RECT 87.865 180.860 88.990 181.080 ;
        RECT 87.275 180.130 88.370 180.690 ;
        RECT 88.540 180.400 88.990 180.860 ;
        RECT 89.160 180.570 89.545 181.540 ;
        RECT 86.150 179.330 86.435 179.790 ;
        RECT 86.605 179.160 86.875 179.620 ;
        RECT 87.275 179.330 87.675 180.130 ;
        RECT 88.540 180.070 89.095 180.400 ;
        RECT 88.540 179.960 88.990 180.070 ;
        RECT 87.865 179.790 88.990 179.960 ;
        RECT 89.265 179.900 89.545 180.570 ;
        RECT 89.715 180.545 90.005 181.710 ;
        RECT 90.180 180.570 90.515 181.540 ;
        RECT 90.685 180.570 90.855 181.710 ;
        RECT 91.025 181.370 93.055 181.540 ;
        RECT 87.865 179.330 88.145 179.790 ;
        RECT 88.665 179.160 88.990 179.620 ;
        RECT 89.160 179.330 89.545 179.900 ;
        RECT 90.180 179.900 90.350 180.570 ;
        RECT 91.025 180.400 91.195 181.370 ;
        RECT 90.520 180.070 90.775 180.400 ;
        RECT 91.000 180.070 91.195 180.400 ;
        RECT 91.365 181.030 92.490 181.200 ;
        RECT 90.605 179.900 90.775 180.070 ;
        RECT 91.365 179.900 91.535 181.030 ;
        RECT 89.715 179.160 90.005 179.885 ;
        RECT 90.180 179.330 90.435 179.900 ;
        RECT 90.605 179.730 91.535 179.900 ;
        RECT 91.705 180.690 92.715 180.860 ;
        RECT 91.705 179.890 91.875 180.690 ;
        RECT 92.080 180.350 92.355 180.490 ;
        RECT 92.075 180.180 92.355 180.350 ;
        RECT 91.360 179.695 91.535 179.730 ;
        RECT 90.605 179.160 90.935 179.560 ;
        RECT 91.360 179.330 91.890 179.695 ;
        RECT 92.080 179.330 92.355 180.180 ;
        RECT 92.525 179.330 92.715 180.690 ;
        RECT 92.885 180.705 93.055 181.370 ;
        RECT 93.225 180.950 93.395 181.710 ;
        RECT 93.630 180.950 94.145 181.360 ;
        RECT 92.885 180.515 93.635 180.705 ;
        RECT 93.805 180.140 94.145 180.950 ;
        RECT 92.915 179.970 94.145 180.140 ;
        RECT 95.235 180.570 95.575 181.540 ;
        RECT 95.745 180.570 95.915 181.710 ;
        RECT 96.185 180.910 96.435 181.710 ;
        RECT 97.080 180.740 97.410 181.540 ;
        RECT 97.710 180.910 98.040 181.710 ;
        RECT 98.210 180.740 98.540 181.540 ;
        RECT 96.105 180.570 98.540 180.740 ;
        RECT 98.915 180.635 99.185 181.540 ;
        RECT 99.355 180.950 99.685 181.710 ;
        RECT 99.865 180.780 100.035 181.540 ;
        RECT 92.895 179.160 93.405 179.695 ;
        RECT 93.625 179.365 93.870 179.970 ;
        RECT 95.235 179.960 95.410 180.570 ;
        RECT 96.105 180.320 96.275 180.570 ;
        RECT 95.580 180.150 96.275 180.320 ;
        RECT 96.450 180.150 96.870 180.350 ;
        RECT 97.040 180.150 97.370 180.350 ;
        RECT 97.540 180.150 97.870 180.350 ;
        RECT 95.235 179.330 95.575 179.960 ;
        RECT 95.745 179.160 95.995 179.960 ;
        RECT 96.185 179.810 97.410 179.980 ;
        RECT 96.185 179.330 96.515 179.810 ;
        RECT 96.685 179.160 96.910 179.620 ;
        RECT 97.080 179.330 97.410 179.810 ;
        RECT 98.040 179.940 98.210 180.570 ;
        RECT 98.395 180.150 98.745 180.400 ;
        RECT 98.040 179.330 98.540 179.940 ;
        RECT 98.915 179.835 99.085 180.635 ;
        RECT 99.370 180.610 100.035 180.780 ;
        RECT 100.295 180.620 101.965 181.710 ;
        RECT 102.135 180.950 102.650 181.360 ;
        RECT 102.885 180.950 103.055 181.710 ;
        RECT 103.225 181.370 105.255 181.540 ;
        RECT 99.370 180.465 99.540 180.610 ;
        RECT 99.255 180.135 99.540 180.465 ;
        RECT 99.370 179.880 99.540 180.135 ;
        RECT 99.775 180.060 100.105 180.430 ;
        RECT 100.295 180.100 101.045 180.620 ;
        RECT 101.215 179.930 101.965 180.450 ;
        RECT 102.135 180.140 102.475 180.950 ;
        RECT 103.225 180.705 103.395 181.370 ;
        RECT 103.790 181.030 104.915 181.200 ;
        RECT 102.645 180.515 103.395 180.705 ;
        RECT 103.565 180.690 104.575 180.860 ;
        RECT 102.135 179.970 103.365 180.140 ;
        RECT 98.915 179.330 99.175 179.835 ;
        RECT 99.370 179.710 100.035 179.880 ;
        RECT 99.355 179.160 99.685 179.540 ;
        RECT 99.865 179.330 100.035 179.710 ;
        RECT 100.295 179.160 101.965 179.930 ;
        RECT 102.410 179.365 102.655 179.970 ;
        RECT 102.875 179.160 103.385 179.695 ;
        RECT 103.565 179.330 103.755 180.690 ;
        RECT 103.925 179.670 104.200 180.490 ;
        RECT 104.405 179.890 104.575 180.690 ;
        RECT 104.745 179.900 104.915 181.030 ;
        RECT 105.085 180.400 105.255 181.370 ;
        RECT 105.425 180.570 105.595 181.710 ;
        RECT 105.765 180.570 106.100 181.540 ;
        RECT 106.480 180.740 106.810 181.540 ;
        RECT 106.980 180.910 107.310 181.710 ;
        RECT 107.610 180.740 107.940 181.540 ;
        RECT 108.585 180.910 108.835 181.710 ;
        RECT 106.480 180.570 108.915 180.740 ;
        RECT 109.105 180.570 109.275 181.710 ;
        RECT 109.445 180.570 109.785 181.540 ;
        RECT 110.045 180.780 110.215 181.540 ;
        RECT 110.395 180.950 110.725 181.710 ;
        RECT 110.045 180.610 110.710 180.780 ;
        RECT 110.895 180.635 111.165 181.540 ;
        RECT 105.085 180.070 105.280 180.400 ;
        RECT 105.505 180.070 105.760 180.400 ;
        RECT 105.505 179.900 105.675 180.070 ;
        RECT 105.930 179.900 106.100 180.570 ;
        RECT 106.275 180.150 106.625 180.400 ;
        RECT 106.810 179.940 106.980 180.570 ;
        RECT 107.150 180.150 107.480 180.350 ;
        RECT 107.650 180.150 107.980 180.350 ;
        RECT 108.150 180.150 108.570 180.350 ;
        RECT 108.745 180.320 108.915 180.570 ;
        RECT 108.745 180.150 109.440 180.320 ;
        RECT 104.745 179.730 105.675 179.900 ;
        RECT 104.745 179.695 104.920 179.730 ;
        RECT 103.925 179.500 104.205 179.670 ;
        RECT 103.925 179.330 104.200 179.500 ;
        RECT 104.390 179.330 104.920 179.695 ;
        RECT 105.345 179.160 105.675 179.560 ;
        RECT 105.845 179.330 106.100 179.900 ;
        RECT 106.480 179.330 106.980 179.940 ;
        RECT 107.610 179.810 108.835 179.980 ;
        RECT 109.610 179.960 109.785 180.570 ;
        RECT 110.540 180.465 110.710 180.610 ;
        RECT 109.975 180.060 110.305 180.430 ;
        RECT 110.540 180.135 110.825 180.465 ;
        RECT 107.610 179.330 107.940 179.810 ;
        RECT 108.110 179.160 108.335 179.620 ;
        RECT 108.505 179.330 108.835 179.810 ;
        RECT 109.025 179.160 109.275 179.960 ;
        RECT 109.445 179.330 109.785 179.960 ;
        RECT 110.540 179.880 110.710 180.135 ;
        RECT 110.045 179.710 110.710 179.880 ;
        RECT 110.995 179.835 111.165 180.635 ;
        RECT 110.045 179.330 110.215 179.710 ;
        RECT 110.395 179.160 110.725 179.540 ;
        RECT 110.905 179.330 111.165 179.835 ;
        RECT 111.335 180.635 111.605 181.540 ;
        RECT 111.775 180.950 112.105 181.710 ;
        RECT 112.285 180.780 112.455 181.540 ;
        RECT 111.335 179.835 111.505 180.635 ;
        RECT 111.790 180.610 112.455 180.780 ;
        RECT 112.715 180.620 114.385 181.710 ;
        RECT 114.555 180.620 115.765 181.710 ;
        RECT 111.790 180.465 111.960 180.610 ;
        RECT 111.675 180.135 111.960 180.465 ;
        RECT 111.790 179.880 111.960 180.135 ;
        RECT 112.195 180.060 112.525 180.430 ;
        RECT 112.715 180.100 113.465 180.620 ;
        RECT 113.635 179.930 114.385 180.450 ;
        RECT 114.555 180.080 115.075 180.620 ;
        RECT 111.335 179.330 111.595 179.835 ;
        RECT 111.790 179.710 112.455 179.880 ;
        RECT 111.775 179.160 112.105 179.540 ;
        RECT 112.285 179.330 112.455 179.710 ;
        RECT 112.715 179.160 114.385 179.930 ;
        RECT 115.245 179.910 115.765 180.450 ;
        RECT 114.555 179.160 115.765 179.910 ;
        RECT 14.650 178.990 115.850 179.160 ;
        RECT 14.735 178.240 15.945 178.990 ;
        RECT 16.120 178.445 21.465 178.990 ;
        RECT 14.735 177.700 15.255 178.240 ;
        RECT 15.425 177.530 15.945 178.070 ;
        RECT 14.735 176.440 15.945 177.530 ;
        RECT 17.710 176.875 18.060 178.125 ;
        RECT 19.540 177.615 19.880 178.445 ;
        RECT 21.750 178.360 22.035 178.820 ;
        RECT 22.205 178.530 22.475 178.990 ;
        RECT 21.750 178.190 22.705 178.360 ;
        RECT 21.635 177.460 22.325 178.020 ;
        RECT 22.495 177.290 22.705 178.190 ;
        RECT 21.750 177.070 22.705 177.290 ;
        RECT 22.875 178.020 23.275 178.820 ;
        RECT 23.465 178.360 23.745 178.820 ;
        RECT 24.265 178.530 24.590 178.990 ;
        RECT 23.465 178.190 24.590 178.360 ;
        RECT 24.760 178.250 25.145 178.820 ;
        RECT 25.315 178.265 25.605 178.990 ;
        RECT 25.865 178.440 26.035 178.820 ;
        RECT 26.215 178.610 26.545 178.990 ;
        RECT 25.865 178.270 26.530 178.440 ;
        RECT 26.725 178.315 26.985 178.820 ;
        RECT 24.140 178.080 24.590 178.190 ;
        RECT 22.875 177.460 23.970 178.020 ;
        RECT 24.140 177.750 24.695 178.080 ;
        RECT 16.120 176.440 21.465 176.875 ;
        RECT 21.750 176.610 22.035 177.070 ;
        RECT 22.205 176.440 22.475 176.900 ;
        RECT 22.875 176.610 23.275 177.460 ;
        RECT 24.140 177.290 24.590 177.750 ;
        RECT 24.865 177.580 25.145 178.250 ;
        RECT 25.795 177.720 26.125 178.090 ;
        RECT 26.360 178.015 26.530 178.270 ;
        RECT 26.360 177.685 26.645 178.015 ;
        RECT 23.465 177.070 24.590 177.290 ;
        RECT 23.465 176.610 23.745 177.070 ;
        RECT 24.265 176.440 24.590 176.900 ;
        RECT 24.760 176.610 25.145 177.580 ;
        RECT 25.315 176.440 25.605 177.605 ;
        RECT 26.360 177.540 26.530 177.685 ;
        RECT 25.865 177.370 26.530 177.540 ;
        RECT 26.815 177.515 26.985 178.315 ;
        RECT 27.195 178.170 27.425 178.990 ;
        RECT 27.595 178.190 27.925 178.820 ;
        RECT 27.175 177.750 27.505 178.000 ;
        RECT 27.675 177.590 27.925 178.190 ;
        RECT 28.095 178.170 28.305 178.990 ;
        RECT 28.540 178.250 28.795 178.820 ;
        RECT 28.965 178.590 29.295 178.990 ;
        RECT 29.720 178.455 30.250 178.820 ;
        RECT 29.720 178.420 29.895 178.455 ;
        RECT 28.965 178.250 29.895 178.420 ;
        RECT 25.865 176.610 26.035 177.370 ;
        RECT 26.215 176.440 26.545 177.200 ;
        RECT 26.715 176.610 26.985 177.515 ;
        RECT 27.195 176.440 27.425 177.580 ;
        RECT 27.595 176.610 27.925 177.590 ;
        RECT 28.540 177.580 28.710 178.250 ;
        RECT 28.965 178.080 29.135 178.250 ;
        RECT 28.880 177.750 29.135 178.080 ;
        RECT 29.360 177.750 29.555 178.080 ;
        RECT 28.095 176.440 28.305 177.580 ;
        RECT 28.540 176.610 28.875 177.580 ;
        RECT 29.045 176.440 29.215 177.580 ;
        RECT 29.385 176.780 29.555 177.750 ;
        RECT 29.725 177.120 29.895 178.250 ;
        RECT 30.065 177.460 30.235 178.260 ;
        RECT 30.440 177.970 30.715 178.820 ;
        RECT 30.435 177.800 30.715 177.970 ;
        RECT 30.440 177.660 30.715 177.800 ;
        RECT 30.885 177.460 31.075 178.820 ;
        RECT 31.255 178.455 31.765 178.990 ;
        RECT 31.985 178.180 32.230 178.785 ;
        RECT 33.410 178.180 33.655 178.785 ;
        RECT 33.875 178.455 34.385 178.990 ;
        RECT 31.275 178.010 32.505 178.180 ;
        RECT 30.065 177.290 31.075 177.460 ;
        RECT 31.245 177.445 31.995 177.635 ;
        RECT 29.725 176.950 30.850 177.120 ;
        RECT 31.245 176.780 31.415 177.445 ;
        RECT 32.165 177.200 32.505 178.010 ;
        RECT 29.385 176.610 31.415 176.780 ;
        RECT 31.585 176.440 31.755 177.200 ;
        RECT 31.990 176.790 32.505 177.200 ;
        RECT 33.135 178.010 34.365 178.180 ;
        RECT 33.135 177.200 33.475 178.010 ;
        RECT 33.645 177.445 34.395 177.635 ;
        RECT 33.135 176.790 33.650 177.200 ;
        RECT 33.885 176.440 34.055 177.200 ;
        RECT 34.225 176.780 34.395 177.445 ;
        RECT 34.565 177.460 34.755 178.820 ;
        RECT 34.925 178.310 35.200 178.820 ;
        RECT 35.390 178.455 35.920 178.820 ;
        RECT 36.345 178.590 36.675 178.990 ;
        RECT 35.745 178.420 35.920 178.455 ;
        RECT 34.925 178.140 35.205 178.310 ;
        RECT 34.925 177.660 35.200 178.140 ;
        RECT 35.405 177.460 35.575 178.260 ;
        RECT 34.565 177.290 35.575 177.460 ;
        RECT 35.745 178.250 36.675 178.420 ;
        RECT 36.845 178.250 37.100 178.820 ;
        RECT 35.745 177.120 35.915 178.250 ;
        RECT 36.505 178.080 36.675 178.250 ;
        RECT 34.790 176.950 35.915 177.120 ;
        RECT 36.085 177.750 36.280 178.080 ;
        RECT 36.505 177.750 36.760 178.080 ;
        RECT 36.085 176.780 36.255 177.750 ;
        RECT 36.930 177.580 37.100 178.250 ;
        RECT 37.735 178.220 40.325 178.990 ;
        RECT 34.225 176.610 36.255 176.780 ;
        RECT 36.425 176.440 36.595 177.580 ;
        RECT 36.765 176.610 37.100 177.580 ;
        RECT 37.735 177.530 38.945 178.050 ;
        RECT 39.115 177.700 40.325 178.220 ;
        RECT 40.495 178.190 40.835 178.820 ;
        RECT 41.005 178.190 41.255 178.990 ;
        RECT 41.445 178.340 41.775 178.820 ;
        RECT 41.945 178.530 42.170 178.990 ;
        RECT 42.340 178.340 42.670 178.820 ;
        RECT 40.495 177.580 40.670 178.190 ;
        RECT 41.445 178.170 42.670 178.340 ;
        RECT 43.300 178.210 43.800 178.820 ;
        RECT 44.175 178.220 46.765 178.990 ;
        RECT 40.840 177.830 41.535 178.000 ;
        RECT 41.365 177.580 41.535 177.830 ;
        RECT 41.710 177.800 42.130 178.000 ;
        RECT 42.300 177.800 42.630 178.000 ;
        RECT 42.800 177.800 43.130 178.000 ;
        RECT 43.300 177.580 43.470 178.210 ;
        RECT 43.655 177.750 44.005 178.000 ;
        RECT 37.735 176.440 40.325 177.530 ;
        RECT 40.495 176.610 40.835 177.580 ;
        RECT 41.005 176.440 41.175 177.580 ;
        RECT 41.365 177.410 43.800 177.580 ;
        RECT 41.445 176.440 41.695 177.240 ;
        RECT 42.340 176.610 42.670 177.410 ;
        RECT 42.970 176.440 43.300 177.240 ;
        RECT 43.470 176.610 43.800 177.410 ;
        RECT 44.175 177.530 45.385 178.050 ;
        RECT 45.555 177.700 46.765 178.220 ;
        RECT 47.210 178.180 47.455 178.785 ;
        RECT 47.675 178.455 48.185 178.990 ;
        RECT 46.935 178.010 48.165 178.180 ;
        RECT 44.175 176.440 46.765 177.530 ;
        RECT 46.935 177.200 47.275 178.010 ;
        RECT 47.445 177.445 48.195 177.635 ;
        RECT 46.935 176.790 47.450 177.200 ;
        RECT 47.685 176.440 47.855 177.200 ;
        RECT 48.025 176.780 48.195 177.445 ;
        RECT 48.365 177.460 48.555 178.820 ;
        RECT 48.725 177.970 49.000 178.820 ;
        RECT 49.190 178.455 49.720 178.820 ;
        RECT 50.145 178.590 50.475 178.990 ;
        RECT 49.545 178.420 49.720 178.455 ;
        RECT 48.725 177.800 49.005 177.970 ;
        RECT 48.725 177.660 49.000 177.800 ;
        RECT 49.205 177.460 49.375 178.260 ;
        RECT 48.365 177.290 49.375 177.460 ;
        RECT 49.545 178.250 50.475 178.420 ;
        RECT 50.645 178.250 50.900 178.820 ;
        RECT 51.075 178.265 51.365 178.990 ;
        RECT 51.650 178.360 51.935 178.820 ;
        RECT 52.105 178.530 52.375 178.990 ;
        RECT 49.545 177.120 49.715 178.250 ;
        RECT 50.305 178.080 50.475 178.250 ;
        RECT 48.590 176.950 49.715 177.120 ;
        RECT 49.885 177.750 50.080 178.080 ;
        RECT 50.305 177.750 50.560 178.080 ;
        RECT 49.885 176.780 50.055 177.750 ;
        RECT 50.730 177.580 50.900 178.250 ;
        RECT 51.650 178.190 52.605 178.360 ;
        RECT 48.025 176.610 50.055 176.780 ;
        RECT 50.225 176.440 50.395 177.580 ;
        RECT 50.565 176.610 50.900 177.580 ;
        RECT 51.075 176.440 51.365 177.605 ;
        RECT 51.535 177.460 52.225 178.020 ;
        RECT 52.395 177.290 52.605 178.190 ;
        RECT 51.650 177.070 52.605 177.290 ;
        RECT 52.775 178.020 53.175 178.820 ;
        RECT 53.365 178.360 53.645 178.820 ;
        RECT 54.165 178.530 54.490 178.990 ;
        RECT 53.365 178.190 54.490 178.360 ;
        RECT 54.660 178.250 55.045 178.820 ;
        RECT 55.275 178.510 55.555 178.990 ;
        RECT 55.725 178.340 55.985 178.730 ;
        RECT 56.160 178.510 56.415 178.990 ;
        RECT 56.585 178.340 56.880 178.730 ;
        RECT 57.060 178.510 57.335 178.990 ;
        RECT 57.505 178.490 57.805 178.820 ;
        RECT 54.040 178.080 54.490 178.190 ;
        RECT 52.775 177.460 53.870 178.020 ;
        RECT 54.040 177.750 54.595 178.080 ;
        RECT 51.650 176.610 51.935 177.070 ;
        RECT 52.105 176.440 52.375 176.900 ;
        RECT 52.775 176.610 53.175 177.460 ;
        RECT 54.040 177.290 54.490 177.750 ;
        RECT 54.765 177.580 55.045 178.250 ;
        RECT 53.365 177.070 54.490 177.290 ;
        RECT 53.365 176.610 53.645 177.070 ;
        RECT 54.165 176.440 54.490 176.900 ;
        RECT 54.660 176.610 55.045 177.580 ;
        RECT 55.230 178.170 56.880 178.340 ;
        RECT 55.230 177.660 55.635 178.170 ;
        RECT 55.805 177.830 56.945 178.000 ;
        RECT 55.230 177.490 55.985 177.660 ;
        RECT 55.270 176.440 55.555 177.310 ;
        RECT 55.725 177.240 55.985 177.490 ;
        RECT 56.775 177.580 56.945 177.830 ;
        RECT 57.115 177.750 57.465 178.320 ;
        RECT 57.635 177.580 57.805 178.490 ;
        RECT 56.775 177.410 57.805 177.580 ;
        RECT 55.725 177.070 56.845 177.240 ;
        RECT 55.725 176.610 55.985 177.070 ;
        RECT 56.160 176.440 56.415 176.900 ;
        RECT 56.585 176.610 56.845 177.070 ;
        RECT 57.015 176.440 57.325 177.240 ;
        RECT 57.495 176.610 57.805 177.410 ;
        RECT 57.975 178.315 58.235 178.820 ;
        RECT 58.415 178.610 58.745 178.990 ;
        RECT 58.925 178.440 59.095 178.820 ;
        RECT 57.975 177.515 58.145 178.315 ;
        RECT 58.430 178.270 59.095 178.440 ;
        RECT 58.430 178.015 58.600 178.270 ;
        RECT 59.815 178.220 62.405 178.990 ;
        RECT 58.315 177.685 58.600 178.015 ;
        RECT 58.835 177.720 59.165 178.090 ;
        RECT 58.430 177.540 58.600 177.685 ;
        RECT 57.975 176.610 58.245 177.515 ;
        RECT 58.430 177.370 59.095 177.540 ;
        RECT 58.415 176.440 58.745 177.200 ;
        RECT 58.925 176.610 59.095 177.370 ;
        RECT 59.815 177.530 61.025 178.050 ;
        RECT 61.195 177.700 62.405 178.220 ;
        RECT 62.615 178.170 62.845 178.990 ;
        RECT 63.015 178.190 63.345 178.820 ;
        RECT 62.595 177.750 62.925 178.000 ;
        RECT 63.095 177.590 63.345 178.190 ;
        RECT 63.515 178.170 63.725 178.990 ;
        RECT 63.960 178.150 64.220 178.990 ;
        RECT 64.395 178.245 64.650 178.820 ;
        RECT 64.820 178.610 65.150 178.990 ;
        RECT 65.365 178.440 65.535 178.820 ;
        RECT 66.065 178.595 66.395 178.990 ;
        RECT 64.820 178.270 65.535 178.440 ;
        RECT 66.565 178.420 66.765 178.775 ;
        RECT 66.935 178.590 67.265 178.990 ;
        RECT 67.435 178.420 67.635 178.765 ;
        RECT 59.815 176.440 62.405 177.530 ;
        RECT 62.615 176.440 62.845 177.580 ;
        RECT 63.015 176.610 63.345 177.590 ;
        RECT 63.515 176.440 63.725 177.580 ;
        RECT 63.960 176.440 64.220 177.590 ;
        RECT 64.395 177.515 64.565 178.245 ;
        RECT 64.820 178.080 64.990 178.270 ;
        RECT 65.795 178.250 67.635 178.420 ;
        RECT 67.805 178.250 68.135 178.990 ;
        RECT 68.370 178.420 68.540 178.670 ;
        RECT 70.205 178.595 70.535 178.990 ;
        RECT 70.705 178.420 70.905 178.775 ;
        RECT 71.075 178.590 71.405 178.990 ;
        RECT 71.575 178.420 71.775 178.765 ;
        RECT 68.370 178.250 68.845 178.420 ;
        RECT 64.735 177.750 64.990 178.080 ;
        RECT 64.820 177.540 64.990 177.750 ;
        RECT 65.270 177.720 65.625 178.090 ;
        RECT 64.395 176.610 64.650 177.515 ;
        RECT 64.820 177.370 65.535 177.540 ;
        RECT 64.820 176.440 65.150 177.200 ;
        RECT 65.365 176.610 65.535 177.370 ;
        RECT 65.795 176.625 66.055 178.250 ;
        RECT 66.235 177.280 66.455 178.080 ;
        RECT 66.695 177.460 66.995 178.080 ;
        RECT 67.165 177.460 67.495 178.080 ;
        RECT 67.665 177.460 67.985 178.080 ;
        RECT 68.155 177.460 68.505 178.080 ;
        RECT 68.675 177.280 68.845 178.250 ;
        RECT 66.235 177.070 68.845 177.280 ;
        RECT 69.935 178.250 71.775 178.420 ;
        RECT 71.945 178.250 72.275 178.990 ;
        RECT 72.510 178.420 72.680 178.670 ;
        RECT 72.510 178.250 72.985 178.420 ;
        RECT 67.805 176.440 68.135 176.890 ;
        RECT 69.935 176.625 70.195 178.250 ;
        RECT 70.375 177.280 70.595 178.080 ;
        RECT 70.835 177.460 71.135 178.080 ;
        RECT 71.305 177.460 71.635 178.080 ;
        RECT 71.805 177.460 72.125 178.080 ;
        RECT 72.295 177.460 72.645 178.080 ;
        RECT 72.815 177.280 72.985 178.250 ;
        RECT 70.375 177.070 72.985 177.280 ;
        RECT 73.155 178.190 73.495 178.820 ;
        RECT 73.665 178.190 73.915 178.990 ;
        RECT 74.105 178.340 74.435 178.820 ;
        RECT 74.605 178.530 74.830 178.990 ;
        RECT 75.000 178.340 75.330 178.820 ;
        RECT 73.155 177.580 73.330 178.190 ;
        RECT 74.105 178.170 75.330 178.340 ;
        RECT 75.960 178.210 76.460 178.820 ;
        RECT 76.835 178.265 77.125 178.990 ;
        RECT 77.295 178.220 78.965 178.990 ;
        RECT 73.500 177.830 74.195 178.000 ;
        RECT 74.025 177.580 74.195 177.830 ;
        RECT 74.370 177.800 74.790 178.000 ;
        RECT 74.960 177.800 75.290 178.000 ;
        RECT 75.460 177.800 75.790 178.000 ;
        RECT 75.960 177.580 76.130 178.210 ;
        RECT 76.315 177.750 76.665 178.000 ;
        RECT 71.945 176.440 72.275 176.890 ;
        RECT 73.155 176.610 73.495 177.580 ;
        RECT 73.665 176.440 73.835 177.580 ;
        RECT 74.025 177.410 76.460 177.580 ;
        RECT 74.105 176.440 74.355 177.240 ;
        RECT 75.000 176.610 75.330 177.410 ;
        RECT 75.630 176.440 75.960 177.240 ;
        RECT 76.130 176.610 76.460 177.410 ;
        RECT 76.835 176.440 77.125 177.605 ;
        RECT 77.295 177.530 78.045 178.050 ;
        RECT 78.215 177.700 78.965 178.220 ;
        RECT 79.250 178.360 79.535 178.820 ;
        RECT 79.705 178.530 79.975 178.990 ;
        RECT 79.250 178.190 80.205 178.360 ;
        RECT 77.295 176.440 78.965 177.530 ;
        RECT 79.135 177.460 79.825 178.020 ;
        RECT 79.995 177.290 80.205 178.190 ;
        RECT 79.250 177.070 80.205 177.290 ;
        RECT 80.375 178.020 80.775 178.820 ;
        RECT 80.965 178.360 81.245 178.820 ;
        RECT 81.765 178.530 82.090 178.990 ;
        RECT 80.965 178.190 82.090 178.360 ;
        RECT 82.260 178.250 82.645 178.820 ;
        RECT 81.640 178.080 82.090 178.190 ;
        RECT 80.375 177.460 81.470 178.020 ;
        RECT 81.640 177.750 82.195 178.080 ;
        RECT 79.250 176.610 79.535 177.070 ;
        RECT 79.705 176.440 79.975 176.900 ;
        RECT 80.375 176.610 80.775 177.460 ;
        RECT 81.640 177.290 82.090 177.750 ;
        RECT 82.365 177.580 82.645 178.250 ;
        RECT 82.905 178.340 83.075 178.820 ;
        RECT 83.255 178.510 83.495 178.990 ;
        RECT 83.745 178.340 83.915 178.820 ;
        RECT 84.085 178.510 84.415 178.990 ;
        RECT 84.585 178.340 84.755 178.820 ;
        RECT 82.905 178.170 83.540 178.340 ;
        RECT 83.745 178.170 84.755 178.340 ;
        RECT 84.925 178.190 85.255 178.990 ;
        RECT 85.665 178.440 85.835 178.820 ;
        RECT 86.015 178.610 86.345 178.990 ;
        RECT 85.665 178.270 86.330 178.440 ;
        RECT 86.525 178.315 86.785 178.820 ;
        RECT 83.370 178.000 83.540 178.170 ;
        RECT 82.820 177.760 83.200 178.000 ;
        RECT 83.370 177.830 83.870 178.000 ;
        RECT 83.370 177.590 83.540 177.830 ;
        RECT 84.260 177.630 84.755 178.170 ;
        RECT 85.595 177.720 85.925 178.090 ;
        RECT 86.160 178.015 86.330 178.270 ;
        RECT 80.965 177.070 82.090 177.290 ;
        RECT 80.965 176.610 81.245 177.070 ;
        RECT 81.765 176.440 82.090 176.900 ;
        RECT 82.260 176.610 82.645 177.580 ;
        RECT 82.825 177.420 83.540 177.590 ;
        RECT 83.745 177.460 84.755 177.630 ;
        RECT 86.160 177.685 86.445 178.015 ;
        RECT 82.825 176.610 83.155 177.420 ;
        RECT 83.325 176.440 83.565 177.240 ;
        RECT 83.745 176.610 83.915 177.460 ;
        RECT 84.085 176.440 84.415 177.240 ;
        RECT 84.585 176.610 84.755 177.460 ;
        RECT 84.925 176.440 85.255 177.590 ;
        RECT 86.160 177.540 86.330 177.685 ;
        RECT 85.665 177.370 86.330 177.540 ;
        RECT 86.615 177.515 86.785 178.315 ;
        RECT 85.665 176.610 85.835 177.370 ;
        RECT 86.015 176.440 86.345 177.200 ;
        RECT 86.515 176.610 86.785 177.515 ;
        RECT 86.955 178.250 87.340 178.820 ;
        RECT 87.510 178.530 87.835 178.990 ;
        RECT 88.355 178.360 88.635 178.820 ;
        RECT 86.955 177.580 87.235 178.250 ;
        RECT 87.510 178.190 88.635 178.360 ;
        RECT 87.510 178.080 87.960 178.190 ;
        RECT 87.405 177.750 87.960 178.080 ;
        RECT 88.825 178.020 89.225 178.820 ;
        RECT 89.625 178.530 89.895 178.990 ;
        RECT 90.065 178.360 90.350 178.820 ;
        RECT 86.955 176.610 87.340 177.580 ;
        RECT 87.510 177.290 87.960 177.750 ;
        RECT 88.130 177.460 89.225 178.020 ;
        RECT 87.510 177.070 88.635 177.290 ;
        RECT 87.510 176.440 87.835 176.900 ;
        RECT 88.355 176.610 88.635 177.070 ;
        RECT 88.825 176.610 89.225 177.460 ;
        RECT 89.395 178.190 90.350 178.360 ;
        RECT 90.635 178.190 90.975 178.820 ;
        RECT 91.145 178.190 91.395 178.990 ;
        RECT 91.585 178.340 91.915 178.820 ;
        RECT 92.085 178.530 92.310 178.990 ;
        RECT 92.480 178.340 92.810 178.820 ;
        RECT 89.395 177.290 89.605 178.190 ;
        RECT 89.775 177.460 90.465 178.020 ;
        RECT 90.635 177.580 90.810 178.190 ;
        RECT 91.585 178.170 92.810 178.340 ;
        RECT 93.440 178.210 93.940 178.820 ;
        RECT 90.980 177.830 91.675 178.000 ;
        RECT 91.505 177.580 91.675 177.830 ;
        RECT 91.850 177.800 92.270 178.000 ;
        RECT 92.440 177.800 92.770 178.000 ;
        RECT 92.940 177.800 93.270 178.000 ;
        RECT 93.440 177.580 93.610 178.210 ;
        RECT 94.315 178.190 94.655 178.820 ;
        RECT 94.825 178.190 95.075 178.990 ;
        RECT 95.265 178.340 95.595 178.820 ;
        RECT 95.765 178.530 95.990 178.990 ;
        RECT 96.160 178.340 96.490 178.820 ;
        RECT 93.795 177.750 94.145 178.000 ;
        RECT 94.315 177.580 94.490 178.190 ;
        RECT 95.265 178.170 96.490 178.340 ;
        RECT 97.120 178.210 97.620 178.820 ;
        RECT 99.120 178.210 99.620 178.820 ;
        RECT 94.660 177.830 95.355 178.000 ;
        RECT 95.185 177.580 95.355 177.830 ;
        RECT 95.530 177.800 95.950 178.000 ;
        RECT 96.120 177.800 96.450 178.000 ;
        RECT 96.620 177.800 96.950 178.000 ;
        RECT 97.120 177.580 97.290 178.210 ;
        RECT 97.475 177.750 97.825 178.000 ;
        RECT 98.915 177.750 99.265 178.000 ;
        RECT 99.450 177.580 99.620 178.210 ;
        RECT 100.250 178.340 100.580 178.820 ;
        RECT 100.750 178.530 100.975 178.990 ;
        RECT 101.145 178.340 101.475 178.820 ;
        RECT 100.250 178.170 101.475 178.340 ;
        RECT 101.665 178.190 101.915 178.990 ;
        RECT 102.085 178.190 102.425 178.820 ;
        RECT 102.595 178.265 102.885 178.990 ;
        RECT 104.090 178.360 104.375 178.820 ;
        RECT 104.545 178.530 104.815 178.990 ;
        RECT 104.090 178.190 105.045 178.360 ;
        RECT 99.790 177.800 100.120 178.000 ;
        RECT 100.290 177.800 100.620 178.000 ;
        RECT 100.790 177.800 101.210 178.000 ;
        RECT 101.385 177.830 102.080 178.000 ;
        RECT 101.385 177.580 101.555 177.830 ;
        RECT 102.250 177.580 102.425 178.190 ;
        RECT 89.395 177.070 90.350 177.290 ;
        RECT 89.625 176.440 89.895 176.900 ;
        RECT 90.065 176.610 90.350 177.070 ;
        RECT 90.635 176.610 90.975 177.580 ;
        RECT 91.145 176.440 91.315 177.580 ;
        RECT 91.505 177.410 93.940 177.580 ;
        RECT 91.585 176.440 91.835 177.240 ;
        RECT 92.480 176.610 92.810 177.410 ;
        RECT 93.110 176.440 93.440 177.240 ;
        RECT 93.610 176.610 93.940 177.410 ;
        RECT 94.315 176.610 94.655 177.580 ;
        RECT 94.825 176.440 94.995 177.580 ;
        RECT 95.185 177.410 97.620 177.580 ;
        RECT 95.265 176.440 95.515 177.240 ;
        RECT 96.160 176.610 96.490 177.410 ;
        RECT 96.790 176.440 97.120 177.240 ;
        RECT 97.290 176.610 97.620 177.410 ;
        RECT 99.120 177.410 101.555 177.580 ;
        RECT 99.120 176.610 99.450 177.410 ;
        RECT 99.620 176.440 99.950 177.240 ;
        RECT 100.250 176.610 100.580 177.410 ;
        RECT 101.225 176.440 101.475 177.240 ;
        RECT 101.745 176.440 101.915 177.580 ;
        RECT 102.085 176.610 102.425 177.580 ;
        RECT 102.595 176.440 102.885 177.605 ;
        RECT 103.975 177.460 104.665 178.020 ;
        RECT 104.835 177.290 105.045 178.190 ;
        RECT 104.090 177.070 105.045 177.290 ;
        RECT 105.215 178.020 105.615 178.820 ;
        RECT 105.805 178.360 106.085 178.820 ;
        RECT 106.605 178.530 106.930 178.990 ;
        RECT 105.805 178.190 106.930 178.360 ;
        RECT 107.100 178.250 107.485 178.820 ;
        RECT 106.480 178.080 106.930 178.190 ;
        RECT 105.215 177.460 106.310 178.020 ;
        RECT 106.480 177.750 107.035 178.080 ;
        RECT 104.090 176.610 104.375 177.070 ;
        RECT 104.545 176.440 104.815 176.900 ;
        RECT 105.215 176.610 105.615 177.460 ;
        RECT 106.480 177.290 106.930 177.750 ;
        RECT 107.205 177.580 107.485 178.250 ;
        RECT 107.655 178.240 108.865 178.990 ;
        RECT 109.125 178.440 109.295 178.820 ;
        RECT 109.475 178.610 109.805 178.990 ;
        RECT 109.125 178.270 109.790 178.440 ;
        RECT 109.985 178.315 110.245 178.820 ;
        RECT 105.805 177.070 106.930 177.290 ;
        RECT 105.805 176.610 106.085 177.070 ;
        RECT 106.605 176.440 106.930 176.900 ;
        RECT 107.100 176.610 107.485 177.580 ;
        RECT 107.655 177.530 108.175 178.070 ;
        RECT 108.345 177.700 108.865 178.240 ;
        RECT 109.055 177.720 109.385 178.090 ;
        RECT 109.620 178.015 109.790 178.270 ;
        RECT 109.620 177.685 109.905 178.015 ;
        RECT 109.620 177.540 109.790 177.685 ;
        RECT 107.655 176.440 108.865 177.530 ;
        RECT 109.125 177.370 109.790 177.540 ;
        RECT 110.075 177.515 110.245 178.315 ;
        RECT 110.875 178.220 114.385 178.990 ;
        RECT 114.555 178.240 115.765 178.990 ;
        RECT 109.125 176.610 109.295 177.370 ;
        RECT 109.475 176.440 109.805 177.200 ;
        RECT 109.975 176.610 110.245 177.515 ;
        RECT 110.875 177.530 112.565 178.050 ;
        RECT 112.735 177.700 114.385 178.220 ;
        RECT 114.555 177.530 115.075 178.070 ;
        RECT 115.245 177.700 115.765 178.240 ;
        RECT 110.875 176.440 114.385 177.530 ;
        RECT 114.555 176.440 115.765 177.530 ;
        RECT 14.650 176.270 115.850 176.440 ;
        RECT 14.735 175.180 15.945 176.270 ;
        RECT 14.735 174.470 15.255 175.010 ;
        RECT 15.425 174.640 15.945 175.180 ;
        RECT 17.035 175.180 20.545 176.270 ;
        RECT 20.920 175.300 21.250 176.100 ;
        RECT 21.420 175.470 21.750 176.270 ;
        RECT 22.050 175.300 22.380 176.100 ;
        RECT 23.025 175.470 23.275 176.270 ;
        RECT 17.035 174.660 18.725 175.180 ;
        RECT 20.920 175.130 23.355 175.300 ;
        RECT 23.545 175.130 23.715 176.270 ;
        RECT 23.885 175.130 24.225 176.100 ;
        RECT 24.510 175.640 24.795 176.100 ;
        RECT 24.965 175.810 25.235 176.270 ;
        RECT 24.510 175.420 25.465 175.640 ;
        RECT 18.895 174.490 20.545 175.010 ;
        RECT 20.715 174.710 21.065 174.960 ;
        RECT 21.250 174.500 21.420 175.130 ;
        RECT 21.590 174.710 21.920 174.910 ;
        RECT 22.090 174.710 22.420 174.910 ;
        RECT 22.590 174.710 23.010 174.910 ;
        RECT 23.185 174.880 23.355 175.130 ;
        RECT 23.185 174.710 23.880 174.880 ;
        RECT 14.735 173.720 15.945 174.470 ;
        RECT 17.035 173.720 20.545 174.490 ;
        RECT 20.920 173.890 21.420 174.500 ;
        RECT 22.050 174.370 23.275 174.540 ;
        RECT 24.050 174.520 24.225 175.130 ;
        RECT 24.395 174.690 25.085 175.250 ;
        RECT 25.255 174.520 25.465 175.420 ;
        RECT 22.050 173.890 22.380 174.370 ;
        RECT 22.550 173.720 22.775 174.180 ;
        RECT 22.945 173.890 23.275 174.370 ;
        RECT 23.465 173.720 23.715 174.520 ;
        RECT 23.885 173.890 24.225 174.520 ;
        RECT 24.510 174.350 25.465 174.520 ;
        RECT 25.635 175.250 26.035 176.100 ;
        RECT 26.225 175.640 26.505 176.100 ;
        RECT 27.025 175.810 27.350 176.270 ;
        RECT 26.225 175.420 27.350 175.640 ;
        RECT 25.635 174.690 26.730 175.250 ;
        RECT 26.900 174.960 27.350 175.420 ;
        RECT 27.520 175.130 27.905 176.100 ;
        RECT 24.510 173.890 24.795 174.350 ;
        RECT 24.965 173.720 25.235 174.180 ;
        RECT 25.635 173.890 26.035 174.690 ;
        RECT 26.900 174.630 27.455 174.960 ;
        RECT 26.900 174.520 27.350 174.630 ;
        RECT 26.225 174.350 27.350 174.520 ;
        RECT 27.625 174.460 27.905 175.130 ;
        RECT 26.225 173.890 26.505 174.350 ;
        RECT 27.025 173.720 27.350 174.180 ;
        RECT 27.520 173.890 27.905 174.460 ;
        RECT 28.080 175.080 28.335 175.960 ;
        RECT 28.505 175.130 28.810 176.270 ;
        RECT 29.150 175.890 29.480 176.270 ;
        RECT 29.660 175.720 29.830 176.010 ;
        RECT 30.000 175.810 30.250 176.270 ;
        RECT 29.030 175.550 29.830 175.720 ;
        RECT 30.420 175.760 31.290 176.100 ;
        RECT 28.080 174.430 28.290 175.080 ;
        RECT 29.030 174.960 29.200 175.550 ;
        RECT 30.420 175.380 30.590 175.760 ;
        RECT 31.525 175.640 31.695 176.100 ;
        RECT 31.865 175.810 32.235 176.270 ;
        RECT 32.530 175.670 32.700 176.010 ;
        RECT 32.870 175.840 33.200 176.270 ;
        RECT 33.435 175.670 33.605 176.010 ;
        RECT 29.370 175.210 30.590 175.380 ;
        RECT 30.760 175.300 31.220 175.590 ;
        RECT 31.525 175.470 32.085 175.640 ;
        RECT 32.530 175.500 33.605 175.670 ;
        RECT 33.775 175.770 34.455 176.100 ;
        RECT 34.670 175.770 34.920 176.100 ;
        RECT 35.090 175.810 35.340 176.270 ;
        RECT 31.915 175.330 32.085 175.470 ;
        RECT 30.760 175.290 31.725 175.300 ;
        RECT 30.420 175.120 30.590 175.210 ;
        RECT 31.050 175.130 31.725 175.290 ;
        RECT 28.460 174.930 29.200 174.960 ;
        RECT 28.460 174.630 29.375 174.930 ;
        RECT 29.050 174.455 29.375 174.630 ;
        RECT 28.080 173.900 28.335 174.430 ;
        RECT 28.505 173.720 28.810 174.180 ;
        RECT 29.055 174.100 29.375 174.455 ;
        RECT 29.545 174.670 30.085 175.040 ;
        RECT 30.420 174.950 30.825 175.120 ;
        RECT 29.545 174.270 29.785 174.670 ;
        RECT 30.265 174.500 30.485 174.780 ;
        RECT 29.955 174.330 30.485 174.500 ;
        RECT 29.955 174.100 30.125 174.330 ;
        RECT 30.655 174.170 30.825 174.950 ;
        RECT 30.995 174.340 31.345 174.960 ;
        RECT 31.515 174.340 31.725 175.130 ;
        RECT 31.915 175.160 33.415 175.330 ;
        RECT 31.915 174.470 32.085 175.160 ;
        RECT 33.775 174.990 33.945 175.770 ;
        RECT 34.750 175.640 34.920 175.770 ;
        RECT 32.255 174.820 33.945 174.990 ;
        RECT 34.115 175.210 34.580 175.600 ;
        RECT 34.750 175.470 35.145 175.640 ;
        RECT 32.255 174.640 32.425 174.820 ;
        RECT 29.055 173.930 30.125 174.100 ;
        RECT 30.295 173.720 30.485 174.160 ;
        RECT 30.655 173.890 31.605 174.170 ;
        RECT 31.915 174.080 32.175 174.470 ;
        RECT 32.595 174.400 33.385 174.650 ;
        RECT 31.825 173.910 32.175 174.080 ;
        RECT 32.385 173.720 32.715 174.180 ;
        RECT 33.590 174.110 33.760 174.820 ;
        RECT 34.115 174.620 34.285 175.210 ;
        RECT 33.930 174.400 34.285 174.620 ;
        RECT 34.455 174.400 34.805 175.020 ;
        RECT 34.975 174.110 35.145 175.470 ;
        RECT 35.510 175.300 35.835 176.085 ;
        RECT 35.315 174.250 35.775 175.300 ;
        RECT 33.590 173.940 34.445 174.110 ;
        RECT 34.650 173.940 35.145 174.110 ;
        RECT 35.315 173.720 35.645 174.080 ;
        RECT 36.005 173.980 36.175 176.100 ;
        RECT 36.345 175.770 36.675 176.270 ;
        RECT 36.845 175.600 37.100 176.100 ;
        RECT 36.350 175.430 37.100 175.600 ;
        RECT 36.350 174.440 36.580 175.430 ;
        RECT 36.750 174.610 37.100 175.260 ;
        RECT 38.195 175.105 38.485 176.270 ;
        RECT 38.655 175.195 38.925 176.100 ;
        RECT 39.095 175.510 39.425 176.270 ;
        RECT 39.605 175.340 39.775 176.100 ;
        RECT 36.350 174.270 37.100 174.440 ;
        RECT 36.345 173.720 36.675 174.100 ;
        RECT 36.845 173.980 37.100 174.270 ;
        RECT 38.195 173.720 38.485 174.445 ;
        RECT 38.655 174.395 38.825 175.195 ;
        RECT 39.110 175.170 39.775 175.340 ;
        RECT 40.700 175.300 41.030 176.100 ;
        RECT 41.200 175.470 41.530 176.270 ;
        RECT 41.830 175.300 42.160 176.100 ;
        RECT 42.805 175.470 43.055 176.270 ;
        RECT 39.110 175.025 39.280 175.170 ;
        RECT 40.700 175.130 43.135 175.300 ;
        RECT 43.325 175.130 43.495 176.270 ;
        RECT 43.665 175.130 44.005 176.100 ;
        RECT 44.290 175.640 44.575 176.100 ;
        RECT 44.745 175.810 45.015 176.270 ;
        RECT 44.290 175.420 45.245 175.640 ;
        RECT 38.995 174.695 39.280 175.025 ;
        RECT 39.110 174.440 39.280 174.695 ;
        RECT 39.515 174.620 39.845 174.990 ;
        RECT 40.495 174.710 40.845 174.960 ;
        RECT 41.030 174.500 41.200 175.130 ;
        RECT 41.370 174.710 41.700 174.910 ;
        RECT 41.870 174.710 42.200 174.910 ;
        RECT 42.370 174.710 42.790 174.910 ;
        RECT 42.965 174.880 43.135 175.130 ;
        RECT 42.965 174.710 43.660 174.880 ;
        RECT 38.655 173.890 38.915 174.395 ;
        RECT 39.110 174.270 39.775 174.440 ;
        RECT 39.095 173.720 39.425 174.100 ;
        RECT 39.605 173.890 39.775 174.270 ;
        RECT 40.700 173.890 41.200 174.500 ;
        RECT 41.830 174.370 43.055 174.540 ;
        RECT 43.830 174.520 44.005 175.130 ;
        RECT 44.175 174.690 44.865 175.250 ;
        RECT 45.035 174.520 45.245 175.420 ;
        RECT 41.830 173.890 42.160 174.370 ;
        RECT 42.330 173.720 42.555 174.180 ;
        RECT 42.725 173.890 43.055 174.370 ;
        RECT 43.245 173.720 43.495 174.520 ;
        RECT 43.665 173.890 44.005 174.520 ;
        RECT 44.290 174.350 45.245 174.520 ;
        RECT 45.415 175.250 45.815 176.100 ;
        RECT 46.005 175.640 46.285 176.100 ;
        RECT 46.805 175.810 47.130 176.270 ;
        RECT 46.005 175.420 47.130 175.640 ;
        RECT 45.415 174.690 46.510 175.250 ;
        RECT 46.680 174.960 47.130 175.420 ;
        RECT 47.300 175.130 47.685 176.100 ;
        RECT 44.290 173.890 44.575 174.350 ;
        RECT 44.745 173.720 45.015 174.180 ;
        RECT 45.415 173.890 45.815 174.690 ;
        RECT 46.680 174.630 47.235 174.960 ;
        RECT 46.680 174.520 47.130 174.630 ;
        RECT 46.005 174.350 47.130 174.520 ;
        RECT 47.405 174.460 47.685 175.130 ;
        RECT 47.855 175.510 48.370 175.920 ;
        RECT 48.605 175.510 48.775 176.270 ;
        RECT 48.945 175.930 50.975 176.100 ;
        RECT 47.855 174.700 48.195 175.510 ;
        RECT 48.945 175.265 49.115 175.930 ;
        RECT 49.510 175.590 50.635 175.760 ;
        RECT 48.365 175.075 49.115 175.265 ;
        RECT 49.285 175.250 50.295 175.420 ;
        RECT 47.855 174.530 49.085 174.700 ;
        RECT 46.005 173.890 46.285 174.350 ;
        RECT 46.805 173.720 47.130 174.180 ;
        RECT 47.300 173.890 47.685 174.460 ;
        RECT 48.130 173.925 48.375 174.530 ;
        RECT 48.595 173.720 49.105 174.255 ;
        RECT 49.285 173.890 49.475 175.250 ;
        RECT 49.645 174.570 49.920 175.050 ;
        RECT 49.645 174.400 49.925 174.570 ;
        RECT 50.125 174.450 50.295 175.250 ;
        RECT 50.465 174.460 50.635 175.590 ;
        RECT 50.805 174.960 50.975 175.930 ;
        RECT 51.145 175.130 51.315 176.270 ;
        RECT 51.485 175.130 51.820 176.100 ;
        RECT 50.805 174.630 51.000 174.960 ;
        RECT 51.225 174.630 51.480 174.960 ;
        RECT 51.225 174.460 51.395 174.630 ;
        RECT 51.650 174.460 51.820 175.130 ;
        RECT 49.645 173.890 49.920 174.400 ;
        RECT 50.465 174.290 51.395 174.460 ;
        RECT 50.465 174.255 50.640 174.290 ;
        RECT 50.110 173.890 50.640 174.255 ;
        RECT 51.065 173.720 51.395 174.120 ;
        RECT 51.565 173.890 51.820 174.460 ;
        RECT 52.000 175.080 52.255 175.960 ;
        RECT 52.425 175.130 52.730 176.270 ;
        RECT 53.070 175.890 53.400 176.270 ;
        RECT 53.580 175.720 53.750 176.010 ;
        RECT 53.920 175.810 54.170 176.270 ;
        RECT 52.950 175.550 53.750 175.720 ;
        RECT 54.340 175.760 55.210 176.100 ;
        RECT 52.000 174.430 52.210 175.080 ;
        RECT 52.950 174.960 53.120 175.550 ;
        RECT 54.340 175.380 54.510 175.760 ;
        RECT 55.445 175.640 55.615 176.100 ;
        RECT 55.785 175.810 56.155 176.270 ;
        RECT 56.450 175.670 56.620 176.010 ;
        RECT 56.790 175.840 57.120 176.270 ;
        RECT 57.355 175.670 57.525 176.010 ;
        RECT 53.290 175.210 54.510 175.380 ;
        RECT 54.680 175.300 55.140 175.590 ;
        RECT 55.445 175.470 56.005 175.640 ;
        RECT 56.450 175.500 57.525 175.670 ;
        RECT 57.695 175.770 58.375 176.100 ;
        RECT 58.590 175.770 58.840 176.100 ;
        RECT 59.010 175.810 59.260 176.270 ;
        RECT 55.835 175.330 56.005 175.470 ;
        RECT 54.680 175.290 55.645 175.300 ;
        RECT 54.340 175.120 54.510 175.210 ;
        RECT 54.970 175.130 55.645 175.290 ;
        RECT 52.380 174.930 53.120 174.960 ;
        RECT 52.380 174.630 53.295 174.930 ;
        RECT 52.970 174.455 53.295 174.630 ;
        RECT 52.000 173.900 52.255 174.430 ;
        RECT 52.425 173.720 52.730 174.180 ;
        RECT 52.975 174.100 53.295 174.455 ;
        RECT 53.465 174.670 54.005 175.040 ;
        RECT 54.340 174.950 54.745 175.120 ;
        RECT 53.465 174.270 53.705 174.670 ;
        RECT 54.185 174.500 54.405 174.780 ;
        RECT 53.875 174.330 54.405 174.500 ;
        RECT 53.875 174.100 54.045 174.330 ;
        RECT 54.575 174.170 54.745 174.950 ;
        RECT 54.915 174.340 55.265 174.960 ;
        RECT 55.435 174.340 55.645 175.130 ;
        RECT 55.835 175.160 57.335 175.330 ;
        RECT 55.835 174.470 56.005 175.160 ;
        RECT 57.695 174.990 57.865 175.770 ;
        RECT 58.670 175.640 58.840 175.770 ;
        RECT 56.175 174.820 57.865 174.990 ;
        RECT 58.035 175.210 58.500 175.600 ;
        RECT 58.670 175.470 59.065 175.640 ;
        RECT 56.175 174.640 56.345 174.820 ;
        RECT 52.975 173.930 54.045 174.100 ;
        RECT 54.215 173.720 54.405 174.160 ;
        RECT 54.575 173.890 55.525 174.170 ;
        RECT 55.835 174.080 56.095 174.470 ;
        RECT 56.515 174.400 57.305 174.650 ;
        RECT 55.745 173.910 56.095 174.080 ;
        RECT 56.305 173.720 56.635 174.180 ;
        RECT 57.510 174.110 57.680 174.820 ;
        RECT 58.035 174.620 58.205 175.210 ;
        RECT 57.850 174.400 58.205 174.620 ;
        RECT 58.375 174.400 58.725 175.020 ;
        RECT 58.895 174.110 59.065 175.470 ;
        RECT 59.430 175.300 59.755 176.085 ;
        RECT 59.235 174.250 59.695 175.300 ;
        RECT 57.510 173.940 58.365 174.110 ;
        RECT 58.570 173.940 59.065 174.110 ;
        RECT 59.235 173.720 59.565 174.080 ;
        RECT 59.925 173.980 60.095 176.100 ;
        RECT 60.265 175.770 60.595 176.270 ;
        RECT 60.765 175.600 61.020 176.100 ;
        RECT 60.270 175.430 61.020 175.600 ;
        RECT 60.270 174.440 60.500 175.430 ;
        RECT 60.670 174.610 61.020 175.260 ;
        RECT 62.120 175.120 62.380 176.270 ;
        RECT 62.555 175.195 62.810 176.100 ;
        RECT 62.980 175.510 63.310 176.270 ;
        RECT 63.525 175.340 63.695 176.100 ;
        RECT 60.270 174.270 61.020 174.440 ;
        RECT 60.265 173.720 60.595 174.100 ;
        RECT 60.765 173.980 61.020 174.270 ;
        RECT 62.120 173.720 62.380 174.560 ;
        RECT 62.555 174.465 62.725 175.195 ;
        RECT 62.980 175.170 63.695 175.340 ;
        RECT 62.980 174.960 63.150 175.170 ;
        RECT 63.955 175.105 64.245 176.270 ;
        RECT 64.880 175.120 65.140 176.270 ;
        RECT 65.315 175.195 65.570 176.100 ;
        RECT 65.740 175.510 66.070 176.270 ;
        RECT 66.285 175.340 66.455 176.100 ;
        RECT 62.895 174.630 63.150 174.960 ;
        RECT 62.555 173.890 62.810 174.465 ;
        RECT 62.980 174.440 63.150 174.630 ;
        RECT 63.430 174.620 63.785 174.990 ;
        RECT 62.980 174.270 63.695 174.440 ;
        RECT 62.980 173.720 63.310 174.100 ;
        RECT 63.525 173.890 63.695 174.270 ;
        RECT 63.955 173.720 64.245 174.445 ;
        RECT 64.880 173.720 65.140 174.560 ;
        RECT 65.315 174.465 65.485 175.195 ;
        RECT 65.740 175.170 66.455 175.340 ;
        RECT 66.725 175.210 67.055 176.270 ;
        RECT 65.740 174.960 65.910 175.170 ;
        RECT 65.655 174.630 65.910 174.960 ;
        RECT 65.315 173.890 65.570 174.465 ;
        RECT 65.740 174.440 65.910 174.630 ;
        RECT 66.190 174.620 66.545 174.990 ;
        RECT 67.235 174.960 67.405 175.885 ;
        RECT 67.575 175.680 67.905 176.080 ;
        RECT 68.075 175.910 68.405 176.270 ;
        RECT 68.605 175.680 69.305 176.100 ;
        RECT 67.575 175.450 69.305 175.680 ;
        RECT 67.575 175.230 67.905 175.450 ;
        RECT 68.100 174.960 68.425 175.250 ;
        RECT 66.715 174.630 67.025 174.960 ;
        RECT 67.235 174.630 67.610 174.960 ;
        RECT 67.930 174.630 68.425 174.960 ;
        RECT 68.600 174.710 68.930 175.250 ;
        RECT 69.100 174.480 69.305 175.450 ;
        RECT 65.740 174.270 66.455 174.440 ;
        RECT 65.740 173.720 66.070 174.100 ;
        RECT 66.285 173.890 66.455 174.270 ;
        RECT 66.725 174.250 68.085 174.460 ;
        RECT 66.725 173.890 67.055 174.250 ;
        RECT 67.225 173.720 67.555 174.080 ;
        RECT 67.755 173.890 68.085 174.250 ;
        RECT 68.595 173.890 69.305 174.480 ;
        RECT 69.475 175.130 69.815 176.100 ;
        RECT 69.985 175.130 70.155 176.270 ;
        RECT 70.425 175.470 70.675 176.270 ;
        RECT 71.320 175.300 71.650 176.100 ;
        RECT 71.950 175.470 72.280 176.270 ;
        RECT 72.450 175.300 72.780 176.100 ;
        RECT 70.345 175.130 72.780 175.300 ;
        RECT 73.155 175.130 73.495 176.100 ;
        RECT 73.665 175.130 73.835 176.270 ;
        RECT 74.105 175.470 74.355 176.270 ;
        RECT 75.000 175.300 75.330 176.100 ;
        RECT 75.630 175.470 75.960 176.270 ;
        RECT 76.130 175.300 76.460 176.100 ;
        RECT 74.025 175.130 76.460 175.300 ;
        RECT 76.835 175.130 77.175 176.100 ;
        RECT 77.345 175.130 77.515 176.270 ;
        RECT 77.785 175.470 78.035 176.270 ;
        RECT 78.680 175.300 79.010 176.100 ;
        RECT 79.310 175.470 79.640 176.270 ;
        RECT 79.810 175.300 80.140 176.100 ;
        RECT 77.705 175.130 80.140 175.300 ;
        RECT 80.515 175.180 82.185 176.270 ;
        RECT 82.360 175.835 87.705 176.270 ;
        RECT 69.475 174.520 69.650 175.130 ;
        RECT 70.345 174.880 70.515 175.130 ;
        RECT 69.820 174.710 70.515 174.880 ;
        RECT 70.690 174.710 71.110 174.910 ;
        RECT 71.280 174.710 71.610 174.910 ;
        RECT 71.780 174.710 72.110 174.910 ;
        RECT 69.475 173.890 69.815 174.520 ;
        RECT 69.985 173.720 70.235 174.520 ;
        RECT 70.425 174.370 71.650 174.540 ;
        RECT 70.425 173.890 70.755 174.370 ;
        RECT 70.925 173.720 71.150 174.180 ;
        RECT 71.320 173.890 71.650 174.370 ;
        RECT 72.280 174.500 72.450 175.130 ;
        RECT 72.635 174.710 72.985 174.960 ;
        RECT 73.155 174.520 73.330 175.130 ;
        RECT 74.025 174.880 74.195 175.130 ;
        RECT 73.500 174.710 74.195 174.880 ;
        RECT 74.370 174.710 74.790 174.910 ;
        RECT 74.960 174.710 75.290 174.910 ;
        RECT 75.460 174.710 75.790 174.910 ;
        RECT 72.280 173.890 72.780 174.500 ;
        RECT 73.155 173.890 73.495 174.520 ;
        RECT 73.665 173.720 73.915 174.520 ;
        RECT 74.105 174.370 75.330 174.540 ;
        RECT 74.105 173.890 74.435 174.370 ;
        RECT 74.605 173.720 74.830 174.180 ;
        RECT 75.000 173.890 75.330 174.370 ;
        RECT 75.960 174.500 76.130 175.130 ;
        RECT 76.315 174.710 76.665 174.960 ;
        RECT 76.835 174.520 77.010 175.130 ;
        RECT 77.705 174.880 77.875 175.130 ;
        RECT 77.180 174.710 77.875 174.880 ;
        RECT 78.050 174.710 78.470 174.910 ;
        RECT 78.640 174.710 78.970 174.910 ;
        RECT 79.140 174.710 79.470 174.910 ;
        RECT 75.960 173.890 76.460 174.500 ;
        RECT 76.835 173.890 77.175 174.520 ;
        RECT 77.345 173.720 77.595 174.520 ;
        RECT 77.785 174.370 79.010 174.540 ;
        RECT 77.785 173.890 78.115 174.370 ;
        RECT 78.285 173.720 78.510 174.180 ;
        RECT 78.680 173.890 79.010 174.370 ;
        RECT 79.640 174.500 79.810 175.130 ;
        RECT 79.995 174.710 80.345 174.960 ;
        RECT 80.515 174.660 81.265 175.180 ;
        RECT 79.640 173.890 80.140 174.500 ;
        RECT 81.435 174.490 82.185 175.010 ;
        RECT 83.950 174.585 84.300 175.835 ;
        RECT 87.915 175.130 88.145 176.270 ;
        RECT 88.315 175.120 88.645 176.100 ;
        RECT 88.815 175.130 89.025 176.270 ;
        RECT 80.515 173.720 82.185 174.490 ;
        RECT 85.780 174.265 86.120 175.095 ;
        RECT 87.895 174.710 88.225 174.960 ;
        RECT 82.360 173.720 87.705 174.265 ;
        RECT 87.915 173.720 88.145 174.540 ;
        RECT 88.395 174.520 88.645 175.120 ;
        RECT 89.715 175.105 90.005 176.270 ;
        RECT 90.750 175.640 91.035 176.100 ;
        RECT 91.205 175.810 91.475 176.270 ;
        RECT 90.750 175.420 91.705 175.640 ;
        RECT 90.635 174.690 91.325 175.250 ;
        RECT 88.315 173.890 88.645 174.520 ;
        RECT 88.815 173.720 89.025 174.540 ;
        RECT 91.495 174.520 91.705 175.420 ;
        RECT 89.715 173.720 90.005 174.445 ;
        RECT 90.750 174.350 91.705 174.520 ;
        RECT 91.875 175.250 92.275 176.100 ;
        RECT 92.465 175.640 92.745 176.100 ;
        RECT 93.265 175.810 93.590 176.270 ;
        RECT 92.465 175.420 93.590 175.640 ;
        RECT 91.875 174.690 92.970 175.250 ;
        RECT 93.140 174.960 93.590 175.420 ;
        RECT 93.760 175.130 94.145 176.100 ;
        RECT 90.750 173.890 91.035 174.350 ;
        RECT 91.205 173.720 91.475 174.180 ;
        RECT 91.875 173.890 92.275 174.690 ;
        RECT 93.140 174.630 93.695 174.960 ;
        RECT 93.140 174.520 93.590 174.630 ;
        RECT 92.465 174.350 93.590 174.520 ;
        RECT 93.865 174.460 94.145 175.130 ;
        RECT 94.315 175.180 95.525 176.270 ;
        RECT 94.315 174.640 94.835 175.180 ;
        RECT 95.735 175.130 95.965 176.270 ;
        RECT 96.135 175.120 96.465 176.100 ;
        RECT 96.635 175.130 96.845 176.270 ;
        RECT 97.280 175.300 97.610 176.100 ;
        RECT 97.780 175.470 98.110 176.270 ;
        RECT 98.410 175.300 98.740 176.100 ;
        RECT 99.385 175.470 99.635 176.270 ;
        RECT 97.280 175.130 99.715 175.300 ;
        RECT 99.905 175.130 100.075 176.270 ;
        RECT 100.245 175.130 100.585 176.100 ;
        RECT 100.870 175.640 101.155 176.100 ;
        RECT 101.325 175.810 101.595 176.270 ;
        RECT 100.870 175.420 101.825 175.640 ;
        RECT 95.005 174.470 95.525 175.010 ;
        RECT 95.715 174.710 96.045 174.960 ;
        RECT 92.465 173.890 92.745 174.350 ;
        RECT 93.265 173.720 93.590 174.180 ;
        RECT 93.760 173.890 94.145 174.460 ;
        RECT 94.315 173.720 95.525 174.470 ;
        RECT 95.735 173.720 95.965 174.540 ;
        RECT 96.215 174.520 96.465 175.120 ;
        RECT 97.075 174.710 97.425 174.960 ;
        RECT 96.135 173.890 96.465 174.520 ;
        RECT 96.635 173.720 96.845 174.540 ;
        RECT 97.610 174.500 97.780 175.130 ;
        RECT 97.950 174.710 98.280 174.910 ;
        RECT 98.450 174.710 98.780 174.910 ;
        RECT 98.950 174.710 99.370 174.910 ;
        RECT 99.545 174.880 99.715 175.130 ;
        RECT 99.545 174.710 100.240 174.880 ;
        RECT 97.280 173.890 97.780 174.500 ;
        RECT 98.410 174.370 99.635 174.540 ;
        RECT 100.410 174.520 100.585 175.130 ;
        RECT 100.755 174.690 101.445 175.250 ;
        RECT 101.615 174.520 101.825 175.420 ;
        RECT 98.410 173.890 98.740 174.370 ;
        RECT 98.910 173.720 99.135 174.180 ;
        RECT 99.305 173.890 99.635 174.370 ;
        RECT 99.825 173.720 100.075 174.520 ;
        RECT 100.245 173.890 100.585 174.520 ;
        RECT 100.870 174.350 101.825 174.520 ;
        RECT 101.995 175.250 102.395 176.100 ;
        RECT 102.585 175.640 102.865 176.100 ;
        RECT 103.385 175.810 103.710 176.270 ;
        RECT 102.585 175.420 103.710 175.640 ;
        RECT 101.995 174.690 103.090 175.250 ;
        RECT 103.260 174.960 103.710 175.420 ;
        RECT 103.880 175.130 104.265 176.100 ;
        RECT 100.870 173.890 101.155 174.350 ;
        RECT 101.325 173.720 101.595 174.180 ;
        RECT 101.995 173.890 102.395 174.690 ;
        RECT 103.260 174.630 103.815 174.960 ;
        RECT 103.260 174.520 103.710 174.630 ;
        RECT 102.585 174.350 103.710 174.520 ;
        RECT 103.985 174.460 104.265 175.130 ;
        RECT 102.585 173.890 102.865 174.350 ;
        RECT 103.385 173.720 103.710 174.180 ;
        RECT 103.880 173.890 104.265 174.460 ;
        RECT 104.440 175.080 104.695 175.960 ;
        RECT 104.865 175.130 105.170 176.270 ;
        RECT 105.510 175.890 105.840 176.270 ;
        RECT 106.020 175.720 106.190 176.010 ;
        RECT 106.360 175.810 106.610 176.270 ;
        RECT 105.390 175.550 106.190 175.720 ;
        RECT 106.780 175.760 107.650 176.100 ;
        RECT 104.440 174.430 104.650 175.080 ;
        RECT 105.390 174.960 105.560 175.550 ;
        RECT 106.780 175.380 106.950 175.760 ;
        RECT 107.885 175.640 108.055 176.100 ;
        RECT 108.225 175.810 108.595 176.270 ;
        RECT 108.890 175.670 109.060 176.010 ;
        RECT 109.230 175.840 109.560 176.270 ;
        RECT 109.795 175.670 109.965 176.010 ;
        RECT 105.730 175.210 106.950 175.380 ;
        RECT 107.120 175.300 107.580 175.590 ;
        RECT 107.885 175.470 108.445 175.640 ;
        RECT 108.890 175.500 109.965 175.670 ;
        RECT 110.135 175.770 110.815 176.100 ;
        RECT 111.030 175.770 111.280 176.100 ;
        RECT 111.450 175.810 111.700 176.270 ;
        RECT 108.275 175.330 108.445 175.470 ;
        RECT 107.120 175.290 108.085 175.300 ;
        RECT 106.780 175.120 106.950 175.210 ;
        RECT 107.410 175.130 108.085 175.290 ;
        RECT 104.820 174.930 105.560 174.960 ;
        RECT 104.820 174.630 105.735 174.930 ;
        RECT 105.410 174.455 105.735 174.630 ;
        RECT 104.440 173.900 104.695 174.430 ;
        RECT 104.865 173.720 105.170 174.180 ;
        RECT 105.415 174.100 105.735 174.455 ;
        RECT 105.905 174.670 106.445 175.040 ;
        RECT 106.780 174.950 107.185 175.120 ;
        RECT 105.905 174.270 106.145 174.670 ;
        RECT 106.625 174.500 106.845 174.780 ;
        RECT 106.315 174.330 106.845 174.500 ;
        RECT 106.315 174.100 106.485 174.330 ;
        RECT 107.015 174.170 107.185 174.950 ;
        RECT 107.355 174.340 107.705 174.960 ;
        RECT 107.875 174.340 108.085 175.130 ;
        RECT 108.275 175.160 109.775 175.330 ;
        RECT 108.275 174.470 108.445 175.160 ;
        RECT 110.135 174.990 110.305 175.770 ;
        RECT 111.110 175.640 111.280 175.770 ;
        RECT 108.615 174.820 110.305 174.990 ;
        RECT 110.475 175.210 110.940 175.600 ;
        RECT 111.110 175.470 111.505 175.640 ;
        RECT 108.615 174.640 108.785 174.820 ;
        RECT 105.415 173.930 106.485 174.100 ;
        RECT 106.655 173.720 106.845 174.160 ;
        RECT 107.015 173.890 107.965 174.170 ;
        RECT 108.275 174.080 108.535 174.470 ;
        RECT 108.955 174.400 109.745 174.650 ;
        RECT 108.185 173.910 108.535 174.080 ;
        RECT 108.745 173.720 109.075 174.180 ;
        RECT 109.950 174.110 110.120 174.820 ;
        RECT 110.475 174.620 110.645 175.210 ;
        RECT 110.290 174.400 110.645 174.620 ;
        RECT 110.815 174.400 111.165 175.020 ;
        RECT 111.335 174.110 111.505 175.470 ;
        RECT 111.870 175.300 112.195 176.085 ;
        RECT 111.675 174.250 112.135 175.300 ;
        RECT 109.950 173.940 110.805 174.110 ;
        RECT 111.010 173.940 111.505 174.110 ;
        RECT 111.675 173.720 112.005 174.080 ;
        RECT 112.365 173.980 112.535 176.100 ;
        RECT 112.705 175.770 113.035 176.270 ;
        RECT 113.205 175.600 113.460 176.100 ;
        RECT 112.710 175.430 113.460 175.600 ;
        RECT 112.710 174.440 112.940 175.430 ;
        RECT 113.110 174.610 113.460 175.260 ;
        RECT 114.555 175.180 115.765 176.270 ;
        RECT 114.555 174.640 115.075 175.180 ;
        RECT 115.245 174.470 115.765 175.010 ;
        RECT 112.710 174.270 113.460 174.440 ;
        RECT 112.705 173.720 113.035 174.100 ;
        RECT 113.205 173.980 113.460 174.270 ;
        RECT 114.555 173.720 115.765 174.470 ;
        RECT 14.650 173.550 115.850 173.720 ;
        RECT 14.735 172.800 15.945 173.550 ;
        RECT 14.735 172.260 15.255 172.800 ;
        RECT 16.575 172.780 20.085 173.550 ;
        RECT 15.425 172.090 15.945 172.630 ;
        RECT 14.735 171.000 15.945 172.090 ;
        RECT 16.575 172.090 18.265 172.610 ;
        RECT 18.435 172.260 20.085 172.780 ;
        RECT 20.255 172.810 20.640 173.380 ;
        RECT 20.810 173.090 21.135 173.550 ;
        RECT 21.655 172.920 21.935 173.380 ;
        RECT 20.255 172.140 20.535 172.810 ;
        RECT 20.810 172.750 21.935 172.920 ;
        RECT 20.810 172.640 21.260 172.750 ;
        RECT 20.705 172.310 21.260 172.640 ;
        RECT 22.125 172.580 22.525 173.380 ;
        RECT 22.925 173.090 23.195 173.550 ;
        RECT 23.365 172.920 23.650 173.380 ;
        RECT 16.575 171.000 20.085 172.090 ;
        RECT 20.255 171.170 20.640 172.140 ;
        RECT 20.810 171.850 21.260 172.310 ;
        RECT 21.430 172.020 22.525 172.580 ;
        RECT 20.810 171.630 21.935 171.850 ;
        RECT 20.810 171.000 21.135 171.460 ;
        RECT 21.655 171.170 21.935 171.630 ;
        RECT 22.125 171.170 22.525 172.020 ;
        RECT 22.695 172.750 23.650 172.920 ;
        RECT 23.935 172.800 25.145 173.550 ;
        RECT 25.315 172.825 25.605 173.550 ;
        RECT 22.695 171.850 22.905 172.750 ;
        RECT 23.075 172.020 23.765 172.580 ;
        RECT 23.935 172.090 24.455 172.630 ;
        RECT 24.625 172.260 25.145 172.800 ;
        RECT 25.835 172.730 26.045 173.550 ;
        RECT 26.215 172.750 26.545 173.380 ;
        RECT 22.695 171.630 23.650 171.850 ;
        RECT 22.925 171.000 23.195 171.460 ;
        RECT 23.365 171.170 23.650 171.630 ;
        RECT 23.935 171.000 25.145 172.090 ;
        RECT 25.315 171.000 25.605 172.165 ;
        RECT 26.215 172.150 26.465 172.750 ;
        RECT 26.715 172.730 26.945 173.550 ;
        RECT 27.360 172.770 27.860 173.380 ;
        RECT 26.635 172.310 26.965 172.560 ;
        RECT 27.155 172.310 27.505 172.560 ;
        RECT 25.835 171.000 26.045 172.140 ;
        RECT 26.215 171.170 26.545 172.150 ;
        RECT 27.690 172.140 27.860 172.770 ;
        RECT 28.490 172.900 28.820 173.380 ;
        RECT 28.990 173.090 29.215 173.550 ;
        RECT 29.385 172.900 29.715 173.380 ;
        RECT 28.490 172.730 29.715 172.900 ;
        RECT 29.905 172.750 30.155 173.550 ;
        RECT 30.325 172.750 30.665 173.380 ;
        RECT 31.040 172.770 31.540 173.380 ;
        RECT 28.030 172.360 28.360 172.560 ;
        RECT 28.530 172.360 28.860 172.560 ;
        RECT 29.030 172.360 29.450 172.560 ;
        RECT 29.625 172.390 30.320 172.560 ;
        RECT 29.625 172.140 29.795 172.390 ;
        RECT 30.490 172.140 30.665 172.750 ;
        RECT 30.835 172.310 31.185 172.560 ;
        RECT 31.370 172.140 31.540 172.770 ;
        RECT 32.170 172.900 32.500 173.380 ;
        RECT 32.670 173.090 32.895 173.550 ;
        RECT 33.065 172.900 33.395 173.380 ;
        RECT 32.170 172.730 33.395 172.900 ;
        RECT 33.585 172.750 33.835 173.550 ;
        RECT 34.005 172.750 34.345 173.380 ;
        RECT 34.720 172.770 35.220 173.380 ;
        RECT 31.710 172.360 32.040 172.560 ;
        RECT 32.210 172.360 32.540 172.560 ;
        RECT 32.710 172.360 33.130 172.560 ;
        RECT 33.305 172.390 34.000 172.560 ;
        RECT 33.305 172.140 33.475 172.390 ;
        RECT 34.170 172.140 34.345 172.750 ;
        RECT 34.515 172.310 34.865 172.560 ;
        RECT 35.050 172.140 35.220 172.770 ;
        RECT 35.850 172.900 36.180 173.380 ;
        RECT 36.350 173.090 36.575 173.550 ;
        RECT 36.745 172.900 37.075 173.380 ;
        RECT 35.850 172.730 37.075 172.900 ;
        RECT 37.265 172.750 37.515 173.550 ;
        RECT 37.685 172.750 38.025 173.380 ;
        RECT 38.310 172.920 38.595 173.380 ;
        RECT 38.765 173.090 39.035 173.550 ;
        RECT 38.310 172.750 39.265 172.920 ;
        RECT 35.390 172.360 35.720 172.560 ;
        RECT 35.890 172.360 36.220 172.560 ;
        RECT 36.390 172.360 36.810 172.560 ;
        RECT 36.985 172.390 37.680 172.560 ;
        RECT 36.985 172.140 37.155 172.390 ;
        RECT 37.850 172.140 38.025 172.750 ;
        RECT 26.715 171.000 26.945 172.140 ;
        RECT 27.360 171.970 29.795 172.140 ;
        RECT 27.360 171.170 27.690 171.970 ;
        RECT 27.860 171.000 28.190 171.800 ;
        RECT 28.490 171.170 28.820 171.970 ;
        RECT 29.465 171.000 29.715 171.800 ;
        RECT 29.985 171.000 30.155 172.140 ;
        RECT 30.325 171.170 30.665 172.140 ;
        RECT 31.040 171.970 33.475 172.140 ;
        RECT 31.040 171.170 31.370 171.970 ;
        RECT 31.540 171.000 31.870 171.800 ;
        RECT 32.170 171.170 32.500 171.970 ;
        RECT 33.145 171.000 33.395 171.800 ;
        RECT 33.665 171.000 33.835 172.140 ;
        RECT 34.005 171.170 34.345 172.140 ;
        RECT 34.720 171.970 37.155 172.140 ;
        RECT 34.720 171.170 35.050 171.970 ;
        RECT 35.220 171.000 35.550 171.800 ;
        RECT 35.850 171.170 36.180 171.970 ;
        RECT 36.825 171.000 37.075 171.800 ;
        RECT 37.345 171.000 37.515 172.140 ;
        RECT 37.685 171.170 38.025 172.140 ;
        RECT 38.195 172.020 38.885 172.580 ;
        RECT 39.055 171.850 39.265 172.750 ;
        RECT 38.310 171.630 39.265 171.850 ;
        RECT 39.435 172.580 39.835 173.380 ;
        RECT 40.025 172.920 40.305 173.380 ;
        RECT 40.825 173.090 41.150 173.550 ;
        RECT 40.025 172.750 41.150 172.920 ;
        RECT 41.320 172.810 41.705 173.380 ;
        RECT 40.700 172.640 41.150 172.750 ;
        RECT 39.435 172.020 40.530 172.580 ;
        RECT 40.700 172.310 41.255 172.640 ;
        RECT 38.310 171.170 38.595 171.630 ;
        RECT 38.765 171.000 39.035 171.460 ;
        RECT 39.435 171.170 39.835 172.020 ;
        RECT 40.700 171.850 41.150 172.310 ;
        RECT 41.425 172.140 41.705 172.810 ;
        RECT 41.875 172.780 43.545 173.550 ;
        RECT 40.025 171.630 41.150 171.850 ;
        RECT 40.025 171.170 40.305 171.630 ;
        RECT 40.825 171.000 41.150 171.460 ;
        RECT 41.320 171.170 41.705 172.140 ;
        RECT 41.875 172.090 42.625 172.610 ;
        RECT 42.795 172.260 43.545 172.780 ;
        RECT 43.715 172.750 44.055 173.380 ;
        RECT 44.225 172.750 44.475 173.550 ;
        RECT 44.665 172.900 44.995 173.380 ;
        RECT 45.165 173.090 45.390 173.550 ;
        RECT 45.560 172.900 45.890 173.380 ;
        RECT 43.715 172.140 43.890 172.750 ;
        RECT 44.665 172.730 45.890 172.900 ;
        RECT 46.520 172.770 47.020 173.380 ;
        RECT 44.060 172.390 44.755 172.560 ;
        RECT 44.585 172.140 44.755 172.390 ;
        RECT 44.930 172.360 45.350 172.560 ;
        RECT 45.520 172.360 45.850 172.560 ;
        RECT 46.020 172.360 46.350 172.560 ;
        RECT 46.520 172.140 46.690 172.770 ;
        RECT 47.395 172.750 47.735 173.380 ;
        RECT 47.905 172.750 48.155 173.550 ;
        RECT 48.345 172.900 48.675 173.380 ;
        RECT 48.845 173.090 49.070 173.550 ;
        RECT 49.240 172.900 49.570 173.380 ;
        RECT 46.875 172.310 47.225 172.560 ;
        RECT 47.395 172.140 47.570 172.750 ;
        RECT 48.345 172.730 49.570 172.900 ;
        RECT 50.200 172.770 50.700 173.380 ;
        RECT 51.075 172.825 51.365 173.550 ;
        RECT 51.535 172.780 55.045 173.550 ;
        RECT 47.740 172.390 48.435 172.560 ;
        RECT 48.265 172.140 48.435 172.390 ;
        RECT 48.610 172.360 49.030 172.560 ;
        RECT 49.200 172.360 49.530 172.560 ;
        RECT 49.700 172.360 50.030 172.560 ;
        RECT 50.200 172.140 50.370 172.770 ;
        RECT 50.555 172.310 50.905 172.560 ;
        RECT 41.875 171.000 43.545 172.090 ;
        RECT 43.715 171.170 44.055 172.140 ;
        RECT 44.225 171.000 44.395 172.140 ;
        RECT 44.585 171.970 47.020 172.140 ;
        RECT 44.665 171.000 44.915 171.800 ;
        RECT 45.560 171.170 45.890 171.970 ;
        RECT 46.190 171.000 46.520 171.800 ;
        RECT 46.690 171.170 47.020 171.970 ;
        RECT 47.395 171.170 47.735 172.140 ;
        RECT 47.905 171.000 48.075 172.140 ;
        RECT 48.265 171.970 50.700 172.140 ;
        RECT 48.345 171.000 48.595 171.800 ;
        RECT 49.240 171.170 49.570 171.970 ;
        RECT 49.870 171.000 50.200 171.800 ;
        RECT 50.370 171.170 50.700 171.970 ;
        RECT 51.075 171.000 51.365 172.165 ;
        RECT 51.535 172.090 53.225 172.610 ;
        RECT 53.395 172.260 55.045 172.780 ;
        RECT 55.275 172.730 55.485 173.550 ;
        RECT 55.655 172.750 55.985 173.380 ;
        RECT 55.655 172.150 55.905 172.750 ;
        RECT 56.155 172.730 56.385 173.550 ;
        RECT 57.145 173.000 57.315 173.380 ;
        RECT 57.495 173.170 57.825 173.550 ;
        RECT 57.145 172.830 57.810 173.000 ;
        RECT 58.005 172.875 58.265 173.380 ;
        RECT 56.075 172.310 56.405 172.560 ;
        RECT 57.075 172.280 57.405 172.650 ;
        RECT 57.640 172.575 57.810 172.830 ;
        RECT 57.640 172.245 57.925 172.575 ;
        RECT 51.535 171.000 55.045 172.090 ;
        RECT 55.275 171.000 55.485 172.140 ;
        RECT 55.655 171.170 55.985 172.150 ;
        RECT 56.155 171.000 56.385 172.140 ;
        RECT 57.640 172.100 57.810 172.245 ;
        RECT 57.145 171.930 57.810 172.100 ;
        RECT 58.095 172.075 58.265 172.875 ;
        RECT 58.895 172.780 62.405 173.550 ;
        RECT 57.145 171.170 57.315 171.930 ;
        RECT 57.495 171.000 57.825 171.760 ;
        RECT 57.995 171.170 58.265 172.075 ;
        RECT 58.895 172.090 60.585 172.610 ;
        RECT 60.755 172.260 62.405 172.780 ;
        RECT 62.580 172.710 62.840 173.550 ;
        RECT 63.015 172.805 63.270 173.380 ;
        RECT 63.440 173.170 63.770 173.550 ;
        RECT 63.985 173.000 64.155 173.380 ;
        RECT 63.440 172.830 64.155 173.000 ;
        RECT 64.505 173.000 64.675 173.380 ;
        RECT 64.890 173.170 65.220 173.550 ;
        RECT 64.505 172.830 65.220 173.000 ;
        RECT 58.895 171.000 62.405 172.090 ;
        RECT 62.580 171.000 62.840 172.150 ;
        RECT 63.015 172.075 63.185 172.805 ;
        RECT 63.440 172.640 63.610 172.830 ;
        RECT 63.355 172.310 63.610 172.640 ;
        RECT 63.440 172.100 63.610 172.310 ;
        RECT 63.890 172.280 64.245 172.650 ;
        RECT 64.415 172.280 64.770 172.650 ;
        RECT 65.050 172.640 65.220 172.830 ;
        RECT 65.390 172.805 65.645 173.380 ;
        RECT 65.050 172.310 65.305 172.640 ;
        RECT 65.050 172.100 65.220 172.310 ;
        RECT 63.015 171.170 63.270 172.075 ;
        RECT 63.440 171.930 64.155 172.100 ;
        RECT 63.440 171.000 63.770 171.760 ;
        RECT 63.985 171.170 64.155 171.930 ;
        RECT 64.505 171.930 65.220 172.100 ;
        RECT 65.475 172.075 65.645 172.805 ;
        RECT 65.820 172.710 66.080 173.550 ;
        RECT 66.255 172.800 67.465 173.550 ;
        RECT 64.505 171.170 64.675 171.930 ;
        RECT 64.890 171.000 65.220 171.760 ;
        RECT 65.390 171.170 65.645 172.075 ;
        RECT 65.820 171.000 66.080 172.150 ;
        RECT 66.255 172.090 66.775 172.630 ;
        RECT 66.945 172.260 67.465 172.800 ;
        RECT 67.635 172.780 71.145 173.550 ;
        RECT 71.320 173.005 76.665 173.550 ;
        RECT 67.635 172.090 69.325 172.610 ;
        RECT 69.495 172.260 71.145 172.780 ;
        RECT 66.255 171.000 67.465 172.090 ;
        RECT 67.635 171.000 71.145 172.090 ;
        RECT 72.910 171.435 73.260 172.685 ;
        RECT 74.740 172.175 75.080 173.005 ;
        RECT 76.835 172.825 77.125 173.550 ;
        RECT 77.670 172.840 77.925 173.370 ;
        RECT 78.105 173.090 78.390 173.550 ;
        RECT 71.320 171.000 76.665 171.435 ;
        RECT 76.835 171.000 77.125 172.165 ;
        RECT 77.670 171.980 77.850 172.840 ;
        RECT 78.570 172.640 78.820 173.290 ;
        RECT 78.020 172.310 78.820 172.640 ;
        RECT 77.670 171.850 77.925 171.980 ;
        RECT 77.585 171.680 77.925 171.850 ;
        RECT 77.670 171.310 77.925 171.680 ;
        RECT 78.105 171.000 78.390 171.800 ;
        RECT 78.570 171.720 78.820 172.310 ;
        RECT 79.020 172.955 79.340 173.285 ;
        RECT 79.520 173.070 80.180 173.550 ;
        RECT 80.380 173.160 81.230 173.330 ;
        RECT 79.020 172.060 79.210 172.955 ;
        RECT 79.530 172.630 80.190 172.900 ;
        RECT 79.860 172.570 80.190 172.630 ;
        RECT 79.380 172.400 79.710 172.460 ;
        RECT 80.380 172.400 80.550 173.160 ;
        RECT 81.790 173.090 82.110 173.550 ;
        RECT 82.310 172.910 82.560 173.340 ;
        RECT 82.850 173.110 83.260 173.550 ;
        RECT 83.430 173.170 84.445 173.370 ;
        RECT 80.720 172.740 81.970 172.910 ;
        RECT 80.720 172.620 81.050 172.740 ;
        RECT 79.380 172.230 81.280 172.400 ;
        RECT 79.020 171.890 80.940 172.060 ;
        RECT 79.020 171.870 79.340 171.890 ;
        RECT 78.570 171.210 78.900 171.720 ;
        RECT 79.170 171.260 79.340 171.870 ;
        RECT 81.110 171.720 81.280 172.230 ;
        RECT 81.450 172.160 81.630 172.570 ;
        RECT 81.800 171.980 81.970 172.740 ;
        RECT 79.510 171.000 79.840 171.690 ;
        RECT 80.070 171.550 81.280 171.720 ;
        RECT 81.450 171.670 81.970 171.980 ;
        RECT 82.140 172.570 82.560 172.910 ;
        RECT 82.850 172.570 83.260 172.900 ;
        RECT 82.140 171.800 82.330 172.570 ;
        RECT 83.430 172.440 83.600 173.170 ;
        RECT 84.745 173.000 84.915 173.330 ;
        RECT 85.085 173.170 85.415 173.550 ;
        RECT 83.770 172.620 84.120 172.990 ;
        RECT 83.430 172.400 83.850 172.440 ;
        RECT 82.500 172.230 83.850 172.400 ;
        RECT 82.500 172.070 82.750 172.230 ;
        RECT 83.260 171.800 83.510 172.060 ;
        RECT 82.140 171.550 83.510 171.800 ;
        RECT 80.070 171.260 80.310 171.550 ;
        RECT 81.110 171.470 81.280 171.550 ;
        RECT 80.510 171.000 80.930 171.380 ;
        RECT 81.110 171.220 81.740 171.470 ;
        RECT 82.210 171.000 82.540 171.380 ;
        RECT 82.710 171.260 82.880 171.550 ;
        RECT 83.680 171.385 83.850 172.230 ;
        RECT 84.300 172.060 84.520 172.930 ;
        RECT 84.745 172.810 85.440 173.000 ;
        RECT 84.020 171.680 84.520 172.060 ;
        RECT 84.690 172.010 85.100 172.630 ;
        RECT 85.270 171.840 85.440 172.810 ;
        RECT 84.745 171.670 85.440 171.840 ;
        RECT 83.060 171.000 83.440 171.380 ;
        RECT 83.680 171.215 84.510 171.385 ;
        RECT 84.745 171.170 84.915 171.670 ;
        RECT 85.085 171.000 85.415 171.500 ;
        RECT 85.630 171.170 85.855 173.290 ;
        RECT 86.025 173.170 86.355 173.550 ;
        RECT 86.525 173.000 86.695 173.290 ;
        RECT 86.030 172.830 86.695 173.000 ;
        RECT 86.960 173.000 87.215 173.290 ;
        RECT 87.385 173.170 87.715 173.550 ;
        RECT 86.960 172.830 87.710 173.000 ;
        RECT 86.030 171.840 86.260 172.830 ;
        RECT 86.430 172.010 86.780 172.660 ;
        RECT 86.960 172.010 87.310 172.660 ;
        RECT 87.480 171.840 87.710 172.830 ;
        RECT 86.030 171.670 86.695 171.840 ;
        RECT 86.025 171.000 86.355 171.500 ;
        RECT 86.525 171.170 86.695 171.670 ;
        RECT 86.960 171.670 87.710 171.840 ;
        RECT 86.960 171.170 87.215 171.670 ;
        RECT 87.385 171.000 87.715 171.500 ;
        RECT 87.885 171.170 88.055 173.290 ;
        RECT 88.415 173.190 88.745 173.550 ;
        RECT 88.915 173.160 89.410 173.330 ;
        RECT 89.615 173.160 90.470 173.330 ;
        RECT 88.285 171.970 88.745 173.020 ;
        RECT 88.225 171.185 88.550 171.970 ;
        RECT 88.915 171.800 89.085 173.160 ;
        RECT 89.255 172.250 89.605 172.870 ;
        RECT 89.775 172.650 90.130 172.870 ;
        RECT 89.775 172.060 89.945 172.650 ;
        RECT 90.300 172.450 90.470 173.160 ;
        RECT 91.345 173.090 91.675 173.550 ;
        RECT 91.885 173.190 92.235 173.360 ;
        RECT 90.675 172.620 91.465 172.870 ;
        RECT 91.885 172.800 92.145 173.190 ;
        RECT 92.455 173.100 93.405 173.380 ;
        RECT 93.575 173.110 93.765 173.550 ;
        RECT 93.935 173.170 95.005 173.340 ;
        RECT 91.635 172.450 91.805 172.630 ;
        RECT 88.915 171.630 89.310 171.800 ;
        RECT 89.480 171.670 89.945 172.060 ;
        RECT 90.115 172.280 91.805 172.450 ;
        RECT 89.140 171.500 89.310 171.630 ;
        RECT 90.115 171.500 90.285 172.280 ;
        RECT 91.975 172.110 92.145 172.800 ;
        RECT 90.645 171.940 92.145 172.110 ;
        RECT 92.335 172.140 92.545 172.930 ;
        RECT 92.715 172.310 93.065 172.930 ;
        RECT 93.235 172.320 93.405 173.100 ;
        RECT 93.935 172.940 94.105 173.170 ;
        RECT 93.575 172.770 94.105 172.940 ;
        RECT 93.575 172.490 93.795 172.770 ;
        RECT 94.275 172.600 94.515 173.000 ;
        RECT 93.235 172.150 93.640 172.320 ;
        RECT 93.975 172.230 94.515 172.600 ;
        RECT 94.685 172.815 95.005 173.170 ;
        RECT 95.250 173.090 95.555 173.550 ;
        RECT 95.725 172.840 95.980 173.370 ;
        RECT 94.685 172.640 95.010 172.815 ;
        RECT 94.685 172.340 95.600 172.640 ;
        RECT 94.860 172.310 95.600 172.340 ;
        RECT 92.335 171.980 93.010 172.140 ;
        RECT 93.470 172.060 93.640 172.150 ;
        RECT 92.335 171.970 93.300 171.980 ;
        RECT 91.975 171.800 92.145 171.940 ;
        RECT 88.720 171.000 88.970 171.460 ;
        RECT 89.140 171.170 89.390 171.500 ;
        RECT 89.605 171.170 90.285 171.500 ;
        RECT 90.455 171.600 91.530 171.770 ;
        RECT 91.975 171.630 92.535 171.800 ;
        RECT 92.840 171.680 93.300 171.970 ;
        RECT 93.470 171.890 94.690 172.060 ;
        RECT 90.455 171.260 90.625 171.600 ;
        RECT 90.860 171.000 91.190 171.430 ;
        RECT 91.360 171.260 91.530 171.600 ;
        RECT 91.825 171.000 92.195 171.460 ;
        RECT 92.365 171.170 92.535 171.630 ;
        RECT 93.470 171.510 93.640 171.890 ;
        RECT 94.860 171.720 95.030 172.310 ;
        RECT 95.770 172.190 95.980 172.840 ;
        RECT 97.115 172.730 97.345 173.550 ;
        RECT 97.515 172.750 97.845 173.380 ;
        RECT 97.095 172.310 97.425 172.560 ;
        RECT 92.770 171.170 93.640 171.510 ;
        RECT 94.230 171.550 95.030 171.720 ;
        RECT 93.810 171.000 94.060 171.460 ;
        RECT 94.230 171.260 94.400 171.550 ;
        RECT 94.580 171.000 94.910 171.380 ;
        RECT 95.250 171.000 95.555 172.140 ;
        RECT 95.725 171.310 95.980 172.190 ;
        RECT 97.595 172.150 97.845 172.750 ;
        RECT 98.015 172.730 98.225 173.550 ;
        RECT 98.730 172.740 98.975 173.345 ;
        RECT 99.195 173.015 99.705 173.550 ;
        RECT 97.115 171.000 97.345 172.140 ;
        RECT 97.515 171.170 97.845 172.150 ;
        RECT 98.455 172.570 99.685 172.740 ;
        RECT 98.015 171.000 98.225 172.140 ;
        RECT 98.455 171.760 98.795 172.570 ;
        RECT 98.965 172.005 99.715 172.195 ;
        RECT 98.455 171.350 98.970 171.760 ;
        RECT 99.205 171.000 99.375 171.760 ;
        RECT 99.545 171.340 99.715 172.005 ;
        RECT 99.885 172.020 100.075 173.380 ;
        RECT 100.245 172.870 100.520 173.380 ;
        RECT 100.710 173.015 101.240 173.380 ;
        RECT 101.665 173.150 101.995 173.550 ;
        RECT 101.065 172.980 101.240 173.015 ;
        RECT 100.245 172.700 100.525 172.870 ;
        RECT 100.245 172.220 100.520 172.700 ;
        RECT 100.725 172.020 100.895 172.820 ;
        RECT 99.885 171.850 100.895 172.020 ;
        RECT 101.065 172.810 101.995 172.980 ;
        RECT 102.165 172.810 102.420 173.380 ;
        RECT 102.595 172.825 102.885 173.550 ;
        RECT 101.065 171.680 101.235 172.810 ;
        RECT 101.825 172.640 101.995 172.810 ;
        RECT 100.110 171.510 101.235 171.680 ;
        RECT 101.405 172.310 101.600 172.640 ;
        RECT 101.825 172.310 102.080 172.640 ;
        RECT 101.405 171.340 101.575 172.310 ;
        RECT 102.250 172.140 102.420 172.810 ;
        RECT 103.095 172.730 103.325 173.550 ;
        RECT 103.495 172.750 103.825 173.380 ;
        RECT 103.075 172.310 103.405 172.560 ;
        RECT 99.545 171.170 101.575 171.340 ;
        RECT 101.745 171.000 101.915 172.140 ;
        RECT 102.085 171.170 102.420 172.140 ;
        RECT 102.595 171.000 102.885 172.165 ;
        RECT 103.575 172.150 103.825 172.750 ;
        RECT 103.995 172.730 104.205 173.550 ;
        RECT 104.440 172.840 104.695 173.370 ;
        RECT 104.865 173.090 105.170 173.550 ;
        RECT 105.415 173.170 106.485 173.340 ;
        RECT 103.095 171.000 103.325 172.140 ;
        RECT 103.495 171.170 103.825 172.150 ;
        RECT 104.440 172.190 104.650 172.840 ;
        RECT 105.415 172.815 105.735 173.170 ;
        RECT 105.410 172.640 105.735 172.815 ;
        RECT 104.820 172.340 105.735 172.640 ;
        RECT 105.905 172.600 106.145 173.000 ;
        RECT 106.315 172.940 106.485 173.170 ;
        RECT 106.655 173.110 106.845 173.550 ;
        RECT 107.015 173.100 107.965 173.380 ;
        RECT 108.185 173.190 108.535 173.360 ;
        RECT 106.315 172.770 106.845 172.940 ;
        RECT 104.820 172.310 105.560 172.340 ;
        RECT 103.995 171.000 104.205 172.140 ;
        RECT 104.440 171.310 104.695 172.190 ;
        RECT 104.865 171.000 105.170 172.140 ;
        RECT 105.390 171.720 105.560 172.310 ;
        RECT 105.905 172.230 106.445 172.600 ;
        RECT 106.625 172.490 106.845 172.770 ;
        RECT 107.015 172.320 107.185 173.100 ;
        RECT 106.780 172.150 107.185 172.320 ;
        RECT 107.355 172.310 107.705 172.930 ;
        RECT 106.780 172.060 106.950 172.150 ;
        RECT 107.875 172.140 108.085 172.930 ;
        RECT 105.730 171.890 106.950 172.060 ;
        RECT 107.410 171.980 108.085 172.140 ;
        RECT 105.390 171.550 106.190 171.720 ;
        RECT 105.510 171.000 105.840 171.380 ;
        RECT 106.020 171.260 106.190 171.550 ;
        RECT 106.780 171.510 106.950 171.890 ;
        RECT 107.120 171.970 108.085 171.980 ;
        RECT 108.275 172.800 108.535 173.190 ;
        RECT 108.745 173.090 109.075 173.550 ;
        RECT 109.950 173.160 110.805 173.330 ;
        RECT 111.010 173.160 111.505 173.330 ;
        RECT 111.675 173.190 112.005 173.550 ;
        RECT 108.275 172.110 108.445 172.800 ;
        RECT 108.615 172.450 108.785 172.630 ;
        RECT 108.955 172.620 109.745 172.870 ;
        RECT 109.950 172.450 110.120 173.160 ;
        RECT 110.290 172.650 110.645 172.870 ;
        RECT 108.615 172.280 110.305 172.450 ;
        RECT 107.120 171.680 107.580 171.970 ;
        RECT 108.275 171.940 109.775 172.110 ;
        RECT 108.275 171.800 108.445 171.940 ;
        RECT 107.885 171.630 108.445 171.800 ;
        RECT 106.360 171.000 106.610 171.460 ;
        RECT 106.780 171.170 107.650 171.510 ;
        RECT 107.885 171.170 108.055 171.630 ;
        RECT 108.890 171.600 109.965 171.770 ;
        RECT 108.225 171.000 108.595 171.460 ;
        RECT 108.890 171.260 109.060 171.600 ;
        RECT 109.230 171.000 109.560 171.430 ;
        RECT 109.795 171.260 109.965 171.600 ;
        RECT 110.135 171.500 110.305 172.280 ;
        RECT 110.475 172.060 110.645 172.650 ;
        RECT 110.815 172.250 111.165 172.870 ;
        RECT 110.475 171.670 110.940 172.060 ;
        RECT 111.335 171.800 111.505 173.160 ;
        RECT 111.675 171.970 112.135 173.020 ;
        RECT 111.110 171.630 111.505 171.800 ;
        RECT 111.110 171.500 111.280 171.630 ;
        RECT 110.135 171.170 110.815 171.500 ;
        RECT 111.030 171.170 111.280 171.500 ;
        RECT 111.450 171.000 111.700 171.460 ;
        RECT 111.870 171.185 112.195 171.970 ;
        RECT 112.365 171.170 112.535 173.290 ;
        RECT 112.705 173.170 113.035 173.550 ;
        RECT 113.205 173.000 113.460 173.290 ;
        RECT 112.710 172.830 113.460 173.000 ;
        RECT 112.710 171.840 112.940 172.830 ;
        RECT 114.555 172.800 115.765 173.550 ;
        RECT 113.110 172.010 113.460 172.660 ;
        RECT 114.555 172.090 115.075 172.630 ;
        RECT 115.245 172.260 115.765 172.800 ;
        RECT 112.710 171.670 113.460 171.840 ;
        RECT 112.705 171.000 113.035 171.500 ;
        RECT 113.205 171.170 113.460 171.670 ;
        RECT 114.555 171.000 115.765 172.090 ;
        RECT 14.650 170.830 115.850 171.000 ;
        RECT 14.735 169.740 15.945 170.830 ;
        RECT 14.735 169.030 15.255 169.570 ;
        RECT 15.425 169.200 15.945 169.740 ;
        RECT 16.635 169.690 16.845 170.830 ;
        RECT 17.015 169.680 17.345 170.660 ;
        RECT 17.515 169.690 17.745 170.830 ;
        RECT 17.955 169.755 18.225 170.660 ;
        RECT 18.395 170.070 18.725 170.830 ;
        RECT 18.905 169.900 19.075 170.660 ;
        RECT 19.450 170.200 19.735 170.660 ;
        RECT 19.905 170.370 20.175 170.830 ;
        RECT 19.450 169.980 20.405 170.200 ;
        RECT 14.735 168.280 15.945 169.030 ;
        RECT 16.635 168.280 16.845 169.100 ;
        RECT 17.015 169.080 17.265 169.680 ;
        RECT 17.435 169.270 17.765 169.520 ;
        RECT 17.015 168.450 17.345 169.080 ;
        RECT 17.515 168.280 17.745 169.100 ;
        RECT 17.955 168.955 18.125 169.755 ;
        RECT 18.410 169.730 19.075 169.900 ;
        RECT 18.410 169.585 18.580 169.730 ;
        RECT 18.295 169.255 18.580 169.585 ;
        RECT 18.410 169.000 18.580 169.255 ;
        RECT 18.815 169.180 19.145 169.550 ;
        RECT 19.335 169.250 20.025 169.810 ;
        RECT 20.195 169.080 20.405 169.980 ;
        RECT 17.955 168.450 18.215 168.955 ;
        RECT 18.410 168.830 19.075 169.000 ;
        RECT 18.395 168.280 18.725 168.660 ;
        RECT 18.905 168.450 19.075 168.830 ;
        RECT 19.450 168.910 20.405 169.080 ;
        RECT 20.575 169.810 20.975 170.660 ;
        RECT 21.165 170.200 21.445 170.660 ;
        RECT 21.965 170.370 22.290 170.830 ;
        RECT 21.165 169.980 22.290 170.200 ;
        RECT 20.575 169.250 21.670 169.810 ;
        RECT 21.840 169.520 22.290 169.980 ;
        RECT 22.460 169.690 22.845 170.660 ;
        RECT 19.450 168.450 19.735 168.910 ;
        RECT 19.905 168.280 20.175 168.740 ;
        RECT 20.575 168.450 20.975 169.250 ;
        RECT 21.840 169.190 22.395 169.520 ;
        RECT 21.840 169.080 22.290 169.190 ;
        RECT 21.165 168.910 22.290 169.080 ;
        RECT 22.565 169.020 22.845 169.690 ;
        RECT 21.165 168.450 21.445 168.910 ;
        RECT 21.965 168.280 22.290 168.740 ;
        RECT 22.460 168.450 22.845 169.020 ;
        RECT 23.020 169.640 23.275 170.520 ;
        RECT 23.445 169.690 23.750 170.830 ;
        RECT 24.090 170.450 24.420 170.830 ;
        RECT 24.600 170.280 24.770 170.570 ;
        RECT 24.940 170.370 25.190 170.830 ;
        RECT 23.970 170.110 24.770 170.280 ;
        RECT 25.360 170.320 26.230 170.660 ;
        RECT 23.020 168.990 23.230 169.640 ;
        RECT 23.970 169.520 24.140 170.110 ;
        RECT 25.360 169.940 25.530 170.320 ;
        RECT 26.465 170.200 26.635 170.660 ;
        RECT 26.805 170.370 27.175 170.830 ;
        RECT 27.470 170.230 27.640 170.570 ;
        RECT 27.810 170.400 28.140 170.830 ;
        RECT 28.375 170.230 28.545 170.570 ;
        RECT 24.310 169.770 25.530 169.940 ;
        RECT 25.700 169.860 26.160 170.150 ;
        RECT 26.465 170.030 27.025 170.200 ;
        RECT 27.470 170.060 28.545 170.230 ;
        RECT 28.715 170.330 29.395 170.660 ;
        RECT 29.610 170.330 29.860 170.660 ;
        RECT 30.030 170.370 30.280 170.830 ;
        RECT 26.855 169.890 27.025 170.030 ;
        RECT 25.700 169.850 26.665 169.860 ;
        RECT 25.360 169.680 25.530 169.770 ;
        RECT 25.990 169.690 26.665 169.850 ;
        RECT 23.400 169.490 24.140 169.520 ;
        RECT 23.400 169.190 24.315 169.490 ;
        RECT 23.990 169.015 24.315 169.190 ;
        RECT 23.020 168.460 23.275 168.990 ;
        RECT 23.445 168.280 23.750 168.740 ;
        RECT 23.995 168.660 24.315 169.015 ;
        RECT 24.485 169.230 25.025 169.600 ;
        RECT 25.360 169.510 25.765 169.680 ;
        RECT 24.485 168.830 24.725 169.230 ;
        RECT 25.205 169.060 25.425 169.340 ;
        RECT 24.895 168.890 25.425 169.060 ;
        RECT 24.895 168.660 25.065 168.890 ;
        RECT 25.595 168.730 25.765 169.510 ;
        RECT 25.935 168.900 26.285 169.520 ;
        RECT 26.455 168.900 26.665 169.690 ;
        RECT 26.855 169.720 28.355 169.890 ;
        RECT 26.855 169.030 27.025 169.720 ;
        RECT 28.715 169.550 28.885 170.330 ;
        RECT 29.690 170.200 29.860 170.330 ;
        RECT 27.195 169.380 28.885 169.550 ;
        RECT 29.055 169.770 29.520 170.160 ;
        RECT 29.690 170.030 30.085 170.200 ;
        RECT 27.195 169.200 27.365 169.380 ;
        RECT 23.995 168.490 25.065 168.660 ;
        RECT 25.235 168.280 25.425 168.720 ;
        RECT 25.595 168.450 26.545 168.730 ;
        RECT 26.855 168.640 27.115 169.030 ;
        RECT 27.535 168.960 28.325 169.210 ;
        RECT 26.765 168.470 27.115 168.640 ;
        RECT 27.325 168.280 27.655 168.740 ;
        RECT 28.530 168.670 28.700 169.380 ;
        RECT 29.055 169.180 29.225 169.770 ;
        RECT 28.870 168.960 29.225 169.180 ;
        RECT 29.395 168.960 29.745 169.580 ;
        RECT 29.915 168.670 30.085 170.030 ;
        RECT 30.450 169.860 30.775 170.645 ;
        RECT 30.255 168.810 30.715 169.860 ;
        RECT 28.530 168.500 29.385 168.670 ;
        RECT 29.590 168.500 30.085 168.670 ;
        RECT 30.255 168.280 30.585 168.640 ;
        RECT 30.945 168.540 31.115 170.660 ;
        RECT 31.285 170.330 31.615 170.830 ;
        RECT 31.785 170.160 32.040 170.660 ;
        RECT 31.290 169.990 32.040 170.160 ;
        RECT 31.290 169.000 31.520 169.990 ;
        RECT 31.690 169.170 32.040 169.820 ;
        RECT 33.175 169.690 33.405 170.830 ;
        RECT 33.575 169.680 33.905 170.660 ;
        RECT 34.075 169.690 34.285 170.830 ;
        RECT 34.630 170.200 34.915 170.660 ;
        RECT 35.085 170.370 35.355 170.830 ;
        RECT 34.630 169.980 35.585 170.200 ;
        RECT 33.155 169.270 33.485 169.520 ;
        RECT 31.290 168.830 32.040 169.000 ;
        RECT 31.285 168.280 31.615 168.660 ;
        RECT 31.785 168.540 32.040 168.830 ;
        RECT 33.175 168.280 33.405 169.100 ;
        RECT 33.655 169.080 33.905 169.680 ;
        RECT 34.515 169.250 35.205 169.810 ;
        RECT 33.575 168.450 33.905 169.080 ;
        RECT 34.075 168.280 34.285 169.100 ;
        RECT 35.375 169.080 35.585 169.980 ;
        RECT 34.630 168.910 35.585 169.080 ;
        RECT 35.755 169.810 36.155 170.660 ;
        RECT 36.345 170.200 36.625 170.660 ;
        RECT 37.145 170.370 37.470 170.830 ;
        RECT 36.345 169.980 37.470 170.200 ;
        RECT 35.755 169.250 36.850 169.810 ;
        RECT 37.020 169.520 37.470 169.980 ;
        RECT 37.640 169.690 38.025 170.660 ;
        RECT 34.630 168.450 34.915 168.910 ;
        RECT 35.085 168.280 35.355 168.740 ;
        RECT 35.755 168.450 36.155 169.250 ;
        RECT 37.020 169.190 37.575 169.520 ;
        RECT 37.020 169.080 37.470 169.190 ;
        RECT 36.345 168.910 37.470 169.080 ;
        RECT 37.745 169.020 38.025 169.690 ;
        RECT 38.195 169.665 38.485 170.830 ;
        RECT 39.115 169.740 41.705 170.830 ;
        RECT 39.115 169.220 40.325 169.740 ;
        RECT 41.880 169.640 42.135 170.520 ;
        RECT 42.305 169.690 42.610 170.830 ;
        RECT 42.950 170.450 43.280 170.830 ;
        RECT 43.460 170.280 43.630 170.570 ;
        RECT 43.800 170.370 44.050 170.830 ;
        RECT 42.830 170.110 43.630 170.280 ;
        RECT 44.220 170.320 45.090 170.660 ;
        RECT 40.495 169.050 41.705 169.570 ;
        RECT 36.345 168.450 36.625 168.910 ;
        RECT 37.145 168.280 37.470 168.740 ;
        RECT 37.640 168.450 38.025 169.020 ;
        RECT 38.195 168.280 38.485 169.005 ;
        RECT 39.115 168.280 41.705 169.050 ;
        RECT 41.880 168.990 42.090 169.640 ;
        RECT 42.830 169.520 43.000 170.110 ;
        RECT 44.220 169.940 44.390 170.320 ;
        RECT 45.325 170.200 45.495 170.660 ;
        RECT 45.665 170.370 46.035 170.830 ;
        RECT 46.330 170.230 46.500 170.570 ;
        RECT 46.670 170.400 47.000 170.830 ;
        RECT 47.235 170.230 47.405 170.570 ;
        RECT 43.170 169.770 44.390 169.940 ;
        RECT 44.560 169.860 45.020 170.150 ;
        RECT 45.325 170.030 45.885 170.200 ;
        RECT 46.330 170.060 47.405 170.230 ;
        RECT 47.575 170.330 48.255 170.660 ;
        RECT 48.470 170.330 48.720 170.660 ;
        RECT 48.890 170.370 49.140 170.830 ;
        RECT 45.715 169.890 45.885 170.030 ;
        RECT 44.560 169.850 45.525 169.860 ;
        RECT 44.220 169.680 44.390 169.770 ;
        RECT 44.850 169.690 45.525 169.850 ;
        RECT 42.260 169.490 43.000 169.520 ;
        RECT 42.260 169.190 43.175 169.490 ;
        RECT 42.850 169.015 43.175 169.190 ;
        RECT 41.880 168.460 42.135 168.990 ;
        RECT 42.305 168.280 42.610 168.740 ;
        RECT 42.855 168.660 43.175 169.015 ;
        RECT 43.345 169.230 43.885 169.600 ;
        RECT 44.220 169.510 44.625 169.680 ;
        RECT 43.345 168.830 43.585 169.230 ;
        RECT 44.065 169.060 44.285 169.340 ;
        RECT 43.755 168.890 44.285 169.060 ;
        RECT 43.755 168.660 43.925 168.890 ;
        RECT 44.455 168.730 44.625 169.510 ;
        RECT 44.795 168.900 45.145 169.520 ;
        RECT 45.315 168.900 45.525 169.690 ;
        RECT 45.715 169.720 47.215 169.890 ;
        RECT 45.715 169.030 45.885 169.720 ;
        RECT 47.575 169.550 47.745 170.330 ;
        RECT 48.550 170.200 48.720 170.330 ;
        RECT 46.055 169.380 47.745 169.550 ;
        RECT 47.915 169.770 48.380 170.160 ;
        RECT 48.550 170.030 48.945 170.200 ;
        RECT 46.055 169.200 46.225 169.380 ;
        RECT 42.855 168.490 43.925 168.660 ;
        RECT 44.095 168.280 44.285 168.720 ;
        RECT 44.455 168.450 45.405 168.730 ;
        RECT 45.715 168.640 45.975 169.030 ;
        RECT 46.395 168.960 47.185 169.210 ;
        RECT 45.625 168.470 45.975 168.640 ;
        RECT 46.185 168.280 46.515 168.740 ;
        RECT 47.390 168.670 47.560 169.380 ;
        RECT 47.915 169.180 48.085 169.770 ;
        RECT 47.730 168.960 48.085 169.180 ;
        RECT 48.255 168.960 48.605 169.580 ;
        RECT 48.775 168.670 48.945 170.030 ;
        RECT 49.310 169.860 49.635 170.645 ;
        RECT 49.115 168.810 49.575 169.860 ;
        RECT 47.390 168.500 48.245 168.670 ;
        RECT 48.450 168.500 48.945 168.670 ;
        RECT 49.115 168.280 49.445 168.640 ;
        RECT 49.805 168.540 49.975 170.660 ;
        RECT 50.145 170.330 50.475 170.830 ;
        RECT 50.645 170.160 50.900 170.660 ;
        RECT 50.150 169.990 50.900 170.160 ;
        RECT 50.150 169.000 50.380 169.990 ;
        RECT 50.550 169.170 50.900 169.820 ;
        RECT 51.135 169.690 51.345 170.830 ;
        RECT 51.515 169.680 51.845 170.660 ;
        RECT 52.015 169.690 52.245 170.830 ;
        RECT 52.495 169.690 52.725 170.830 ;
        RECT 52.895 169.680 53.225 170.660 ;
        RECT 53.395 169.690 53.605 170.830 ;
        RECT 53.985 169.680 54.315 170.830 ;
        RECT 54.485 169.810 54.655 170.660 ;
        RECT 54.825 170.030 55.155 170.830 ;
        RECT 55.325 169.810 55.495 170.660 ;
        RECT 55.675 170.030 55.915 170.830 ;
        RECT 56.085 169.850 56.415 170.660 ;
        RECT 50.150 168.830 50.900 169.000 ;
        RECT 50.145 168.280 50.475 168.660 ;
        RECT 50.645 168.540 50.900 168.830 ;
        RECT 51.135 168.280 51.345 169.100 ;
        RECT 51.515 169.080 51.765 169.680 ;
        RECT 51.935 169.270 52.265 169.520 ;
        RECT 52.475 169.270 52.805 169.520 ;
        RECT 51.515 168.450 51.845 169.080 ;
        RECT 52.015 168.280 52.245 169.100 ;
        RECT 52.495 168.280 52.725 169.100 ;
        RECT 52.975 169.080 53.225 169.680 ;
        RECT 54.485 169.640 55.495 169.810 ;
        RECT 55.700 169.680 56.415 169.850 ;
        RECT 56.595 169.740 58.265 170.830 ;
        RECT 58.440 170.395 63.785 170.830 ;
        RECT 54.485 169.470 54.980 169.640 ;
        RECT 54.485 169.300 54.985 169.470 ;
        RECT 55.700 169.440 55.870 169.680 ;
        RECT 54.485 169.100 54.980 169.300 ;
        RECT 55.370 169.270 55.870 169.440 ;
        RECT 56.040 169.270 56.420 169.510 ;
        RECT 55.700 169.100 55.870 169.270 ;
        RECT 56.595 169.220 57.345 169.740 ;
        RECT 52.895 168.450 53.225 169.080 ;
        RECT 53.395 168.280 53.605 169.100 ;
        RECT 53.985 168.280 54.315 169.080 ;
        RECT 54.485 168.930 55.495 169.100 ;
        RECT 55.700 168.930 56.335 169.100 ;
        RECT 57.515 169.050 58.265 169.570 ;
        RECT 60.030 169.145 60.380 170.395 ;
        RECT 63.955 169.665 64.245 170.830 ;
        RECT 64.420 169.680 64.680 170.830 ;
        RECT 64.855 169.755 65.110 170.660 ;
        RECT 65.280 170.070 65.610 170.830 ;
        RECT 65.825 169.900 65.995 170.660 ;
        RECT 54.485 168.450 54.655 168.930 ;
        RECT 54.825 168.280 55.155 168.760 ;
        RECT 55.325 168.450 55.495 168.930 ;
        RECT 55.745 168.280 55.985 168.760 ;
        RECT 56.165 168.450 56.335 168.930 ;
        RECT 56.595 168.280 58.265 169.050 ;
        RECT 61.860 168.825 62.200 169.655 ;
        RECT 58.440 168.280 63.785 168.825 ;
        RECT 63.955 168.280 64.245 169.005 ;
        RECT 64.420 168.280 64.680 169.120 ;
        RECT 64.855 169.025 65.025 169.755 ;
        RECT 65.280 169.730 65.995 169.900 ;
        RECT 66.255 169.860 66.565 170.660 ;
        RECT 66.735 170.030 67.045 170.830 ;
        RECT 67.215 170.200 67.475 170.660 ;
        RECT 67.645 170.370 67.900 170.830 ;
        RECT 68.075 170.200 68.335 170.660 ;
        RECT 67.215 170.030 68.335 170.200 ;
        RECT 65.280 169.520 65.450 169.730 ;
        RECT 66.255 169.690 67.285 169.860 ;
        RECT 65.195 169.190 65.450 169.520 ;
        RECT 64.855 168.450 65.110 169.025 ;
        RECT 65.280 169.000 65.450 169.190 ;
        RECT 65.730 169.180 66.085 169.550 ;
        RECT 65.280 168.830 65.995 169.000 ;
        RECT 65.280 168.280 65.610 168.660 ;
        RECT 65.825 168.450 65.995 168.830 ;
        RECT 66.255 168.780 66.425 169.690 ;
        RECT 66.595 168.950 66.945 169.520 ;
        RECT 67.115 169.440 67.285 169.690 ;
        RECT 68.075 169.780 68.335 170.030 ;
        RECT 68.505 169.960 68.790 170.830 ;
        RECT 68.075 169.610 68.830 169.780 ;
        RECT 67.115 169.270 68.255 169.440 ;
        RECT 68.425 169.100 68.830 169.610 ;
        RECT 69.475 169.740 72.065 170.830 ;
        RECT 72.610 169.850 72.865 170.520 ;
        RECT 73.045 170.030 73.330 170.830 ;
        RECT 73.510 170.110 73.840 170.620 ;
        RECT 69.475 169.220 70.685 169.740 ;
        RECT 67.180 168.930 68.830 169.100 ;
        RECT 70.855 169.050 72.065 169.570 ;
        RECT 72.610 169.130 72.790 169.850 ;
        RECT 73.510 169.520 73.760 170.110 ;
        RECT 74.110 169.960 74.280 170.570 ;
        RECT 74.450 170.140 74.780 170.830 ;
        RECT 75.010 170.280 75.250 170.570 ;
        RECT 75.450 170.450 75.870 170.830 ;
        RECT 76.050 170.360 76.680 170.610 ;
        RECT 77.150 170.450 77.480 170.830 ;
        RECT 76.050 170.280 76.220 170.360 ;
        RECT 77.650 170.280 77.820 170.570 ;
        RECT 78.000 170.450 78.380 170.830 ;
        RECT 78.620 170.445 79.450 170.615 ;
        RECT 75.010 170.110 76.220 170.280 ;
        RECT 72.960 169.190 73.760 169.520 ;
        RECT 66.255 168.450 66.555 168.780 ;
        RECT 66.725 168.280 67.000 168.760 ;
        RECT 67.180 168.540 67.475 168.930 ;
        RECT 67.645 168.280 67.900 168.760 ;
        RECT 68.075 168.540 68.335 168.930 ;
        RECT 68.505 168.280 68.785 168.760 ;
        RECT 69.475 168.280 72.065 169.050 ;
        RECT 72.525 168.990 72.790 169.130 ;
        RECT 72.525 168.960 72.865 168.990 ;
        RECT 72.610 168.460 72.865 168.960 ;
        RECT 73.045 168.280 73.330 168.740 ;
        RECT 73.510 168.540 73.760 169.190 ;
        RECT 73.960 169.940 74.280 169.960 ;
        RECT 73.960 169.770 75.880 169.940 ;
        RECT 73.960 168.875 74.150 169.770 ;
        RECT 76.050 169.600 76.220 170.110 ;
        RECT 76.390 169.850 76.910 170.160 ;
        RECT 74.320 169.430 76.220 169.600 ;
        RECT 74.320 169.370 74.650 169.430 ;
        RECT 74.800 169.200 75.130 169.260 ;
        RECT 74.470 168.930 75.130 169.200 ;
        RECT 73.960 168.545 74.280 168.875 ;
        RECT 74.460 168.280 75.120 168.760 ;
        RECT 75.320 168.670 75.490 169.430 ;
        RECT 76.390 169.260 76.570 169.670 ;
        RECT 75.660 169.090 75.990 169.210 ;
        RECT 76.740 169.090 76.910 169.850 ;
        RECT 75.660 168.920 76.910 169.090 ;
        RECT 77.080 170.030 78.450 170.280 ;
        RECT 77.080 169.260 77.270 170.030 ;
        RECT 78.200 169.770 78.450 170.030 ;
        RECT 77.440 169.600 77.690 169.760 ;
        RECT 78.620 169.600 78.790 170.445 ;
        RECT 79.685 170.160 79.855 170.660 ;
        RECT 80.025 170.330 80.355 170.830 ;
        RECT 78.960 169.770 79.460 170.150 ;
        RECT 79.685 169.990 80.380 170.160 ;
        RECT 77.440 169.430 78.790 169.600 ;
        RECT 78.370 169.390 78.790 169.430 ;
        RECT 77.080 168.920 77.500 169.260 ;
        RECT 77.790 168.930 78.200 169.260 ;
        RECT 75.320 168.500 76.170 168.670 ;
        RECT 76.730 168.280 77.050 168.740 ;
        RECT 77.250 168.490 77.500 168.920 ;
        RECT 77.790 168.280 78.200 168.720 ;
        RECT 78.370 168.660 78.540 169.390 ;
        RECT 78.710 168.840 79.060 169.210 ;
        RECT 79.240 168.900 79.460 169.770 ;
        RECT 79.630 169.200 80.040 169.820 ;
        RECT 80.210 169.020 80.380 169.990 ;
        RECT 79.685 168.830 80.380 169.020 ;
        RECT 78.370 168.460 79.385 168.660 ;
        RECT 79.685 168.500 79.855 168.830 ;
        RECT 80.025 168.280 80.355 168.660 ;
        RECT 80.570 168.540 80.795 170.660 ;
        RECT 80.965 170.330 81.295 170.830 ;
        RECT 81.465 170.160 81.635 170.660 ;
        RECT 80.970 169.990 81.635 170.160 ;
        RECT 80.970 169.000 81.200 169.990 ;
        RECT 81.985 169.900 82.155 170.660 ;
        RECT 82.335 170.070 82.665 170.830 ;
        RECT 81.370 169.170 81.720 169.820 ;
        RECT 81.985 169.730 82.650 169.900 ;
        RECT 82.835 169.755 83.105 170.660 ;
        RECT 83.525 170.100 83.820 170.830 ;
        RECT 83.990 169.930 84.250 170.655 ;
        RECT 84.420 170.100 84.680 170.830 ;
        RECT 84.850 169.930 85.110 170.655 ;
        RECT 85.280 170.100 85.540 170.830 ;
        RECT 85.710 169.930 85.970 170.655 ;
        RECT 86.140 170.100 86.400 170.830 ;
        RECT 86.570 169.930 86.830 170.655 ;
        RECT 82.480 169.585 82.650 169.730 ;
        RECT 81.915 169.180 82.245 169.550 ;
        RECT 82.480 169.255 82.765 169.585 ;
        RECT 82.480 169.000 82.650 169.255 ;
        RECT 80.970 168.830 81.635 169.000 ;
        RECT 80.965 168.280 81.295 168.660 ;
        RECT 81.465 168.540 81.635 168.830 ;
        RECT 81.985 168.830 82.650 169.000 ;
        RECT 82.935 168.955 83.105 169.755 ;
        RECT 81.985 168.450 82.155 168.830 ;
        RECT 82.335 168.280 82.665 168.660 ;
        RECT 82.845 168.450 83.105 168.955 ;
        RECT 83.520 169.690 86.830 169.930 ;
        RECT 87.000 169.720 87.260 170.830 ;
        RECT 83.520 169.100 84.490 169.690 ;
        RECT 87.430 169.520 87.680 170.655 ;
        RECT 87.860 169.720 88.155 170.830 ;
        RECT 88.335 169.755 88.605 170.660 ;
        RECT 88.775 170.070 89.105 170.830 ;
        RECT 89.285 169.900 89.455 170.660 ;
        RECT 84.660 169.270 87.680 169.520 ;
        RECT 83.520 168.930 86.830 169.100 ;
        RECT 83.520 168.280 83.820 168.760 ;
        RECT 83.990 168.475 84.250 168.930 ;
        RECT 84.420 168.280 84.680 168.760 ;
        RECT 84.850 168.475 85.110 168.930 ;
        RECT 85.280 168.280 85.540 168.760 ;
        RECT 85.710 168.475 85.970 168.930 ;
        RECT 86.140 168.280 86.400 168.760 ;
        RECT 86.570 168.475 86.830 168.930 ;
        RECT 87.000 168.280 87.260 168.805 ;
        RECT 87.430 168.460 87.680 169.270 ;
        RECT 87.850 168.910 88.165 169.520 ;
        RECT 88.335 168.955 88.505 169.755 ;
        RECT 88.790 169.730 89.455 169.900 ;
        RECT 88.790 169.585 88.960 169.730 ;
        RECT 89.715 169.665 90.005 170.830 ;
        RECT 90.180 169.690 90.515 170.660 ;
        RECT 90.685 169.690 90.855 170.830 ;
        RECT 91.025 170.490 93.055 170.660 ;
        RECT 88.675 169.255 88.960 169.585 ;
        RECT 88.790 169.000 88.960 169.255 ;
        RECT 89.195 169.180 89.525 169.550 ;
        RECT 90.180 169.020 90.350 169.690 ;
        RECT 91.025 169.520 91.195 170.490 ;
        RECT 90.520 169.190 90.775 169.520 ;
        RECT 91.000 169.190 91.195 169.520 ;
        RECT 91.365 170.150 92.490 170.320 ;
        RECT 90.605 169.020 90.775 169.190 ;
        RECT 91.365 169.020 91.535 170.150 ;
        RECT 87.860 168.280 88.105 168.740 ;
        RECT 88.335 168.450 88.595 168.955 ;
        RECT 88.790 168.830 89.455 169.000 ;
        RECT 88.775 168.280 89.105 168.660 ;
        RECT 89.285 168.450 89.455 168.830 ;
        RECT 89.715 168.280 90.005 169.005 ;
        RECT 90.180 168.450 90.435 169.020 ;
        RECT 90.605 168.850 91.535 169.020 ;
        RECT 91.705 169.810 92.715 169.980 ;
        RECT 91.705 169.010 91.875 169.810 ;
        RECT 92.080 169.130 92.355 169.610 ;
        RECT 92.075 168.960 92.355 169.130 ;
        RECT 91.360 168.815 91.535 168.850 ;
        RECT 90.605 168.280 90.935 168.680 ;
        RECT 91.360 168.450 91.890 168.815 ;
        RECT 92.080 168.450 92.355 168.960 ;
        RECT 92.525 168.450 92.715 169.810 ;
        RECT 92.885 169.825 93.055 170.490 ;
        RECT 93.225 170.070 93.395 170.830 ;
        RECT 93.630 170.070 94.145 170.480 ;
        RECT 92.885 169.635 93.635 169.825 ;
        RECT 93.805 169.260 94.145 170.070 ;
        RECT 92.915 169.090 94.145 169.260 ;
        RECT 94.320 169.690 94.655 170.660 ;
        RECT 94.825 169.690 94.995 170.830 ;
        RECT 95.165 170.490 97.195 170.660 ;
        RECT 92.895 168.280 93.405 168.815 ;
        RECT 93.625 168.485 93.870 169.090 ;
        RECT 94.320 169.020 94.490 169.690 ;
        RECT 95.165 169.520 95.335 170.490 ;
        RECT 94.660 169.190 94.915 169.520 ;
        RECT 95.140 169.190 95.335 169.520 ;
        RECT 95.505 170.150 96.630 170.320 ;
        RECT 94.745 169.020 94.915 169.190 ;
        RECT 95.505 169.020 95.675 170.150 ;
        RECT 94.320 168.450 94.575 169.020 ;
        RECT 94.745 168.850 95.675 169.020 ;
        RECT 95.845 169.810 96.855 169.980 ;
        RECT 95.845 169.010 96.015 169.810 ;
        RECT 96.220 169.130 96.495 169.610 ;
        RECT 96.215 168.960 96.495 169.130 ;
        RECT 95.500 168.815 95.675 168.850 ;
        RECT 94.745 168.280 95.075 168.680 ;
        RECT 95.500 168.450 96.030 168.815 ;
        RECT 96.220 168.450 96.495 168.960 ;
        RECT 96.665 168.450 96.855 169.810 ;
        RECT 97.025 169.825 97.195 170.490 ;
        RECT 97.365 170.070 97.535 170.830 ;
        RECT 97.770 170.070 98.285 170.480 ;
        RECT 97.025 169.635 97.775 169.825 ;
        RECT 97.945 169.260 98.285 170.070 ;
        RECT 97.055 169.090 98.285 169.260 ;
        RECT 98.455 170.070 98.970 170.480 ;
        RECT 99.205 170.070 99.375 170.830 ;
        RECT 99.545 170.490 101.575 170.660 ;
        RECT 98.455 169.260 98.795 170.070 ;
        RECT 99.545 169.825 99.715 170.490 ;
        RECT 100.110 170.150 101.235 170.320 ;
        RECT 98.965 169.635 99.715 169.825 ;
        RECT 99.885 169.810 100.895 169.980 ;
        RECT 98.455 169.090 99.685 169.260 ;
        RECT 97.035 168.280 97.545 168.815 ;
        RECT 97.765 168.485 98.010 169.090 ;
        RECT 98.730 168.485 98.975 169.090 ;
        RECT 99.195 168.280 99.705 168.815 ;
        RECT 99.885 168.450 100.075 169.810 ;
        RECT 100.245 169.130 100.520 169.610 ;
        RECT 100.245 168.960 100.525 169.130 ;
        RECT 100.725 169.010 100.895 169.810 ;
        RECT 101.065 169.020 101.235 170.150 ;
        RECT 101.405 169.520 101.575 170.490 ;
        RECT 101.745 169.690 101.915 170.830 ;
        RECT 102.085 169.690 102.420 170.660 ;
        RECT 101.405 169.190 101.600 169.520 ;
        RECT 101.825 169.190 102.080 169.520 ;
        RECT 101.825 169.020 101.995 169.190 ;
        RECT 102.250 169.020 102.420 169.690 ;
        RECT 103.515 170.070 104.030 170.480 ;
        RECT 104.265 170.070 104.435 170.830 ;
        RECT 104.605 170.490 106.635 170.660 ;
        RECT 103.515 169.260 103.855 170.070 ;
        RECT 104.605 169.825 104.775 170.490 ;
        RECT 105.170 170.150 106.295 170.320 ;
        RECT 104.025 169.635 104.775 169.825 ;
        RECT 104.945 169.810 105.955 169.980 ;
        RECT 103.515 169.090 104.745 169.260 ;
        RECT 100.245 168.450 100.520 168.960 ;
        RECT 101.065 168.850 101.995 169.020 ;
        RECT 101.065 168.815 101.240 168.850 ;
        RECT 100.710 168.450 101.240 168.815 ;
        RECT 101.665 168.280 101.995 168.680 ;
        RECT 102.165 168.450 102.420 169.020 ;
        RECT 103.790 168.485 104.035 169.090 ;
        RECT 104.255 168.280 104.765 168.815 ;
        RECT 104.945 168.450 105.135 169.810 ;
        RECT 105.305 169.470 105.580 169.610 ;
        RECT 105.305 169.300 105.585 169.470 ;
        RECT 105.305 168.450 105.580 169.300 ;
        RECT 105.785 169.010 105.955 169.810 ;
        RECT 106.125 169.020 106.295 170.150 ;
        RECT 106.465 169.520 106.635 170.490 ;
        RECT 106.805 169.690 106.975 170.830 ;
        RECT 107.145 169.690 107.480 170.660 ;
        RECT 107.770 170.200 108.055 170.660 ;
        RECT 108.225 170.370 108.495 170.830 ;
        RECT 107.770 169.980 108.725 170.200 ;
        RECT 106.465 169.190 106.660 169.520 ;
        RECT 106.885 169.190 107.140 169.520 ;
        RECT 106.885 169.020 107.055 169.190 ;
        RECT 107.310 169.020 107.480 169.690 ;
        RECT 107.655 169.250 108.345 169.810 ;
        RECT 108.515 169.080 108.725 169.980 ;
        RECT 106.125 168.850 107.055 169.020 ;
        RECT 106.125 168.815 106.300 168.850 ;
        RECT 105.770 168.450 106.300 168.815 ;
        RECT 106.725 168.280 107.055 168.680 ;
        RECT 107.225 168.450 107.480 169.020 ;
        RECT 107.770 168.910 108.725 169.080 ;
        RECT 108.895 169.810 109.295 170.660 ;
        RECT 109.485 170.200 109.765 170.660 ;
        RECT 110.285 170.370 110.610 170.830 ;
        RECT 109.485 169.980 110.610 170.200 ;
        RECT 108.895 169.250 109.990 169.810 ;
        RECT 110.160 169.520 110.610 169.980 ;
        RECT 110.780 169.690 111.165 170.660 ;
        RECT 111.340 170.405 111.675 170.830 ;
        RECT 111.845 170.225 112.030 170.630 ;
        RECT 107.770 168.450 108.055 168.910 ;
        RECT 108.225 168.280 108.495 168.740 ;
        RECT 108.895 168.450 109.295 169.250 ;
        RECT 110.160 169.190 110.715 169.520 ;
        RECT 110.160 169.080 110.610 169.190 ;
        RECT 109.485 168.910 110.610 169.080 ;
        RECT 110.885 169.020 111.165 169.690 ;
        RECT 109.485 168.450 109.765 168.910 ;
        RECT 110.285 168.280 110.610 168.740 ;
        RECT 110.780 168.450 111.165 169.020 ;
        RECT 111.365 170.050 112.030 170.225 ;
        RECT 112.235 170.050 112.565 170.830 ;
        RECT 111.365 169.020 111.705 170.050 ;
        RECT 112.735 169.860 113.005 170.630 ;
        RECT 111.875 169.690 113.005 169.860 ;
        RECT 111.875 169.190 112.125 169.690 ;
        RECT 111.365 168.850 112.050 169.020 ;
        RECT 112.305 168.940 112.665 169.520 ;
        RECT 111.340 168.280 111.675 168.680 ;
        RECT 111.845 168.450 112.050 168.850 ;
        RECT 112.835 168.780 113.005 169.690 ;
        RECT 112.260 168.280 112.535 168.760 ;
        RECT 112.745 168.450 113.005 168.780 ;
        RECT 113.175 169.755 113.445 170.660 ;
        RECT 113.615 170.070 113.945 170.830 ;
        RECT 114.125 169.900 114.295 170.660 ;
        RECT 113.175 168.955 113.345 169.755 ;
        RECT 113.630 169.730 114.295 169.900 ;
        RECT 114.555 169.740 115.765 170.830 ;
        RECT 113.630 169.585 113.800 169.730 ;
        RECT 113.515 169.255 113.800 169.585 ;
        RECT 113.630 169.000 113.800 169.255 ;
        RECT 114.035 169.180 114.365 169.550 ;
        RECT 114.555 169.200 115.075 169.740 ;
        RECT 115.245 169.030 115.765 169.570 ;
        RECT 113.175 168.450 113.435 168.955 ;
        RECT 113.630 168.830 114.295 169.000 ;
        RECT 113.615 168.280 113.945 168.660 ;
        RECT 114.125 168.450 114.295 168.830 ;
        RECT 114.555 168.280 115.765 169.030 ;
        RECT 14.650 168.110 115.850 168.280 ;
        RECT 14.735 167.360 15.945 168.110 ;
        RECT 16.120 167.560 16.375 167.850 ;
        RECT 16.545 167.730 16.875 168.110 ;
        RECT 16.120 167.390 16.870 167.560 ;
        RECT 14.735 166.820 15.255 167.360 ;
        RECT 15.425 166.650 15.945 167.190 ;
        RECT 14.735 165.560 15.945 166.650 ;
        RECT 16.120 166.570 16.470 167.220 ;
        RECT 16.640 166.400 16.870 167.390 ;
        RECT 16.120 166.230 16.870 166.400 ;
        RECT 16.120 165.730 16.375 166.230 ;
        RECT 16.545 165.560 16.875 166.060 ;
        RECT 17.045 165.730 17.215 167.850 ;
        RECT 17.575 167.750 17.905 168.110 ;
        RECT 18.075 167.720 18.570 167.890 ;
        RECT 18.775 167.720 19.630 167.890 ;
        RECT 17.445 166.530 17.905 167.580 ;
        RECT 17.385 165.745 17.710 166.530 ;
        RECT 18.075 166.360 18.245 167.720 ;
        RECT 18.415 166.810 18.765 167.430 ;
        RECT 18.935 167.210 19.290 167.430 ;
        RECT 18.935 166.620 19.105 167.210 ;
        RECT 19.460 167.010 19.630 167.720 ;
        RECT 20.505 167.650 20.835 168.110 ;
        RECT 21.045 167.750 21.395 167.920 ;
        RECT 19.835 167.180 20.625 167.430 ;
        RECT 21.045 167.360 21.305 167.750 ;
        RECT 21.615 167.660 22.565 167.940 ;
        RECT 22.735 167.670 22.925 168.110 ;
        RECT 23.095 167.730 24.165 167.900 ;
        RECT 20.795 167.010 20.965 167.190 ;
        RECT 18.075 166.190 18.470 166.360 ;
        RECT 18.640 166.230 19.105 166.620 ;
        RECT 19.275 166.840 20.965 167.010 ;
        RECT 18.300 166.060 18.470 166.190 ;
        RECT 19.275 166.060 19.445 166.840 ;
        RECT 21.135 166.670 21.305 167.360 ;
        RECT 19.805 166.500 21.305 166.670 ;
        RECT 21.495 166.700 21.705 167.490 ;
        RECT 21.875 166.870 22.225 167.490 ;
        RECT 22.395 166.880 22.565 167.660 ;
        RECT 23.095 167.500 23.265 167.730 ;
        RECT 22.735 167.330 23.265 167.500 ;
        RECT 22.735 167.050 22.955 167.330 ;
        RECT 23.435 167.160 23.675 167.560 ;
        RECT 22.395 166.710 22.800 166.880 ;
        RECT 23.135 166.790 23.675 167.160 ;
        RECT 23.845 167.375 24.165 167.730 ;
        RECT 24.410 167.650 24.715 168.110 ;
        RECT 24.885 167.400 25.140 167.930 ;
        RECT 23.845 167.200 24.170 167.375 ;
        RECT 23.845 166.900 24.760 167.200 ;
        RECT 24.020 166.870 24.760 166.900 ;
        RECT 21.495 166.540 22.170 166.700 ;
        RECT 22.630 166.620 22.800 166.710 ;
        RECT 21.495 166.530 22.460 166.540 ;
        RECT 21.135 166.360 21.305 166.500 ;
        RECT 17.880 165.560 18.130 166.020 ;
        RECT 18.300 165.730 18.550 166.060 ;
        RECT 18.765 165.730 19.445 166.060 ;
        RECT 19.615 166.160 20.690 166.330 ;
        RECT 21.135 166.190 21.695 166.360 ;
        RECT 22.000 166.240 22.460 166.530 ;
        RECT 22.630 166.450 23.850 166.620 ;
        RECT 19.615 165.820 19.785 166.160 ;
        RECT 20.020 165.560 20.350 165.990 ;
        RECT 20.520 165.820 20.690 166.160 ;
        RECT 20.985 165.560 21.355 166.020 ;
        RECT 21.525 165.730 21.695 166.190 ;
        RECT 22.630 166.070 22.800 166.450 ;
        RECT 24.020 166.280 24.190 166.870 ;
        RECT 24.930 166.750 25.140 167.400 ;
        RECT 25.315 167.385 25.605 168.110 ;
        RECT 21.930 165.730 22.800 166.070 ;
        RECT 23.390 166.110 24.190 166.280 ;
        RECT 22.970 165.560 23.220 166.020 ;
        RECT 23.390 165.820 23.560 166.110 ;
        RECT 23.740 165.560 24.070 165.940 ;
        RECT 24.410 165.560 24.715 166.700 ;
        RECT 24.885 165.870 25.140 166.750 ;
        RECT 25.780 167.370 26.035 167.940 ;
        RECT 26.205 167.710 26.535 168.110 ;
        RECT 26.960 167.575 27.490 167.940 ;
        RECT 26.960 167.540 27.135 167.575 ;
        RECT 26.205 167.370 27.135 167.540 ;
        RECT 25.315 165.560 25.605 166.725 ;
        RECT 25.780 166.700 25.950 167.370 ;
        RECT 26.205 167.200 26.375 167.370 ;
        RECT 26.120 166.870 26.375 167.200 ;
        RECT 26.600 166.870 26.795 167.200 ;
        RECT 25.780 165.730 26.115 166.700 ;
        RECT 26.285 165.560 26.455 166.700 ;
        RECT 26.625 165.900 26.795 166.870 ;
        RECT 26.965 166.240 27.135 167.370 ;
        RECT 27.305 166.580 27.475 167.380 ;
        RECT 27.680 167.090 27.955 167.940 ;
        RECT 27.675 166.920 27.955 167.090 ;
        RECT 27.680 166.780 27.955 166.920 ;
        RECT 28.125 166.580 28.315 167.940 ;
        RECT 28.495 167.575 29.005 168.110 ;
        RECT 29.225 167.300 29.470 167.905 ;
        RECT 29.915 167.435 30.175 167.940 ;
        RECT 30.355 167.730 30.685 168.110 ;
        RECT 30.865 167.560 31.035 167.940 ;
        RECT 28.515 167.130 29.745 167.300 ;
        RECT 27.305 166.410 28.315 166.580 ;
        RECT 28.485 166.565 29.235 166.755 ;
        RECT 26.965 166.070 28.090 166.240 ;
        RECT 28.485 165.900 28.655 166.565 ;
        RECT 29.405 166.320 29.745 167.130 ;
        RECT 26.625 165.730 28.655 165.900 ;
        RECT 28.825 165.560 28.995 166.320 ;
        RECT 29.230 165.910 29.745 166.320 ;
        RECT 29.915 166.635 30.085 167.435 ;
        RECT 30.370 167.390 31.035 167.560 ;
        RECT 31.760 167.400 32.015 167.930 ;
        RECT 32.185 167.650 32.490 168.110 ;
        RECT 32.735 167.730 33.805 167.900 ;
        RECT 30.370 167.135 30.540 167.390 ;
        RECT 30.255 166.805 30.540 167.135 ;
        RECT 30.775 166.840 31.105 167.210 ;
        RECT 30.370 166.660 30.540 166.805 ;
        RECT 31.760 166.750 31.970 167.400 ;
        RECT 32.735 167.375 33.055 167.730 ;
        RECT 32.730 167.200 33.055 167.375 ;
        RECT 32.140 166.900 33.055 167.200 ;
        RECT 33.225 167.160 33.465 167.560 ;
        RECT 33.635 167.500 33.805 167.730 ;
        RECT 33.975 167.670 34.165 168.110 ;
        RECT 34.335 167.660 35.285 167.940 ;
        RECT 35.505 167.750 35.855 167.920 ;
        RECT 33.635 167.330 34.165 167.500 ;
        RECT 32.140 166.870 32.880 166.900 ;
        RECT 29.915 165.730 30.185 166.635 ;
        RECT 30.370 166.490 31.035 166.660 ;
        RECT 30.355 165.560 30.685 166.320 ;
        RECT 30.865 165.730 31.035 166.490 ;
        RECT 31.760 165.870 32.015 166.750 ;
        RECT 32.185 165.560 32.490 166.700 ;
        RECT 32.710 166.280 32.880 166.870 ;
        RECT 33.225 166.790 33.765 167.160 ;
        RECT 33.945 167.050 34.165 167.330 ;
        RECT 34.335 166.880 34.505 167.660 ;
        RECT 34.100 166.710 34.505 166.880 ;
        RECT 34.675 166.870 35.025 167.490 ;
        RECT 34.100 166.620 34.270 166.710 ;
        RECT 35.195 166.700 35.405 167.490 ;
        RECT 33.050 166.450 34.270 166.620 ;
        RECT 34.730 166.540 35.405 166.700 ;
        RECT 32.710 166.110 33.510 166.280 ;
        RECT 32.830 165.560 33.160 165.940 ;
        RECT 33.340 165.820 33.510 166.110 ;
        RECT 34.100 166.070 34.270 166.450 ;
        RECT 34.440 166.530 35.405 166.540 ;
        RECT 35.595 167.360 35.855 167.750 ;
        RECT 36.065 167.650 36.395 168.110 ;
        RECT 37.270 167.720 38.125 167.890 ;
        RECT 38.330 167.720 38.825 167.890 ;
        RECT 38.995 167.750 39.325 168.110 ;
        RECT 35.595 166.670 35.765 167.360 ;
        RECT 35.935 167.010 36.105 167.190 ;
        RECT 36.275 167.180 37.065 167.430 ;
        RECT 37.270 167.010 37.440 167.720 ;
        RECT 37.610 167.210 37.965 167.430 ;
        RECT 35.935 166.840 37.625 167.010 ;
        RECT 34.440 166.240 34.900 166.530 ;
        RECT 35.595 166.500 37.095 166.670 ;
        RECT 35.595 166.360 35.765 166.500 ;
        RECT 35.205 166.190 35.765 166.360 ;
        RECT 33.680 165.560 33.930 166.020 ;
        RECT 34.100 165.730 34.970 166.070 ;
        RECT 35.205 165.730 35.375 166.190 ;
        RECT 36.210 166.160 37.285 166.330 ;
        RECT 35.545 165.560 35.915 166.020 ;
        RECT 36.210 165.820 36.380 166.160 ;
        RECT 36.550 165.560 36.880 165.990 ;
        RECT 37.115 165.820 37.285 166.160 ;
        RECT 37.455 166.060 37.625 166.840 ;
        RECT 37.795 166.620 37.965 167.210 ;
        RECT 38.135 166.810 38.485 167.430 ;
        RECT 37.795 166.230 38.260 166.620 ;
        RECT 38.655 166.360 38.825 167.720 ;
        RECT 38.995 166.530 39.455 167.580 ;
        RECT 38.430 166.190 38.825 166.360 ;
        RECT 38.430 166.060 38.600 166.190 ;
        RECT 37.455 165.730 38.135 166.060 ;
        RECT 38.350 165.730 38.600 166.060 ;
        RECT 38.770 165.560 39.020 166.020 ;
        RECT 39.190 165.745 39.515 166.530 ;
        RECT 39.685 165.730 39.855 167.850 ;
        RECT 40.025 167.730 40.355 168.110 ;
        RECT 40.525 167.560 40.780 167.850 ;
        RECT 40.955 167.600 41.260 168.110 ;
        RECT 40.030 167.390 40.780 167.560 ;
        RECT 40.030 166.400 40.260 167.390 ;
        RECT 40.430 166.570 40.780 167.220 ;
        RECT 40.955 166.870 41.270 167.430 ;
        RECT 41.440 167.120 41.690 167.930 ;
        RECT 41.860 167.585 42.120 168.110 ;
        RECT 42.300 167.120 42.550 167.930 ;
        RECT 42.720 167.550 42.980 168.110 ;
        RECT 43.150 167.460 43.410 167.915 ;
        RECT 43.580 167.630 43.840 168.110 ;
        RECT 44.010 167.460 44.270 167.915 ;
        RECT 44.440 167.630 44.700 168.110 ;
        RECT 44.870 167.460 45.130 167.915 ;
        RECT 45.300 167.630 45.545 168.110 ;
        RECT 45.715 167.460 45.990 167.915 ;
        RECT 46.160 167.630 46.405 168.110 ;
        RECT 46.575 167.460 46.835 167.915 ;
        RECT 47.015 167.630 47.265 168.110 ;
        RECT 47.435 167.460 47.695 167.915 ;
        RECT 47.875 167.630 48.125 168.110 ;
        RECT 48.295 167.460 48.555 167.915 ;
        RECT 48.735 167.630 48.995 168.110 ;
        RECT 49.165 167.460 49.425 167.915 ;
        RECT 49.595 167.630 49.895 168.110 ;
        RECT 43.150 167.290 49.895 167.460 ;
        RECT 51.075 167.385 51.365 168.110 ;
        RECT 51.540 167.400 51.795 167.930 ;
        RECT 51.965 167.650 52.270 168.110 ;
        RECT 52.515 167.730 53.585 167.900 ;
        RECT 41.440 166.870 48.560 167.120 ;
        RECT 40.030 166.230 40.780 166.400 ;
        RECT 40.025 165.560 40.355 166.060 ;
        RECT 40.525 165.730 40.780 166.230 ;
        RECT 40.965 165.560 41.260 166.370 ;
        RECT 41.440 165.730 41.685 166.870 ;
        RECT 41.860 165.560 42.120 166.370 ;
        RECT 42.300 165.735 42.550 166.870 ;
        RECT 48.730 166.700 49.895 167.290 ;
        RECT 51.540 166.750 51.750 167.400 ;
        RECT 52.515 167.375 52.835 167.730 ;
        RECT 52.510 167.200 52.835 167.375 ;
        RECT 51.920 166.900 52.835 167.200 ;
        RECT 53.005 167.160 53.245 167.560 ;
        RECT 53.415 167.500 53.585 167.730 ;
        RECT 53.755 167.670 53.945 168.110 ;
        RECT 54.115 167.660 55.065 167.940 ;
        RECT 55.285 167.750 55.635 167.920 ;
        RECT 53.415 167.330 53.945 167.500 ;
        RECT 51.920 166.870 52.660 166.900 ;
        RECT 43.150 166.475 49.895 166.700 ;
        RECT 43.150 166.460 48.555 166.475 ;
        RECT 42.720 165.565 42.980 166.360 ;
        RECT 43.150 165.735 43.410 166.460 ;
        RECT 43.580 165.565 43.840 166.290 ;
        RECT 44.010 165.735 44.270 166.460 ;
        RECT 44.440 165.565 44.700 166.290 ;
        RECT 44.870 165.735 45.130 166.460 ;
        RECT 45.300 165.565 45.560 166.290 ;
        RECT 45.730 165.735 45.990 166.460 ;
        RECT 46.160 165.565 46.405 166.290 ;
        RECT 46.575 165.735 46.835 166.460 ;
        RECT 47.020 165.565 47.265 166.290 ;
        RECT 47.435 165.735 47.695 166.460 ;
        RECT 47.880 165.565 48.125 166.290 ;
        RECT 48.295 165.735 48.555 166.460 ;
        RECT 48.740 165.565 48.995 166.290 ;
        RECT 49.165 165.735 49.455 166.475 ;
        RECT 42.720 165.560 48.995 165.565 ;
        RECT 49.625 165.560 49.895 166.305 ;
        RECT 51.075 165.560 51.365 166.725 ;
        RECT 51.540 165.870 51.795 166.750 ;
        RECT 51.965 165.560 52.270 166.700 ;
        RECT 52.490 166.280 52.660 166.870 ;
        RECT 53.005 166.790 53.545 167.160 ;
        RECT 53.725 167.050 53.945 167.330 ;
        RECT 54.115 166.880 54.285 167.660 ;
        RECT 53.880 166.710 54.285 166.880 ;
        RECT 54.455 166.870 54.805 167.490 ;
        RECT 53.880 166.620 54.050 166.710 ;
        RECT 54.975 166.700 55.185 167.490 ;
        RECT 52.830 166.450 54.050 166.620 ;
        RECT 54.510 166.540 55.185 166.700 ;
        RECT 52.490 166.110 53.290 166.280 ;
        RECT 52.610 165.560 52.940 165.940 ;
        RECT 53.120 165.820 53.290 166.110 ;
        RECT 53.880 166.070 54.050 166.450 ;
        RECT 54.220 166.530 55.185 166.540 ;
        RECT 55.375 167.360 55.635 167.750 ;
        RECT 55.845 167.650 56.175 168.110 ;
        RECT 57.050 167.720 57.905 167.890 ;
        RECT 58.110 167.720 58.605 167.890 ;
        RECT 58.775 167.750 59.105 168.110 ;
        RECT 55.375 166.670 55.545 167.360 ;
        RECT 55.715 167.010 55.885 167.190 ;
        RECT 56.055 167.180 56.845 167.430 ;
        RECT 57.050 167.010 57.220 167.720 ;
        RECT 57.390 167.210 57.745 167.430 ;
        RECT 55.715 166.840 57.405 167.010 ;
        RECT 54.220 166.240 54.680 166.530 ;
        RECT 55.375 166.500 56.875 166.670 ;
        RECT 55.375 166.360 55.545 166.500 ;
        RECT 54.985 166.190 55.545 166.360 ;
        RECT 53.460 165.560 53.710 166.020 ;
        RECT 53.880 165.730 54.750 166.070 ;
        RECT 54.985 165.730 55.155 166.190 ;
        RECT 55.990 166.160 57.065 166.330 ;
        RECT 55.325 165.560 55.695 166.020 ;
        RECT 55.990 165.820 56.160 166.160 ;
        RECT 56.330 165.560 56.660 165.990 ;
        RECT 56.895 165.820 57.065 166.160 ;
        RECT 57.235 166.060 57.405 166.840 ;
        RECT 57.575 166.620 57.745 167.210 ;
        RECT 57.915 166.810 58.265 167.430 ;
        RECT 57.575 166.230 58.040 166.620 ;
        RECT 58.435 166.360 58.605 167.720 ;
        RECT 58.775 166.530 59.235 167.580 ;
        RECT 58.210 166.190 58.605 166.360 ;
        RECT 58.210 166.060 58.380 166.190 ;
        RECT 57.235 165.730 57.915 166.060 ;
        RECT 58.130 165.730 58.380 166.060 ;
        RECT 58.550 165.560 58.800 166.020 ;
        RECT 58.970 165.745 59.295 166.530 ;
        RECT 59.465 165.730 59.635 167.850 ;
        RECT 59.805 167.730 60.135 168.110 ;
        RECT 60.305 167.560 60.560 167.850 ;
        RECT 60.795 167.630 61.075 168.110 ;
        RECT 59.810 167.390 60.560 167.560 ;
        RECT 61.245 167.460 61.505 167.850 ;
        RECT 61.680 167.630 61.935 168.110 ;
        RECT 62.105 167.460 62.400 167.850 ;
        RECT 62.580 167.630 62.855 168.110 ;
        RECT 63.025 167.610 63.325 167.940 ;
        RECT 63.555 167.630 63.835 168.110 ;
        RECT 59.810 166.400 60.040 167.390 ;
        RECT 60.750 167.290 62.400 167.460 ;
        RECT 60.210 166.570 60.560 167.220 ;
        RECT 60.750 166.780 61.155 167.290 ;
        RECT 61.325 166.950 62.465 167.120 ;
        RECT 60.750 166.610 61.505 166.780 ;
        RECT 59.810 166.230 60.560 166.400 ;
        RECT 59.805 165.560 60.135 166.060 ;
        RECT 60.305 165.730 60.560 166.230 ;
        RECT 60.790 165.560 61.075 166.430 ;
        RECT 61.245 166.360 61.505 166.610 ;
        RECT 62.295 166.700 62.465 166.950 ;
        RECT 62.635 166.870 62.985 167.440 ;
        RECT 63.155 166.700 63.325 167.610 ;
        RECT 64.005 167.460 64.265 167.850 ;
        RECT 64.440 167.630 64.695 168.110 ;
        RECT 64.865 167.460 65.160 167.850 ;
        RECT 65.340 167.630 65.615 168.110 ;
        RECT 65.785 167.610 66.085 167.940 ;
        RECT 62.295 166.530 63.325 166.700 ;
        RECT 63.510 167.290 65.160 167.460 ;
        RECT 63.510 166.780 63.915 167.290 ;
        RECT 64.085 166.950 65.225 167.120 ;
        RECT 63.510 166.610 64.265 166.780 ;
        RECT 61.245 166.190 62.365 166.360 ;
        RECT 61.245 165.730 61.505 166.190 ;
        RECT 61.680 165.560 61.935 166.020 ;
        RECT 62.105 165.730 62.365 166.190 ;
        RECT 62.535 165.560 62.845 166.360 ;
        RECT 63.015 165.730 63.325 166.530 ;
        RECT 63.550 165.560 63.835 166.430 ;
        RECT 64.005 166.360 64.265 166.610 ;
        RECT 65.055 166.700 65.225 166.950 ;
        RECT 65.395 166.870 65.745 167.440 ;
        RECT 65.915 166.700 66.085 167.610 ;
        RECT 66.265 167.580 66.595 167.940 ;
        RECT 66.765 167.750 67.095 168.110 ;
        RECT 67.295 167.580 67.625 167.940 ;
        RECT 66.265 167.370 67.625 167.580 ;
        RECT 68.135 167.350 68.845 167.940 ;
        RECT 68.615 167.260 68.845 167.350 ;
        RECT 69.475 167.340 71.145 168.110 ;
        RECT 66.255 166.870 66.565 167.200 ;
        RECT 66.775 166.870 67.150 167.200 ;
        RECT 67.470 166.870 67.965 167.200 ;
        RECT 65.055 166.530 66.085 166.700 ;
        RECT 64.005 166.190 65.125 166.360 ;
        RECT 64.005 165.730 64.265 166.190 ;
        RECT 64.440 165.560 64.695 166.020 ;
        RECT 64.865 165.730 65.125 166.190 ;
        RECT 65.295 165.560 65.605 166.360 ;
        RECT 65.775 165.730 66.085 166.530 ;
        RECT 66.265 165.560 66.595 166.620 ;
        RECT 66.775 165.945 66.945 166.870 ;
        RECT 67.115 166.380 67.445 166.600 ;
        RECT 67.640 166.580 67.965 166.870 ;
        RECT 68.140 166.580 68.470 167.120 ;
        RECT 68.640 166.380 68.845 167.260 ;
        RECT 67.115 166.150 68.845 166.380 ;
        RECT 67.115 165.750 67.445 166.150 ;
        RECT 67.615 165.560 67.945 165.920 ;
        RECT 68.145 165.730 68.845 166.150 ;
        RECT 69.475 166.650 70.225 167.170 ;
        RECT 70.395 166.820 71.145 167.340 ;
        RECT 71.375 167.290 71.585 168.110 ;
        RECT 71.755 167.310 72.085 167.940 ;
        RECT 71.755 166.710 72.005 167.310 ;
        RECT 72.255 167.290 72.485 168.110 ;
        RECT 72.970 167.300 73.215 167.905 ;
        RECT 73.435 167.575 73.945 168.110 ;
        RECT 72.695 167.130 73.925 167.300 ;
        RECT 72.175 166.870 72.505 167.120 ;
        RECT 69.475 165.560 71.145 166.650 ;
        RECT 71.375 165.560 71.585 166.700 ;
        RECT 71.755 165.730 72.085 166.710 ;
        RECT 72.255 165.560 72.485 166.700 ;
        RECT 72.695 166.320 73.035 167.130 ;
        RECT 73.205 166.565 73.955 166.755 ;
        RECT 72.695 165.910 73.210 166.320 ;
        RECT 73.445 165.560 73.615 166.320 ;
        RECT 73.785 165.900 73.955 166.565 ;
        RECT 74.125 166.580 74.315 167.940 ;
        RECT 74.485 167.430 74.760 167.940 ;
        RECT 74.950 167.575 75.480 167.940 ;
        RECT 75.905 167.710 76.235 168.110 ;
        RECT 75.305 167.540 75.480 167.575 ;
        RECT 74.485 167.260 74.765 167.430 ;
        RECT 74.485 166.780 74.760 167.260 ;
        RECT 74.965 166.580 75.135 167.380 ;
        RECT 74.125 166.410 75.135 166.580 ;
        RECT 75.305 167.370 76.235 167.540 ;
        RECT 76.405 167.370 76.660 167.940 ;
        RECT 76.835 167.385 77.125 168.110 ;
        RECT 75.305 166.240 75.475 167.370 ;
        RECT 76.065 167.200 76.235 167.370 ;
        RECT 74.350 166.070 75.475 166.240 ;
        RECT 75.645 166.870 75.840 167.200 ;
        RECT 76.065 166.870 76.320 167.200 ;
        RECT 75.645 165.900 75.815 166.870 ;
        RECT 76.490 166.700 76.660 167.370 ;
        RECT 77.355 167.290 77.565 168.110 ;
        RECT 77.735 167.310 78.065 167.940 ;
        RECT 73.785 165.730 75.815 165.900 ;
        RECT 75.985 165.560 76.155 166.700 ;
        RECT 76.325 165.730 76.660 166.700 ;
        RECT 76.835 165.560 77.125 166.725 ;
        RECT 77.735 166.710 77.985 167.310 ;
        RECT 78.235 167.290 78.465 168.110 ;
        RECT 79.135 167.600 79.440 168.110 ;
        RECT 78.155 166.870 78.485 167.120 ;
        RECT 79.135 166.870 79.450 167.430 ;
        RECT 79.620 167.120 79.870 167.930 ;
        RECT 80.040 167.585 80.300 168.110 ;
        RECT 80.480 167.120 80.730 167.930 ;
        RECT 80.900 167.550 81.160 168.110 ;
        RECT 81.330 167.460 81.590 167.915 ;
        RECT 81.760 167.630 82.020 168.110 ;
        RECT 82.190 167.460 82.450 167.915 ;
        RECT 82.620 167.630 82.880 168.110 ;
        RECT 83.050 167.460 83.310 167.915 ;
        RECT 83.480 167.630 83.725 168.110 ;
        RECT 83.895 167.460 84.170 167.915 ;
        RECT 84.340 167.630 84.585 168.110 ;
        RECT 84.755 167.460 85.015 167.915 ;
        RECT 85.195 167.630 85.445 168.110 ;
        RECT 85.615 167.460 85.875 167.915 ;
        RECT 86.055 167.630 86.305 168.110 ;
        RECT 86.475 167.460 86.735 167.915 ;
        RECT 86.915 167.630 87.175 168.110 ;
        RECT 87.345 167.460 87.605 167.915 ;
        RECT 87.775 167.630 88.075 168.110 ;
        RECT 81.330 167.290 88.075 167.460 ;
        RECT 89.295 167.290 89.525 168.110 ;
        RECT 89.695 167.310 90.025 167.940 ;
        RECT 79.620 166.870 86.740 167.120 ;
        RECT 77.355 165.560 77.565 166.700 ;
        RECT 77.735 165.730 78.065 166.710 ;
        RECT 78.235 165.560 78.465 166.700 ;
        RECT 79.145 165.560 79.440 166.370 ;
        RECT 79.620 165.730 79.865 166.870 ;
        RECT 80.040 165.560 80.300 166.370 ;
        RECT 80.480 165.735 80.730 166.870 ;
        RECT 86.910 166.700 88.075 167.290 ;
        RECT 89.275 166.870 89.605 167.120 ;
        RECT 89.775 166.710 90.025 167.310 ;
        RECT 90.195 167.290 90.405 168.110 ;
        RECT 90.635 167.600 90.940 168.110 ;
        RECT 90.635 166.870 90.950 167.430 ;
        RECT 91.120 167.120 91.370 167.930 ;
        RECT 91.540 167.585 91.800 168.110 ;
        RECT 91.980 167.120 92.230 167.930 ;
        RECT 92.400 167.550 92.660 168.110 ;
        RECT 92.830 167.460 93.090 167.915 ;
        RECT 93.260 167.630 93.520 168.110 ;
        RECT 93.690 167.460 93.950 167.915 ;
        RECT 94.120 167.630 94.380 168.110 ;
        RECT 94.550 167.460 94.810 167.915 ;
        RECT 94.980 167.630 95.225 168.110 ;
        RECT 95.395 167.460 95.670 167.915 ;
        RECT 95.840 167.630 96.085 168.110 ;
        RECT 96.255 167.460 96.515 167.915 ;
        RECT 96.695 167.630 96.945 168.110 ;
        RECT 97.115 167.460 97.375 167.915 ;
        RECT 97.555 167.630 97.805 168.110 ;
        RECT 97.975 167.460 98.235 167.915 ;
        RECT 98.415 167.630 98.675 168.110 ;
        RECT 98.845 167.460 99.105 167.915 ;
        RECT 99.275 167.630 99.575 168.110 ;
        RECT 92.830 167.290 99.575 167.460 ;
        RECT 100.505 167.420 100.835 168.110 ;
        RECT 101.295 167.515 101.915 167.940 ;
        RECT 102.085 167.620 102.415 168.110 ;
        RECT 91.120 166.870 98.240 167.120 ;
        RECT 81.330 166.475 88.075 166.700 ;
        RECT 81.330 166.460 86.735 166.475 ;
        RECT 80.900 165.565 81.160 166.360 ;
        RECT 81.330 165.735 81.590 166.460 ;
        RECT 81.760 165.565 82.020 166.290 ;
        RECT 82.190 165.735 82.450 166.460 ;
        RECT 82.620 165.565 82.880 166.290 ;
        RECT 83.050 165.735 83.310 166.460 ;
        RECT 83.480 165.565 83.740 166.290 ;
        RECT 83.910 165.735 84.170 166.460 ;
        RECT 84.340 165.565 84.585 166.290 ;
        RECT 84.755 165.735 85.015 166.460 ;
        RECT 85.200 165.565 85.445 166.290 ;
        RECT 85.615 165.735 85.875 166.460 ;
        RECT 86.060 165.565 86.305 166.290 ;
        RECT 86.475 165.735 86.735 166.460 ;
        RECT 86.920 165.565 87.175 166.290 ;
        RECT 87.345 165.735 87.635 166.475 ;
        RECT 80.900 165.560 87.175 165.565 ;
        RECT 87.805 165.560 88.075 166.305 ;
        RECT 89.295 165.560 89.525 166.700 ;
        RECT 89.695 165.730 90.025 166.710 ;
        RECT 90.195 165.560 90.405 166.700 ;
        RECT 90.645 165.560 90.940 166.370 ;
        RECT 91.120 165.730 91.365 166.870 ;
        RECT 91.540 165.560 91.800 166.370 ;
        RECT 91.980 165.735 92.230 166.870 ;
        RECT 98.410 166.750 99.575 167.290 ;
        RECT 101.555 167.180 101.915 167.515 ;
        RECT 100.495 166.900 101.915 167.180 ;
        RECT 98.410 166.700 99.605 166.750 ;
        RECT 92.830 166.580 99.605 166.700 ;
        RECT 92.830 166.475 99.575 166.580 ;
        RECT 92.830 166.460 98.235 166.475 ;
        RECT 92.400 165.565 92.660 166.360 ;
        RECT 92.830 165.735 93.090 166.460 ;
        RECT 93.260 165.565 93.520 166.290 ;
        RECT 93.690 165.735 93.950 166.460 ;
        RECT 94.120 165.565 94.380 166.290 ;
        RECT 94.550 165.735 94.810 166.460 ;
        RECT 94.980 165.565 95.240 166.290 ;
        RECT 95.410 165.735 95.670 166.460 ;
        RECT 95.840 165.565 96.085 166.290 ;
        RECT 96.255 165.735 96.515 166.460 ;
        RECT 96.700 165.565 96.945 166.290 ;
        RECT 97.115 165.735 97.375 166.460 ;
        RECT 97.560 165.565 97.805 166.290 ;
        RECT 97.975 165.735 98.235 166.460 ;
        RECT 98.420 165.565 98.675 166.290 ;
        RECT 98.845 165.735 99.135 166.475 ;
        RECT 92.400 165.560 98.675 165.565 ;
        RECT 99.305 165.560 99.575 166.305 ;
        RECT 99.965 165.560 100.295 166.730 ;
        RECT 100.495 165.730 100.825 166.900 ;
        RECT 101.025 165.560 101.355 166.730 ;
        RECT 101.555 165.730 101.915 166.900 ;
        RECT 102.085 166.870 102.425 167.450 ;
        RECT 102.595 167.385 102.885 168.110 ;
        RECT 103.555 167.290 103.785 168.110 ;
        RECT 103.955 167.310 104.285 167.940 ;
        RECT 103.535 166.870 103.865 167.120 ;
        RECT 102.085 165.560 102.415 166.700 ;
        RECT 102.595 165.560 102.885 166.725 ;
        RECT 104.035 166.710 104.285 167.310 ;
        RECT 104.455 167.290 104.665 168.110 ;
        RECT 104.900 167.400 105.155 167.930 ;
        RECT 105.325 167.650 105.630 168.110 ;
        RECT 105.875 167.730 106.945 167.900 ;
        RECT 103.555 165.560 103.785 166.700 ;
        RECT 103.955 165.730 104.285 166.710 ;
        RECT 104.900 166.750 105.110 167.400 ;
        RECT 105.875 167.375 106.195 167.730 ;
        RECT 105.870 167.200 106.195 167.375 ;
        RECT 105.280 166.900 106.195 167.200 ;
        RECT 106.365 167.160 106.605 167.560 ;
        RECT 106.775 167.500 106.945 167.730 ;
        RECT 107.115 167.670 107.305 168.110 ;
        RECT 107.475 167.660 108.425 167.940 ;
        RECT 108.645 167.750 108.995 167.920 ;
        RECT 106.775 167.330 107.305 167.500 ;
        RECT 105.280 166.870 106.020 166.900 ;
        RECT 104.455 165.560 104.665 166.700 ;
        RECT 104.900 165.870 105.155 166.750 ;
        RECT 105.325 165.560 105.630 166.700 ;
        RECT 105.850 166.280 106.020 166.870 ;
        RECT 106.365 166.790 106.905 167.160 ;
        RECT 107.085 167.050 107.305 167.330 ;
        RECT 107.475 166.880 107.645 167.660 ;
        RECT 107.240 166.710 107.645 166.880 ;
        RECT 107.815 166.870 108.165 167.490 ;
        RECT 107.240 166.620 107.410 166.710 ;
        RECT 108.335 166.700 108.545 167.490 ;
        RECT 106.190 166.450 107.410 166.620 ;
        RECT 107.870 166.540 108.545 166.700 ;
        RECT 105.850 166.110 106.650 166.280 ;
        RECT 105.970 165.560 106.300 165.940 ;
        RECT 106.480 165.820 106.650 166.110 ;
        RECT 107.240 166.070 107.410 166.450 ;
        RECT 107.580 166.530 108.545 166.540 ;
        RECT 108.735 167.360 108.995 167.750 ;
        RECT 109.205 167.650 109.535 168.110 ;
        RECT 110.410 167.720 111.265 167.890 ;
        RECT 111.470 167.720 111.965 167.890 ;
        RECT 112.135 167.750 112.465 168.110 ;
        RECT 108.735 166.670 108.905 167.360 ;
        RECT 109.075 167.010 109.245 167.190 ;
        RECT 109.415 167.180 110.205 167.430 ;
        RECT 110.410 167.010 110.580 167.720 ;
        RECT 110.750 167.210 111.105 167.430 ;
        RECT 109.075 166.840 110.765 167.010 ;
        RECT 107.580 166.240 108.040 166.530 ;
        RECT 108.735 166.500 110.235 166.670 ;
        RECT 108.735 166.360 108.905 166.500 ;
        RECT 108.345 166.190 108.905 166.360 ;
        RECT 106.820 165.560 107.070 166.020 ;
        RECT 107.240 165.730 108.110 166.070 ;
        RECT 108.345 165.730 108.515 166.190 ;
        RECT 109.350 166.160 110.425 166.330 ;
        RECT 108.685 165.560 109.055 166.020 ;
        RECT 109.350 165.820 109.520 166.160 ;
        RECT 109.690 165.560 110.020 165.990 ;
        RECT 110.255 165.820 110.425 166.160 ;
        RECT 110.595 166.060 110.765 166.840 ;
        RECT 110.935 166.620 111.105 167.210 ;
        RECT 111.275 166.810 111.625 167.430 ;
        RECT 110.935 166.230 111.400 166.620 ;
        RECT 111.795 166.360 111.965 167.720 ;
        RECT 112.135 166.530 112.595 167.580 ;
        RECT 111.570 166.190 111.965 166.360 ;
        RECT 111.570 166.060 111.740 166.190 ;
        RECT 110.595 165.730 111.275 166.060 ;
        RECT 111.490 165.730 111.740 166.060 ;
        RECT 111.910 165.560 112.160 166.020 ;
        RECT 112.330 165.745 112.655 166.530 ;
        RECT 112.825 165.730 112.995 167.850 ;
        RECT 113.165 167.730 113.495 168.110 ;
        RECT 113.665 167.560 113.920 167.850 ;
        RECT 113.170 167.390 113.920 167.560 ;
        RECT 113.170 166.400 113.400 167.390 ;
        RECT 114.555 167.360 115.765 168.110 ;
        RECT 113.570 166.570 113.920 167.220 ;
        RECT 114.555 166.650 115.075 167.190 ;
        RECT 115.245 166.820 115.765 167.360 ;
        RECT 113.170 166.230 113.920 166.400 ;
        RECT 113.165 165.560 113.495 166.060 ;
        RECT 113.665 165.730 113.920 166.230 ;
        RECT 114.555 165.560 115.765 166.650 ;
        RECT 14.650 165.390 115.850 165.560 ;
        RECT 14.735 164.300 15.945 165.390 ;
        RECT 16.205 164.720 16.375 165.220 ;
        RECT 16.545 164.890 16.875 165.390 ;
        RECT 16.205 164.550 16.870 164.720 ;
        RECT 14.735 163.590 15.255 164.130 ;
        RECT 15.425 163.760 15.945 164.300 ;
        RECT 16.120 163.730 16.470 164.380 ;
        RECT 14.735 162.840 15.945 163.590 ;
        RECT 16.640 163.560 16.870 164.550 ;
        RECT 16.205 163.390 16.870 163.560 ;
        RECT 16.205 163.100 16.375 163.390 ;
        RECT 16.545 162.840 16.875 163.220 ;
        RECT 17.045 163.100 17.270 165.220 ;
        RECT 17.485 164.890 17.815 165.390 ;
        RECT 17.985 164.720 18.155 165.220 ;
        RECT 18.390 165.005 19.220 165.175 ;
        RECT 19.460 165.010 19.840 165.390 ;
        RECT 17.460 164.550 18.155 164.720 ;
        RECT 17.460 163.580 17.630 164.550 ;
        RECT 17.800 163.760 18.210 164.380 ;
        RECT 18.380 164.330 18.880 164.710 ;
        RECT 17.460 163.390 18.155 163.580 ;
        RECT 18.380 163.460 18.600 164.330 ;
        RECT 19.050 164.160 19.220 165.005 ;
        RECT 20.020 164.840 20.190 165.130 ;
        RECT 20.360 165.010 20.690 165.390 ;
        RECT 21.160 164.920 21.790 165.170 ;
        RECT 21.970 165.010 22.390 165.390 ;
        RECT 21.620 164.840 21.790 164.920 ;
        RECT 22.590 164.840 22.830 165.130 ;
        RECT 19.390 164.590 20.760 164.840 ;
        RECT 19.390 164.330 19.640 164.590 ;
        RECT 20.150 164.160 20.400 164.320 ;
        RECT 19.050 163.990 20.400 164.160 ;
        RECT 19.050 163.950 19.470 163.990 ;
        RECT 18.780 163.400 19.130 163.770 ;
        RECT 17.485 162.840 17.815 163.220 ;
        RECT 17.985 163.060 18.155 163.390 ;
        RECT 19.300 163.220 19.470 163.950 ;
        RECT 20.570 163.820 20.760 164.590 ;
        RECT 19.640 163.490 20.050 163.820 ;
        RECT 20.340 163.480 20.760 163.820 ;
        RECT 20.930 164.410 21.450 164.720 ;
        RECT 21.620 164.670 22.830 164.840 ;
        RECT 23.060 164.700 23.390 165.390 ;
        RECT 20.930 163.650 21.100 164.410 ;
        RECT 21.270 163.820 21.450 164.230 ;
        RECT 21.620 164.160 21.790 164.670 ;
        RECT 23.560 164.520 23.730 165.130 ;
        RECT 24.000 164.670 24.330 165.180 ;
        RECT 23.560 164.500 23.880 164.520 ;
        RECT 21.960 164.330 23.880 164.500 ;
        RECT 21.620 163.990 23.520 164.160 ;
        RECT 21.850 163.650 22.180 163.770 ;
        RECT 20.930 163.480 22.180 163.650 ;
        RECT 18.455 163.020 19.470 163.220 ;
        RECT 19.640 162.840 20.050 163.280 ;
        RECT 20.340 163.050 20.590 163.480 ;
        RECT 20.790 162.840 21.110 163.300 ;
        RECT 22.350 163.230 22.520 163.990 ;
        RECT 23.190 163.930 23.520 163.990 ;
        RECT 22.710 163.760 23.040 163.820 ;
        RECT 22.710 163.490 23.370 163.760 ;
        RECT 23.690 163.435 23.880 164.330 ;
        RECT 21.670 163.060 22.520 163.230 ;
        RECT 22.720 162.840 23.380 163.320 ;
        RECT 23.560 163.105 23.880 163.435 ;
        RECT 24.080 164.080 24.330 164.670 ;
        RECT 24.510 164.590 24.795 165.390 ;
        RECT 24.975 164.410 25.230 165.080 ;
        RECT 26.785 164.645 27.055 165.390 ;
        RECT 27.685 165.385 33.960 165.390 ;
        RECT 27.225 164.475 27.515 165.215 ;
        RECT 27.685 164.660 27.940 165.385 ;
        RECT 28.125 164.490 28.385 165.215 ;
        RECT 28.555 164.660 28.800 165.385 ;
        RECT 28.985 164.490 29.245 165.215 ;
        RECT 29.415 164.660 29.660 165.385 ;
        RECT 29.845 164.490 30.105 165.215 ;
        RECT 30.275 164.660 30.520 165.385 ;
        RECT 30.690 164.490 30.950 165.215 ;
        RECT 31.120 164.660 31.380 165.385 ;
        RECT 31.550 164.490 31.810 165.215 ;
        RECT 31.980 164.660 32.240 165.385 ;
        RECT 32.410 164.490 32.670 165.215 ;
        RECT 32.840 164.660 33.100 165.385 ;
        RECT 33.270 164.490 33.530 165.215 ;
        RECT 33.700 164.590 33.960 165.385 ;
        RECT 28.125 164.475 33.530 164.490 ;
        RECT 24.080 163.750 24.880 164.080 ;
        RECT 24.080 163.100 24.330 163.750 ;
        RECT 25.050 163.550 25.230 164.410 ;
        RECT 24.975 163.350 25.230 163.550 ;
        RECT 26.785 164.250 33.530 164.475 ;
        RECT 26.785 163.660 27.950 164.250 ;
        RECT 34.130 164.080 34.380 165.215 ;
        RECT 34.560 164.580 34.820 165.390 ;
        RECT 34.995 164.080 35.240 165.220 ;
        RECT 35.420 164.580 35.715 165.390 ;
        RECT 35.955 164.555 36.210 165.390 ;
        RECT 36.380 164.385 36.640 165.190 ;
        RECT 36.810 164.555 37.070 165.390 ;
        RECT 37.240 164.385 37.495 165.190 ;
        RECT 35.895 164.215 37.495 164.385 ;
        RECT 38.195 164.225 38.485 165.390 ;
        RECT 39.115 164.315 39.385 165.220 ;
        RECT 39.555 164.630 39.885 165.390 ;
        RECT 40.065 164.460 40.235 165.220 ;
        RECT 28.120 163.830 35.240 164.080 ;
        RECT 26.785 163.490 33.530 163.660 ;
        RECT 24.510 162.840 24.795 163.300 ;
        RECT 24.975 163.180 25.315 163.350 ;
        RECT 24.975 163.020 25.230 163.180 ;
        RECT 26.785 162.840 27.085 163.320 ;
        RECT 27.255 163.035 27.515 163.490 ;
        RECT 27.685 162.840 27.945 163.320 ;
        RECT 28.125 163.035 28.385 163.490 ;
        RECT 28.555 162.840 28.805 163.320 ;
        RECT 28.985 163.035 29.245 163.490 ;
        RECT 29.415 162.840 29.665 163.320 ;
        RECT 29.845 163.035 30.105 163.490 ;
        RECT 30.275 162.840 30.520 163.320 ;
        RECT 30.690 163.035 30.965 163.490 ;
        RECT 31.135 162.840 31.380 163.320 ;
        RECT 31.550 163.035 31.810 163.490 ;
        RECT 31.980 162.840 32.240 163.320 ;
        RECT 32.410 163.035 32.670 163.490 ;
        RECT 32.840 162.840 33.100 163.320 ;
        RECT 33.270 163.035 33.530 163.490 ;
        RECT 33.700 162.840 33.960 163.400 ;
        RECT 34.130 163.020 34.380 163.830 ;
        RECT 34.560 162.840 34.820 163.365 ;
        RECT 34.990 163.020 35.240 163.830 ;
        RECT 35.410 163.520 35.725 164.080 ;
        RECT 35.895 163.650 36.175 164.215 ;
        RECT 36.345 163.820 37.565 164.045 ;
        RECT 35.895 163.480 36.625 163.650 ;
        RECT 35.420 162.840 35.725 163.350 ;
        RECT 35.900 162.840 36.230 163.310 ;
        RECT 36.400 163.035 36.625 163.480 ;
        RECT 36.795 162.840 37.090 163.365 ;
        RECT 38.195 162.840 38.485 163.565 ;
        RECT 39.115 163.515 39.285 164.315 ;
        RECT 39.570 164.290 40.235 164.460 ;
        RECT 39.570 164.145 39.740 164.290 ;
        RECT 39.455 163.815 39.740 164.145 ;
        RECT 40.500 164.250 40.835 165.220 ;
        RECT 41.005 164.250 41.175 165.390 ;
        RECT 41.345 165.050 43.375 165.220 ;
        RECT 39.570 163.560 39.740 163.815 ;
        RECT 39.975 163.740 40.305 164.110 ;
        RECT 40.500 163.580 40.670 164.250 ;
        RECT 41.345 164.080 41.515 165.050 ;
        RECT 40.840 163.750 41.095 164.080 ;
        RECT 41.320 163.750 41.515 164.080 ;
        RECT 41.685 164.710 42.810 164.880 ;
        RECT 40.925 163.580 41.095 163.750 ;
        RECT 41.685 163.580 41.855 164.710 ;
        RECT 39.115 163.010 39.375 163.515 ;
        RECT 39.570 163.390 40.235 163.560 ;
        RECT 39.555 162.840 39.885 163.220 ;
        RECT 40.065 163.010 40.235 163.390 ;
        RECT 40.500 163.010 40.755 163.580 ;
        RECT 40.925 163.410 41.855 163.580 ;
        RECT 42.025 164.370 43.035 164.540 ;
        RECT 42.025 163.570 42.195 164.370 ;
        RECT 42.400 164.030 42.675 164.170 ;
        RECT 42.395 163.860 42.675 164.030 ;
        RECT 41.680 163.375 41.855 163.410 ;
        RECT 40.925 162.840 41.255 163.240 ;
        RECT 41.680 163.010 42.210 163.375 ;
        RECT 42.400 163.010 42.675 163.860 ;
        RECT 42.845 163.010 43.035 164.370 ;
        RECT 43.205 164.385 43.375 165.050 ;
        RECT 43.545 164.630 43.715 165.390 ;
        RECT 43.950 164.630 44.465 165.040 ;
        RECT 43.205 164.195 43.955 164.385 ;
        RECT 44.125 163.820 44.465 164.630 ;
        RECT 43.235 163.650 44.465 163.820 ;
        RECT 44.635 164.300 46.305 165.390 ;
        RECT 46.475 164.630 46.990 165.040 ;
        RECT 47.225 164.630 47.395 165.390 ;
        RECT 47.565 165.050 49.595 165.220 ;
        RECT 44.635 163.780 45.385 164.300 ;
        RECT 43.215 162.840 43.725 163.375 ;
        RECT 43.945 163.045 44.190 163.650 ;
        RECT 45.555 163.610 46.305 164.130 ;
        RECT 46.475 163.820 46.815 164.630 ;
        RECT 47.565 164.385 47.735 165.050 ;
        RECT 48.130 164.710 49.255 164.880 ;
        RECT 46.985 164.195 47.735 164.385 ;
        RECT 47.905 164.370 48.915 164.540 ;
        RECT 46.475 163.650 47.705 163.820 ;
        RECT 44.635 162.840 46.305 163.610 ;
        RECT 46.750 163.045 46.995 163.650 ;
        RECT 47.215 162.840 47.725 163.375 ;
        RECT 47.905 163.010 48.095 164.370 ;
        RECT 48.265 163.350 48.540 164.170 ;
        RECT 48.745 163.570 48.915 164.370 ;
        RECT 49.085 163.580 49.255 164.710 ;
        RECT 49.425 164.080 49.595 165.050 ;
        RECT 49.765 164.250 49.935 165.390 ;
        RECT 50.105 164.250 50.440 165.220 ;
        RECT 49.425 163.750 49.620 164.080 ;
        RECT 49.845 163.750 50.100 164.080 ;
        RECT 49.845 163.580 50.015 163.750 ;
        RECT 50.270 163.580 50.440 164.250 ;
        RECT 50.615 164.630 51.130 165.040 ;
        RECT 51.365 164.630 51.535 165.390 ;
        RECT 51.705 165.050 53.735 165.220 ;
        RECT 50.615 163.820 50.955 164.630 ;
        RECT 51.705 164.385 51.875 165.050 ;
        RECT 52.270 164.710 53.395 164.880 ;
        RECT 51.125 164.195 51.875 164.385 ;
        RECT 52.045 164.370 53.055 164.540 ;
        RECT 50.615 163.650 51.845 163.820 ;
        RECT 49.085 163.410 50.015 163.580 ;
        RECT 49.085 163.375 49.260 163.410 ;
        RECT 48.265 163.180 48.545 163.350 ;
        RECT 48.265 163.010 48.540 163.180 ;
        RECT 48.730 163.010 49.260 163.375 ;
        RECT 49.685 162.840 50.015 163.240 ;
        RECT 50.185 163.010 50.440 163.580 ;
        RECT 50.890 163.045 51.135 163.650 ;
        RECT 51.355 162.840 51.865 163.375 ;
        RECT 52.045 163.010 52.235 164.370 ;
        RECT 52.405 163.690 52.680 164.170 ;
        RECT 52.405 163.520 52.685 163.690 ;
        RECT 52.885 163.570 53.055 164.370 ;
        RECT 53.225 163.580 53.395 164.710 ;
        RECT 53.565 164.080 53.735 165.050 ;
        RECT 53.905 164.250 54.075 165.390 ;
        RECT 54.245 164.250 54.580 165.220 ;
        RECT 53.565 163.750 53.760 164.080 ;
        RECT 53.985 163.750 54.240 164.080 ;
        RECT 53.985 163.580 54.155 163.750 ;
        RECT 54.410 163.580 54.580 164.250 ;
        RECT 52.405 163.010 52.680 163.520 ;
        RECT 53.225 163.410 54.155 163.580 ;
        RECT 53.225 163.375 53.400 163.410 ;
        RECT 52.870 163.010 53.400 163.375 ;
        RECT 53.825 162.840 54.155 163.240 ;
        RECT 54.325 163.010 54.580 163.580 ;
        RECT 54.755 164.315 55.025 165.220 ;
        RECT 55.195 164.630 55.525 165.390 ;
        RECT 55.705 164.460 55.875 165.220 ;
        RECT 54.755 163.515 54.925 164.315 ;
        RECT 55.210 164.290 55.875 164.460 ;
        RECT 56.225 164.460 56.395 165.220 ;
        RECT 56.575 164.630 56.905 165.390 ;
        RECT 56.225 164.290 56.890 164.460 ;
        RECT 57.075 164.315 57.345 165.220 ;
        RECT 55.210 164.145 55.380 164.290 ;
        RECT 55.095 163.815 55.380 164.145 ;
        RECT 56.720 164.145 56.890 164.290 ;
        RECT 55.210 163.560 55.380 163.815 ;
        RECT 55.615 163.740 55.945 164.110 ;
        RECT 56.155 163.740 56.485 164.110 ;
        RECT 56.720 163.815 57.005 164.145 ;
        RECT 56.720 163.560 56.890 163.815 ;
        RECT 54.755 163.010 55.015 163.515 ;
        RECT 55.210 163.390 55.875 163.560 ;
        RECT 55.195 162.840 55.525 163.220 ;
        RECT 55.705 163.010 55.875 163.390 ;
        RECT 56.225 163.390 56.890 163.560 ;
        RECT 57.175 163.515 57.345 164.315 ;
        RECT 58.015 164.250 58.245 165.390 ;
        RECT 58.415 164.240 58.745 165.220 ;
        RECT 58.915 164.250 59.125 165.390 ;
        RECT 60.425 164.240 60.755 165.390 ;
        RECT 60.925 164.370 61.095 165.220 ;
        RECT 61.265 164.590 61.595 165.390 ;
        RECT 61.765 164.370 61.935 165.220 ;
        RECT 62.115 164.590 62.355 165.390 ;
        RECT 62.525 164.410 62.855 165.220 ;
        RECT 57.995 163.830 58.325 164.080 ;
        RECT 56.225 163.010 56.395 163.390 ;
        RECT 56.575 162.840 56.905 163.220 ;
        RECT 57.085 163.010 57.345 163.515 ;
        RECT 58.015 162.840 58.245 163.660 ;
        RECT 58.495 163.640 58.745 164.240 ;
        RECT 60.925 164.200 61.935 164.370 ;
        RECT 62.140 164.240 62.855 164.410 ;
        RECT 60.925 163.660 61.420 164.200 ;
        RECT 62.140 164.000 62.310 164.240 ;
        RECT 63.955 164.225 64.245 165.390 ;
        RECT 65.340 164.240 65.600 165.390 ;
        RECT 65.775 164.315 66.030 165.220 ;
        RECT 66.200 164.630 66.530 165.390 ;
        RECT 66.745 164.460 66.915 165.220 ;
        RECT 61.810 163.830 62.310 164.000 ;
        RECT 62.480 163.830 62.860 164.070 ;
        RECT 62.140 163.660 62.310 163.830 ;
        RECT 58.415 163.010 58.745 163.640 ;
        RECT 58.915 162.840 59.125 163.660 ;
        RECT 60.425 162.840 60.755 163.640 ;
        RECT 60.925 163.490 61.935 163.660 ;
        RECT 62.140 163.490 62.775 163.660 ;
        RECT 60.925 163.010 61.095 163.490 ;
        RECT 61.265 162.840 61.595 163.320 ;
        RECT 61.765 163.010 61.935 163.490 ;
        RECT 62.185 162.840 62.425 163.320 ;
        RECT 62.605 163.010 62.775 163.490 ;
        RECT 63.955 162.840 64.245 163.565 ;
        RECT 65.340 162.840 65.600 163.680 ;
        RECT 65.775 163.585 65.945 164.315 ;
        RECT 66.200 164.290 66.915 164.460 ;
        RECT 67.265 164.460 67.435 165.220 ;
        RECT 67.650 164.630 67.980 165.390 ;
        RECT 67.265 164.290 67.980 164.460 ;
        RECT 68.150 164.315 68.405 165.220 ;
        RECT 66.200 164.080 66.370 164.290 ;
        RECT 66.115 163.750 66.370 164.080 ;
        RECT 65.775 163.010 66.030 163.585 ;
        RECT 66.200 163.560 66.370 163.750 ;
        RECT 66.650 163.740 67.005 164.110 ;
        RECT 67.175 163.740 67.530 164.110 ;
        RECT 67.810 164.080 67.980 164.290 ;
        RECT 67.810 163.750 68.065 164.080 ;
        RECT 67.810 163.560 67.980 163.750 ;
        RECT 68.235 163.585 68.405 164.315 ;
        RECT 68.580 164.240 68.840 165.390 ;
        RECT 69.935 164.300 73.445 165.390 ;
        RECT 73.615 164.630 74.130 165.040 ;
        RECT 74.365 164.630 74.535 165.390 ;
        RECT 74.705 165.050 76.735 165.220 ;
        RECT 69.935 163.780 71.625 164.300 ;
        RECT 66.200 163.390 66.915 163.560 ;
        RECT 66.200 162.840 66.530 163.220 ;
        RECT 66.745 163.010 66.915 163.390 ;
        RECT 67.265 163.390 67.980 163.560 ;
        RECT 67.265 163.010 67.435 163.390 ;
        RECT 67.650 162.840 67.980 163.220 ;
        RECT 68.150 163.010 68.405 163.585 ;
        RECT 68.580 162.840 68.840 163.680 ;
        RECT 71.795 163.610 73.445 164.130 ;
        RECT 73.615 163.820 73.955 164.630 ;
        RECT 74.705 164.385 74.875 165.050 ;
        RECT 75.270 164.710 76.395 164.880 ;
        RECT 74.125 164.195 74.875 164.385 ;
        RECT 75.045 164.370 76.055 164.540 ;
        RECT 73.615 163.650 74.845 163.820 ;
        RECT 69.935 162.840 73.445 163.610 ;
        RECT 73.890 163.045 74.135 163.650 ;
        RECT 74.355 162.840 74.865 163.375 ;
        RECT 75.045 163.010 75.235 164.370 ;
        RECT 75.405 163.350 75.680 164.170 ;
        RECT 75.885 163.570 76.055 164.370 ;
        RECT 76.225 163.580 76.395 164.710 ;
        RECT 76.565 164.080 76.735 165.050 ;
        RECT 76.905 164.250 77.075 165.390 ;
        RECT 77.245 164.250 77.580 165.220 ;
        RECT 77.845 164.460 78.015 165.220 ;
        RECT 78.195 164.630 78.525 165.390 ;
        RECT 77.845 164.290 78.510 164.460 ;
        RECT 78.695 164.315 78.965 165.220 ;
        RECT 80.060 164.955 85.405 165.390 ;
        RECT 76.565 163.750 76.760 164.080 ;
        RECT 76.985 163.750 77.240 164.080 ;
        RECT 76.985 163.580 77.155 163.750 ;
        RECT 77.410 163.580 77.580 164.250 ;
        RECT 78.340 164.145 78.510 164.290 ;
        RECT 77.775 163.740 78.105 164.110 ;
        RECT 78.340 163.815 78.625 164.145 ;
        RECT 76.225 163.410 77.155 163.580 ;
        RECT 76.225 163.375 76.400 163.410 ;
        RECT 75.405 163.180 75.685 163.350 ;
        RECT 75.405 163.010 75.680 163.180 ;
        RECT 75.870 163.010 76.400 163.375 ;
        RECT 76.825 162.840 77.155 163.240 ;
        RECT 77.325 163.010 77.580 163.580 ;
        RECT 78.340 163.560 78.510 163.815 ;
        RECT 77.845 163.390 78.510 163.560 ;
        RECT 78.795 163.515 78.965 164.315 ;
        RECT 81.650 163.705 82.000 164.955 ;
        RECT 85.575 164.630 86.090 165.040 ;
        RECT 86.325 164.630 86.495 165.390 ;
        RECT 86.665 165.050 88.695 165.220 ;
        RECT 77.845 163.010 78.015 163.390 ;
        RECT 78.195 162.840 78.525 163.220 ;
        RECT 78.705 163.010 78.965 163.515 ;
        RECT 83.480 163.385 83.820 164.215 ;
        RECT 85.575 163.820 85.915 164.630 ;
        RECT 86.665 164.385 86.835 165.050 ;
        RECT 87.230 164.710 88.355 164.880 ;
        RECT 86.085 164.195 86.835 164.385 ;
        RECT 87.005 164.370 88.015 164.540 ;
        RECT 85.575 163.650 86.805 163.820 ;
        RECT 80.060 162.840 85.405 163.385 ;
        RECT 85.850 163.045 86.095 163.650 ;
        RECT 86.315 162.840 86.825 163.375 ;
        RECT 87.005 163.010 87.195 164.370 ;
        RECT 87.365 164.030 87.640 164.170 ;
        RECT 87.365 163.860 87.645 164.030 ;
        RECT 87.365 163.010 87.640 163.860 ;
        RECT 87.845 163.570 88.015 164.370 ;
        RECT 88.185 163.580 88.355 164.710 ;
        RECT 88.525 164.080 88.695 165.050 ;
        RECT 88.865 164.250 89.035 165.390 ;
        RECT 89.205 164.250 89.540 165.220 ;
        RECT 88.525 163.750 88.720 164.080 ;
        RECT 88.945 163.750 89.200 164.080 ;
        RECT 88.945 163.580 89.115 163.750 ;
        RECT 89.370 163.580 89.540 164.250 ;
        RECT 89.715 164.225 90.005 165.390 ;
        RECT 90.550 165.050 90.805 165.080 ;
        RECT 90.465 164.880 90.805 165.050 ;
        RECT 90.550 164.410 90.805 164.880 ;
        RECT 90.985 164.590 91.270 165.390 ;
        RECT 91.450 164.670 91.780 165.180 ;
        RECT 88.185 163.410 89.115 163.580 ;
        RECT 88.185 163.375 88.360 163.410 ;
        RECT 87.830 163.010 88.360 163.375 ;
        RECT 88.785 162.840 89.115 163.240 ;
        RECT 89.285 163.010 89.540 163.580 ;
        RECT 89.715 162.840 90.005 163.565 ;
        RECT 90.550 163.550 90.730 164.410 ;
        RECT 91.450 164.080 91.700 164.670 ;
        RECT 92.050 164.520 92.220 165.130 ;
        RECT 92.390 164.700 92.720 165.390 ;
        RECT 92.950 164.840 93.190 165.130 ;
        RECT 93.390 165.010 93.810 165.390 ;
        RECT 93.990 164.920 94.620 165.170 ;
        RECT 95.090 165.010 95.420 165.390 ;
        RECT 93.990 164.840 94.160 164.920 ;
        RECT 95.590 164.840 95.760 165.130 ;
        RECT 95.940 165.010 96.320 165.390 ;
        RECT 96.560 165.005 97.390 165.175 ;
        RECT 92.950 164.670 94.160 164.840 ;
        RECT 90.900 163.750 91.700 164.080 ;
        RECT 90.550 163.020 90.805 163.550 ;
        RECT 90.985 162.840 91.270 163.300 ;
        RECT 91.450 163.100 91.700 163.750 ;
        RECT 91.900 164.500 92.220 164.520 ;
        RECT 91.900 164.330 93.820 164.500 ;
        RECT 91.900 163.435 92.090 164.330 ;
        RECT 93.990 164.160 94.160 164.670 ;
        RECT 94.330 164.410 94.850 164.720 ;
        RECT 92.260 163.990 94.160 164.160 ;
        RECT 92.260 163.930 92.590 163.990 ;
        RECT 92.740 163.760 93.070 163.820 ;
        RECT 92.410 163.490 93.070 163.760 ;
        RECT 91.900 163.105 92.220 163.435 ;
        RECT 92.400 162.840 93.060 163.320 ;
        RECT 93.260 163.230 93.430 163.990 ;
        RECT 94.330 163.820 94.510 164.230 ;
        RECT 93.600 163.650 93.930 163.770 ;
        RECT 94.680 163.650 94.850 164.410 ;
        RECT 93.600 163.480 94.850 163.650 ;
        RECT 95.020 164.590 96.390 164.840 ;
        RECT 95.020 163.820 95.210 164.590 ;
        RECT 96.140 164.330 96.390 164.590 ;
        RECT 95.380 164.160 95.630 164.320 ;
        RECT 96.560 164.160 96.730 165.005 ;
        RECT 97.625 164.720 97.795 165.220 ;
        RECT 97.965 164.890 98.295 165.390 ;
        RECT 96.900 164.330 97.400 164.710 ;
        RECT 97.625 164.550 98.320 164.720 ;
        RECT 95.380 163.990 96.730 164.160 ;
        RECT 96.310 163.950 96.730 163.990 ;
        RECT 95.020 163.480 95.440 163.820 ;
        RECT 95.730 163.490 96.140 163.820 ;
        RECT 93.260 163.060 94.110 163.230 ;
        RECT 94.670 162.840 94.990 163.300 ;
        RECT 95.190 163.050 95.440 163.480 ;
        RECT 95.730 162.840 96.140 163.280 ;
        RECT 96.310 163.220 96.480 163.950 ;
        RECT 96.650 163.400 97.000 163.770 ;
        RECT 97.180 163.460 97.400 164.330 ;
        RECT 97.570 163.760 97.980 164.380 ;
        RECT 98.150 163.580 98.320 164.550 ;
        RECT 97.625 163.390 98.320 163.580 ;
        RECT 96.310 163.020 97.325 163.220 ;
        RECT 97.625 163.060 97.795 163.390 ;
        RECT 97.965 162.840 98.295 163.220 ;
        RECT 98.510 163.100 98.735 165.220 ;
        RECT 98.905 164.890 99.235 165.390 ;
        RECT 99.405 164.720 99.575 165.220 ;
        RECT 98.910 164.550 99.575 164.720 ;
        RECT 98.910 163.560 99.140 164.550 ;
        RECT 99.310 163.730 99.660 164.380 ;
        RECT 99.840 164.200 100.095 165.080 ;
        RECT 100.265 164.250 100.570 165.390 ;
        RECT 100.910 165.010 101.240 165.390 ;
        RECT 101.420 164.840 101.590 165.130 ;
        RECT 101.760 164.930 102.010 165.390 ;
        RECT 100.790 164.670 101.590 164.840 ;
        RECT 102.180 164.880 103.050 165.220 ;
        RECT 98.910 163.390 99.575 163.560 ;
        RECT 98.905 162.840 99.235 163.220 ;
        RECT 99.405 163.100 99.575 163.390 ;
        RECT 99.840 163.550 100.050 164.200 ;
        RECT 100.790 164.080 100.960 164.670 ;
        RECT 102.180 164.500 102.350 164.880 ;
        RECT 103.285 164.760 103.455 165.220 ;
        RECT 103.625 164.930 103.995 165.390 ;
        RECT 104.290 164.790 104.460 165.130 ;
        RECT 104.630 164.960 104.960 165.390 ;
        RECT 105.195 164.790 105.365 165.130 ;
        RECT 101.130 164.330 102.350 164.500 ;
        RECT 102.520 164.420 102.980 164.710 ;
        RECT 103.285 164.590 103.845 164.760 ;
        RECT 104.290 164.620 105.365 164.790 ;
        RECT 105.535 164.890 106.215 165.220 ;
        RECT 106.430 164.890 106.680 165.220 ;
        RECT 106.850 164.930 107.100 165.390 ;
        RECT 103.675 164.450 103.845 164.590 ;
        RECT 102.520 164.410 103.485 164.420 ;
        RECT 102.180 164.240 102.350 164.330 ;
        RECT 102.810 164.250 103.485 164.410 ;
        RECT 100.220 164.050 100.960 164.080 ;
        RECT 100.220 163.750 101.135 164.050 ;
        RECT 100.810 163.575 101.135 163.750 ;
        RECT 99.840 163.020 100.095 163.550 ;
        RECT 100.265 162.840 100.570 163.300 ;
        RECT 100.815 163.220 101.135 163.575 ;
        RECT 101.305 163.790 101.845 164.160 ;
        RECT 102.180 164.070 102.585 164.240 ;
        RECT 101.305 163.390 101.545 163.790 ;
        RECT 102.025 163.620 102.245 163.900 ;
        RECT 101.715 163.450 102.245 163.620 ;
        RECT 101.715 163.220 101.885 163.450 ;
        RECT 102.415 163.290 102.585 164.070 ;
        RECT 102.755 163.460 103.105 164.080 ;
        RECT 103.275 163.460 103.485 164.250 ;
        RECT 103.675 164.280 105.175 164.450 ;
        RECT 103.675 163.590 103.845 164.280 ;
        RECT 105.535 164.110 105.705 164.890 ;
        RECT 106.510 164.760 106.680 164.890 ;
        RECT 104.015 163.940 105.705 164.110 ;
        RECT 105.875 164.330 106.340 164.720 ;
        RECT 106.510 164.590 106.905 164.760 ;
        RECT 104.015 163.760 104.185 163.940 ;
        RECT 100.815 163.050 101.885 163.220 ;
        RECT 102.055 162.840 102.245 163.280 ;
        RECT 102.415 163.010 103.365 163.290 ;
        RECT 103.675 163.200 103.935 163.590 ;
        RECT 104.355 163.520 105.145 163.770 ;
        RECT 103.585 163.030 103.935 163.200 ;
        RECT 104.145 162.840 104.475 163.300 ;
        RECT 105.350 163.230 105.520 163.940 ;
        RECT 105.875 163.740 106.045 164.330 ;
        RECT 105.690 163.520 106.045 163.740 ;
        RECT 106.215 163.520 106.565 164.140 ;
        RECT 106.735 163.230 106.905 164.590 ;
        RECT 107.270 164.420 107.595 165.205 ;
        RECT 107.075 163.370 107.535 164.420 ;
        RECT 105.350 163.060 106.205 163.230 ;
        RECT 106.410 163.060 106.905 163.230 ;
        RECT 107.075 162.840 107.405 163.200 ;
        RECT 107.765 163.100 107.935 165.220 ;
        RECT 108.105 164.890 108.435 165.390 ;
        RECT 108.605 164.720 108.860 165.220 ;
        RECT 108.110 164.550 108.860 164.720 ;
        RECT 108.110 163.560 108.340 164.550 ;
        RECT 108.510 163.730 108.860 164.380 ;
        RECT 109.035 164.250 109.420 165.220 ;
        RECT 109.590 164.930 109.915 165.390 ;
        RECT 110.435 164.760 110.715 165.220 ;
        RECT 109.590 164.540 110.715 164.760 ;
        RECT 109.035 163.580 109.315 164.250 ;
        RECT 109.590 164.080 110.040 164.540 ;
        RECT 110.905 164.370 111.305 165.220 ;
        RECT 111.705 164.930 111.975 165.390 ;
        RECT 112.145 164.760 112.430 165.220 ;
        RECT 109.485 163.750 110.040 164.080 ;
        RECT 110.210 163.810 111.305 164.370 ;
        RECT 109.590 163.640 110.040 163.750 ;
        RECT 108.110 163.390 108.860 163.560 ;
        RECT 108.105 162.840 108.435 163.220 ;
        RECT 108.605 163.100 108.860 163.390 ;
        RECT 109.035 163.010 109.420 163.580 ;
        RECT 109.590 163.470 110.715 163.640 ;
        RECT 109.590 162.840 109.915 163.300 ;
        RECT 110.435 163.010 110.715 163.470 ;
        RECT 110.905 163.010 111.305 163.810 ;
        RECT 111.475 164.540 112.430 164.760 ;
        RECT 111.475 163.640 111.685 164.540 ;
        RECT 111.855 163.810 112.545 164.370 ;
        RECT 112.715 164.300 114.385 165.390 ;
        RECT 114.555 164.300 115.765 165.390 ;
        RECT 112.715 163.780 113.465 164.300 ;
        RECT 111.475 163.470 112.430 163.640 ;
        RECT 113.635 163.610 114.385 164.130 ;
        RECT 114.555 163.760 115.075 164.300 ;
        RECT 111.705 162.840 111.975 163.300 ;
        RECT 112.145 163.010 112.430 163.470 ;
        RECT 112.715 162.840 114.385 163.610 ;
        RECT 115.245 163.590 115.765 164.130 ;
        RECT 114.555 162.840 115.765 163.590 ;
        RECT 14.650 162.670 115.850 162.840 ;
        RECT 14.735 161.920 15.945 162.670 ;
        RECT 14.735 161.380 15.255 161.920 ;
        RECT 16.115 161.900 17.785 162.670 ;
        RECT 15.425 161.210 15.945 161.750 ;
        RECT 14.735 160.120 15.945 161.210 ;
        RECT 16.115 161.210 16.865 161.730 ;
        RECT 17.035 161.380 17.785 161.900 ;
        RECT 18.015 161.850 18.225 162.670 ;
        RECT 18.395 161.870 18.725 162.500 ;
        RECT 18.395 161.270 18.645 161.870 ;
        RECT 18.895 161.850 19.125 162.670 ;
        RECT 19.340 161.930 19.595 162.500 ;
        RECT 19.765 162.270 20.095 162.670 ;
        RECT 20.520 162.135 21.050 162.500 ;
        RECT 20.520 162.100 20.695 162.135 ;
        RECT 19.765 161.930 20.695 162.100 ;
        RECT 21.240 161.990 21.515 162.500 ;
        RECT 18.815 161.430 19.145 161.680 ;
        RECT 16.115 160.120 17.785 161.210 ;
        RECT 18.015 160.120 18.225 161.260 ;
        RECT 18.395 160.290 18.725 161.270 ;
        RECT 19.340 161.260 19.510 161.930 ;
        RECT 19.765 161.760 19.935 161.930 ;
        RECT 19.680 161.430 19.935 161.760 ;
        RECT 20.160 161.430 20.355 161.760 ;
        RECT 18.895 160.120 19.125 161.260 ;
        RECT 19.340 160.290 19.675 161.260 ;
        RECT 19.845 160.120 20.015 161.260 ;
        RECT 20.185 160.460 20.355 161.430 ;
        RECT 20.525 160.800 20.695 161.930 ;
        RECT 20.865 161.140 21.035 161.940 ;
        RECT 21.235 161.820 21.515 161.990 ;
        RECT 21.240 161.340 21.515 161.820 ;
        RECT 21.685 161.140 21.875 162.500 ;
        RECT 22.055 162.135 22.565 162.670 ;
        RECT 22.785 161.860 23.030 162.465 ;
        RECT 23.475 161.900 25.145 162.670 ;
        RECT 25.315 161.945 25.605 162.670 ;
        RECT 25.775 161.900 27.445 162.670 ;
        RECT 22.075 161.690 23.305 161.860 ;
        RECT 20.865 160.970 21.875 161.140 ;
        RECT 22.045 161.125 22.795 161.315 ;
        RECT 20.525 160.630 21.650 160.800 ;
        RECT 22.045 160.460 22.215 161.125 ;
        RECT 22.965 160.880 23.305 161.690 ;
        RECT 20.185 160.290 22.215 160.460 ;
        RECT 22.385 160.120 22.555 160.880 ;
        RECT 22.790 160.470 23.305 160.880 ;
        RECT 23.475 161.210 24.225 161.730 ;
        RECT 24.395 161.380 25.145 161.900 ;
        RECT 23.475 160.120 25.145 161.210 ;
        RECT 25.315 160.120 25.605 161.285 ;
        RECT 25.775 161.210 26.525 161.730 ;
        RECT 26.695 161.380 27.445 161.900 ;
        RECT 27.890 161.860 28.135 162.465 ;
        RECT 28.355 162.135 28.865 162.670 ;
        RECT 27.615 161.690 28.845 161.860 ;
        RECT 25.775 160.120 27.445 161.210 ;
        RECT 27.615 160.880 27.955 161.690 ;
        RECT 28.125 161.125 28.875 161.315 ;
        RECT 27.615 160.470 28.130 160.880 ;
        RECT 28.365 160.120 28.535 160.880 ;
        RECT 28.705 160.460 28.875 161.125 ;
        RECT 29.045 161.140 29.235 162.500 ;
        RECT 29.405 161.650 29.680 162.500 ;
        RECT 29.870 162.135 30.400 162.500 ;
        RECT 30.825 162.270 31.155 162.670 ;
        RECT 30.225 162.100 30.400 162.135 ;
        RECT 29.405 161.480 29.685 161.650 ;
        RECT 29.405 161.340 29.680 161.480 ;
        RECT 29.885 161.140 30.055 161.940 ;
        RECT 29.045 160.970 30.055 161.140 ;
        RECT 30.225 161.930 31.155 162.100 ;
        RECT 31.325 161.930 31.580 162.500 ;
        RECT 32.765 162.120 32.935 162.500 ;
        RECT 33.115 162.290 33.445 162.670 ;
        RECT 32.765 161.950 33.430 162.120 ;
        RECT 33.625 161.995 33.885 162.500 ;
        RECT 30.225 160.800 30.395 161.930 ;
        RECT 30.985 161.760 31.155 161.930 ;
        RECT 29.270 160.630 30.395 160.800 ;
        RECT 30.565 161.430 30.760 161.760 ;
        RECT 30.985 161.430 31.240 161.760 ;
        RECT 30.565 160.460 30.735 161.430 ;
        RECT 31.410 161.260 31.580 161.930 ;
        RECT 32.695 161.400 33.025 161.770 ;
        RECT 33.260 161.695 33.430 161.950 ;
        RECT 28.705 160.290 30.735 160.460 ;
        RECT 30.905 160.120 31.075 161.260 ;
        RECT 31.245 160.290 31.580 161.260 ;
        RECT 33.260 161.365 33.545 161.695 ;
        RECT 33.260 161.220 33.430 161.365 ;
        RECT 32.765 161.050 33.430 161.220 ;
        RECT 33.715 161.195 33.885 161.995 ;
        RECT 32.765 160.290 32.935 161.050 ;
        RECT 33.115 160.120 33.445 160.880 ;
        RECT 33.615 160.290 33.885 161.195 ;
        RECT 34.060 161.930 34.315 162.500 ;
        RECT 34.485 162.270 34.815 162.670 ;
        RECT 35.240 162.135 35.770 162.500 ;
        RECT 35.240 162.100 35.415 162.135 ;
        RECT 34.485 161.930 35.415 162.100 ;
        RECT 35.960 161.990 36.235 162.500 ;
        RECT 34.060 161.260 34.230 161.930 ;
        RECT 34.485 161.760 34.655 161.930 ;
        RECT 34.400 161.430 34.655 161.760 ;
        RECT 34.880 161.430 35.075 161.760 ;
        RECT 34.060 160.290 34.395 161.260 ;
        RECT 34.565 160.120 34.735 161.260 ;
        RECT 34.905 160.460 35.075 161.430 ;
        RECT 35.245 160.800 35.415 161.930 ;
        RECT 35.585 161.140 35.755 161.940 ;
        RECT 35.955 161.820 36.235 161.990 ;
        RECT 35.960 161.340 36.235 161.820 ;
        RECT 36.405 161.140 36.595 162.500 ;
        RECT 36.775 162.135 37.285 162.670 ;
        RECT 37.505 161.860 37.750 162.465 ;
        RECT 38.195 161.900 39.865 162.670 ;
        RECT 36.795 161.690 38.025 161.860 ;
        RECT 35.585 160.970 36.595 161.140 ;
        RECT 36.765 161.125 37.515 161.315 ;
        RECT 35.245 160.630 36.370 160.800 ;
        RECT 36.765 160.460 36.935 161.125 ;
        RECT 37.685 160.880 38.025 161.690 ;
        RECT 34.905 160.290 36.935 160.460 ;
        RECT 37.105 160.120 37.275 160.880 ;
        RECT 37.510 160.470 38.025 160.880 ;
        RECT 38.195 161.210 38.945 161.730 ;
        RECT 39.115 161.380 39.865 161.900 ;
        RECT 40.035 161.870 40.375 162.500 ;
        RECT 40.545 161.870 40.795 162.670 ;
        RECT 40.985 162.020 41.315 162.500 ;
        RECT 41.485 162.210 41.710 162.670 ;
        RECT 41.880 162.020 42.210 162.500 ;
        RECT 40.035 161.260 40.210 161.870 ;
        RECT 40.985 161.850 42.210 162.020 ;
        RECT 42.840 161.890 43.340 162.500 ;
        RECT 43.830 162.040 44.115 162.500 ;
        RECT 44.285 162.210 44.555 162.670 ;
        RECT 40.380 161.510 41.075 161.680 ;
        RECT 40.905 161.260 41.075 161.510 ;
        RECT 41.250 161.480 41.670 161.680 ;
        RECT 41.840 161.480 42.170 161.680 ;
        RECT 42.340 161.480 42.670 161.680 ;
        RECT 42.840 161.260 43.010 161.890 ;
        RECT 43.830 161.870 44.785 162.040 ;
        RECT 43.195 161.430 43.545 161.680 ;
        RECT 38.195 160.120 39.865 161.210 ;
        RECT 40.035 160.290 40.375 161.260 ;
        RECT 40.545 160.120 40.715 161.260 ;
        RECT 40.905 161.090 43.340 161.260 ;
        RECT 43.715 161.140 44.405 161.700 ;
        RECT 40.985 160.120 41.235 160.920 ;
        RECT 41.880 160.290 42.210 161.090 ;
        RECT 42.510 160.120 42.840 160.920 ;
        RECT 43.010 160.290 43.340 161.090 ;
        RECT 44.575 160.970 44.785 161.870 ;
        RECT 43.830 160.750 44.785 160.970 ;
        RECT 44.955 161.700 45.355 162.500 ;
        RECT 45.545 162.040 45.825 162.500 ;
        RECT 46.345 162.210 46.670 162.670 ;
        RECT 45.545 161.870 46.670 162.040 ;
        RECT 46.840 161.930 47.225 162.500 ;
        RECT 46.220 161.760 46.670 161.870 ;
        RECT 44.955 161.140 46.050 161.700 ;
        RECT 46.220 161.430 46.775 161.760 ;
        RECT 43.830 160.290 44.115 160.750 ;
        RECT 44.285 160.120 44.555 160.580 ;
        RECT 44.955 160.290 45.355 161.140 ;
        RECT 46.220 160.970 46.670 161.430 ;
        RECT 46.945 161.260 47.225 161.930 ;
        RECT 45.545 160.750 46.670 160.970 ;
        RECT 45.545 160.290 45.825 160.750 ;
        RECT 46.345 160.120 46.670 160.580 ;
        RECT 46.840 160.290 47.225 161.260 ;
        RECT 47.395 161.930 47.780 162.500 ;
        RECT 47.950 162.210 48.275 162.670 ;
        RECT 48.795 162.040 49.075 162.500 ;
        RECT 47.395 161.260 47.675 161.930 ;
        RECT 47.950 161.870 49.075 162.040 ;
        RECT 47.950 161.760 48.400 161.870 ;
        RECT 47.845 161.430 48.400 161.760 ;
        RECT 49.265 161.700 49.665 162.500 ;
        RECT 50.065 162.210 50.335 162.670 ;
        RECT 50.505 162.040 50.790 162.500 ;
        RECT 47.395 160.290 47.780 161.260 ;
        RECT 47.950 160.970 48.400 161.430 ;
        RECT 48.570 161.140 49.665 161.700 ;
        RECT 47.950 160.750 49.075 160.970 ;
        RECT 47.950 160.120 48.275 160.580 ;
        RECT 48.795 160.290 49.075 160.750 ;
        RECT 49.265 160.290 49.665 161.140 ;
        RECT 49.835 161.870 50.790 162.040 ;
        RECT 51.075 161.945 51.365 162.670 ;
        RECT 52.110 162.040 52.395 162.500 ;
        RECT 52.565 162.210 52.835 162.670 ;
        RECT 52.110 161.870 53.065 162.040 ;
        RECT 49.835 160.970 50.045 161.870 ;
        RECT 50.215 161.140 50.905 161.700 ;
        RECT 49.835 160.750 50.790 160.970 ;
        RECT 50.065 160.120 50.335 160.580 ;
        RECT 50.505 160.290 50.790 160.750 ;
        RECT 51.075 160.120 51.365 161.285 ;
        RECT 51.995 161.140 52.685 161.700 ;
        RECT 52.855 160.970 53.065 161.870 ;
        RECT 52.110 160.750 53.065 160.970 ;
        RECT 53.235 161.700 53.635 162.500 ;
        RECT 53.825 162.040 54.105 162.500 ;
        RECT 54.625 162.210 54.950 162.670 ;
        RECT 53.825 161.870 54.950 162.040 ;
        RECT 55.120 161.930 55.505 162.500 ;
        RECT 54.500 161.760 54.950 161.870 ;
        RECT 53.235 161.140 54.330 161.700 ;
        RECT 54.500 161.430 55.055 161.760 ;
        RECT 52.110 160.290 52.395 160.750 ;
        RECT 52.565 160.120 52.835 160.580 ;
        RECT 53.235 160.290 53.635 161.140 ;
        RECT 54.500 160.970 54.950 161.430 ;
        RECT 55.225 161.260 55.505 161.930 ;
        RECT 55.825 161.870 56.155 162.670 ;
        RECT 56.325 162.020 56.495 162.500 ;
        RECT 56.665 162.190 56.995 162.670 ;
        RECT 57.165 162.020 57.335 162.500 ;
        RECT 57.585 162.190 57.825 162.670 ;
        RECT 58.005 162.020 58.175 162.500 ;
        RECT 56.325 161.850 57.335 162.020 ;
        RECT 57.540 161.850 58.175 162.020 ;
        RECT 56.325 161.310 56.820 161.850 ;
        RECT 57.540 161.680 57.710 161.850 ;
        RECT 59.360 161.830 59.620 162.670 ;
        RECT 59.795 161.925 60.050 162.500 ;
        RECT 60.220 162.290 60.550 162.670 ;
        RECT 60.765 162.120 60.935 162.500 ;
        RECT 60.220 161.950 60.935 162.120 ;
        RECT 57.210 161.510 57.710 161.680 ;
        RECT 53.825 160.750 54.950 160.970 ;
        RECT 53.825 160.290 54.105 160.750 ;
        RECT 54.625 160.120 54.950 160.580 ;
        RECT 55.120 160.290 55.505 161.260 ;
        RECT 55.825 160.120 56.155 161.270 ;
        RECT 56.325 161.140 57.335 161.310 ;
        RECT 56.325 160.290 56.495 161.140 ;
        RECT 56.665 160.120 56.995 160.920 ;
        RECT 57.165 160.290 57.335 161.140 ;
        RECT 57.540 161.270 57.710 161.510 ;
        RECT 57.880 161.440 58.260 161.680 ;
        RECT 57.540 161.100 58.255 161.270 ;
        RECT 57.515 160.120 57.755 160.920 ;
        RECT 57.925 160.290 58.255 161.100 ;
        RECT 59.360 160.120 59.620 161.270 ;
        RECT 59.795 161.195 59.965 161.925 ;
        RECT 60.220 161.760 60.390 161.950 ;
        RECT 61.200 161.830 61.460 162.670 ;
        RECT 61.635 161.925 61.890 162.500 ;
        RECT 62.060 162.290 62.390 162.670 ;
        RECT 62.605 162.120 62.775 162.500 ;
        RECT 62.060 161.950 62.775 162.120 ;
        RECT 63.125 162.120 63.295 162.500 ;
        RECT 63.510 162.290 63.840 162.670 ;
        RECT 63.125 161.950 63.840 162.120 ;
        RECT 60.135 161.430 60.390 161.760 ;
        RECT 60.220 161.220 60.390 161.430 ;
        RECT 60.670 161.400 61.025 161.770 ;
        RECT 59.795 160.290 60.050 161.195 ;
        RECT 60.220 161.050 60.935 161.220 ;
        RECT 60.220 160.120 60.550 160.880 ;
        RECT 60.765 160.290 60.935 161.050 ;
        RECT 61.200 160.120 61.460 161.270 ;
        RECT 61.635 161.195 61.805 161.925 ;
        RECT 62.060 161.760 62.230 161.950 ;
        RECT 61.975 161.430 62.230 161.760 ;
        RECT 62.060 161.220 62.230 161.430 ;
        RECT 62.510 161.400 62.865 161.770 ;
        RECT 63.035 161.400 63.390 161.770 ;
        RECT 63.670 161.760 63.840 161.950 ;
        RECT 64.010 161.925 64.265 162.500 ;
        RECT 63.670 161.430 63.925 161.760 ;
        RECT 63.670 161.220 63.840 161.430 ;
        RECT 61.635 160.290 61.890 161.195 ;
        RECT 62.060 161.050 62.775 161.220 ;
        RECT 62.060 160.120 62.390 160.880 ;
        RECT 62.605 160.290 62.775 161.050 ;
        RECT 63.125 161.050 63.840 161.220 ;
        RECT 64.095 161.195 64.265 161.925 ;
        RECT 64.440 161.830 64.700 162.670 ;
        RECT 65.340 161.830 65.600 162.670 ;
        RECT 65.775 161.925 66.030 162.500 ;
        RECT 66.200 162.290 66.530 162.670 ;
        RECT 66.745 162.120 66.915 162.500 ;
        RECT 66.200 161.950 66.915 162.120 ;
        RECT 67.265 162.120 67.435 162.500 ;
        RECT 67.650 162.290 67.980 162.670 ;
        RECT 67.265 161.950 67.980 162.120 ;
        RECT 63.125 160.290 63.295 161.050 ;
        RECT 63.510 160.120 63.840 160.880 ;
        RECT 64.010 160.290 64.265 161.195 ;
        RECT 64.440 160.120 64.700 161.270 ;
        RECT 65.340 160.120 65.600 161.270 ;
        RECT 65.775 161.195 65.945 161.925 ;
        RECT 66.200 161.760 66.370 161.950 ;
        RECT 66.115 161.430 66.370 161.760 ;
        RECT 66.200 161.220 66.370 161.430 ;
        RECT 66.650 161.400 67.005 161.770 ;
        RECT 67.175 161.400 67.530 161.770 ;
        RECT 67.810 161.760 67.980 161.950 ;
        RECT 68.150 161.925 68.405 162.500 ;
        RECT 67.810 161.430 68.065 161.760 ;
        RECT 67.810 161.220 67.980 161.430 ;
        RECT 65.775 160.290 66.030 161.195 ;
        RECT 66.200 161.050 66.915 161.220 ;
        RECT 66.200 160.120 66.530 160.880 ;
        RECT 66.745 160.290 66.915 161.050 ;
        RECT 67.265 161.050 67.980 161.220 ;
        RECT 68.235 161.195 68.405 161.925 ;
        RECT 68.580 161.830 68.840 162.670 ;
        RECT 69.015 161.870 69.355 162.500 ;
        RECT 69.525 161.870 69.775 162.670 ;
        RECT 69.965 162.020 70.295 162.500 ;
        RECT 70.465 162.210 70.690 162.670 ;
        RECT 70.860 162.020 71.190 162.500 ;
        RECT 67.265 160.290 67.435 161.050 ;
        RECT 67.650 160.120 67.980 160.880 ;
        RECT 68.150 160.290 68.405 161.195 ;
        RECT 68.580 160.120 68.840 161.270 ;
        RECT 69.015 161.260 69.190 161.870 ;
        RECT 69.965 161.850 71.190 162.020 ;
        RECT 71.820 161.890 72.320 162.500 ;
        RECT 69.360 161.510 70.055 161.680 ;
        RECT 69.885 161.260 70.055 161.510 ;
        RECT 70.230 161.480 70.650 161.680 ;
        RECT 70.820 161.480 71.150 161.680 ;
        RECT 71.320 161.480 71.650 161.680 ;
        RECT 71.820 161.260 71.990 161.890 ;
        RECT 72.970 161.860 73.215 162.465 ;
        RECT 73.435 162.135 73.945 162.670 ;
        RECT 72.695 161.690 73.925 161.860 ;
        RECT 72.175 161.430 72.525 161.680 ;
        RECT 69.015 160.290 69.355 161.260 ;
        RECT 69.525 160.120 69.695 161.260 ;
        RECT 69.885 161.090 72.320 161.260 ;
        RECT 69.965 160.120 70.215 160.920 ;
        RECT 70.860 160.290 71.190 161.090 ;
        RECT 71.490 160.120 71.820 160.920 ;
        RECT 71.990 160.290 72.320 161.090 ;
        RECT 72.695 160.880 73.035 161.690 ;
        RECT 73.205 161.125 73.955 161.315 ;
        RECT 72.695 160.470 73.210 160.880 ;
        RECT 73.445 160.120 73.615 160.880 ;
        RECT 73.785 160.460 73.955 161.125 ;
        RECT 74.125 161.140 74.315 162.500 ;
        RECT 74.485 161.990 74.760 162.500 ;
        RECT 74.950 162.135 75.480 162.500 ;
        RECT 75.905 162.270 76.235 162.670 ;
        RECT 75.305 162.100 75.480 162.135 ;
        RECT 74.485 161.820 74.765 161.990 ;
        RECT 74.485 161.340 74.760 161.820 ;
        RECT 74.965 161.140 75.135 161.940 ;
        RECT 74.125 160.970 75.135 161.140 ;
        RECT 75.305 161.930 76.235 162.100 ;
        RECT 76.405 161.930 76.660 162.500 ;
        RECT 76.835 161.945 77.125 162.670 ;
        RECT 75.305 160.800 75.475 161.930 ;
        RECT 76.065 161.760 76.235 161.930 ;
        RECT 74.350 160.630 75.475 160.800 ;
        RECT 75.645 161.430 75.840 161.760 ;
        RECT 76.065 161.430 76.320 161.760 ;
        RECT 75.645 160.460 75.815 161.430 ;
        RECT 76.490 161.260 76.660 161.930 ;
        RECT 77.295 161.900 78.965 162.670 ;
        RECT 73.785 160.290 75.815 160.460 ;
        RECT 75.985 160.120 76.155 161.260 ;
        RECT 76.325 160.290 76.660 161.260 ;
        RECT 76.835 160.120 77.125 161.285 ;
        RECT 77.295 161.210 78.045 161.730 ;
        RECT 78.215 161.380 78.965 161.900 ;
        RECT 79.195 161.850 79.405 162.670 ;
        RECT 79.575 161.870 79.905 162.500 ;
        RECT 79.575 161.270 79.825 161.870 ;
        RECT 80.075 161.850 80.305 162.670 ;
        RECT 80.605 162.120 80.775 162.500 ;
        RECT 80.955 162.290 81.285 162.670 ;
        RECT 80.605 161.950 81.270 162.120 ;
        RECT 81.465 161.995 81.725 162.500 ;
        RECT 79.995 161.430 80.325 161.680 ;
        RECT 80.535 161.400 80.865 161.770 ;
        RECT 81.100 161.695 81.270 161.950 ;
        RECT 81.100 161.365 81.385 161.695 ;
        RECT 77.295 160.120 78.965 161.210 ;
        RECT 79.195 160.120 79.405 161.260 ;
        RECT 79.575 160.290 79.905 161.270 ;
        RECT 80.075 160.120 80.305 161.260 ;
        RECT 81.100 161.220 81.270 161.365 ;
        RECT 80.605 161.050 81.270 161.220 ;
        RECT 81.555 161.195 81.725 161.995 ;
        RECT 83.190 161.990 83.445 162.490 ;
        RECT 83.625 162.210 83.910 162.670 ;
        RECT 83.105 161.960 83.445 161.990 ;
        RECT 83.105 161.820 83.370 161.960 ;
        RECT 80.605 160.290 80.775 161.050 ;
        RECT 80.955 160.120 81.285 160.880 ;
        RECT 81.455 160.290 81.725 161.195 ;
        RECT 83.190 161.100 83.370 161.820 ;
        RECT 84.090 161.760 84.340 162.410 ;
        RECT 83.540 161.430 84.340 161.760 ;
        RECT 83.190 160.430 83.445 161.100 ;
        RECT 83.625 160.120 83.910 160.920 ;
        RECT 84.090 160.840 84.340 161.430 ;
        RECT 84.540 162.075 84.860 162.405 ;
        RECT 85.040 162.190 85.700 162.670 ;
        RECT 85.900 162.280 86.750 162.450 ;
        RECT 84.540 161.180 84.730 162.075 ;
        RECT 85.050 161.750 85.710 162.020 ;
        RECT 85.380 161.690 85.710 161.750 ;
        RECT 84.900 161.520 85.230 161.580 ;
        RECT 85.900 161.520 86.070 162.280 ;
        RECT 87.310 162.210 87.630 162.670 ;
        RECT 87.830 162.030 88.080 162.460 ;
        RECT 88.370 162.230 88.780 162.670 ;
        RECT 88.950 162.290 89.965 162.490 ;
        RECT 86.240 161.860 87.490 162.030 ;
        RECT 86.240 161.740 86.570 161.860 ;
        RECT 84.900 161.350 86.800 161.520 ;
        RECT 84.540 161.010 86.460 161.180 ;
        RECT 84.540 160.990 84.860 161.010 ;
        RECT 84.090 160.330 84.420 160.840 ;
        RECT 84.690 160.380 84.860 160.990 ;
        RECT 86.630 160.840 86.800 161.350 ;
        RECT 86.970 161.280 87.150 161.690 ;
        RECT 87.320 161.100 87.490 161.860 ;
        RECT 85.030 160.120 85.360 160.810 ;
        RECT 85.590 160.670 86.800 160.840 ;
        RECT 86.970 160.790 87.490 161.100 ;
        RECT 87.660 161.690 88.080 162.030 ;
        RECT 88.370 161.690 88.780 162.020 ;
        RECT 87.660 160.920 87.850 161.690 ;
        RECT 88.950 161.560 89.120 162.290 ;
        RECT 90.265 162.120 90.435 162.450 ;
        RECT 90.605 162.290 90.935 162.670 ;
        RECT 89.290 161.740 89.640 162.110 ;
        RECT 88.950 161.520 89.370 161.560 ;
        RECT 88.020 161.350 89.370 161.520 ;
        RECT 88.020 161.190 88.270 161.350 ;
        RECT 88.780 160.920 89.030 161.180 ;
        RECT 87.660 160.670 89.030 160.920 ;
        RECT 85.590 160.380 85.830 160.670 ;
        RECT 86.630 160.590 86.800 160.670 ;
        RECT 86.030 160.120 86.450 160.500 ;
        RECT 86.630 160.340 87.260 160.590 ;
        RECT 87.730 160.120 88.060 160.500 ;
        RECT 88.230 160.380 88.400 160.670 ;
        RECT 89.200 160.505 89.370 161.350 ;
        RECT 89.820 161.180 90.040 162.050 ;
        RECT 90.265 161.930 90.960 162.120 ;
        RECT 89.540 160.800 90.040 161.180 ;
        RECT 90.210 161.130 90.620 161.750 ;
        RECT 90.790 160.960 90.960 161.930 ;
        RECT 90.265 160.790 90.960 160.960 ;
        RECT 88.580 160.120 88.960 160.500 ;
        RECT 89.200 160.335 90.030 160.505 ;
        RECT 90.265 160.290 90.435 160.790 ;
        RECT 90.605 160.120 90.935 160.620 ;
        RECT 91.150 160.290 91.375 162.410 ;
        RECT 91.545 162.290 91.875 162.670 ;
        RECT 92.045 162.120 92.215 162.410 ;
        RECT 91.550 161.950 92.215 162.120 ;
        RECT 92.475 161.995 92.735 162.500 ;
        RECT 92.915 162.290 93.245 162.670 ;
        RECT 93.425 162.120 93.595 162.500 ;
        RECT 91.550 160.960 91.780 161.950 ;
        RECT 91.950 161.130 92.300 161.780 ;
        RECT 92.475 161.195 92.645 161.995 ;
        RECT 92.930 161.950 93.595 162.120 ;
        RECT 92.930 161.695 93.100 161.950 ;
        RECT 94.775 161.930 95.160 162.500 ;
        RECT 95.330 162.210 95.655 162.670 ;
        RECT 96.175 162.040 96.455 162.500 ;
        RECT 92.815 161.365 93.100 161.695 ;
        RECT 93.335 161.400 93.665 161.770 ;
        RECT 92.930 161.220 93.100 161.365 ;
        RECT 94.775 161.260 95.055 161.930 ;
        RECT 95.330 161.870 96.455 162.040 ;
        RECT 95.330 161.760 95.780 161.870 ;
        RECT 95.225 161.430 95.780 161.760 ;
        RECT 96.645 161.700 97.045 162.500 ;
        RECT 97.445 162.210 97.715 162.670 ;
        RECT 97.885 162.040 98.170 162.500 ;
        RECT 91.550 160.790 92.215 160.960 ;
        RECT 91.545 160.120 91.875 160.620 ;
        RECT 92.045 160.290 92.215 160.790 ;
        RECT 92.475 160.290 92.745 161.195 ;
        RECT 92.930 161.050 93.595 161.220 ;
        RECT 92.915 160.120 93.245 160.880 ;
        RECT 93.425 160.290 93.595 161.050 ;
        RECT 94.775 160.290 95.160 161.260 ;
        RECT 95.330 160.970 95.780 161.430 ;
        RECT 95.950 161.140 97.045 161.700 ;
        RECT 95.330 160.750 96.455 160.970 ;
        RECT 95.330 160.120 95.655 160.580 ;
        RECT 96.175 160.290 96.455 160.750 ;
        RECT 96.645 160.290 97.045 161.140 ;
        RECT 97.215 161.870 98.170 162.040 ;
        RECT 98.660 161.890 99.160 162.500 ;
        RECT 97.215 160.970 97.425 161.870 ;
        RECT 97.595 161.140 98.285 161.700 ;
        RECT 98.455 161.430 98.805 161.680 ;
        RECT 98.990 161.260 99.160 161.890 ;
        RECT 99.790 162.020 100.120 162.500 ;
        RECT 100.290 162.210 100.515 162.670 ;
        RECT 100.685 162.020 101.015 162.500 ;
        RECT 99.790 161.850 101.015 162.020 ;
        RECT 101.205 161.870 101.455 162.670 ;
        RECT 101.625 161.870 101.965 162.500 ;
        RECT 102.595 161.945 102.885 162.670 ;
        RECT 99.330 161.480 99.660 161.680 ;
        RECT 99.830 161.480 100.160 161.680 ;
        RECT 100.330 161.480 100.750 161.680 ;
        RECT 100.925 161.510 101.620 161.680 ;
        RECT 100.925 161.260 101.095 161.510 ;
        RECT 101.790 161.260 101.965 161.870 ;
        RECT 104.250 161.860 104.495 162.465 ;
        RECT 104.715 162.135 105.225 162.670 ;
        RECT 103.975 161.690 105.205 161.860 ;
        RECT 98.660 161.090 101.095 161.260 ;
        RECT 97.215 160.750 98.170 160.970 ;
        RECT 97.445 160.120 97.715 160.580 ;
        RECT 97.885 160.290 98.170 160.750 ;
        RECT 98.660 160.290 98.990 161.090 ;
        RECT 99.160 160.120 99.490 160.920 ;
        RECT 99.790 160.290 100.120 161.090 ;
        RECT 100.765 160.120 101.015 160.920 ;
        RECT 101.285 160.120 101.455 161.260 ;
        RECT 101.625 160.290 101.965 161.260 ;
        RECT 102.595 160.120 102.885 161.285 ;
        RECT 103.975 160.880 104.315 161.690 ;
        RECT 104.485 161.125 105.235 161.315 ;
        RECT 103.975 160.470 104.490 160.880 ;
        RECT 104.725 160.120 104.895 160.880 ;
        RECT 105.065 160.460 105.235 161.125 ;
        RECT 105.405 161.140 105.595 162.500 ;
        RECT 105.765 161.650 106.040 162.500 ;
        RECT 106.230 162.135 106.760 162.500 ;
        RECT 107.185 162.270 107.515 162.670 ;
        RECT 106.585 162.100 106.760 162.135 ;
        RECT 105.765 161.480 106.045 161.650 ;
        RECT 105.765 161.340 106.040 161.480 ;
        RECT 106.245 161.140 106.415 161.940 ;
        RECT 105.405 160.970 106.415 161.140 ;
        RECT 106.585 161.930 107.515 162.100 ;
        RECT 107.685 161.930 107.940 162.500 ;
        RECT 106.585 160.800 106.755 161.930 ;
        RECT 107.345 161.760 107.515 161.930 ;
        RECT 105.630 160.630 106.755 160.800 ;
        RECT 106.925 161.430 107.120 161.760 ;
        RECT 107.345 161.430 107.600 161.760 ;
        RECT 106.925 160.460 107.095 161.430 ;
        RECT 107.770 161.260 107.940 161.930 ;
        RECT 109.185 161.870 109.515 162.670 ;
        RECT 109.685 162.020 109.855 162.500 ;
        RECT 110.025 162.190 110.355 162.670 ;
        RECT 110.525 162.020 110.695 162.500 ;
        RECT 110.945 162.190 111.185 162.670 ;
        RECT 111.365 162.020 111.535 162.500 ;
        RECT 109.685 161.850 110.695 162.020 ;
        RECT 110.900 161.850 111.535 162.020 ;
        RECT 111.885 162.120 112.055 162.500 ;
        RECT 112.235 162.290 112.565 162.670 ;
        RECT 111.885 161.950 112.550 162.120 ;
        RECT 112.745 161.995 113.005 162.500 ;
        RECT 109.685 161.820 110.185 161.850 ;
        RECT 109.685 161.310 110.180 161.820 ;
        RECT 110.900 161.680 111.070 161.850 ;
        RECT 110.570 161.510 111.070 161.680 ;
        RECT 105.065 160.290 107.095 160.460 ;
        RECT 107.265 160.120 107.435 161.260 ;
        RECT 107.605 160.290 107.940 161.260 ;
        RECT 109.185 160.120 109.515 161.270 ;
        RECT 109.685 161.140 110.695 161.310 ;
        RECT 109.685 160.290 109.855 161.140 ;
        RECT 110.025 160.120 110.355 160.920 ;
        RECT 110.525 160.290 110.695 161.140 ;
        RECT 110.900 161.270 111.070 161.510 ;
        RECT 111.240 161.440 111.620 161.680 ;
        RECT 111.815 161.400 112.145 161.770 ;
        RECT 112.380 161.695 112.550 161.950 ;
        RECT 112.380 161.365 112.665 161.695 ;
        RECT 110.900 161.100 111.615 161.270 ;
        RECT 112.380 161.220 112.550 161.365 ;
        RECT 110.875 160.120 111.115 160.920 ;
        RECT 111.285 160.290 111.615 161.100 ;
        RECT 111.885 161.050 112.550 161.220 ;
        RECT 112.835 161.195 113.005 161.995 ;
        RECT 113.175 161.920 114.385 162.670 ;
        RECT 114.555 161.920 115.765 162.670 ;
        RECT 111.885 160.290 112.055 161.050 ;
        RECT 112.235 160.120 112.565 160.880 ;
        RECT 112.735 160.290 113.005 161.195 ;
        RECT 113.175 161.210 113.695 161.750 ;
        RECT 113.865 161.380 114.385 161.920 ;
        RECT 114.555 161.210 115.075 161.750 ;
        RECT 115.245 161.380 115.765 161.920 ;
        RECT 113.175 160.120 114.385 161.210 ;
        RECT 114.555 160.120 115.765 161.210 ;
        RECT 14.650 159.950 115.850 160.120 ;
        RECT 14.735 158.860 15.945 159.950 ;
        RECT 16.950 158.970 17.205 159.640 ;
        RECT 17.385 159.150 17.670 159.950 ;
        RECT 17.850 159.230 18.180 159.740 ;
        RECT 16.950 158.930 17.130 158.970 ;
        RECT 14.735 158.150 15.255 158.690 ;
        RECT 15.425 158.320 15.945 158.860 ;
        RECT 16.865 158.760 17.130 158.930 ;
        RECT 14.735 157.400 15.945 158.150 ;
        RECT 16.950 158.110 17.130 158.760 ;
        RECT 17.850 158.640 18.100 159.230 ;
        RECT 18.450 159.080 18.620 159.690 ;
        RECT 18.790 159.260 19.120 159.950 ;
        RECT 19.350 159.400 19.590 159.690 ;
        RECT 19.790 159.570 20.210 159.950 ;
        RECT 20.390 159.480 21.020 159.730 ;
        RECT 21.490 159.570 21.820 159.950 ;
        RECT 20.390 159.400 20.560 159.480 ;
        RECT 21.990 159.400 22.160 159.690 ;
        RECT 22.340 159.570 22.720 159.950 ;
        RECT 22.960 159.565 23.790 159.735 ;
        RECT 19.350 159.230 20.560 159.400 ;
        RECT 17.300 158.310 18.100 158.640 ;
        RECT 16.950 157.580 17.205 158.110 ;
        RECT 17.385 157.400 17.670 157.860 ;
        RECT 17.850 157.660 18.100 158.310 ;
        RECT 18.300 159.060 18.620 159.080 ;
        RECT 18.300 158.890 20.220 159.060 ;
        RECT 18.300 157.995 18.490 158.890 ;
        RECT 20.390 158.720 20.560 159.230 ;
        RECT 20.730 158.970 21.250 159.280 ;
        RECT 18.660 158.550 20.560 158.720 ;
        RECT 18.660 158.490 18.990 158.550 ;
        RECT 19.140 158.320 19.470 158.380 ;
        RECT 18.810 158.050 19.470 158.320 ;
        RECT 18.300 157.665 18.620 157.995 ;
        RECT 18.800 157.400 19.460 157.880 ;
        RECT 19.660 157.790 19.830 158.550 ;
        RECT 20.730 158.380 20.910 158.790 ;
        RECT 20.000 158.210 20.330 158.330 ;
        RECT 21.080 158.210 21.250 158.970 ;
        RECT 20.000 158.040 21.250 158.210 ;
        RECT 21.420 159.150 22.790 159.400 ;
        RECT 21.420 158.380 21.610 159.150 ;
        RECT 22.540 158.890 22.790 159.150 ;
        RECT 21.780 158.720 22.030 158.880 ;
        RECT 22.960 158.720 23.130 159.565 ;
        RECT 24.025 159.280 24.195 159.780 ;
        RECT 24.365 159.450 24.695 159.950 ;
        RECT 23.300 158.890 23.800 159.270 ;
        RECT 24.025 159.110 24.720 159.280 ;
        RECT 21.780 158.550 23.130 158.720 ;
        RECT 22.710 158.510 23.130 158.550 ;
        RECT 21.420 158.040 21.840 158.380 ;
        RECT 22.130 158.050 22.540 158.380 ;
        RECT 19.660 157.620 20.510 157.790 ;
        RECT 21.070 157.400 21.390 157.860 ;
        RECT 21.590 157.610 21.840 158.040 ;
        RECT 22.130 157.400 22.540 157.840 ;
        RECT 22.710 157.780 22.880 158.510 ;
        RECT 23.050 157.960 23.400 158.330 ;
        RECT 23.580 158.020 23.800 158.890 ;
        RECT 23.970 158.320 24.380 158.940 ;
        RECT 24.550 158.140 24.720 159.110 ;
        RECT 24.025 157.950 24.720 158.140 ;
        RECT 22.710 157.580 23.725 157.780 ;
        RECT 24.025 157.620 24.195 157.950 ;
        RECT 24.365 157.400 24.695 157.780 ;
        RECT 24.910 157.660 25.135 159.780 ;
        RECT 25.305 159.450 25.635 159.950 ;
        RECT 25.805 159.280 25.975 159.780 ;
        RECT 25.310 159.110 25.975 159.280 ;
        RECT 25.310 158.120 25.540 159.110 ;
        RECT 25.710 158.290 26.060 158.940 ;
        RECT 27.195 158.810 27.425 159.950 ;
        RECT 27.595 158.800 27.925 159.780 ;
        RECT 28.095 158.810 28.305 159.950 ;
        RECT 28.910 159.610 29.165 159.640 ;
        RECT 28.825 159.440 29.165 159.610 ;
        RECT 28.910 158.970 29.165 159.440 ;
        RECT 29.345 159.150 29.630 159.950 ;
        RECT 29.810 159.230 30.140 159.740 ;
        RECT 27.175 158.390 27.505 158.640 ;
        RECT 25.310 157.950 25.975 158.120 ;
        RECT 25.305 157.400 25.635 157.780 ;
        RECT 25.805 157.660 25.975 157.950 ;
        RECT 27.195 157.400 27.425 158.220 ;
        RECT 27.675 158.200 27.925 158.800 ;
        RECT 27.595 157.570 27.925 158.200 ;
        RECT 28.095 157.400 28.305 158.220 ;
        RECT 28.910 158.110 29.090 158.970 ;
        RECT 29.810 158.640 30.060 159.230 ;
        RECT 30.410 159.080 30.580 159.690 ;
        RECT 30.750 159.260 31.080 159.950 ;
        RECT 31.310 159.400 31.550 159.690 ;
        RECT 31.750 159.570 32.170 159.950 ;
        RECT 32.350 159.480 32.980 159.730 ;
        RECT 33.450 159.570 33.780 159.950 ;
        RECT 32.350 159.400 32.520 159.480 ;
        RECT 33.950 159.400 34.120 159.690 ;
        RECT 34.300 159.570 34.680 159.950 ;
        RECT 34.920 159.565 35.750 159.735 ;
        RECT 31.310 159.230 32.520 159.400 ;
        RECT 29.260 158.310 30.060 158.640 ;
        RECT 28.910 157.580 29.165 158.110 ;
        RECT 29.345 157.400 29.630 157.860 ;
        RECT 29.810 157.660 30.060 158.310 ;
        RECT 30.260 159.060 30.580 159.080 ;
        RECT 30.260 158.890 32.180 159.060 ;
        RECT 30.260 157.995 30.450 158.890 ;
        RECT 32.350 158.720 32.520 159.230 ;
        RECT 32.690 158.970 33.210 159.280 ;
        RECT 30.620 158.550 32.520 158.720 ;
        RECT 30.620 158.490 30.950 158.550 ;
        RECT 31.100 158.320 31.430 158.380 ;
        RECT 30.770 158.050 31.430 158.320 ;
        RECT 30.260 157.665 30.580 157.995 ;
        RECT 30.760 157.400 31.420 157.880 ;
        RECT 31.620 157.790 31.790 158.550 ;
        RECT 32.690 158.380 32.870 158.790 ;
        RECT 31.960 158.210 32.290 158.330 ;
        RECT 33.040 158.210 33.210 158.970 ;
        RECT 31.960 158.040 33.210 158.210 ;
        RECT 33.380 159.150 34.750 159.400 ;
        RECT 33.380 158.380 33.570 159.150 ;
        RECT 34.500 158.890 34.750 159.150 ;
        RECT 33.740 158.720 33.990 158.880 ;
        RECT 34.920 158.720 35.090 159.565 ;
        RECT 35.985 159.280 36.155 159.780 ;
        RECT 36.325 159.450 36.655 159.950 ;
        RECT 35.260 158.890 35.760 159.270 ;
        RECT 35.985 159.110 36.680 159.280 ;
        RECT 33.740 158.550 35.090 158.720 ;
        RECT 34.670 158.510 35.090 158.550 ;
        RECT 33.380 158.040 33.800 158.380 ;
        RECT 34.090 158.050 34.500 158.380 ;
        RECT 31.620 157.620 32.470 157.790 ;
        RECT 33.030 157.400 33.350 157.860 ;
        RECT 33.550 157.610 33.800 158.040 ;
        RECT 34.090 157.400 34.500 157.840 ;
        RECT 34.670 157.780 34.840 158.510 ;
        RECT 35.010 157.960 35.360 158.330 ;
        RECT 35.540 158.020 35.760 158.890 ;
        RECT 35.930 158.320 36.340 158.940 ;
        RECT 36.510 158.140 36.680 159.110 ;
        RECT 35.985 157.950 36.680 158.140 ;
        RECT 34.670 157.580 35.685 157.780 ;
        RECT 35.985 157.620 36.155 157.950 ;
        RECT 36.325 157.400 36.655 157.780 ;
        RECT 36.870 157.660 37.095 159.780 ;
        RECT 37.265 159.450 37.595 159.950 ;
        RECT 37.765 159.280 37.935 159.780 ;
        RECT 37.270 159.110 37.935 159.280 ;
        RECT 37.270 158.120 37.500 159.110 ;
        RECT 37.670 158.290 38.020 158.940 ;
        RECT 38.195 158.785 38.485 159.950 ;
        RECT 39.115 158.860 41.705 159.950 ;
        RECT 39.115 158.340 40.325 158.860 ;
        RECT 41.875 158.810 42.215 159.780 ;
        RECT 42.385 158.810 42.555 159.950 ;
        RECT 42.825 159.150 43.075 159.950 ;
        RECT 43.720 158.980 44.050 159.780 ;
        RECT 44.350 159.150 44.680 159.950 ;
        RECT 44.850 158.980 45.180 159.780 ;
        RECT 42.745 158.810 45.180 158.980 ;
        RECT 45.555 158.810 45.895 159.780 ;
        RECT 46.065 158.810 46.235 159.950 ;
        RECT 46.505 159.150 46.755 159.950 ;
        RECT 47.400 158.980 47.730 159.780 ;
        RECT 48.030 159.150 48.360 159.950 ;
        RECT 48.530 158.980 48.860 159.780 ;
        RECT 46.425 158.810 48.860 158.980 ;
        RECT 49.235 158.810 49.575 159.780 ;
        RECT 49.745 158.810 49.915 159.950 ;
        RECT 50.185 159.150 50.435 159.950 ;
        RECT 51.080 158.980 51.410 159.780 ;
        RECT 51.710 159.150 52.040 159.950 ;
        RECT 52.210 158.980 52.540 159.780 ;
        RECT 50.105 158.810 52.540 158.980 ;
        RECT 52.915 158.860 54.585 159.950 ;
        RECT 54.845 159.205 55.115 159.950 ;
        RECT 55.745 159.945 62.020 159.950 ;
        RECT 55.285 159.035 55.575 159.775 ;
        RECT 55.745 159.220 56.000 159.945 ;
        RECT 56.185 159.050 56.445 159.775 ;
        RECT 56.615 159.220 56.860 159.945 ;
        RECT 57.045 159.050 57.305 159.775 ;
        RECT 57.475 159.220 57.720 159.945 ;
        RECT 57.905 159.050 58.165 159.775 ;
        RECT 58.335 159.220 58.580 159.945 ;
        RECT 58.750 159.050 59.010 159.775 ;
        RECT 59.180 159.220 59.440 159.945 ;
        RECT 59.610 159.050 59.870 159.775 ;
        RECT 60.040 159.220 60.300 159.945 ;
        RECT 60.470 159.050 60.730 159.775 ;
        RECT 60.900 159.220 61.160 159.945 ;
        RECT 61.330 159.050 61.590 159.775 ;
        RECT 61.760 159.150 62.020 159.945 ;
        RECT 56.185 159.035 61.590 159.050 ;
        RECT 54.845 158.930 61.590 159.035 ;
        RECT 40.495 158.170 41.705 158.690 ;
        RECT 37.270 157.950 37.935 158.120 ;
        RECT 37.265 157.400 37.595 157.780 ;
        RECT 37.765 157.660 37.935 157.950 ;
        RECT 38.195 157.400 38.485 158.125 ;
        RECT 39.115 157.400 41.705 158.170 ;
        RECT 41.875 158.200 42.050 158.810 ;
        RECT 42.745 158.560 42.915 158.810 ;
        RECT 42.220 158.390 42.915 158.560 ;
        RECT 43.090 158.390 43.510 158.590 ;
        RECT 43.680 158.390 44.010 158.590 ;
        RECT 44.180 158.390 44.510 158.590 ;
        RECT 41.875 157.570 42.215 158.200 ;
        RECT 42.385 157.400 42.635 158.200 ;
        RECT 42.825 158.050 44.050 158.220 ;
        RECT 42.825 157.570 43.155 158.050 ;
        RECT 43.325 157.400 43.550 157.860 ;
        RECT 43.720 157.570 44.050 158.050 ;
        RECT 44.680 158.180 44.850 158.810 ;
        RECT 45.035 158.390 45.385 158.640 ;
        RECT 45.555 158.200 45.730 158.810 ;
        RECT 46.425 158.560 46.595 158.810 ;
        RECT 45.900 158.390 46.595 158.560 ;
        RECT 46.770 158.390 47.190 158.590 ;
        RECT 47.360 158.390 47.690 158.590 ;
        RECT 47.860 158.390 48.190 158.590 ;
        RECT 44.680 157.570 45.180 158.180 ;
        RECT 45.555 157.570 45.895 158.200 ;
        RECT 46.065 157.400 46.315 158.200 ;
        RECT 46.505 158.050 47.730 158.220 ;
        RECT 46.505 157.570 46.835 158.050 ;
        RECT 47.005 157.400 47.230 157.860 ;
        RECT 47.400 157.570 47.730 158.050 ;
        RECT 48.360 158.180 48.530 158.810 ;
        RECT 48.715 158.390 49.065 158.640 ;
        RECT 49.235 158.200 49.410 158.810 ;
        RECT 50.105 158.560 50.275 158.810 ;
        RECT 49.580 158.390 50.275 158.560 ;
        RECT 50.450 158.390 50.870 158.590 ;
        RECT 51.040 158.390 51.370 158.590 ;
        RECT 51.540 158.390 51.870 158.590 ;
        RECT 48.360 157.570 48.860 158.180 ;
        RECT 49.235 157.570 49.575 158.200 ;
        RECT 49.745 157.400 49.995 158.200 ;
        RECT 50.185 158.050 51.410 158.220 ;
        RECT 50.185 157.570 50.515 158.050 ;
        RECT 50.685 157.400 50.910 157.860 ;
        RECT 51.080 157.570 51.410 158.050 ;
        RECT 52.040 158.180 52.210 158.810 ;
        RECT 52.395 158.390 52.745 158.640 ;
        RECT 52.915 158.340 53.665 158.860 ;
        RECT 54.815 158.810 61.590 158.930 ;
        RECT 54.815 158.760 56.010 158.810 ;
        RECT 52.040 157.570 52.540 158.180 ;
        RECT 53.835 158.170 54.585 158.690 ;
        RECT 52.915 157.400 54.585 158.170 ;
        RECT 54.845 158.220 56.010 158.760 ;
        RECT 62.190 158.640 62.440 159.775 ;
        RECT 62.620 159.140 62.880 159.950 ;
        RECT 63.055 158.640 63.300 159.780 ;
        RECT 63.480 159.140 63.775 159.950 ;
        RECT 63.955 158.785 64.245 159.950 ;
        RECT 65.425 159.020 65.595 159.780 ;
        RECT 65.810 159.190 66.140 159.950 ;
        RECT 65.425 158.850 66.140 159.020 ;
        RECT 66.310 158.875 66.565 159.780 ;
        RECT 56.180 158.390 63.300 158.640 ;
        RECT 54.845 158.050 61.590 158.220 ;
        RECT 54.845 157.400 55.145 157.880 ;
        RECT 55.315 157.595 55.575 158.050 ;
        RECT 55.745 157.400 56.005 157.880 ;
        RECT 56.185 157.595 56.445 158.050 ;
        RECT 56.615 157.400 56.865 157.880 ;
        RECT 57.045 157.595 57.305 158.050 ;
        RECT 57.475 157.400 57.725 157.880 ;
        RECT 57.905 157.595 58.165 158.050 ;
        RECT 58.335 157.400 58.580 157.880 ;
        RECT 58.750 157.595 59.025 158.050 ;
        RECT 59.195 157.400 59.440 157.880 ;
        RECT 59.610 157.595 59.870 158.050 ;
        RECT 60.040 157.400 60.300 157.880 ;
        RECT 60.470 157.595 60.730 158.050 ;
        RECT 60.900 157.400 61.160 157.880 ;
        RECT 61.330 157.595 61.590 158.050 ;
        RECT 61.760 157.400 62.020 157.960 ;
        RECT 62.190 157.580 62.440 158.390 ;
        RECT 62.620 157.400 62.880 157.925 ;
        RECT 63.050 157.580 63.300 158.390 ;
        RECT 63.470 158.080 63.785 158.640 ;
        RECT 65.335 158.300 65.690 158.670 ;
        RECT 65.970 158.640 66.140 158.850 ;
        RECT 65.970 158.310 66.225 158.640 ;
        RECT 63.480 157.400 63.785 157.910 ;
        RECT 63.955 157.400 64.245 158.125 ;
        RECT 65.970 158.120 66.140 158.310 ;
        RECT 66.395 158.145 66.565 158.875 ;
        RECT 66.740 158.800 67.000 159.950 ;
        RECT 67.380 158.980 67.710 159.780 ;
        RECT 67.880 159.150 68.210 159.950 ;
        RECT 68.510 158.980 68.840 159.780 ;
        RECT 69.485 159.150 69.735 159.950 ;
        RECT 67.380 158.810 69.815 158.980 ;
        RECT 70.005 158.810 70.175 159.950 ;
        RECT 70.345 158.810 70.685 159.780 ;
        RECT 67.175 158.390 67.525 158.640 ;
        RECT 65.425 157.950 66.140 158.120 ;
        RECT 65.425 157.570 65.595 157.950 ;
        RECT 65.810 157.400 66.140 157.780 ;
        RECT 66.310 157.570 66.565 158.145 ;
        RECT 66.740 157.400 67.000 158.240 ;
        RECT 67.710 158.180 67.880 158.810 ;
        RECT 68.050 158.390 68.380 158.590 ;
        RECT 68.550 158.390 68.880 158.590 ;
        RECT 69.050 158.390 69.470 158.590 ;
        RECT 69.645 158.560 69.815 158.810 ;
        RECT 69.645 158.390 70.340 158.560 ;
        RECT 67.380 157.570 67.880 158.180 ;
        RECT 68.510 158.050 69.735 158.220 ;
        RECT 70.510 158.200 70.685 158.810 ;
        RECT 68.510 157.570 68.840 158.050 ;
        RECT 69.010 157.400 69.235 157.860 ;
        RECT 69.405 157.570 69.735 158.050 ;
        RECT 69.925 157.400 70.175 158.200 ;
        RECT 70.345 157.570 70.685 158.200 ;
        RECT 70.855 158.810 71.195 159.780 ;
        RECT 71.365 158.810 71.535 159.950 ;
        RECT 71.805 159.150 72.055 159.950 ;
        RECT 72.700 158.980 73.030 159.780 ;
        RECT 73.330 159.150 73.660 159.950 ;
        RECT 73.830 158.980 74.160 159.780 ;
        RECT 71.725 158.810 74.160 158.980 ;
        RECT 75.370 158.970 75.625 159.640 ;
        RECT 75.805 159.150 76.090 159.950 ;
        RECT 76.270 159.230 76.600 159.740 ;
        RECT 70.855 158.760 71.085 158.810 ;
        RECT 70.855 158.200 71.030 158.760 ;
        RECT 71.725 158.560 71.895 158.810 ;
        RECT 71.200 158.390 71.895 158.560 ;
        RECT 72.070 158.390 72.490 158.590 ;
        RECT 72.660 158.390 72.990 158.590 ;
        RECT 73.160 158.390 73.490 158.590 ;
        RECT 70.855 157.570 71.195 158.200 ;
        RECT 71.365 157.400 71.615 158.200 ;
        RECT 71.805 158.050 73.030 158.220 ;
        RECT 71.805 157.570 72.135 158.050 ;
        RECT 72.305 157.400 72.530 157.860 ;
        RECT 72.700 157.570 73.030 158.050 ;
        RECT 73.660 158.180 73.830 158.810 ;
        RECT 74.015 158.390 74.365 158.640 ;
        RECT 75.370 158.250 75.550 158.970 ;
        RECT 76.270 158.640 76.520 159.230 ;
        RECT 76.870 159.080 77.040 159.690 ;
        RECT 77.210 159.260 77.540 159.950 ;
        RECT 77.770 159.400 78.010 159.690 ;
        RECT 78.210 159.570 78.630 159.950 ;
        RECT 78.810 159.480 79.440 159.730 ;
        RECT 79.910 159.570 80.240 159.950 ;
        RECT 78.810 159.400 78.980 159.480 ;
        RECT 80.410 159.400 80.580 159.690 ;
        RECT 80.760 159.570 81.140 159.950 ;
        RECT 81.380 159.565 82.210 159.735 ;
        RECT 77.770 159.230 78.980 159.400 ;
        RECT 75.720 158.310 76.520 158.640 ;
        RECT 73.660 157.570 74.160 158.180 ;
        RECT 75.285 158.110 75.550 158.250 ;
        RECT 75.285 158.080 75.625 158.110 ;
        RECT 75.370 157.580 75.625 158.080 ;
        RECT 75.805 157.400 76.090 157.860 ;
        RECT 76.270 157.660 76.520 158.310 ;
        RECT 76.720 159.060 77.040 159.080 ;
        RECT 76.720 158.890 78.640 159.060 ;
        RECT 76.720 157.995 76.910 158.890 ;
        RECT 78.810 158.720 78.980 159.230 ;
        RECT 79.150 158.970 79.670 159.280 ;
        RECT 77.080 158.550 78.980 158.720 ;
        RECT 77.080 158.490 77.410 158.550 ;
        RECT 77.560 158.320 77.890 158.380 ;
        RECT 77.230 158.050 77.890 158.320 ;
        RECT 76.720 157.665 77.040 157.995 ;
        RECT 77.220 157.400 77.880 157.880 ;
        RECT 78.080 157.790 78.250 158.550 ;
        RECT 79.150 158.380 79.330 158.790 ;
        RECT 78.420 158.210 78.750 158.330 ;
        RECT 79.500 158.210 79.670 158.970 ;
        RECT 78.420 158.040 79.670 158.210 ;
        RECT 79.840 159.150 81.210 159.400 ;
        RECT 79.840 158.380 80.030 159.150 ;
        RECT 80.960 158.890 81.210 159.150 ;
        RECT 80.200 158.720 80.450 158.880 ;
        RECT 81.380 158.720 81.550 159.565 ;
        RECT 82.445 159.280 82.615 159.780 ;
        RECT 82.785 159.450 83.115 159.950 ;
        RECT 81.720 158.890 82.220 159.270 ;
        RECT 82.445 159.110 83.140 159.280 ;
        RECT 80.200 158.550 81.550 158.720 ;
        RECT 81.130 158.510 81.550 158.550 ;
        RECT 79.840 158.040 80.260 158.380 ;
        RECT 80.550 158.050 80.960 158.380 ;
        RECT 78.080 157.620 78.930 157.790 ;
        RECT 79.490 157.400 79.810 157.860 ;
        RECT 80.010 157.610 80.260 158.040 ;
        RECT 80.550 157.400 80.960 157.840 ;
        RECT 81.130 157.780 81.300 158.510 ;
        RECT 81.470 157.960 81.820 158.330 ;
        RECT 82.000 158.020 82.220 158.890 ;
        RECT 82.390 158.320 82.800 158.940 ;
        RECT 82.970 158.140 83.140 159.110 ;
        RECT 82.445 157.950 83.140 158.140 ;
        RECT 81.130 157.580 82.145 157.780 ;
        RECT 82.445 157.620 82.615 157.950 ;
        RECT 82.785 157.400 83.115 157.780 ;
        RECT 83.330 157.660 83.555 159.780 ;
        RECT 83.725 159.450 84.055 159.950 ;
        RECT 84.225 159.280 84.395 159.780 ;
        RECT 83.730 159.110 84.395 159.280 ;
        RECT 83.730 158.120 83.960 159.110 ;
        RECT 84.130 158.290 84.480 158.940 ;
        RECT 84.655 158.860 85.865 159.950 ;
        RECT 84.655 158.320 85.175 158.860 ;
        RECT 86.075 158.810 86.305 159.950 ;
        RECT 86.475 158.800 86.805 159.780 ;
        RECT 86.975 158.810 87.185 159.950 ;
        RECT 88.425 159.020 88.595 159.780 ;
        RECT 88.775 159.190 89.105 159.950 ;
        RECT 88.425 158.850 89.090 159.020 ;
        RECT 89.275 158.875 89.545 159.780 ;
        RECT 85.345 158.150 85.865 158.690 ;
        RECT 86.055 158.390 86.385 158.640 ;
        RECT 83.730 157.950 84.395 158.120 ;
        RECT 83.725 157.400 84.055 157.780 ;
        RECT 84.225 157.660 84.395 157.950 ;
        RECT 84.655 157.400 85.865 158.150 ;
        RECT 86.075 157.400 86.305 158.220 ;
        RECT 86.555 158.200 86.805 158.800 ;
        RECT 88.920 158.705 89.090 158.850 ;
        RECT 88.355 158.300 88.685 158.670 ;
        RECT 88.920 158.375 89.205 158.705 ;
        RECT 86.475 157.570 86.805 158.200 ;
        RECT 86.975 157.400 87.185 158.220 ;
        RECT 88.920 158.120 89.090 158.375 ;
        RECT 88.425 157.950 89.090 158.120 ;
        RECT 89.375 158.075 89.545 158.875 ;
        RECT 89.715 158.785 90.005 159.950 ;
        RECT 91.095 158.810 91.365 159.780 ;
        RECT 91.575 159.150 91.855 159.950 ;
        RECT 92.025 159.440 93.680 159.730 ;
        RECT 92.090 159.100 93.680 159.270 ;
        RECT 92.090 158.980 92.260 159.100 ;
        RECT 91.535 158.810 92.260 158.980 ;
        RECT 88.425 157.570 88.595 157.950 ;
        RECT 88.775 157.400 89.105 157.780 ;
        RECT 89.285 157.570 89.545 158.075 ;
        RECT 89.715 157.400 90.005 158.125 ;
        RECT 91.095 158.075 91.265 158.810 ;
        RECT 91.535 158.640 91.705 158.810 ;
        RECT 92.450 158.760 93.165 158.930 ;
        RECT 93.360 158.810 93.680 159.100 ;
        RECT 94.775 158.810 95.115 159.780 ;
        RECT 95.285 158.810 95.455 159.950 ;
        RECT 95.725 159.150 95.975 159.950 ;
        RECT 96.620 158.980 96.950 159.780 ;
        RECT 97.250 159.150 97.580 159.950 ;
        RECT 97.750 158.980 98.080 159.780 ;
        RECT 95.645 158.810 98.080 158.980 ;
        RECT 99.120 158.980 99.450 159.780 ;
        RECT 99.620 159.150 99.950 159.950 ;
        RECT 100.250 158.980 100.580 159.780 ;
        RECT 101.225 159.150 101.475 159.950 ;
        RECT 99.120 158.810 101.555 158.980 ;
        RECT 101.745 158.810 101.915 159.950 ;
        RECT 102.085 158.810 102.425 159.780 ;
        RECT 91.435 158.310 91.705 158.640 ;
        RECT 91.875 158.310 92.280 158.640 ;
        RECT 92.450 158.310 93.160 158.760 ;
        RECT 91.535 158.140 91.705 158.310 ;
        RECT 91.095 157.730 91.365 158.075 ;
        RECT 91.535 157.970 93.145 158.140 ;
        RECT 93.330 158.070 93.680 158.640 ;
        RECT 94.775 158.200 94.950 158.810 ;
        RECT 95.645 158.560 95.815 158.810 ;
        RECT 95.120 158.390 95.815 158.560 ;
        RECT 95.990 158.390 96.410 158.590 ;
        RECT 96.580 158.390 96.910 158.590 ;
        RECT 97.080 158.390 97.410 158.590 ;
        RECT 91.555 157.400 91.935 157.800 ;
        RECT 92.105 157.620 92.275 157.970 ;
        RECT 92.445 157.400 92.775 157.800 ;
        RECT 92.975 157.620 93.145 157.970 ;
        RECT 93.345 157.400 93.675 157.900 ;
        RECT 94.775 157.570 95.115 158.200 ;
        RECT 95.285 157.400 95.535 158.200 ;
        RECT 95.725 158.050 96.950 158.220 ;
        RECT 95.725 157.570 96.055 158.050 ;
        RECT 96.225 157.400 96.450 157.860 ;
        RECT 96.620 157.570 96.950 158.050 ;
        RECT 97.580 158.180 97.750 158.810 ;
        RECT 97.935 158.390 98.285 158.640 ;
        RECT 98.915 158.390 99.265 158.640 ;
        RECT 99.450 158.180 99.620 158.810 ;
        RECT 99.790 158.390 100.120 158.590 ;
        RECT 100.290 158.390 100.620 158.590 ;
        RECT 100.790 158.390 101.210 158.590 ;
        RECT 101.385 158.560 101.555 158.810 ;
        RECT 101.385 158.390 102.080 158.560 ;
        RECT 97.580 157.570 98.080 158.180 ;
        RECT 99.120 157.570 99.620 158.180 ;
        RECT 100.250 158.050 101.475 158.220 ;
        RECT 102.250 158.200 102.425 158.810 ;
        RECT 102.605 158.970 102.935 159.780 ;
        RECT 103.105 159.150 103.345 159.950 ;
        RECT 102.605 158.800 103.320 158.970 ;
        RECT 102.600 158.390 102.980 158.630 ;
        RECT 103.150 158.560 103.320 158.800 ;
        RECT 103.525 158.930 103.695 159.780 ;
        RECT 103.865 159.150 104.195 159.950 ;
        RECT 104.365 158.930 104.535 159.780 ;
        RECT 103.525 158.760 104.535 158.930 ;
        RECT 104.705 158.800 105.035 159.950 ;
        RECT 105.470 159.320 105.755 159.780 ;
        RECT 105.925 159.490 106.195 159.950 ;
        RECT 105.470 159.100 106.425 159.320 ;
        RECT 103.150 158.390 103.650 158.560 ;
        RECT 103.150 158.220 103.320 158.390 ;
        RECT 104.040 158.250 104.535 158.760 ;
        RECT 105.355 158.370 106.045 158.930 ;
        RECT 104.035 158.220 104.535 158.250 ;
        RECT 100.250 157.570 100.580 158.050 ;
        RECT 100.750 157.400 100.975 157.860 ;
        RECT 101.145 157.570 101.475 158.050 ;
        RECT 101.665 157.400 101.915 158.200 ;
        RECT 102.085 157.570 102.425 158.200 ;
        RECT 102.685 158.050 103.320 158.220 ;
        RECT 103.525 158.050 104.535 158.220 ;
        RECT 106.215 158.200 106.425 159.100 ;
        RECT 102.685 157.570 102.855 158.050 ;
        RECT 103.035 157.400 103.275 157.880 ;
        RECT 103.525 157.570 103.695 158.050 ;
        RECT 103.865 157.400 104.195 157.880 ;
        RECT 104.365 157.570 104.535 158.050 ;
        RECT 104.705 157.400 105.035 158.200 ;
        RECT 105.470 158.030 106.425 158.200 ;
        RECT 106.595 158.930 106.995 159.780 ;
        RECT 107.185 159.320 107.465 159.780 ;
        RECT 107.985 159.490 108.310 159.950 ;
        RECT 107.185 159.100 108.310 159.320 ;
        RECT 106.595 158.370 107.690 158.930 ;
        RECT 107.860 158.640 108.310 159.100 ;
        RECT 108.480 158.810 108.865 159.780 ;
        RECT 109.040 159.515 114.385 159.950 ;
        RECT 105.470 157.570 105.755 158.030 ;
        RECT 105.925 157.400 106.195 157.860 ;
        RECT 106.595 157.570 106.995 158.370 ;
        RECT 107.860 158.310 108.415 158.640 ;
        RECT 107.860 158.200 108.310 158.310 ;
        RECT 107.185 158.030 108.310 158.200 ;
        RECT 108.585 158.140 108.865 158.810 ;
        RECT 110.630 158.265 110.980 159.515 ;
        RECT 114.555 158.860 115.765 159.950 ;
        RECT 107.185 157.570 107.465 158.030 ;
        RECT 107.985 157.400 108.310 157.860 ;
        RECT 108.480 157.570 108.865 158.140 ;
        RECT 112.460 157.945 112.800 158.775 ;
        RECT 114.555 158.320 115.075 158.860 ;
        RECT 115.245 158.150 115.765 158.690 ;
        RECT 109.040 157.400 114.385 157.945 ;
        RECT 114.555 157.400 115.765 158.150 ;
        RECT 14.650 157.230 115.850 157.400 ;
        RECT 14.735 156.480 15.945 157.230 ;
        RECT 14.735 155.940 15.255 156.480 ;
        RECT 16.115 156.460 18.705 157.230 ;
        RECT 15.425 155.770 15.945 156.310 ;
        RECT 14.735 154.680 15.945 155.770 ;
        RECT 16.115 155.770 17.325 156.290 ;
        RECT 17.495 155.940 18.705 156.460 ;
        RECT 18.875 156.555 19.135 157.060 ;
        RECT 19.315 156.850 19.645 157.230 ;
        RECT 19.825 156.680 19.995 157.060 ;
        RECT 16.115 154.680 18.705 155.770 ;
        RECT 18.875 155.755 19.045 156.555 ;
        RECT 19.330 156.510 19.995 156.680 ;
        RECT 19.330 156.255 19.500 156.510 ;
        RECT 20.530 156.420 20.775 157.025 ;
        RECT 20.995 156.695 21.505 157.230 ;
        RECT 19.215 155.925 19.500 156.255 ;
        RECT 19.735 155.960 20.065 156.330 ;
        RECT 20.255 156.250 21.485 156.420 ;
        RECT 19.330 155.780 19.500 155.925 ;
        RECT 18.875 154.850 19.145 155.755 ;
        RECT 19.330 155.610 19.995 155.780 ;
        RECT 19.315 154.680 19.645 155.440 ;
        RECT 19.825 154.850 19.995 155.610 ;
        RECT 20.255 155.440 20.595 156.250 ;
        RECT 20.765 155.685 21.515 155.875 ;
        RECT 20.255 155.030 20.770 155.440 ;
        RECT 21.005 154.680 21.175 155.440 ;
        RECT 21.345 155.020 21.515 155.685 ;
        RECT 21.685 155.700 21.875 157.060 ;
        RECT 22.045 156.210 22.320 157.060 ;
        RECT 22.510 156.695 23.040 157.060 ;
        RECT 23.465 156.830 23.795 157.230 ;
        RECT 22.865 156.660 23.040 156.695 ;
        RECT 22.045 156.040 22.325 156.210 ;
        RECT 22.045 155.900 22.320 156.040 ;
        RECT 22.525 155.700 22.695 156.500 ;
        RECT 21.685 155.530 22.695 155.700 ;
        RECT 22.865 156.490 23.795 156.660 ;
        RECT 23.965 156.490 24.220 157.060 ;
        RECT 25.315 156.505 25.605 157.230 ;
        RECT 22.865 155.360 23.035 156.490 ;
        RECT 23.625 156.320 23.795 156.490 ;
        RECT 21.910 155.190 23.035 155.360 ;
        RECT 23.205 155.990 23.400 156.320 ;
        RECT 23.625 155.990 23.880 156.320 ;
        RECT 23.205 155.020 23.375 155.990 ;
        RECT 24.050 155.820 24.220 156.490 ;
        RECT 26.695 156.460 30.205 157.230 ;
        RECT 21.345 154.850 23.375 155.020 ;
        RECT 23.545 154.680 23.715 155.820 ;
        RECT 23.885 154.850 24.220 155.820 ;
        RECT 25.315 154.680 25.605 155.845 ;
        RECT 26.695 155.770 28.385 156.290 ;
        RECT 28.555 155.940 30.205 156.460 ;
        RECT 30.375 156.430 30.715 157.060 ;
        RECT 30.885 156.430 31.135 157.230 ;
        RECT 31.325 156.580 31.655 157.060 ;
        RECT 31.825 156.770 32.050 157.230 ;
        RECT 32.220 156.580 32.550 157.060 ;
        RECT 30.375 155.820 30.550 156.430 ;
        RECT 31.325 156.410 32.550 156.580 ;
        RECT 33.180 156.450 33.680 157.060 ;
        RECT 34.055 156.460 35.725 157.230 ;
        RECT 30.720 156.070 31.415 156.240 ;
        RECT 31.245 155.820 31.415 156.070 ;
        RECT 31.590 156.040 32.010 156.240 ;
        RECT 32.180 156.040 32.510 156.240 ;
        RECT 32.680 156.040 33.010 156.240 ;
        RECT 33.180 155.820 33.350 156.450 ;
        RECT 33.535 155.990 33.885 156.240 ;
        RECT 26.695 154.680 30.205 155.770 ;
        RECT 30.375 154.850 30.715 155.820 ;
        RECT 30.885 154.680 31.055 155.820 ;
        RECT 31.245 155.650 33.680 155.820 ;
        RECT 31.325 154.680 31.575 155.480 ;
        RECT 32.220 154.850 32.550 155.650 ;
        RECT 32.850 154.680 33.180 155.480 ;
        RECT 33.350 154.850 33.680 155.650 ;
        RECT 34.055 155.770 34.805 156.290 ;
        RECT 34.975 155.940 35.725 156.460 ;
        RECT 36.100 156.450 36.600 157.060 ;
        RECT 35.895 155.990 36.245 156.240 ;
        RECT 36.430 155.820 36.600 156.450 ;
        RECT 37.230 156.580 37.560 157.060 ;
        RECT 37.730 156.770 37.955 157.230 ;
        RECT 38.125 156.580 38.455 157.060 ;
        RECT 37.230 156.410 38.455 156.580 ;
        RECT 38.645 156.430 38.895 157.230 ;
        RECT 39.065 156.430 39.405 157.060 ;
        RECT 39.780 156.450 40.280 157.060 ;
        RECT 36.770 156.040 37.100 156.240 ;
        RECT 37.270 156.040 37.600 156.240 ;
        RECT 37.770 156.040 38.190 156.240 ;
        RECT 38.365 156.070 39.060 156.240 ;
        RECT 38.365 155.820 38.535 156.070 ;
        RECT 39.230 155.820 39.405 156.430 ;
        RECT 39.575 155.990 39.925 156.240 ;
        RECT 40.110 155.820 40.280 156.450 ;
        RECT 40.910 156.580 41.240 157.060 ;
        RECT 41.410 156.770 41.635 157.230 ;
        RECT 41.805 156.580 42.135 157.060 ;
        RECT 40.910 156.410 42.135 156.580 ;
        RECT 42.325 156.430 42.575 157.230 ;
        RECT 42.745 156.430 43.085 157.060 ;
        RECT 43.255 156.460 45.845 157.230 ;
        RECT 40.450 156.040 40.780 156.240 ;
        RECT 40.950 156.040 41.280 156.240 ;
        RECT 41.450 156.040 41.870 156.240 ;
        RECT 42.045 156.070 42.740 156.240 ;
        RECT 42.045 155.820 42.215 156.070 ;
        RECT 42.910 155.820 43.085 156.430 ;
        RECT 34.055 154.680 35.725 155.770 ;
        RECT 36.100 155.650 38.535 155.820 ;
        RECT 36.100 154.850 36.430 155.650 ;
        RECT 36.600 154.680 36.930 155.480 ;
        RECT 37.230 154.850 37.560 155.650 ;
        RECT 38.205 154.680 38.455 155.480 ;
        RECT 38.725 154.680 38.895 155.820 ;
        RECT 39.065 154.850 39.405 155.820 ;
        RECT 39.780 155.650 42.215 155.820 ;
        RECT 39.780 154.850 40.110 155.650 ;
        RECT 40.280 154.680 40.610 155.480 ;
        RECT 40.910 154.850 41.240 155.650 ;
        RECT 41.885 154.680 42.135 155.480 ;
        RECT 42.405 154.680 42.575 155.820 ;
        RECT 42.745 154.850 43.085 155.820 ;
        RECT 43.255 155.770 44.465 156.290 ;
        RECT 44.635 155.940 45.845 156.460 ;
        RECT 46.055 156.410 46.285 157.230 ;
        RECT 46.455 156.430 46.785 157.060 ;
        RECT 46.035 155.990 46.365 156.240 ;
        RECT 46.535 155.830 46.785 156.430 ;
        RECT 46.955 156.410 47.165 157.230 ;
        RECT 48.065 156.540 48.395 157.230 ;
        RECT 48.855 156.635 49.475 157.060 ;
        RECT 49.645 156.740 49.975 157.230 ;
        RECT 49.115 156.300 49.475 156.635 ;
        RECT 48.055 156.020 49.475 156.300 ;
        RECT 43.255 154.680 45.845 155.770 ;
        RECT 46.055 154.680 46.285 155.820 ;
        RECT 46.455 154.850 46.785 155.830 ;
        RECT 46.955 154.680 47.165 155.820 ;
        RECT 47.525 154.680 47.855 155.850 ;
        RECT 48.055 154.850 48.385 156.020 ;
        RECT 48.585 154.680 48.915 155.850 ;
        RECT 49.115 154.850 49.475 156.020 ;
        RECT 49.645 155.990 49.985 156.570 ;
        RECT 51.075 156.505 51.365 157.230 ;
        RECT 51.995 156.460 53.665 157.230 ;
        RECT 53.925 156.680 54.095 157.060 ;
        RECT 54.275 156.850 54.605 157.230 ;
        RECT 53.925 156.510 54.590 156.680 ;
        RECT 54.785 156.555 55.045 157.060 ;
        RECT 49.645 154.680 49.975 155.820 ;
        RECT 51.075 154.680 51.365 155.845 ;
        RECT 51.995 155.770 52.745 156.290 ;
        RECT 52.915 155.940 53.665 156.460 ;
        RECT 53.855 155.960 54.185 156.330 ;
        RECT 54.420 156.255 54.590 156.510 ;
        RECT 54.420 155.925 54.705 156.255 ;
        RECT 54.420 155.780 54.590 155.925 ;
        RECT 51.995 154.680 53.665 155.770 ;
        RECT 53.925 155.610 54.590 155.780 ;
        RECT 54.875 155.755 55.045 156.555 ;
        RECT 53.925 154.850 54.095 155.610 ;
        RECT 54.275 154.680 54.605 155.440 ;
        RECT 54.775 154.850 55.045 155.755 ;
        RECT 55.590 156.520 55.845 157.050 ;
        RECT 56.025 156.770 56.310 157.230 ;
        RECT 55.590 155.660 55.770 156.520 ;
        RECT 56.490 156.320 56.740 156.970 ;
        RECT 55.940 155.990 56.740 156.320 ;
        RECT 55.590 155.530 55.845 155.660 ;
        RECT 55.505 155.360 55.845 155.530 ;
        RECT 55.590 154.990 55.845 155.360 ;
        RECT 56.025 154.680 56.310 155.480 ;
        RECT 56.490 155.400 56.740 155.990 ;
        RECT 56.940 156.635 57.260 156.965 ;
        RECT 57.440 156.750 58.100 157.230 ;
        RECT 58.300 156.840 59.150 157.010 ;
        RECT 56.940 155.740 57.130 156.635 ;
        RECT 57.450 156.310 58.110 156.580 ;
        RECT 57.780 156.250 58.110 156.310 ;
        RECT 57.300 156.080 57.630 156.140 ;
        RECT 58.300 156.080 58.470 156.840 ;
        RECT 59.710 156.770 60.030 157.230 ;
        RECT 60.230 156.590 60.480 157.020 ;
        RECT 60.770 156.790 61.180 157.230 ;
        RECT 61.350 156.850 62.365 157.050 ;
        RECT 58.640 156.420 59.890 156.590 ;
        RECT 58.640 156.300 58.970 156.420 ;
        RECT 57.300 155.910 59.200 156.080 ;
        RECT 56.940 155.570 58.860 155.740 ;
        RECT 56.940 155.550 57.260 155.570 ;
        RECT 56.490 154.890 56.820 155.400 ;
        RECT 57.090 154.940 57.260 155.550 ;
        RECT 59.030 155.400 59.200 155.910 ;
        RECT 59.370 155.840 59.550 156.250 ;
        RECT 59.720 155.660 59.890 156.420 ;
        RECT 57.430 154.680 57.760 155.370 ;
        RECT 57.990 155.230 59.200 155.400 ;
        RECT 59.370 155.350 59.890 155.660 ;
        RECT 60.060 156.250 60.480 156.590 ;
        RECT 60.770 156.250 61.180 156.580 ;
        RECT 60.060 155.480 60.250 156.250 ;
        RECT 61.350 156.120 61.520 156.850 ;
        RECT 62.665 156.680 62.835 157.010 ;
        RECT 63.005 156.850 63.335 157.230 ;
        RECT 61.690 156.300 62.040 156.670 ;
        RECT 61.350 156.080 61.770 156.120 ;
        RECT 60.420 155.910 61.770 156.080 ;
        RECT 60.420 155.750 60.670 155.910 ;
        RECT 61.180 155.480 61.430 155.740 ;
        RECT 60.060 155.230 61.430 155.480 ;
        RECT 57.990 154.940 58.230 155.230 ;
        RECT 59.030 155.150 59.200 155.230 ;
        RECT 58.430 154.680 58.850 155.060 ;
        RECT 59.030 154.900 59.660 155.150 ;
        RECT 60.130 154.680 60.460 155.060 ;
        RECT 60.630 154.940 60.800 155.230 ;
        RECT 61.600 155.065 61.770 155.910 ;
        RECT 62.220 155.740 62.440 156.610 ;
        RECT 62.665 156.490 63.360 156.680 ;
        RECT 61.940 155.360 62.440 155.740 ;
        RECT 62.610 155.690 63.020 156.310 ;
        RECT 63.190 155.520 63.360 156.490 ;
        RECT 62.665 155.350 63.360 155.520 ;
        RECT 60.980 154.680 61.360 155.060 ;
        RECT 61.600 154.895 62.430 155.065 ;
        RECT 62.665 154.850 62.835 155.350 ;
        RECT 63.005 154.680 63.335 155.180 ;
        RECT 63.550 154.850 63.775 156.970 ;
        RECT 63.945 156.850 64.275 157.230 ;
        RECT 64.445 156.680 64.615 156.970 ;
        RECT 63.950 156.510 64.615 156.680 ;
        RECT 63.950 155.520 64.180 156.510 ;
        RECT 64.875 156.480 66.085 157.230 ;
        RECT 66.345 156.680 66.515 157.060 ;
        RECT 66.730 156.850 67.060 157.230 ;
        RECT 66.345 156.510 67.060 156.680 ;
        RECT 64.350 155.690 64.700 156.340 ;
        RECT 64.875 155.770 65.395 156.310 ;
        RECT 65.565 155.940 66.085 156.480 ;
        RECT 66.255 155.960 66.610 156.330 ;
        RECT 66.890 156.320 67.060 156.510 ;
        RECT 67.230 156.485 67.485 157.060 ;
        RECT 66.890 155.990 67.145 156.320 ;
        RECT 66.890 155.780 67.060 155.990 ;
        RECT 63.950 155.350 64.615 155.520 ;
        RECT 63.945 154.680 64.275 155.180 ;
        RECT 64.445 154.850 64.615 155.350 ;
        RECT 64.875 154.680 66.085 155.770 ;
        RECT 66.345 155.610 67.060 155.780 ;
        RECT 67.315 155.755 67.485 156.485 ;
        RECT 67.660 156.390 67.920 157.230 ;
        RECT 68.105 156.700 68.435 157.060 ;
        RECT 68.605 156.870 68.935 157.230 ;
        RECT 69.135 156.700 69.465 157.060 ;
        RECT 68.105 156.490 69.465 156.700 ;
        RECT 69.975 156.470 70.685 157.060 ;
        RECT 68.095 155.990 68.405 156.320 ;
        RECT 68.615 155.990 68.990 156.320 ;
        RECT 69.310 155.990 69.805 156.320 ;
        RECT 66.345 154.850 66.515 155.610 ;
        RECT 66.730 154.680 67.060 155.440 ;
        RECT 67.230 154.850 67.485 155.755 ;
        RECT 67.660 154.680 67.920 155.830 ;
        RECT 68.105 154.680 68.435 155.740 ;
        RECT 68.615 155.065 68.785 155.990 ;
        RECT 68.955 155.500 69.285 155.720 ;
        RECT 69.480 155.700 69.805 155.990 ;
        RECT 69.980 155.700 70.310 156.240 ;
        RECT 70.480 155.500 70.685 156.470 ;
        RECT 71.980 156.450 72.480 157.060 ;
        RECT 71.775 155.990 72.125 156.240 ;
        RECT 72.310 155.820 72.480 156.450 ;
        RECT 73.110 156.580 73.440 157.060 ;
        RECT 73.610 156.770 73.835 157.230 ;
        RECT 74.005 156.580 74.335 157.060 ;
        RECT 73.110 156.410 74.335 156.580 ;
        RECT 74.525 156.430 74.775 157.230 ;
        RECT 74.945 156.430 75.285 157.060 ;
        RECT 75.455 156.480 76.665 157.230 ;
        RECT 76.835 156.505 77.125 157.230 ;
        RECT 78.220 156.685 83.565 157.230 ;
        RECT 83.740 156.685 89.085 157.230 ;
        RECT 72.650 156.040 72.980 156.240 ;
        RECT 73.150 156.040 73.480 156.240 ;
        RECT 73.650 156.040 74.070 156.240 ;
        RECT 74.245 156.070 74.940 156.240 ;
        RECT 74.245 155.820 74.415 156.070 ;
        RECT 75.110 155.820 75.285 156.430 ;
        RECT 68.955 155.270 70.685 155.500 ;
        RECT 68.955 154.870 69.285 155.270 ;
        RECT 69.455 154.680 69.785 155.040 ;
        RECT 69.985 154.850 70.685 155.270 ;
        RECT 71.980 155.650 74.415 155.820 ;
        RECT 71.980 154.850 72.310 155.650 ;
        RECT 72.480 154.680 72.810 155.480 ;
        RECT 73.110 154.850 73.440 155.650 ;
        RECT 74.085 154.680 74.335 155.480 ;
        RECT 74.605 154.680 74.775 155.820 ;
        RECT 74.945 154.850 75.285 155.820 ;
        RECT 75.455 155.770 75.975 156.310 ;
        RECT 76.145 155.940 76.665 156.480 ;
        RECT 75.455 154.680 76.665 155.770 ;
        RECT 76.835 154.680 77.125 155.845 ;
        RECT 79.810 155.115 80.160 156.365 ;
        RECT 81.640 155.855 81.980 156.685 ;
        RECT 85.330 155.115 85.680 156.365 ;
        RECT 87.160 155.855 87.500 156.685 ;
        RECT 89.255 156.430 89.595 157.060 ;
        RECT 89.765 156.430 90.015 157.230 ;
        RECT 90.205 156.580 90.535 157.060 ;
        RECT 90.705 156.770 90.930 157.230 ;
        RECT 91.100 156.580 91.430 157.060 ;
        RECT 89.255 155.820 89.430 156.430 ;
        RECT 90.205 156.410 91.430 156.580 ;
        RECT 92.060 156.450 92.560 157.060 ;
        RECT 89.600 156.070 90.295 156.240 ;
        RECT 90.125 155.820 90.295 156.070 ;
        RECT 90.470 156.040 90.890 156.240 ;
        RECT 91.060 156.040 91.390 156.240 ;
        RECT 91.560 156.040 91.890 156.240 ;
        RECT 92.060 155.820 92.230 156.450 ;
        RECT 93.855 156.430 94.195 157.060 ;
        RECT 94.365 156.430 94.615 157.230 ;
        RECT 94.805 156.580 95.135 157.060 ;
        RECT 95.305 156.770 95.530 157.230 ;
        RECT 95.700 156.580 96.030 157.060 ;
        RECT 92.415 155.990 92.765 156.240 ;
        RECT 93.855 155.820 94.030 156.430 ;
        RECT 94.805 156.410 96.030 156.580 ;
        RECT 96.660 156.450 97.160 157.060 ;
        RECT 97.740 156.450 98.240 157.060 ;
        RECT 94.200 156.070 94.895 156.240 ;
        RECT 94.725 155.820 94.895 156.070 ;
        RECT 95.070 156.040 95.490 156.240 ;
        RECT 95.660 156.040 95.990 156.240 ;
        RECT 96.160 156.040 96.490 156.240 ;
        RECT 96.660 155.820 96.830 156.450 ;
        RECT 97.015 155.990 97.365 156.240 ;
        RECT 97.535 155.990 97.885 156.240 ;
        RECT 98.070 155.820 98.240 156.450 ;
        RECT 98.870 156.580 99.200 157.060 ;
        RECT 99.370 156.770 99.595 157.230 ;
        RECT 99.765 156.580 100.095 157.060 ;
        RECT 98.870 156.410 100.095 156.580 ;
        RECT 100.285 156.430 100.535 157.230 ;
        RECT 100.705 156.430 101.045 157.060 ;
        RECT 101.305 156.680 101.475 157.060 ;
        RECT 101.655 156.850 101.985 157.230 ;
        RECT 101.305 156.510 101.970 156.680 ;
        RECT 102.165 156.555 102.425 157.060 ;
        RECT 98.410 156.040 98.740 156.240 ;
        RECT 98.910 156.040 99.240 156.240 ;
        RECT 99.410 156.040 99.830 156.240 ;
        RECT 100.005 156.070 100.700 156.240 ;
        RECT 100.005 155.820 100.175 156.070 ;
        RECT 100.870 155.820 101.045 156.430 ;
        RECT 101.235 155.960 101.565 156.330 ;
        RECT 101.800 156.255 101.970 156.510 ;
        RECT 78.220 154.680 83.565 155.115 ;
        RECT 83.740 154.680 89.085 155.115 ;
        RECT 89.255 154.850 89.595 155.820 ;
        RECT 89.765 154.680 89.935 155.820 ;
        RECT 90.125 155.650 92.560 155.820 ;
        RECT 90.205 154.680 90.455 155.480 ;
        RECT 91.100 154.850 91.430 155.650 ;
        RECT 91.730 154.680 92.060 155.480 ;
        RECT 92.230 154.850 92.560 155.650 ;
        RECT 93.855 154.850 94.195 155.820 ;
        RECT 94.365 154.680 94.535 155.820 ;
        RECT 94.725 155.650 97.160 155.820 ;
        RECT 94.805 154.680 95.055 155.480 ;
        RECT 95.700 154.850 96.030 155.650 ;
        RECT 96.330 154.680 96.660 155.480 ;
        RECT 96.830 154.850 97.160 155.650 ;
        RECT 97.740 155.650 100.175 155.820 ;
        RECT 97.740 154.850 98.070 155.650 ;
        RECT 98.240 154.680 98.570 155.480 ;
        RECT 98.870 154.850 99.200 155.650 ;
        RECT 99.845 154.680 100.095 155.480 ;
        RECT 100.365 154.680 100.535 155.820 ;
        RECT 100.705 154.850 101.045 155.820 ;
        RECT 101.800 155.925 102.085 156.255 ;
        RECT 101.800 155.780 101.970 155.925 ;
        RECT 101.305 155.610 101.970 155.780 ;
        RECT 102.255 155.755 102.425 156.555 ;
        RECT 102.595 156.505 102.885 157.230 ;
        RECT 103.055 156.480 104.265 157.230 ;
        RECT 101.305 154.850 101.475 155.610 ;
        RECT 101.655 154.680 101.985 155.440 ;
        RECT 102.155 154.850 102.425 155.755 ;
        RECT 102.595 154.680 102.885 155.845 ;
        RECT 103.055 155.770 103.575 156.310 ;
        RECT 103.745 155.940 104.265 156.480 ;
        RECT 104.435 156.460 107.945 157.230 ;
        RECT 104.435 155.770 106.125 156.290 ;
        RECT 106.295 155.940 107.945 156.460 ;
        RECT 108.175 156.410 108.385 157.230 ;
        RECT 108.555 156.430 108.885 157.060 ;
        RECT 108.555 155.830 108.805 156.430 ;
        RECT 109.055 156.410 109.285 157.230 ;
        RECT 110.505 156.680 110.675 157.060 ;
        RECT 110.855 156.850 111.185 157.230 ;
        RECT 110.505 156.510 111.170 156.680 ;
        RECT 111.365 156.555 111.625 157.060 ;
        RECT 108.975 155.990 109.305 156.240 ;
        RECT 110.435 155.960 110.765 156.330 ;
        RECT 111.000 156.255 111.170 156.510 ;
        RECT 111.000 155.925 111.285 156.255 ;
        RECT 103.055 154.680 104.265 155.770 ;
        RECT 104.435 154.680 107.945 155.770 ;
        RECT 108.175 154.680 108.385 155.820 ;
        RECT 108.555 154.850 108.885 155.830 ;
        RECT 109.055 154.680 109.285 155.820 ;
        RECT 111.000 155.780 111.170 155.925 ;
        RECT 110.505 155.610 111.170 155.780 ;
        RECT 111.455 155.755 111.625 156.555 ;
        RECT 111.795 156.460 114.385 157.230 ;
        RECT 114.555 156.480 115.765 157.230 ;
        RECT 110.505 154.850 110.675 155.610 ;
        RECT 110.855 154.680 111.185 155.440 ;
        RECT 111.355 154.850 111.625 155.755 ;
        RECT 111.795 155.770 113.005 156.290 ;
        RECT 113.175 155.940 114.385 156.460 ;
        RECT 114.555 155.770 115.075 156.310 ;
        RECT 115.245 155.940 115.765 156.480 ;
        RECT 111.795 154.680 114.385 155.770 ;
        RECT 114.555 154.680 115.765 155.770 ;
        RECT 14.650 154.510 115.850 154.680 ;
        RECT 14.735 153.420 15.945 154.510 ;
        RECT 14.735 152.710 15.255 153.250 ;
        RECT 15.425 152.880 15.945 153.420 ;
        RECT 16.490 153.530 16.745 154.200 ;
        RECT 16.925 153.710 17.210 154.510 ;
        RECT 17.390 153.790 17.720 154.300 ;
        RECT 14.735 151.960 15.945 152.710 ;
        RECT 16.490 152.670 16.670 153.530 ;
        RECT 17.390 153.200 17.640 153.790 ;
        RECT 17.990 153.640 18.160 154.250 ;
        RECT 18.330 153.820 18.660 154.510 ;
        RECT 18.890 153.960 19.130 154.250 ;
        RECT 19.330 154.130 19.750 154.510 ;
        RECT 19.930 154.040 20.560 154.290 ;
        RECT 21.030 154.130 21.360 154.510 ;
        RECT 19.930 153.960 20.100 154.040 ;
        RECT 21.530 153.960 21.700 154.250 ;
        RECT 21.880 154.130 22.260 154.510 ;
        RECT 22.500 154.125 23.330 154.295 ;
        RECT 18.890 153.790 20.100 153.960 ;
        RECT 16.840 152.870 17.640 153.200 ;
        RECT 16.490 152.470 16.745 152.670 ;
        RECT 16.405 152.300 16.745 152.470 ;
        RECT 16.490 152.140 16.745 152.300 ;
        RECT 16.925 151.960 17.210 152.420 ;
        RECT 17.390 152.220 17.640 152.870 ;
        RECT 17.840 153.620 18.160 153.640 ;
        RECT 17.840 153.450 19.760 153.620 ;
        RECT 17.840 152.555 18.030 153.450 ;
        RECT 19.930 153.280 20.100 153.790 ;
        RECT 20.270 153.530 20.790 153.840 ;
        RECT 18.200 153.110 20.100 153.280 ;
        RECT 18.200 153.050 18.530 153.110 ;
        RECT 18.680 152.880 19.010 152.940 ;
        RECT 18.350 152.610 19.010 152.880 ;
        RECT 17.840 152.225 18.160 152.555 ;
        RECT 18.340 151.960 19.000 152.440 ;
        RECT 19.200 152.350 19.370 153.110 ;
        RECT 20.270 152.940 20.450 153.350 ;
        RECT 19.540 152.770 19.870 152.890 ;
        RECT 20.620 152.770 20.790 153.530 ;
        RECT 19.540 152.600 20.790 152.770 ;
        RECT 20.960 153.710 22.330 153.960 ;
        RECT 20.960 152.940 21.150 153.710 ;
        RECT 22.080 153.450 22.330 153.710 ;
        RECT 21.320 153.280 21.570 153.440 ;
        RECT 22.500 153.280 22.670 154.125 ;
        RECT 23.565 153.840 23.735 154.340 ;
        RECT 23.905 154.010 24.235 154.510 ;
        RECT 22.840 153.450 23.340 153.830 ;
        RECT 23.565 153.670 24.260 153.840 ;
        RECT 21.320 153.110 22.670 153.280 ;
        RECT 22.250 153.070 22.670 153.110 ;
        RECT 20.960 152.600 21.380 152.940 ;
        RECT 21.670 152.610 22.080 152.940 ;
        RECT 19.200 152.180 20.050 152.350 ;
        RECT 20.610 151.960 20.930 152.420 ;
        RECT 21.130 152.170 21.380 152.600 ;
        RECT 21.670 151.960 22.080 152.400 ;
        RECT 22.250 152.340 22.420 153.070 ;
        RECT 22.590 152.520 22.940 152.890 ;
        RECT 23.120 152.580 23.340 153.450 ;
        RECT 23.510 152.880 23.920 153.500 ;
        RECT 24.090 152.700 24.260 153.670 ;
        RECT 23.565 152.510 24.260 152.700 ;
        RECT 22.250 152.140 23.265 152.340 ;
        RECT 23.565 152.180 23.735 152.510 ;
        RECT 23.905 151.960 24.235 152.340 ;
        RECT 24.450 152.220 24.675 154.340 ;
        RECT 24.845 154.010 25.175 154.510 ;
        RECT 25.345 153.840 25.515 154.340 ;
        RECT 24.850 153.670 25.515 153.840 ;
        RECT 24.850 152.680 25.080 153.670 ;
        RECT 25.250 152.850 25.600 153.500 ;
        RECT 25.775 153.435 26.045 154.340 ;
        RECT 26.215 153.750 26.545 154.510 ;
        RECT 26.725 153.580 26.895 154.340 ;
        RECT 24.850 152.510 25.515 152.680 ;
        RECT 24.845 151.960 25.175 152.340 ;
        RECT 25.345 152.220 25.515 152.510 ;
        RECT 25.775 152.635 25.945 153.435 ;
        RECT 26.230 153.410 26.895 153.580 ;
        RECT 26.230 153.265 26.400 153.410 ;
        RECT 26.115 152.935 26.400 153.265 ;
        RECT 28.075 153.370 28.345 154.340 ;
        RECT 28.555 153.710 28.835 154.510 ;
        RECT 29.005 154.000 30.660 154.290 ;
        RECT 29.070 153.660 30.660 153.830 ;
        RECT 29.070 153.540 29.240 153.660 ;
        RECT 28.515 153.370 29.240 153.540 ;
        RECT 26.230 152.680 26.400 152.935 ;
        RECT 26.635 152.860 26.965 153.230 ;
        RECT 25.775 152.130 26.035 152.635 ;
        RECT 26.230 152.510 26.895 152.680 ;
        RECT 26.215 151.960 26.545 152.340 ;
        RECT 26.725 152.130 26.895 152.510 ;
        RECT 28.075 152.635 28.245 153.370 ;
        RECT 28.515 153.200 28.685 153.370 ;
        RECT 28.415 152.870 28.685 153.200 ;
        RECT 28.855 152.870 29.260 153.200 ;
        RECT 29.430 152.870 30.140 153.490 ;
        RECT 30.340 153.370 30.660 153.660 ;
        RECT 30.835 153.370 31.175 154.340 ;
        RECT 31.345 153.370 31.515 154.510 ;
        RECT 31.785 153.710 32.035 154.510 ;
        RECT 32.680 153.540 33.010 154.340 ;
        RECT 33.310 153.710 33.640 154.510 ;
        RECT 33.810 153.540 34.140 154.340 ;
        RECT 31.705 153.370 34.140 153.540 ;
        RECT 34.720 153.540 35.050 154.340 ;
        RECT 35.220 153.710 35.550 154.510 ;
        RECT 35.850 153.540 36.180 154.340 ;
        RECT 36.825 153.710 37.075 154.510 ;
        RECT 34.720 153.370 37.155 153.540 ;
        RECT 37.345 153.370 37.515 154.510 ;
        RECT 37.685 153.370 38.025 154.340 ;
        RECT 28.515 152.700 28.685 152.870 ;
        RECT 28.075 152.290 28.345 152.635 ;
        RECT 28.515 152.530 30.125 152.700 ;
        RECT 30.310 152.630 30.660 153.200 ;
        RECT 30.835 152.760 31.010 153.370 ;
        RECT 31.705 153.120 31.875 153.370 ;
        RECT 31.180 152.950 31.875 153.120 ;
        RECT 32.050 152.950 32.470 153.150 ;
        RECT 32.640 152.950 32.970 153.150 ;
        RECT 33.140 152.950 33.470 153.150 ;
        RECT 28.535 151.960 28.915 152.360 ;
        RECT 29.085 152.180 29.255 152.530 ;
        RECT 29.425 151.960 29.755 152.360 ;
        RECT 29.955 152.180 30.125 152.530 ;
        RECT 30.325 151.960 30.655 152.460 ;
        RECT 30.835 152.130 31.175 152.760 ;
        RECT 31.345 151.960 31.595 152.760 ;
        RECT 31.785 152.610 33.010 152.780 ;
        RECT 31.785 152.130 32.115 152.610 ;
        RECT 32.285 151.960 32.510 152.420 ;
        RECT 32.680 152.130 33.010 152.610 ;
        RECT 33.640 152.740 33.810 153.370 ;
        RECT 33.995 152.950 34.345 153.200 ;
        RECT 34.515 152.950 34.865 153.200 ;
        RECT 35.050 152.740 35.220 153.370 ;
        RECT 35.390 152.950 35.720 153.150 ;
        RECT 35.890 152.950 36.220 153.150 ;
        RECT 36.390 152.950 36.810 153.150 ;
        RECT 36.985 153.120 37.155 153.370 ;
        RECT 36.985 152.950 37.680 153.120 ;
        RECT 33.640 152.130 34.140 152.740 ;
        RECT 34.720 152.130 35.220 152.740 ;
        RECT 35.850 152.610 37.075 152.780 ;
        RECT 37.850 152.760 38.025 153.370 ;
        RECT 38.195 153.345 38.485 154.510 ;
        RECT 38.660 154.000 40.315 154.290 ;
        RECT 38.660 153.660 40.250 153.830 ;
        RECT 40.485 153.710 40.765 154.510 ;
        RECT 38.660 153.370 38.980 153.660 ;
        RECT 40.080 153.540 40.250 153.660 ;
        RECT 39.175 153.320 39.890 153.490 ;
        RECT 40.080 153.370 40.805 153.540 ;
        RECT 40.975 153.370 41.245 154.340 ;
        RECT 35.850 152.130 36.180 152.610 ;
        RECT 36.350 151.960 36.575 152.420 ;
        RECT 36.745 152.130 37.075 152.610 ;
        RECT 37.265 151.960 37.515 152.760 ;
        RECT 37.685 152.130 38.025 152.760 ;
        RECT 38.195 151.960 38.485 152.685 ;
        RECT 38.660 152.630 39.010 153.200 ;
        RECT 39.180 152.870 39.890 153.320 ;
        RECT 40.635 153.200 40.805 153.370 ;
        RECT 40.060 152.870 40.465 153.200 ;
        RECT 40.635 152.870 40.905 153.200 ;
        RECT 40.635 152.700 40.805 152.870 ;
        RECT 39.195 152.530 40.805 152.700 ;
        RECT 41.075 152.635 41.245 153.370 ;
        RECT 38.665 151.960 38.995 152.460 ;
        RECT 39.195 152.180 39.365 152.530 ;
        RECT 39.565 151.960 39.895 152.360 ;
        RECT 40.065 152.180 40.235 152.530 ;
        RECT 40.405 151.960 40.785 152.360 ;
        RECT 40.975 152.290 41.245 152.635 ;
        RECT 41.875 153.370 42.145 154.340 ;
        RECT 42.355 153.710 42.635 154.510 ;
        RECT 42.805 154.000 44.460 154.290 ;
        RECT 44.750 153.880 45.035 154.340 ;
        RECT 45.205 154.050 45.475 154.510 ;
        RECT 42.870 153.660 44.460 153.830 ;
        RECT 44.750 153.660 45.705 153.880 ;
        RECT 42.870 153.540 43.040 153.660 ;
        RECT 42.315 153.370 43.040 153.540 ;
        RECT 41.875 152.635 42.045 153.370 ;
        RECT 42.315 153.200 42.485 153.370 ;
        RECT 43.230 153.320 43.945 153.490 ;
        RECT 44.140 153.370 44.460 153.660 ;
        RECT 42.215 152.870 42.485 153.200 ;
        RECT 42.655 152.870 43.060 153.200 ;
        RECT 43.230 152.870 43.940 153.320 ;
        RECT 42.315 152.700 42.485 152.870 ;
        RECT 41.875 152.290 42.145 152.635 ;
        RECT 42.315 152.530 43.925 152.700 ;
        RECT 44.110 152.630 44.460 153.200 ;
        RECT 44.635 152.930 45.325 153.490 ;
        RECT 45.495 152.760 45.705 153.660 ;
        RECT 42.335 151.960 42.715 152.360 ;
        RECT 42.885 152.180 43.055 152.530 ;
        RECT 43.225 151.960 43.555 152.360 ;
        RECT 43.755 152.180 43.925 152.530 ;
        RECT 44.750 152.590 45.705 152.760 ;
        RECT 45.875 153.490 46.275 154.340 ;
        RECT 46.465 153.880 46.745 154.340 ;
        RECT 47.265 154.050 47.590 154.510 ;
        RECT 46.465 153.660 47.590 153.880 ;
        RECT 45.875 152.930 46.970 153.490 ;
        RECT 47.140 153.200 47.590 153.660 ;
        RECT 47.760 153.370 48.145 154.340 ;
        RECT 44.125 151.960 44.455 152.460 ;
        RECT 44.750 152.130 45.035 152.590 ;
        RECT 45.205 151.960 45.475 152.420 ;
        RECT 45.875 152.130 46.275 152.930 ;
        RECT 47.140 152.870 47.695 153.200 ;
        RECT 47.140 152.760 47.590 152.870 ;
        RECT 46.465 152.590 47.590 152.760 ;
        RECT 47.865 152.700 48.145 153.370 ;
        RECT 46.465 152.130 46.745 152.590 ;
        RECT 47.265 151.960 47.590 152.420 ;
        RECT 47.760 152.130 48.145 152.700 ;
        RECT 48.320 153.320 48.575 154.200 ;
        RECT 48.745 153.370 49.050 154.510 ;
        RECT 49.390 154.130 49.720 154.510 ;
        RECT 49.900 153.960 50.070 154.250 ;
        RECT 50.240 154.050 50.490 154.510 ;
        RECT 49.270 153.790 50.070 153.960 ;
        RECT 50.660 154.000 51.530 154.340 ;
        RECT 48.320 152.670 48.530 153.320 ;
        RECT 49.270 153.200 49.440 153.790 ;
        RECT 50.660 153.620 50.830 154.000 ;
        RECT 51.765 153.880 51.935 154.340 ;
        RECT 52.105 154.050 52.475 154.510 ;
        RECT 52.770 153.910 52.940 154.250 ;
        RECT 53.110 154.080 53.440 154.510 ;
        RECT 53.675 153.910 53.845 154.250 ;
        RECT 49.610 153.450 50.830 153.620 ;
        RECT 51.000 153.540 51.460 153.830 ;
        RECT 51.765 153.710 52.325 153.880 ;
        RECT 52.770 153.740 53.845 153.910 ;
        RECT 54.015 154.010 54.695 154.340 ;
        RECT 54.910 154.010 55.160 154.340 ;
        RECT 55.330 154.050 55.580 154.510 ;
        RECT 52.155 153.570 52.325 153.710 ;
        RECT 51.000 153.530 51.965 153.540 ;
        RECT 50.660 153.360 50.830 153.450 ;
        RECT 51.290 153.370 51.965 153.530 ;
        RECT 48.700 153.170 49.440 153.200 ;
        RECT 48.700 152.870 49.615 153.170 ;
        RECT 49.290 152.695 49.615 152.870 ;
        RECT 48.320 152.140 48.575 152.670 ;
        RECT 48.745 151.960 49.050 152.420 ;
        RECT 49.295 152.340 49.615 152.695 ;
        RECT 49.785 152.910 50.325 153.280 ;
        RECT 50.660 153.190 51.065 153.360 ;
        RECT 49.785 152.510 50.025 152.910 ;
        RECT 50.505 152.740 50.725 153.020 ;
        RECT 50.195 152.570 50.725 152.740 ;
        RECT 50.195 152.340 50.365 152.570 ;
        RECT 50.895 152.410 51.065 153.190 ;
        RECT 51.235 152.580 51.585 153.200 ;
        RECT 51.755 152.580 51.965 153.370 ;
        RECT 52.155 153.400 53.655 153.570 ;
        RECT 52.155 152.710 52.325 153.400 ;
        RECT 54.015 153.230 54.185 154.010 ;
        RECT 54.990 153.880 55.160 154.010 ;
        RECT 52.495 153.060 54.185 153.230 ;
        RECT 54.355 153.450 54.820 153.840 ;
        RECT 54.990 153.710 55.385 153.880 ;
        RECT 52.495 152.880 52.665 153.060 ;
        RECT 49.295 152.170 50.365 152.340 ;
        RECT 50.535 151.960 50.725 152.400 ;
        RECT 50.895 152.130 51.845 152.410 ;
        RECT 52.155 152.320 52.415 152.710 ;
        RECT 52.835 152.640 53.625 152.890 ;
        RECT 52.065 152.150 52.415 152.320 ;
        RECT 52.625 151.960 52.955 152.420 ;
        RECT 53.830 152.350 54.000 153.060 ;
        RECT 54.355 152.860 54.525 153.450 ;
        RECT 54.170 152.640 54.525 152.860 ;
        RECT 54.695 152.640 55.045 153.260 ;
        RECT 55.215 152.350 55.385 153.710 ;
        RECT 55.750 153.540 56.075 154.325 ;
        RECT 55.555 152.490 56.015 153.540 ;
        RECT 53.830 152.180 54.685 152.350 ;
        RECT 54.890 152.180 55.385 152.350 ;
        RECT 55.555 151.960 55.885 152.320 ;
        RECT 56.245 152.220 56.415 154.340 ;
        RECT 56.585 154.010 56.915 154.510 ;
        RECT 57.085 153.840 57.340 154.340 ;
        RECT 56.590 153.670 57.340 153.840 ;
        RECT 56.590 152.680 56.820 153.670 ;
        RECT 56.990 152.850 57.340 153.500 ;
        RECT 57.515 153.370 57.855 154.340 ;
        RECT 58.025 153.370 58.195 154.510 ;
        RECT 58.465 153.710 58.715 154.510 ;
        RECT 59.360 153.540 59.690 154.340 ;
        RECT 59.990 153.710 60.320 154.510 ;
        RECT 60.490 153.540 60.820 154.340 ;
        RECT 61.250 153.640 61.535 154.510 ;
        RECT 61.705 153.880 61.965 154.340 ;
        RECT 62.140 154.050 62.395 154.510 ;
        RECT 62.565 153.880 62.825 154.340 ;
        RECT 61.705 153.710 62.825 153.880 ;
        RECT 62.995 153.710 63.305 154.510 ;
        RECT 58.385 153.370 60.820 153.540 ;
        RECT 61.705 153.460 61.965 153.710 ;
        RECT 62.175 153.660 62.345 153.710 ;
        RECT 63.475 153.540 63.785 154.340 ;
        RECT 57.515 152.760 57.690 153.370 ;
        RECT 58.385 153.120 58.555 153.370 ;
        RECT 57.860 152.950 58.555 153.120 ;
        RECT 58.730 152.950 59.150 153.150 ;
        RECT 59.320 152.950 59.650 153.150 ;
        RECT 59.820 152.950 60.150 153.150 ;
        RECT 56.590 152.510 57.340 152.680 ;
        RECT 56.585 151.960 56.915 152.340 ;
        RECT 57.085 152.220 57.340 152.510 ;
        RECT 57.515 152.130 57.855 152.760 ;
        RECT 58.025 151.960 58.275 152.760 ;
        RECT 58.465 152.610 59.690 152.780 ;
        RECT 58.465 152.130 58.795 152.610 ;
        RECT 58.965 151.960 59.190 152.420 ;
        RECT 59.360 152.130 59.690 152.610 ;
        RECT 60.320 152.740 60.490 153.370 ;
        RECT 61.210 153.290 61.965 153.460 ;
        RECT 62.755 153.370 63.785 153.540 ;
        RECT 60.675 152.950 61.025 153.200 ;
        RECT 61.210 152.780 61.615 153.290 ;
        RECT 62.755 153.120 62.925 153.370 ;
        RECT 61.785 152.950 62.925 153.120 ;
        RECT 60.320 152.130 60.820 152.740 ;
        RECT 61.210 152.610 62.860 152.780 ;
        RECT 63.095 152.630 63.445 153.200 ;
        RECT 61.255 151.960 61.535 152.440 ;
        RECT 61.705 152.220 61.965 152.610 ;
        RECT 62.140 151.960 62.395 152.440 ;
        RECT 62.565 152.220 62.860 152.610 ;
        RECT 63.615 152.460 63.785 153.370 ;
        RECT 63.955 153.345 64.245 154.510 ;
        RECT 64.530 153.880 64.815 154.340 ;
        RECT 64.985 154.050 65.255 154.510 ;
        RECT 64.530 153.660 65.485 153.880 ;
        RECT 64.415 152.930 65.105 153.490 ;
        RECT 65.275 152.760 65.485 153.660 ;
        RECT 63.040 151.960 63.315 152.440 ;
        RECT 63.485 152.130 63.785 152.460 ;
        RECT 63.955 151.960 64.245 152.685 ;
        RECT 64.530 152.590 65.485 152.760 ;
        RECT 65.655 153.490 66.055 154.340 ;
        RECT 66.245 153.880 66.525 154.340 ;
        RECT 67.045 154.050 67.370 154.510 ;
        RECT 66.245 153.660 67.370 153.880 ;
        RECT 65.655 152.930 66.750 153.490 ;
        RECT 66.920 153.200 67.370 153.660 ;
        RECT 67.540 153.370 67.925 154.340 ;
        RECT 64.530 152.130 64.815 152.590 ;
        RECT 64.985 151.960 65.255 152.420 ;
        RECT 65.655 152.130 66.055 152.930 ;
        RECT 66.920 152.870 67.475 153.200 ;
        RECT 66.920 152.760 67.370 152.870 ;
        RECT 66.245 152.590 67.370 152.760 ;
        RECT 67.645 152.700 67.925 153.370 ;
        RECT 66.245 152.130 66.525 152.590 ;
        RECT 67.045 151.960 67.370 152.420 ;
        RECT 67.540 152.130 67.925 152.700 ;
        RECT 68.095 153.660 68.355 154.340 ;
        RECT 68.525 153.730 68.775 154.510 ;
        RECT 69.025 153.960 69.275 154.340 ;
        RECT 69.445 154.130 69.800 154.510 ;
        RECT 70.805 154.120 71.140 154.340 ;
        RECT 70.405 153.960 70.635 154.000 ;
        RECT 69.025 153.760 70.635 153.960 ;
        RECT 69.025 153.750 69.860 153.760 ;
        RECT 70.450 153.670 70.635 153.760 ;
        RECT 68.095 152.460 68.265 153.660 ;
        RECT 69.965 153.560 70.295 153.590 ;
        RECT 68.495 153.500 70.295 153.560 ;
        RECT 70.885 153.500 71.140 154.120 ;
        RECT 68.435 153.390 71.140 153.500 ;
        RECT 68.435 153.355 68.635 153.390 ;
        RECT 68.435 152.780 68.605 153.355 ;
        RECT 69.965 153.330 71.140 153.390 ;
        RECT 71.315 153.540 71.625 154.340 ;
        RECT 71.795 153.710 72.105 154.510 ;
        RECT 72.275 153.880 72.535 154.340 ;
        RECT 72.705 154.050 72.960 154.510 ;
        RECT 73.135 153.880 73.395 154.340 ;
        RECT 72.275 153.710 73.395 153.880 ;
        RECT 71.315 153.370 72.345 153.540 ;
        RECT 68.835 152.915 69.245 153.220 ;
        RECT 69.415 152.950 69.745 153.160 ;
        RECT 68.435 152.660 68.705 152.780 ;
        RECT 68.435 152.615 69.280 152.660 ;
        RECT 68.525 152.490 69.280 152.615 ;
        RECT 69.535 152.550 69.745 152.950 ;
        RECT 69.990 152.950 70.465 153.160 ;
        RECT 70.655 152.950 71.145 153.150 ;
        RECT 69.990 152.550 70.210 152.950 ;
        RECT 68.095 152.130 68.355 152.460 ;
        RECT 69.110 152.340 69.280 152.490 ;
        RECT 68.525 151.960 68.855 152.320 ;
        RECT 69.110 152.130 70.410 152.340 ;
        RECT 70.685 151.960 71.140 152.725 ;
        RECT 71.315 152.460 71.485 153.370 ;
        RECT 71.655 152.630 72.005 153.200 ;
        RECT 72.175 153.120 72.345 153.370 ;
        RECT 73.135 153.460 73.395 153.710 ;
        RECT 73.565 153.640 73.850 154.510 ;
        RECT 74.165 153.580 74.335 154.340 ;
        RECT 74.550 153.750 74.880 154.510 ;
        RECT 73.135 153.290 73.890 153.460 ;
        RECT 74.165 153.410 74.880 153.580 ;
        RECT 75.050 153.435 75.305 154.340 ;
        RECT 72.175 152.950 73.315 153.120 ;
        RECT 73.485 152.780 73.890 153.290 ;
        RECT 74.075 152.860 74.430 153.230 ;
        RECT 74.710 153.200 74.880 153.410 ;
        RECT 74.710 152.870 74.965 153.200 ;
        RECT 72.240 152.610 73.890 152.780 ;
        RECT 74.710 152.680 74.880 152.870 ;
        RECT 75.135 152.705 75.305 153.435 ;
        RECT 75.480 153.360 75.740 154.510 ;
        RECT 76.435 153.370 76.645 154.510 ;
        RECT 76.815 153.360 77.145 154.340 ;
        RECT 77.315 153.370 77.545 154.510 ;
        RECT 77.755 153.750 78.270 154.160 ;
        RECT 78.505 153.750 78.675 154.510 ;
        RECT 78.845 154.170 80.875 154.340 ;
        RECT 71.315 152.130 71.615 152.460 ;
        RECT 71.785 151.960 72.060 152.440 ;
        RECT 72.240 152.220 72.535 152.610 ;
        RECT 72.705 151.960 72.960 152.440 ;
        RECT 73.135 152.220 73.395 152.610 ;
        RECT 74.165 152.510 74.880 152.680 ;
        RECT 73.565 151.960 73.845 152.440 ;
        RECT 74.165 152.130 74.335 152.510 ;
        RECT 74.550 151.960 74.880 152.340 ;
        RECT 75.050 152.130 75.305 152.705 ;
        RECT 75.480 151.960 75.740 152.800 ;
        RECT 76.435 151.960 76.645 152.780 ;
        RECT 76.815 152.760 77.065 153.360 ;
        RECT 77.235 152.950 77.565 153.200 ;
        RECT 77.755 152.940 78.095 153.750 ;
        RECT 78.845 153.505 79.015 154.170 ;
        RECT 79.410 153.830 80.535 154.000 ;
        RECT 78.265 153.315 79.015 153.505 ;
        RECT 79.185 153.490 80.195 153.660 ;
        RECT 76.815 152.130 77.145 152.760 ;
        RECT 77.315 151.960 77.545 152.780 ;
        RECT 77.755 152.770 78.985 152.940 ;
        RECT 78.030 152.165 78.275 152.770 ;
        RECT 78.495 151.960 79.005 152.495 ;
        RECT 79.185 152.130 79.375 153.490 ;
        RECT 79.545 152.470 79.820 153.290 ;
        RECT 80.025 152.690 80.195 153.490 ;
        RECT 80.365 152.700 80.535 153.830 ;
        RECT 80.705 153.200 80.875 154.170 ;
        RECT 81.045 153.370 81.215 154.510 ;
        RECT 81.385 153.370 81.720 154.340 ;
        RECT 82.445 153.580 82.615 154.340 ;
        RECT 82.795 153.750 83.125 154.510 ;
        RECT 82.445 153.410 83.110 153.580 ;
        RECT 83.295 153.435 83.565 154.340 ;
        RECT 80.705 152.870 80.900 153.200 ;
        RECT 81.125 152.870 81.380 153.200 ;
        RECT 81.125 152.700 81.295 152.870 ;
        RECT 81.550 152.700 81.720 153.370 ;
        RECT 82.940 153.265 83.110 153.410 ;
        RECT 82.375 152.860 82.705 153.230 ;
        RECT 82.940 152.935 83.225 153.265 ;
        RECT 80.365 152.530 81.295 152.700 ;
        RECT 80.365 152.495 80.540 152.530 ;
        RECT 79.545 152.300 79.825 152.470 ;
        RECT 79.545 152.130 79.820 152.300 ;
        RECT 80.010 152.130 80.540 152.495 ;
        RECT 80.965 151.960 81.295 152.360 ;
        RECT 81.465 152.130 81.720 152.700 ;
        RECT 82.940 152.680 83.110 152.935 ;
        RECT 82.445 152.510 83.110 152.680 ;
        RECT 83.395 152.635 83.565 153.435 ;
        RECT 84.655 153.750 85.170 154.160 ;
        RECT 85.405 153.750 85.575 154.510 ;
        RECT 85.745 154.170 87.775 154.340 ;
        RECT 84.655 152.940 84.995 153.750 ;
        RECT 85.745 153.505 85.915 154.170 ;
        RECT 86.310 153.830 87.435 154.000 ;
        RECT 85.165 153.315 85.915 153.505 ;
        RECT 86.085 153.490 87.095 153.660 ;
        RECT 84.655 152.770 85.885 152.940 ;
        RECT 82.445 152.130 82.615 152.510 ;
        RECT 82.795 151.960 83.125 152.340 ;
        RECT 83.305 152.130 83.565 152.635 ;
        RECT 84.930 152.165 85.175 152.770 ;
        RECT 85.395 151.960 85.905 152.495 ;
        RECT 86.085 152.130 86.275 153.490 ;
        RECT 86.445 153.150 86.720 153.290 ;
        RECT 86.445 152.980 86.725 153.150 ;
        RECT 86.445 152.130 86.720 152.980 ;
        RECT 86.925 152.690 87.095 153.490 ;
        RECT 87.265 152.700 87.435 153.830 ;
        RECT 87.605 153.200 87.775 154.170 ;
        RECT 87.945 153.370 88.115 154.510 ;
        RECT 88.285 153.370 88.620 154.340 ;
        RECT 87.605 152.870 87.800 153.200 ;
        RECT 88.025 152.870 88.280 153.200 ;
        RECT 88.025 152.700 88.195 152.870 ;
        RECT 88.450 152.700 88.620 153.370 ;
        RECT 89.715 153.345 90.005 154.510 ;
        RECT 90.635 153.420 92.305 154.510 ;
        RECT 90.635 152.900 91.385 153.420 ;
        RECT 92.475 153.370 92.815 154.340 ;
        RECT 92.985 153.370 93.155 154.510 ;
        RECT 93.425 153.710 93.675 154.510 ;
        RECT 94.320 153.540 94.650 154.340 ;
        RECT 94.950 153.710 95.280 154.510 ;
        RECT 95.450 153.540 95.780 154.340 ;
        RECT 93.345 153.370 95.780 153.540 ;
        RECT 96.155 153.370 96.495 154.340 ;
        RECT 96.665 153.370 96.835 154.510 ;
        RECT 97.105 153.710 97.355 154.510 ;
        RECT 98.000 153.540 98.330 154.340 ;
        RECT 98.630 153.710 98.960 154.510 ;
        RECT 99.130 153.540 99.460 154.340 ;
        RECT 97.025 153.370 99.460 153.540 ;
        RECT 99.835 153.420 101.045 154.510 ;
        RECT 101.215 153.750 101.730 154.160 ;
        RECT 101.965 153.750 102.135 154.510 ;
        RECT 102.305 154.170 104.335 154.340 ;
        RECT 91.555 152.730 92.305 153.250 ;
        RECT 87.265 152.530 88.195 152.700 ;
        RECT 87.265 152.495 87.440 152.530 ;
        RECT 86.910 152.130 87.440 152.495 ;
        RECT 87.865 151.960 88.195 152.360 ;
        RECT 88.365 152.130 88.620 152.700 ;
        RECT 89.715 151.960 90.005 152.685 ;
        RECT 90.635 151.960 92.305 152.730 ;
        RECT 92.475 152.760 92.650 153.370 ;
        RECT 93.345 153.120 93.515 153.370 ;
        RECT 92.820 152.950 93.515 153.120 ;
        RECT 93.690 152.950 94.110 153.150 ;
        RECT 94.280 152.950 94.610 153.150 ;
        RECT 94.780 152.950 95.110 153.150 ;
        RECT 92.475 152.130 92.815 152.760 ;
        RECT 92.985 151.960 93.235 152.760 ;
        RECT 93.425 152.610 94.650 152.780 ;
        RECT 93.425 152.130 93.755 152.610 ;
        RECT 93.925 151.960 94.150 152.420 ;
        RECT 94.320 152.130 94.650 152.610 ;
        RECT 95.280 152.740 95.450 153.370 ;
        RECT 95.635 152.950 95.985 153.200 ;
        RECT 96.155 152.760 96.330 153.370 ;
        RECT 97.025 153.120 97.195 153.370 ;
        RECT 96.500 152.950 97.195 153.120 ;
        RECT 97.370 152.950 97.790 153.150 ;
        RECT 97.960 152.950 98.290 153.150 ;
        RECT 98.460 152.950 98.790 153.150 ;
        RECT 95.280 152.130 95.780 152.740 ;
        RECT 96.155 152.130 96.495 152.760 ;
        RECT 96.665 151.960 96.915 152.760 ;
        RECT 97.105 152.610 98.330 152.780 ;
        RECT 97.105 152.130 97.435 152.610 ;
        RECT 97.605 151.960 97.830 152.420 ;
        RECT 98.000 152.130 98.330 152.610 ;
        RECT 98.960 152.740 99.130 153.370 ;
        RECT 99.315 152.950 99.665 153.200 ;
        RECT 99.835 152.880 100.355 153.420 ;
        RECT 98.960 152.130 99.460 152.740 ;
        RECT 100.525 152.710 101.045 153.250 ;
        RECT 101.215 152.940 101.555 153.750 ;
        RECT 102.305 153.505 102.475 154.170 ;
        RECT 102.870 153.830 103.995 154.000 ;
        RECT 101.725 153.315 102.475 153.505 ;
        RECT 102.645 153.490 103.655 153.660 ;
        RECT 101.215 152.770 102.445 152.940 ;
        RECT 99.835 151.960 101.045 152.710 ;
        RECT 101.490 152.165 101.735 152.770 ;
        RECT 101.955 151.960 102.465 152.495 ;
        RECT 102.645 152.130 102.835 153.490 ;
        RECT 103.005 152.810 103.280 153.290 ;
        RECT 103.005 152.640 103.285 152.810 ;
        RECT 103.485 152.690 103.655 153.490 ;
        RECT 103.825 152.700 103.995 153.830 ;
        RECT 104.165 153.200 104.335 154.170 ;
        RECT 104.505 153.370 104.675 154.510 ;
        RECT 104.845 153.370 105.180 154.340 ;
        RECT 104.165 152.870 104.360 153.200 ;
        RECT 104.585 152.870 104.840 153.200 ;
        RECT 104.585 152.700 104.755 152.870 ;
        RECT 105.010 152.700 105.180 153.370 ;
        RECT 103.005 152.130 103.280 152.640 ;
        RECT 103.825 152.530 104.755 152.700 ;
        RECT 103.825 152.495 104.000 152.530 ;
        RECT 103.470 152.130 104.000 152.495 ;
        RECT 104.425 151.960 104.755 152.360 ;
        RECT 104.925 152.130 105.180 152.700 ;
        RECT 105.360 153.320 105.615 154.200 ;
        RECT 105.785 153.370 106.090 154.510 ;
        RECT 106.430 154.130 106.760 154.510 ;
        RECT 106.940 153.960 107.110 154.250 ;
        RECT 107.280 154.050 107.530 154.510 ;
        RECT 106.310 153.790 107.110 153.960 ;
        RECT 107.700 154.000 108.570 154.340 ;
        RECT 105.360 152.670 105.570 153.320 ;
        RECT 106.310 153.200 106.480 153.790 ;
        RECT 107.700 153.620 107.870 154.000 ;
        RECT 108.805 153.880 108.975 154.340 ;
        RECT 109.145 154.050 109.515 154.510 ;
        RECT 109.810 153.910 109.980 154.250 ;
        RECT 110.150 154.080 110.480 154.510 ;
        RECT 110.715 153.910 110.885 154.250 ;
        RECT 106.650 153.450 107.870 153.620 ;
        RECT 108.040 153.540 108.500 153.830 ;
        RECT 108.805 153.710 109.365 153.880 ;
        RECT 109.810 153.740 110.885 153.910 ;
        RECT 111.055 154.010 111.735 154.340 ;
        RECT 111.950 154.010 112.200 154.340 ;
        RECT 112.370 154.050 112.620 154.510 ;
        RECT 109.195 153.570 109.365 153.710 ;
        RECT 108.040 153.530 109.005 153.540 ;
        RECT 107.700 153.360 107.870 153.450 ;
        RECT 108.330 153.370 109.005 153.530 ;
        RECT 105.740 153.170 106.480 153.200 ;
        RECT 105.740 152.870 106.655 153.170 ;
        RECT 106.330 152.695 106.655 152.870 ;
        RECT 105.360 152.140 105.615 152.670 ;
        RECT 105.785 151.960 106.090 152.420 ;
        RECT 106.335 152.340 106.655 152.695 ;
        RECT 106.825 152.910 107.365 153.280 ;
        RECT 107.700 153.190 108.105 153.360 ;
        RECT 106.825 152.510 107.065 152.910 ;
        RECT 107.545 152.740 107.765 153.020 ;
        RECT 107.235 152.570 107.765 152.740 ;
        RECT 107.235 152.340 107.405 152.570 ;
        RECT 107.935 152.410 108.105 153.190 ;
        RECT 108.275 152.580 108.625 153.200 ;
        RECT 108.795 152.580 109.005 153.370 ;
        RECT 109.195 153.400 110.695 153.570 ;
        RECT 109.195 152.710 109.365 153.400 ;
        RECT 111.055 153.230 111.225 154.010 ;
        RECT 112.030 153.880 112.200 154.010 ;
        RECT 109.535 153.060 111.225 153.230 ;
        RECT 111.395 153.450 111.860 153.840 ;
        RECT 112.030 153.710 112.425 153.880 ;
        RECT 109.535 152.880 109.705 153.060 ;
        RECT 106.335 152.170 107.405 152.340 ;
        RECT 107.575 151.960 107.765 152.400 ;
        RECT 107.935 152.130 108.885 152.410 ;
        RECT 109.195 152.320 109.455 152.710 ;
        RECT 109.875 152.640 110.665 152.890 ;
        RECT 109.105 152.150 109.455 152.320 ;
        RECT 109.665 151.960 109.995 152.420 ;
        RECT 110.870 152.350 111.040 153.060 ;
        RECT 111.395 152.860 111.565 153.450 ;
        RECT 111.210 152.640 111.565 152.860 ;
        RECT 111.735 152.640 112.085 153.260 ;
        RECT 112.255 152.350 112.425 153.710 ;
        RECT 112.790 153.540 113.115 154.325 ;
        RECT 112.595 152.490 113.055 153.540 ;
        RECT 110.870 152.180 111.725 152.350 ;
        RECT 111.930 152.180 112.425 152.350 ;
        RECT 112.595 151.960 112.925 152.320 ;
        RECT 113.285 152.220 113.455 154.340 ;
        RECT 113.625 154.010 113.955 154.510 ;
        RECT 114.125 153.840 114.380 154.340 ;
        RECT 113.630 153.670 114.380 153.840 ;
        RECT 113.630 152.680 113.860 153.670 ;
        RECT 114.030 152.850 114.380 153.500 ;
        RECT 114.555 153.420 115.765 154.510 ;
        RECT 114.555 152.880 115.075 153.420 ;
        RECT 115.245 152.710 115.765 153.250 ;
        RECT 113.630 152.510 114.380 152.680 ;
        RECT 113.625 151.960 113.955 152.340 ;
        RECT 114.125 152.220 114.380 152.510 ;
        RECT 114.555 151.960 115.765 152.710 ;
        RECT 14.650 151.790 115.850 151.960 ;
        RECT 14.735 151.040 15.945 151.790 ;
        RECT 14.735 150.500 15.255 151.040 ;
        RECT 16.115 151.020 19.625 151.790 ;
        RECT 15.425 150.330 15.945 150.870 ;
        RECT 14.735 149.240 15.945 150.330 ;
        RECT 16.115 150.330 17.805 150.850 ;
        RECT 17.975 150.500 19.625 151.020 ;
        RECT 19.835 150.970 20.065 151.790 ;
        RECT 20.235 150.990 20.565 151.620 ;
        RECT 19.815 150.550 20.145 150.800 ;
        RECT 20.315 150.390 20.565 150.990 ;
        RECT 20.735 150.970 20.945 151.790 ;
        RECT 21.180 151.050 21.435 151.620 ;
        RECT 21.605 151.390 21.935 151.790 ;
        RECT 22.360 151.255 22.890 151.620 ;
        RECT 22.360 151.220 22.535 151.255 ;
        RECT 21.605 151.050 22.535 151.220 ;
        RECT 16.115 149.240 19.625 150.330 ;
        RECT 19.835 149.240 20.065 150.380 ;
        RECT 20.235 149.410 20.565 150.390 ;
        RECT 21.180 150.380 21.350 151.050 ;
        RECT 21.605 150.880 21.775 151.050 ;
        RECT 21.520 150.550 21.775 150.880 ;
        RECT 22.000 150.550 22.195 150.880 ;
        RECT 20.735 149.240 20.945 150.380 ;
        RECT 21.180 149.410 21.515 150.380 ;
        RECT 21.685 149.240 21.855 150.380 ;
        RECT 22.025 149.580 22.195 150.550 ;
        RECT 22.365 149.920 22.535 151.050 ;
        RECT 22.705 150.260 22.875 151.060 ;
        RECT 23.080 150.770 23.355 151.620 ;
        RECT 23.075 150.600 23.355 150.770 ;
        RECT 23.080 150.460 23.355 150.600 ;
        RECT 23.525 150.260 23.715 151.620 ;
        RECT 23.895 151.255 24.405 151.790 ;
        RECT 24.625 150.980 24.870 151.585 ;
        RECT 25.315 151.065 25.605 151.790 ;
        RECT 25.775 151.040 26.985 151.790 ;
        RECT 23.915 150.810 25.145 150.980 ;
        RECT 22.705 150.090 23.715 150.260 ;
        RECT 23.885 150.245 24.635 150.435 ;
        RECT 22.365 149.750 23.490 149.920 ;
        RECT 23.885 149.580 24.055 150.245 ;
        RECT 24.805 150.000 25.145 150.810 ;
        RECT 22.025 149.410 24.055 149.580 ;
        RECT 24.225 149.240 24.395 150.000 ;
        RECT 24.630 149.590 25.145 150.000 ;
        RECT 25.315 149.240 25.605 150.405 ;
        RECT 25.775 150.330 26.295 150.870 ;
        RECT 26.465 150.500 26.985 151.040 ;
        RECT 27.195 150.970 27.425 151.790 ;
        RECT 27.595 150.990 27.925 151.620 ;
        RECT 27.175 150.550 27.505 150.800 ;
        RECT 27.675 150.390 27.925 150.990 ;
        RECT 28.095 150.970 28.305 151.790 ;
        RECT 29.730 150.980 29.975 151.585 ;
        RECT 30.195 151.255 30.705 151.790 ;
        RECT 25.775 149.240 26.985 150.330 ;
        RECT 27.195 149.240 27.425 150.380 ;
        RECT 27.595 149.410 27.925 150.390 ;
        RECT 29.455 150.810 30.685 150.980 ;
        RECT 28.095 149.240 28.305 150.380 ;
        RECT 29.455 150.000 29.795 150.810 ;
        RECT 29.965 150.245 30.715 150.435 ;
        RECT 29.455 149.590 29.970 150.000 ;
        RECT 30.205 149.240 30.375 150.000 ;
        RECT 30.545 149.580 30.715 150.245 ;
        RECT 30.885 150.260 31.075 151.620 ;
        RECT 31.245 151.110 31.520 151.620 ;
        RECT 31.710 151.255 32.240 151.620 ;
        RECT 32.665 151.390 32.995 151.790 ;
        RECT 32.065 151.220 32.240 151.255 ;
        RECT 31.245 150.940 31.525 151.110 ;
        RECT 31.245 150.460 31.520 150.940 ;
        RECT 31.725 150.260 31.895 151.060 ;
        RECT 30.885 150.090 31.895 150.260 ;
        RECT 32.065 151.050 32.995 151.220 ;
        RECT 33.165 151.050 33.420 151.620 ;
        RECT 32.065 149.920 32.235 151.050 ;
        RECT 32.825 150.880 32.995 151.050 ;
        RECT 31.110 149.750 32.235 149.920 ;
        RECT 32.405 150.550 32.600 150.880 ;
        RECT 32.825 150.550 33.080 150.880 ;
        RECT 32.405 149.580 32.575 150.550 ;
        RECT 33.250 150.380 33.420 151.050 ;
        RECT 30.545 149.410 32.575 149.580 ;
        RECT 32.745 149.240 32.915 150.380 ;
        RECT 33.085 149.410 33.420 150.380 ;
        RECT 33.595 150.990 33.935 151.620 ;
        RECT 34.105 150.990 34.355 151.790 ;
        RECT 34.545 151.140 34.875 151.620 ;
        RECT 35.045 151.330 35.270 151.790 ;
        RECT 35.440 151.140 35.770 151.620 ;
        RECT 33.595 150.380 33.770 150.990 ;
        RECT 34.545 150.970 35.770 151.140 ;
        RECT 36.400 151.010 36.900 151.620 ;
        RECT 37.275 151.020 38.945 151.790 ;
        RECT 39.125 151.290 39.455 151.790 ;
        RECT 39.655 151.220 39.825 151.570 ;
        RECT 40.025 151.390 40.355 151.790 ;
        RECT 40.525 151.220 40.695 151.570 ;
        RECT 40.865 151.390 41.245 151.790 ;
        RECT 33.940 150.630 34.635 150.800 ;
        RECT 34.465 150.380 34.635 150.630 ;
        RECT 34.810 150.600 35.230 150.800 ;
        RECT 35.400 150.600 35.730 150.800 ;
        RECT 35.900 150.600 36.230 150.800 ;
        RECT 36.400 150.380 36.570 151.010 ;
        RECT 36.755 150.550 37.105 150.800 ;
        RECT 33.595 149.410 33.935 150.380 ;
        RECT 34.105 149.240 34.275 150.380 ;
        RECT 34.465 150.210 36.900 150.380 ;
        RECT 34.545 149.240 34.795 150.040 ;
        RECT 35.440 149.410 35.770 150.210 ;
        RECT 36.070 149.240 36.400 150.040 ;
        RECT 36.570 149.410 36.900 150.210 ;
        RECT 37.275 150.330 38.025 150.850 ;
        RECT 38.195 150.500 38.945 151.020 ;
        RECT 39.120 150.550 39.470 151.120 ;
        RECT 39.655 151.050 41.265 151.220 ;
        RECT 41.435 151.115 41.705 151.460 ;
        RECT 41.095 150.880 41.265 151.050 ;
        RECT 37.275 149.240 38.945 150.330 ;
        RECT 39.120 150.090 39.440 150.380 ;
        RECT 39.640 150.260 40.350 150.880 ;
        RECT 40.520 150.550 40.925 150.880 ;
        RECT 41.095 150.550 41.365 150.880 ;
        RECT 41.095 150.380 41.265 150.550 ;
        RECT 41.535 150.380 41.705 151.115 ;
        RECT 40.540 150.210 41.265 150.380 ;
        RECT 40.540 150.090 40.710 150.210 ;
        RECT 39.120 149.920 40.710 150.090 ;
        RECT 39.120 149.460 40.775 149.750 ;
        RECT 40.945 149.240 41.225 150.040 ;
        RECT 41.435 149.410 41.705 150.380 ;
        RECT 41.875 150.990 42.215 151.620 ;
        RECT 42.385 150.990 42.635 151.790 ;
        RECT 42.825 151.140 43.155 151.620 ;
        RECT 43.325 151.330 43.550 151.790 ;
        RECT 43.720 151.140 44.050 151.620 ;
        RECT 41.875 150.940 42.105 150.990 ;
        RECT 42.825 150.970 44.050 151.140 ;
        RECT 44.680 151.010 45.180 151.620 ;
        RECT 41.875 150.380 42.050 150.940 ;
        RECT 42.220 150.630 42.915 150.800 ;
        RECT 42.745 150.380 42.915 150.630 ;
        RECT 43.090 150.600 43.510 150.800 ;
        RECT 43.680 150.600 44.010 150.800 ;
        RECT 44.180 150.600 44.510 150.800 ;
        RECT 44.680 150.380 44.850 151.010 ;
        RECT 45.830 150.980 46.075 151.585 ;
        RECT 46.295 151.255 46.805 151.790 ;
        RECT 45.555 150.810 46.785 150.980 ;
        RECT 45.035 150.550 45.385 150.800 ;
        RECT 41.875 149.410 42.215 150.380 ;
        RECT 42.385 149.240 42.555 150.380 ;
        RECT 42.745 150.210 45.180 150.380 ;
        RECT 42.825 149.240 43.075 150.040 ;
        RECT 43.720 149.410 44.050 150.210 ;
        RECT 44.350 149.240 44.680 150.040 ;
        RECT 44.850 149.410 45.180 150.210 ;
        RECT 45.555 150.000 45.895 150.810 ;
        RECT 46.065 150.245 46.815 150.435 ;
        RECT 45.555 149.590 46.070 150.000 ;
        RECT 46.305 149.240 46.475 150.000 ;
        RECT 46.645 149.580 46.815 150.245 ;
        RECT 46.985 150.260 47.175 151.620 ;
        RECT 47.345 151.110 47.620 151.620 ;
        RECT 47.810 151.255 48.340 151.620 ;
        RECT 48.765 151.390 49.095 151.790 ;
        RECT 48.165 151.220 48.340 151.255 ;
        RECT 47.345 150.940 47.625 151.110 ;
        RECT 47.345 150.460 47.620 150.940 ;
        RECT 47.825 150.260 47.995 151.060 ;
        RECT 46.985 150.090 47.995 150.260 ;
        RECT 48.165 151.050 49.095 151.220 ;
        RECT 49.265 151.050 49.520 151.620 ;
        RECT 48.165 149.920 48.335 151.050 ;
        RECT 48.925 150.880 49.095 151.050 ;
        RECT 47.210 149.750 48.335 149.920 ;
        RECT 48.505 150.550 48.700 150.880 ;
        RECT 48.925 150.550 49.180 150.880 ;
        RECT 48.505 149.580 48.675 150.550 ;
        RECT 49.350 150.380 49.520 151.050 ;
        RECT 49.695 151.040 50.905 151.790 ;
        RECT 51.075 151.065 51.365 151.790 ;
        RECT 46.645 149.410 48.675 149.580 ;
        RECT 48.845 149.240 49.015 150.380 ;
        RECT 49.185 149.410 49.520 150.380 ;
        RECT 49.695 150.330 50.215 150.870 ;
        RECT 50.385 150.500 50.905 151.040 ;
        RECT 52.460 151.050 52.715 151.620 ;
        RECT 52.885 151.390 53.215 151.790 ;
        RECT 53.640 151.255 54.170 151.620 ;
        RECT 54.360 151.450 54.635 151.620 ;
        RECT 54.355 151.280 54.635 151.450 ;
        RECT 53.640 151.220 53.815 151.255 ;
        RECT 52.885 151.050 53.815 151.220 ;
        RECT 49.695 149.240 50.905 150.330 ;
        RECT 51.075 149.240 51.365 150.405 ;
        RECT 52.460 150.380 52.630 151.050 ;
        RECT 52.885 150.880 53.055 151.050 ;
        RECT 52.800 150.550 53.055 150.880 ;
        RECT 53.280 150.550 53.475 150.880 ;
        RECT 52.460 149.410 52.795 150.380 ;
        RECT 52.965 149.240 53.135 150.380 ;
        RECT 53.305 149.580 53.475 150.550 ;
        RECT 53.645 149.920 53.815 151.050 ;
        RECT 53.985 150.260 54.155 151.060 ;
        RECT 54.360 150.460 54.635 151.280 ;
        RECT 54.805 150.260 54.995 151.620 ;
        RECT 55.175 151.255 55.685 151.790 ;
        RECT 55.905 150.980 56.150 151.585 ;
        RECT 56.595 151.020 59.185 151.790 ;
        RECT 55.195 150.810 56.425 150.980 ;
        RECT 53.985 150.090 54.995 150.260 ;
        RECT 55.165 150.245 55.915 150.435 ;
        RECT 53.645 149.750 54.770 149.920 ;
        RECT 55.165 149.580 55.335 150.245 ;
        RECT 56.085 150.000 56.425 150.810 ;
        RECT 53.305 149.410 55.335 149.580 ;
        RECT 55.505 149.240 55.675 150.000 ;
        RECT 55.910 149.590 56.425 150.000 ;
        RECT 56.595 150.330 57.805 150.850 ;
        RECT 57.975 150.500 59.185 151.020 ;
        RECT 59.730 151.080 59.985 151.610 ;
        RECT 60.165 151.330 60.450 151.790 ;
        RECT 56.595 149.240 59.185 150.330 ;
        RECT 59.730 150.220 59.910 151.080 ;
        RECT 60.630 150.880 60.880 151.530 ;
        RECT 60.080 150.550 60.880 150.880 ;
        RECT 59.730 149.750 59.985 150.220 ;
        RECT 59.645 149.580 59.985 149.750 ;
        RECT 59.730 149.550 59.985 149.580 ;
        RECT 60.165 149.240 60.450 150.040 ;
        RECT 60.630 149.960 60.880 150.550 ;
        RECT 61.080 151.195 61.400 151.525 ;
        RECT 61.580 151.310 62.240 151.790 ;
        RECT 62.440 151.400 63.290 151.570 ;
        RECT 61.080 150.300 61.270 151.195 ;
        RECT 61.590 150.870 62.250 151.140 ;
        RECT 61.920 150.810 62.250 150.870 ;
        RECT 61.440 150.640 61.770 150.700 ;
        RECT 62.440 150.640 62.610 151.400 ;
        RECT 63.850 151.330 64.170 151.790 ;
        RECT 64.370 151.150 64.620 151.580 ;
        RECT 64.910 151.350 65.320 151.790 ;
        RECT 65.490 151.410 66.505 151.610 ;
        RECT 62.780 150.980 64.030 151.150 ;
        RECT 62.780 150.860 63.110 150.980 ;
        RECT 61.440 150.470 63.340 150.640 ;
        RECT 61.080 150.130 63.000 150.300 ;
        RECT 61.080 150.110 61.400 150.130 ;
        RECT 60.630 149.450 60.960 149.960 ;
        RECT 61.230 149.500 61.400 150.110 ;
        RECT 63.170 149.960 63.340 150.470 ;
        RECT 63.510 150.400 63.690 150.810 ;
        RECT 63.860 150.220 64.030 150.980 ;
        RECT 61.570 149.240 61.900 149.930 ;
        RECT 62.130 149.790 63.340 149.960 ;
        RECT 63.510 149.910 64.030 150.220 ;
        RECT 64.200 150.810 64.620 151.150 ;
        RECT 64.910 150.810 65.320 151.140 ;
        RECT 64.200 150.040 64.390 150.810 ;
        RECT 65.490 150.680 65.660 151.410 ;
        RECT 66.805 151.240 66.975 151.570 ;
        RECT 67.145 151.410 67.475 151.790 ;
        RECT 65.830 150.860 66.180 151.230 ;
        RECT 65.490 150.640 65.910 150.680 ;
        RECT 64.560 150.470 65.910 150.640 ;
        RECT 64.560 150.310 64.810 150.470 ;
        RECT 65.320 150.040 65.570 150.300 ;
        RECT 64.200 149.790 65.570 150.040 ;
        RECT 62.130 149.500 62.370 149.790 ;
        RECT 63.170 149.710 63.340 149.790 ;
        RECT 62.570 149.240 62.990 149.620 ;
        RECT 63.170 149.460 63.800 149.710 ;
        RECT 64.270 149.240 64.600 149.620 ;
        RECT 64.770 149.500 64.940 149.790 ;
        RECT 65.740 149.625 65.910 150.470 ;
        RECT 66.360 150.300 66.580 151.170 ;
        RECT 66.805 151.050 67.500 151.240 ;
        RECT 66.080 149.920 66.580 150.300 ;
        RECT 66.750 150.250 67.160 150.870 ;
        RECT 67.330 150.080 67.500 151.050 ;
        RECT 66.805 149.910 67.500 150.080 ;
        RECT 65.120 149.240 65.500 149.620 ;
        RECT 65.740 149.455 66.570 149.625 ;
        RECT 66.805 149.410 66.975 149.910 ;
        RECT 67.145 149.240 67.475 149.740 ;
        RECT 67.690 149.410 67.915 151.530 ;
        RECT 68.085 151.410 68.415 151.790 ;
        RECT 68.585 151.240 68.755 151.530 ;
        RECT 68.090 151.070 68.755 151.240 ;
        RECT 69.935 151.115 70.205 151.460 ;
        RECT 70.395 151.390 70.775 151.790 ;
        RECT 70.945 151.220 71.115 151.570 ;
        RECT 71.285 151.390 71.615 151.790 ;
        RECT 71.815 151.220 71.985 151.570 ;
        RECT 72.185 151.290 72.515 151.790 ;
        RECT 68.090 150.080 68.320 151.070 ;
        RECT 68.490 150.250 68.840 150.900 ;
        RECT 69.935 150.380 70.105 151.115 ;
        RECT 70.375 151.050 71.985 151.220 ;
        RECT 70.375 150.880 70.545 151.050 ;
        RECT 70.275 150.550 70.545 150.880 ;
        RECT 70.715 150.550 71.120 150.880 ;
        RECT 70.375 150.380 70.545 150.550 ;
        RECT 68.090 149.910 68.755 150.080 ;
        RECT 68.085 149.240 68.415 149.740 ;
        RECT 68.585 149.410 68.755 149.910 ;
        RECT 69.935 149.410 70.205 150.380 ;
        RECT 70.375 150.210 71.100 150.380 ;
        RECT 71.290 150.260 72.000 150.880 ;
        RECT 72.170 150.550 72.520 151.120 ;
        RECT 72.695 150.990 73.035 151.620 ;
        RECT 73.205 150.990 73.455 151.790 ;
        RECT 73.645 151.140 73.975 151.620 ;
        RECT 74.145 151.330 74.370 151.790 ;
        RECT 74.540 151.140 74.870 151.620 ;
        RECT 72.695 150.940 72.925 150.990 ;
        RECT 73.645 150.970 74.870 151.140 ;
        RECT 75.500 151.010 76.000 151.620 ;
        RECT 76.835 151.065 77.125 151.790 ;
        RECT 77.670 151.450 77.925 151.610 ;
        RECT 77.585 151.280 77.925 151.450 ;
        RECT 78.105 151.330 78.390 151.790 ;
        RECT 77.670 151.080 77.925 151.280 ;
        RECT 72.695 150.380 72.870 150.940 ;
        RECT 73.040 150.630 73.735 150.800 ;
        RECT 73.565 150.380 73.735 150.630 ;
        RECT 73.910 150.600 74.330 150.800 ;
        RECT 74.500 150.600 74.830 150.800 ;
        RECT 75.000 150.600 75.330 150.800 ;
        RECT 75.500 150.380 75.670 151.010 ;
        RECT 75.855 150.550 76.205 150.800 ;
        RECT 70.930 150.090 71.100 150.210 ;
        RECT 72.200 150.090 72.520 150.380 ;
        RECT 70.415 149.240 70.695 150.040 ;
        RECT 70.930 149.920 72.520 150.090 ;
        RECT 70.865 149.460 72.520 149.750 ;
        RECT 72.695 149.410 73.035 150.380 ;
        RECT 73.205 149.240 73.375 150.380 ;
        RECT 73.565 150.210 76.000 150.380 ;
        RECT 73.645 149.240 73.895 150.040 ;
        RECT 74.540 149.410 74.870 150.210 ;
        RECT 75.170 149.240 75.500 150.040 ;
        RECT 75.670 149.410 76.000 150.210 ;
        RECT 76.835 149.240 77.125 150.405 ;
        RECT 77.670 150.220 77.850 151.080 ;
        RECT 78.570 150.880 78.820 151.530 ;
        RECT 78.020 150.550 78.820 150.880 ;
        RECT 77.670 149.550 77.925 150.220 ;
        RECT 78.105 149.240 78.390 150.040 ;
        RECT 78.570 149.960 78.820 150.550 ;
        RECT 79.020 151.195 79.340 151.525 ;
        RECT 79.520 151.310 80.180 151.790 ;
        RECT 80.380 151.400 81.230 151.570 ;
        RECT 79.020 150.300 79.210 151.195 ;
        RECT 79.530 150.870 80.190 151.140 ;
        RECT 79.860 150.810 80.190 150.870 ;
        RECT 79.380 150.640 79.710 150.700 ;
        RECT 80.380 150.640 80.550 151.400 ;
        RECT 81.790 151.330 82.110 151.790 ;
        RECT 82.310 151.150 82.560 151.580 ;
        RECT 82.850 151.350 83.260 151.790 ;
        RECT 83.430 151.410 84.445 151.610 ;
        RECT 80.720 150.980 81.970 151.150 ;
        RECT 80.720 150.860 81.050 150.980 ;
        RECT 79.380 150.470 81.280 150.640 ;
        RECT 79.020 150.130 80.940 150.300 ;
        RECT 79.020 150.110 79.340 150.130 ;
        RECT 78.570 149.450 78.900 149.960 ;
        RECT 79.170 149.500 79.340 150.110 ;
        RECT 81.110 149.960 81.280 150.470 ;
        RECT 81.450 150.400 81.630 150.810 ;
        RECT 81.800 150.220 81.970 150.980 ;
        RECT 79.510 149.240 79.840 149.930 ;
        RECT 80.070 149.790 81.280 149.960 ;
        RECT 81.450 149.910 81.970 150.220 ;
        RECT 82.140 150.810 82.560 151.150 ;
        RECT 82.850 150.810 83.260 151.140 ;
        RECT 82.140 150.040 82.330 150.810 ;
        RECT 83.430 150.680 83.600 151.410 ;
        RECT 84.745 151.240 84.915 151.570 ;
        RECT 85.085 151.410 85.415 151.790 ;
        RECT 83.770 150.860 84.120 151.230 ;
        RECT 83.430 150.640 83.850 150.680 ;
        RECT 82.500 150.470 83.850 150.640 ;
        RECT 82.500 150.310 82.750 150.470 ;
        RECT 83.260 150.040 83.510 150.300 ;
        RECT 82.140 149.790 83.510 150.040 ;
        RECT 80.070 149.500 80.310 149.790 ;
        RECT 81.110 149.710 81.280 149.790 ;
        RECT 80.510 149.240 80.930 149.620 ;
        RECT 81.110 149.460 81.740 149.710 ;
        RECT 82.210 149.240 82.540 149.620 ;
        RECT 82.710 149.500 82.880 149.790 ;
        RECT 83.680 149.625 83.850 150.470 ;
        RECT 84.300 150.300 84.520 151.170 ;
        RECT 84.745 151.050 85.440 151.240 ;
        RECT 84.020 149.920 84.520 150.300 ;
        RECT 84.690 150.250 85.100 150.870 ;
        RECT 85.270 150.080 85.440 151.050 ;
        RECT 84.745 149.910 85.440 150.080 ;
        RECT 83.060 149.240 83.440 149.620 ;
        RECT 83.680 149.455 84.510 149.625 ;
        RECT 84.745 149.410 84.915 149.910 ;
        RECT 85.085 149.240 85.415 149.740 ;
        RECT 85.630 149.410 85.855 151.530 ;
        RECT 86.025 151.410 86.355 151.790 ;
        RECT 86.525 151.240 86.695 151.530 ;
        RECT 86.030 151.070 86.695 151.240 ;
        RECT 86.960 151.240 87.215 151.530 ;
        RECT 87.385 151.410 87.715 151.790 ;
        RECT 86.960 151.070 87.710 151.240 ;
        RECT 86.030 150.080 86.260 151.070 ;
        RECT 86.430 150.250 86.780 150.900 ;
        RECT 86.960 150.250 87.310 150.900 ;
        RECT 87.480 150.080 87.710 151.070 ;
        RECT 86.030 149.910 86.695 150.080 ;
        RECT 86.025 149.240 86.355 149.740 ;
        RECT 86.525 149.410 86.695 149.910 ;
        RECT 86.960 149.910 87.710 150.080 ;
        RECT 86.960 149.410 87.215 149.910 ;
        RECT 87.385 149.240 87.715 149.740 ;
        RECT 87.885 149.410 88.055 151.530 ;
        RECT 88.415 151.430 88.745 151.790 ;
        RECT 88.915 151.400 89.410 151.570 ;
        RECT 89.615 151.400 90.470 151.570 ;
        RECT 88.285 150.210 88.745 151.260 ;
        RECT 88.225 149.425 88.550 150.210 ;
        RECT 88.915 150.040 89.085 151.400 ;
        RECT 89.255 150.490 89.605 151.110 ;
        RECT 89.775 150.890 90.130 151.110 ;
        RECT 89.775 150.300 89.945 150.890 ;
        RECT 90.300 150.690 90.470 151.400 ;
        RECT 91.345 151.330 91.675 151.790 ;
        RECT 91.885 151.430 92.235 151.600 ;
        RECT 90.675 150.860 91.465 151.110 ;
        RECT 91.885 151.040 92.145 151.430 ;
        RECT 92.455 151.340 93.405 151.620 ;
        RECT 93.575 151.350 93.765 151.790 ;
        RECT 93.935 151.410 95.005 151.580 ;
        RECT 91.635 150.690 91.805 150.870 ;
        RECT 88.915 149.870 89.310 150.040 ;
        RECT 89.480 149.910 89.945 150.300 ;
        RECT 90.115 150.520 91.805 150.690 ;
        RECT 89.140 149.740 89.310 149.870 ;
        RECT 90.115 149.740 90.285 150.520 ;
        RECT 91.975 150.350 92.145 151.040 ;
        RECT 90.645 150.180 92.145 150.350 ;
        RECT 92.335 150.380 92.545 151.170 ;
        RECT 92.715 150.550 93.065 151.170 ;
        RECT 93.235 150.560 93.405 151.340 ;
        RECT 93.935 151.180 94.105 151.410 ;
        RECT 93.575 151.010 94.105 151.180 ;
        RECT 93.575 150.730 93.795 151.010 ;
        RECT 94.275 150.840 94.515 151.240 ;
        RECT 93.235 150.390 93.640 150.560 ;
        RECT 93.975 150.470 94.515 150.840 ;
        RECT 94.685 151.055 95.005 151.410 ;
        RECT 95.250 151.330 95.555 151.790 ;
        RECT 95.725 151.080 95.980 151.610 ;
        RECT 94.685 150.880 95.010 151.055 ;
        RECT 94.685 150.580 95.600 150.880 ;
        RECT 94.860 150.550 95.600 150.580 ;
        RECT 92.335 150.220 93.010 150.380 ;
        RECT 93.470 150.300 93.640 150.390 ;
        RECT 92.335 150.210 93.300 150.220 ;
        RECT 91.975 150.040 92.145 150.180 ;
        RECT 88.720 149.240 88.970 149.700 ;
        RECT 89.140 149.410 89.390 149.740 ;
        RECT 89.605 149.410 90.285 149.740 ;
        RECT 90.455 149.840 91.530 150.010 ;
        RECT 91.975 149.870 92.535 150.040 ;
        RECT 92.840 149.920 93.300 150.210 ;
        RECT 93.470 150.130 94.690 150.300 ;
        RECT 90.455 149.500 90.625 149.840 ;
        RECT 90.860 149.240 91.190 149.670 ;
        RECT 91.360 149.500 91.530 149.840 ;
        RECT 91.825 149.240 92.195 149.700 ;
        RECT 92.365 149.410 92.535 149.870 ;
        RECT 93.470 149.750 93.640 150.130 ;
        RECT 94.860 149.960 95.030 150.550 ;
        RECT 95.770 150.430 95.980 151.080 ;
        RECT 96.270 151.160 96.555 151.620 ;
        RECT 96.725 151.330 96.995 151.790 ;
        RECT 96.270 150.990 97.225 151.160 ;
        RECT 92.770 149.410 93.640 149.750 ;
        RECT 94.230 149.790 95.030 149.960 ;
        RECT 93.810 149.240 94.060 149.700 ;
        RECT 94.230 149.500 94.400 149.790 ;
        RECT 94.580 149.240 94.910 149.620 ;
        RECT 95.250 149.240 95.555 150.380 ;
        RECT 95.725 149.550 95.980 150.430 ;
        RECT 96.155 150.260 96.845 150.820 ;
        RECT 97.015 150.090 97.225 150.990 ;
        RECT 96.270 149.870 97.225 150.090 ;
        RECT 97.395 150.820 97.795 151.620 ;
        RECT 97.985 151.160 98.265 151.620 ;
        RECT 98.785 151.330 99.110 151.790 ;
        RECT 97.985 150.990 99.110 151.160 ;
        RECT 99.280 151.050 99.665 151.620 ;
        RECT 99.845 151.290 100.175 151.790 ;
        RECT 100.375 151.220 100.545 151.570 ;
        RECT 100.745 151.390 101.075 151.790 ;
        RECT 101.245 151.220 101.415 151.570 ;
        RECT 101.585 151.390 101.965 151.790 ;
        RECT 98.660 150.880 99.110 150.990 ;
        RECT 97.395 150.260 98.490 150.820 ;
        RECT 98.660 150.550 99.215 150.880 ;
        RECT 96.270 149.410 96.555 149.870 ;
        RECT 96.725 149.240 96.995 149.700 ;
        RECT 97.395 149.410 97.795 150.260 ;
        RECT 98.660 150.090 99.110 150.550 ;
        RECT 99.385 150.380 99.665 151.050 ;
        RECT 99.840 150.550 100.190 151.120 ;
        RECT 100.375 151.050 101.985 151.220 ;
        RECT 102.155 151.115 102.425 151.460 ;
        RECT 101.815 150.880 101.985 151.050 ;
        RECT 97.985 149.870 99.110 150.090 ;
        RECT 97.985 149.410 98.265 149.870 ;
        RECT 98.785 149.240 99.110 149.700 ;
        RECT 99.280 149.410 99.665 150.380 ;
        RECT 99.840 150.090 100.160 150.380 ;
        RECT 100.360 150.260 101.070 150.880 ;
        RECT 101.240 150.550 101.645 150.880 ;
        RECT 101.815 150.550 102.085 150.880 ;
        RECT 101.815 150.380 101.985 150.550 ;
        RECT 102.255 150.380 102.425 151.115 ;
        RECT 102.595 151.065 102.885 151.790 ;
        RECT 103.515 151.020 105.185 151.790 ;
        RECT 101.260 150.210 101.985 150.380 ;
        RECT 101.260 150.090 101.430 150.210 ;
        RECT 99.840 149.920 101.430 150.090 ;
        RECT 99.840 149.460 101.495 149.750 ;
        RECT 101.665 149.240 101.945 150.040 ;
        RECT 102.155 149.410 102.425 150.380 ;
        RECT 102.595 149.240 102.885 150.405 ;
        RECT 103.515 150.330 104.265 150.850 ;
        RECT 104.435 150.500 105.185 151.020 ;
        RECT 105.630 150.980 105.875 151.585 ;
        RECT 106.095 151.255 106.605 151.790 ;
        RECT 105.355 150.810 106.585 150.980 ;
        RECT 103.515 149.240 105.185 150.330 ;
        RECT 105.355 150.000 105.695 150.810 ;
        RECT 105.865 150.245 106.615 150.435 ;
        RECT 105.355 149.590 105.870 150.000 ;
        RECT 106.105 149.240 106.275 150.000 ;
        RECT 106.445 149.580 106.615 150.245 ;
        RECT 106.785 150.260 106.975 151.620 ;
        RECT 107.145 151.450 107.420 151.620 ;
        RECT 107.145 151.280 107.425 151.450 ;
        RECT 107.145 150.460 107.420 151.280 ;
        RECT 107.610 151.255 108.140 151.620 ;
        RECT 108.565 151.390 108.895 151.790 ;
        RECT 107.965 151.220 108.140 151.255 ;
        RECT 107.625 150.260 107.795 151.060 ;
        RECT 106.785 150.090 107.795 150.260 ;
        RECT 107.965 151.050 108.895 151.220 ;
        RECT 109.065 151.050 109.320 151.620 ;
        RECT 107.965 149.920 108.135 151.050 ;
        RECT 108.725 150.880 108.895 151.050 ;
        RECT 107.010 149.750 108.135 149.920 ;
        RECT 108.305 150.550 108.500 150.880 ;
        RECT 108.725 150.550 108.980 150.880 ;
        RECT 108.305 149.580 108.475 150.550 ;
        RECT 109.150 150.380 109.320 151.050 ;
        RECT 106.445 149.410 108.475 149.580 ;
        RECT 108.645 149.240 108.815 150.380 ;
        RECT 108.985 149.410 109.320 150.380 ;
        RECT 109.495 151.050 109.880 151.620 ;
        RECT 110.050 151.330 110.375 151.790 ;
        RECT 110.895 151.160 111.175 151.620 ;
        RECT 109.495 150.380 109.775 151.050 ;
        RECT 110.050 150.990 111.175 151.160 ;
        RECT 110.050 150.880 110.500 150.990 ;
        RECT 109.945 150.550 110.500 150.880 ;
        RECT 111.365 150.820 111.765 151.620 ;
        RECT 112.165 151.330 112.435 151.790 ;
        RECT 112.605 151.160 112.890 151.620 ;
        RECT 109.495 149.410 109.880 150.380 ;
        RECT 110.050 150.090 110.500 150.550 ;
        RECT 110.670 150.260 111.765 150.820 ;
        RECT 110.050 149.870 111.175 150.090 ;
        RECT 110.050 149.240 110.375 149.700 ;
        RECT 110.895 149.410 111.175 149.870 ;
        RECT 111.365 149.410 111.765 150.260 ;
        RECT 111.935 150.990 112.890 151.160 ;
        RECT 113.175 151.115 113.435 151.620 ;
        RECT 113.615 151.410 113.945 151.790 ;
        RECT 114.125 151.240 114.295 151.620 ;
        RECT 111.935 150.090 112.145 150.990 ;
        RECT 112.315 150.260 113.005 150.820 ;
        RECT 113.175 150.315 113.345 151.115 ;
        RECT 113.630 151.070 114.295 151.240 ;
        RECT 113.630 150.815 113.800 151.070 ;
        RECT 114.555 151.040 115.765 151.790 ;
        RECT 113.515 150.485 113.800 150.815 ;
        RECT 114.035 150.520 114.365 150.890 ;
        RECT 113.630 150.340 113.800 150.485 ;
        RECT 111.935 149.870 112.890 150.090 ;
        RECT 112.165 149.240 112.435 149.700 ;
        RECT 112.605 149.410 112.890 149.870 ;
        RECT 113.175 149.410 113.445 150.315 ;
        RECT 113.630 150.170 114.295 150.340 ;
        RECT 113.615 149.240 113.945 150.000 ;
        RECT 114.125 149.410 114.295 150.170 ;
        RECT 114.555 150.330 115.075 150.870 ;
        RECT 115.245 150.500 115.765 151.040 ;
        RECT 114.555 149.240 115.765 150.330 ;
        RECT 14.650 149.070 115.850 149.240 ;
        RECT 14.735 147.980 15.945 149.070 ;
        RECT 14.735 147.270 15.255 147.810 ;
        RECT 15.425 147.440 15.945 147.980 ;
        RECT 16.115 147.980 19.625 149.070 ;
        RECT 16.115 147.460 17.805 147.980 ;
        RECT 19.855 147.930 20.065 149.070 ;
        RECT 20.235 147.920 20.565 148.900 ;
        RECT 20.735 147.930 20.965 149.070 ;
        RECT 21.175 147.980 22.385 149.070 ;
        RECT 22.645 148.140 22.815 148.900 ;
        RECT 22.995 148.310 23.325 149.070 ;
        RECT 17.975 147.290 19.625 147.810 ;
        RECT 14.735 146.520 15.945 147.270 ;
        RECT 16.115 146.520 19.625 147.290 ;
        RECT 19.855 146.520 20.065 147.340 ;
        RECT 20.235 147.320 20.485 147.920 ;
        RECT 20.655 147.510 20.985 147.760 ;
        RECT 21.175 147.440 21.695 147.980 ;
        RECT 22.645 147.970 23.310 148.140 ;
        RECT 23.495 147.995 23.765 148.900 ;
        RECT 24.310 148.730 24.565 148.760 ;
        RECT 24.225 148.560 24.565 148.730 ;
        RECT 23.140 147.825 23.310 147.970 ;
        RECT 20.235 146.690 20.565 147.320 ;
        RECT 20.735 146.520 20.965 147.340 ;
        RECT 21.865 147.270 22.385 147.810 ;
        RECT 22.575 147.420 22.905 147.790 ;
        RECT 23.140 147.495 23.425 147.825 ;
        RECT 21.175 146.520 22.385 147.270 ;
        RECT 23.140 147.240 23.310 147.495 ;
        RECT 22.645 147.070 23.310 147.240 ;
        RECT 23.595 147.195 23.765 147.995 ;
        RECT 22.645 146.690 22.815 147.070 ;
        RECT 22.995 146.520 23.325 146.900 ;
        RECT 23.505 146.690 23.765 147.195 ;
        RECT 24.310 148.090 24.565 148.560 ;
        RECT 24.745 148.270 25.030 149.070 ;
        RECT 25.210 148.350 25.540 148.860 ;
        RECT 24.310 147.230 24.490 148.090 ;
        RECT 25.210 147.760 25.460 148.350 ;
        RECT 25.810 148.200 25.980 148.810 ;
        RECT 26.150 148.380 26.480 149.070 ;
        RECT 26.710 148.520 26.950 148.810 ;
        RECT 27.150 148.690 27.570 149.070 ;
        RECT 27.750 148.600 28.380 148.850 ;
        RECT 28.850 148.690 29.180 149.070 ;
        RECT 27.750 148.520 27.920 148.600 ;
        RECT 29.350 148.520 29.520 148.810 ;
        RECT 29.700 148.690 30.080 149.070 ;
        RECT 30.320 148.685 31.150 148.855 ;
        RECT 26.710 148.350 27.920 148.520 ;
        RECT 24.660 147.430 25.460 147.760 ;
        RECT 24.310 146.700 24.565 147.230 ;
        RECT 24.745 146.520 25.030 146.980 ;
        RECT 25.210 146.780 25.460 147.430 ;
        RECT 25.660 148.180 25.980 148.200 ;
        RECT 25.660 148.010 27.580 148.180 ;
        RECT 25.660 147.115 25.850 148.010 ;
        RECT 27.750 147.840 27.920 148.350 ;
        RECT 28.090 148.090 28.610 148.400 ;
        RECT 26.020 147.670 27.920 147.840 ;
        RECT 26.020 147.610 26.350 147.670 ;
        RECT 26.500 147.440 26.830 147.500 ;
        RECT 26.170 147.170 26.830 147.440 ;
        RECT 25.660 146.785 25.980 147.115 ;
        RECT 26.160 146.520 26.820 147.000 ;
        RECT 27.020 146.910 27.190 147.670 ;
        RECT 28.090 147.500 28.270 147.910 ;
        RECT 27.360 147.330 27.690 147.450 ;
        RECT 28.440 147.330 28.610 148.090 ;
        RECT 27.360 147.160 28.610 147.330 ;
        RECT 28.780 148.270 30.150 148.520 ;
        RECT 28.780 147.500 28.970 148.270 ;
        RECT 29.900 148.010 30.150 148.270 ;
        RECT 29.140 147.840 29.390 148.000 ;
        RECT 30.320 147.840 30.490 148.685 ;
        RECT 31.385 148.400 31.555 148.900 ;
        RECT 31.725 148.570 32.055 149.070 ;
        RECT 30.660 148.010 31.160 148.390 ;
        RECT 31.385 148.230 32.080 148.400 ;
        RECT 29.140 147.670 30.490 147.840 ;
        RECT 30.070 147.630 30.490 147.670 ;
        RECT 28.780 147.160 29.200 147.500 ;
        RECT 29.490 147.170 29.900 147.500 ;
        RECT 27.020 146.740 27.870 146.910 ;
        RECT 28.430 146.520 28.750 146.980 ;
        RECT 28.950 146.730 29.200 147.160 ;
        RECT 29.490 146.520 29.900 146.960 ;
        RECT 30.070 146.900 30.240 147.630 ;
        RECT 30.410 147.080 30.760 147.450 ;
        RECT 30.940 147.140 31.160 148.010 ;
        RECT 31.330 147.440 31.740 148.060 ;
        RECT 31.910 147.260 32.080 148.230 ;
        RECT 31.385 147.070 32.080 147.260 ;
        RECT 30.070 146.700 31.085 146.900 ;
        RECT 31.385 146.740 31.555 147.070 ;
        RECT 31.725 146.520 32.055 146.900 ;
        RECT 32.270 146.780 32.495 148.900 ;
        RECT 32.665 148.570 32.995 149.070 ;
        RECT 33.165 148.400 33.335 148.900 ;
        RECT 32.670 148.230 33.335 148.400 ;
        RECT 32.670 147.240 32.900 148.230 ;
        RECT 33.070 147.410 33.420 148.060 ;
        RECT 33.595 147.995 33.865 148.900 ;
        RECT 34.035 148.310 34.365 149.070 ;
        RECT 34.545 148.140 34.715 148.900 ;
        RECT 32.670 147.070 33.335 147.240 ;
        RECT 32.665 146.520 32.995 146.900 ;
        RECT 33.165 146.780 33.335 147.070 ;
        RECT 33.595 147.195 33.765 147.995 ;
        RECT 34.050 147.970 34.715 148.140 ;
        RECT 34.975 147.980 36.645 149.070 ;
        RECT 34.050 147.825 34.220 147.970 ;
        RECT 33.935 147.495 34.220 147.825 ;
        RECT 34.050 147.240 34.220 147.495 ;
        RECT 34.455 147.420 34.785 147.790 ;
        RECT 34.975 147.460 35.725 147.980 ;
        RECT 36.855 147.930 37.085 149.070 ;
        RECT 37.255 147.920 37.585 148.900 ;
        RECT 37.755 147.930 37.965 149.070 ;
        RECT 35.895 147.290 36.645 147.810 ;
        RECT 36.835 147.510 37.165 147.760 ;
        RECT 33.595 146.690 33.855 147.195 ;
        RECT 34.050 147.070 34.715 147.240 ;
        RECT 34.035 146.520 34.365 146.900 ;
        RECT 34.545 146.690 34.715 147.070 ;
        RECT 34.975 146.520 36.645 147.290 ;
        RECT 36.855 146.520 37.085 147.340 ;
        RECT 37.335 147.320 37.585 147.920 ;
        RECT 38.195 147.905 38.485 149.070 ;
        RECT 39.030 148.090 39.285 148.760 ;
        RECT 39.465 148.270 39.750 149.070 ;
        RECT 39.930 148.350 40.260 148.860 ;
        RECT 39.030 148.050 39.210 148.090 ;
        RECT 38.945 147.880 39.210 148.050 ;
        RECT 37.255 146.690 37.585 147.320 ;
        RECT 37.755 146.520 37.965 147.340 ;
        RECT 38.195 146.520 38.485 147.245 ;
        RECT 39.030 147.230 39.210 147.880 ;
        RECT 39.930 147.760 40.180 148.350 ;
        RECT 40.530 148.200 40.700 148.810 ;
        RECT 40.870 148.380 41.200 149.070 ;
        RECT 41.430 148.520 41.670 148.810 ;
        RECT 41.870 148.690 42.290 149.070 ;
        RECT 42.470 148.600 43.100 148.850 ;
        RECT 43.570 148.690 43.900 149.070 ;
        RECT 42.470 148.520 42.640 148.600 ;
        RECT 44.070 148.520 44.240 148.810 ;
        RECT 44.420 148.690 44.800 149.070 ;
        RECT 45.040 148.685 45.870 148.855 ;
        RECT 41.430 148.350 42.640 148.520 ;
        RECT 39.380 147.430 40.180 147.760 ;
        RECT 39.030 146.700 39.285 147.230 ;
        RECT 39.465 146.520 39.750 146.980 ;
        RECT 39.930 146.780 40.180 147.430 ;
        RECT 40.380 148.180 40.700 148.200 ;
        RECT 40.380 148.010 42.300 148.180 ;
        RECT 40.380 147.115 40.570 148.010 ;
        RECT 42.470 147.840 42.640 148.350 ;
        RECT 42.810 148.090 43.330 148.400 ;
        RECT 40.740 147.670 42.640 147.840 ;
        RECT 40.740 147.610 41.070 147.670 ;
        RECT 41.220 147.440 41.550 147.500 ;
        RECT 40.890 147.170 41.550 147.440 ;
        RECT 40.380 146.785 40.700 147.115 ;
        RECT 40.880 146.520 41.540 147.000 ;
        RECT 41.740 146.910 41.910 147.670 ;
        RECT 42.810 147.500 42.990 147.910 ;
        RECT 42.080 147.330 42.410 147.450 ;
        RECT 43.160 147.330 43.330 148.090 ;
        RECT 42.080 147.160 43.330 147.330 ;
        RECT 43.500 148.270 44.870 148.520 ;
        RECT 43.500 147.500 43.690 148.270 ;
        RECT 44.620 148.010 44.870 148.270 ;
        RECT 43.860 147.840 44.110 148.000 ;
        RECT 45.040 147.840 45.210 148.685 ;
        RECT 46.105 148.400 46.275 148.900 ;
        RECT 46.445 148.570 46.775 149.070 ;
        RECT 45.380 148.010 45.880 148.390 ;
        RECT 46.105 148.230 46.800 148.400 ;
        RECT 43.860 147.670 45.210 147.840 ;
        RECT 44.790 147.630 45.210 147.670 ;
        RECT 43.500 147.160 43.920 147.500 ;
        RECT 44.210 147.170 44.620 147.500 ;
        RECT 41.740 146.740 42.590 146.910 ;
        RECT 43.150 146.520 43.470 146.980 ;
        RECT 43.670 146.730 43.920 147.160 ;
        RECT 44.210 146.520 44.620 146.960 ;
        RECT 44.790 146.900 44.960 147.630 ;
        RECT 45.130 147.080 45.480 147.450 ;
        RECT 45.660 147.140 45.880 148.010 ;
        RECT 46.050 147.440 46.460 148.060 ;
        RECT 46.630 147.260 46.800 148.230 ;
        RECT 46.105 147.070 46.800 147.260 ;
        RECT 44.790 146.700 45.805 146.900 ;
        RECT 46.105 146.740 46.275 147.070 ;
        RECT 46.445 146.520 46.775 146.900 ;
        RECT 46.990 146.780 47.215 148.900 ;
        RECT 47.385 148.570 47.715 149.070 ;
        RECT 47.885 148.400 48.055 148.900 ;
        RECT 47.390 148.230 48.055 148.400 ;
        RECT 47.390 147.240 47.620 148.230 ;
        RECT 47.790 147.410 48.140 148.060 ;
        RECT 48.315 147.930 48.655 148.900 ;
        RECT 48.825 147.930 48.995 149.070 ;
        RECT 49.265 148.270 49.515 149.070 ;
        RECT 50.160 148.100 50.490 148.900 ;
        RECT 50.790 148.270 51.120 149.070 ;
        RECT 51.290 148.100 51.620 148.900 ;
        RECT 49.185 147.930 51.620 148.100 ;
        RECT 51.995 147.995 52.265 148.900 ;
        RECT 52.435 148.310 52.765 149.070 ;
        RECT 52.945 148.140 53.115 148.900 ;
        RECT 48.315 147.320 48.490 147.930 ;
        RECT 49.185 147.680 49.355 147.930 ;
        RECT 48.660 147.510 49.355 147.680 ;
        RECT 49.530 147.510 49.950 147.710 ;
        RECT 50.120 147.510 50.450 147.710 ;
        RECT 50.620 147.510 50.950 147.710 ;
        RECT 47.390 147.070 48.055 147.240 ;
        RECT 47.385 146.520 47.715 146.900 ;
        RECT 47.885 146.780 48.055 147.070 ;
        RECT 48.315 146.690 48.655 147.320 ;
        RECT 48.825 146.520 49.075 147.320 ;
        RECT 49.265 147.170 50.490 147.340 ;
        RECT 49.265 146.690 49.595 147.170 ;
        RECT 49.765 146.520 49.990 146.980 ;
        RECT 50.160 146.690 50.490 147.170 ;
        RECT 51.120 147.300 51.290 147.930 ;
        RECT 51.475 147.510 51.825 147.760 ;
        RECT 51.120 146.690 51.620 147.300 ;
        RECT 51.995 147.195 52.165 147.995 ;
        RECT 52.450 147.970 53.115 148.140 ;
        RECT 54.295 147.980 57.805 149.070 ;
        RECT 58.180 148.100 58.510 148.900 ;
        RECT 58.680 148.270 59.010 149.070 ;
        RECT 59.310 148.100 59.640 148.900 ;
        RECT 60.285 148.270 60.535 149.070 ;
        RECT 52.450 147.825 52.620 147.970 ;
        RECT 52.335 147.495 52.620 147.825 ;
        RECT 52.450 147.240 52.620 147.495 ;
        RECT 52.855 147.420 53.185 147.790 ;
        RECT 54.295 147.460 55.985 147.980 ;
        RECT 58.180 147.930 60.615 148.100 ;
        RECT 60.805 147.930 60.975 149.070 ;
        RECT 61.145 147.930 61.485 148.900 ;
        RECT 62.615 147.930 62.845 149.070 ;
        RECT 56.155 147.290 57.805 147.810 ;
        RECT 57.975 147.510 58.325 147.760 ;
        RECT 58.510 147.300 58.680 147.930 ;
        RECT 58.850 147.510 59.180 147.710 ;
        RECT 59.350 147.510 59.680 147.710 ;
        RECT 59.850 147.510 60.270 147.710 ;
        RECT 60.445 147.680 60.615 147.930 ;
        RECT 61.255 147.880 61.485 147.930 ;
        RECT 63.015 147.920 63.345 148.900 ;
        RECT 63.515 147.930 63.725 149.070 ;
        RECT 60.445 147.510 61.140 147.680 ;
        RECT 51.995 146.690 52.255 147.195 ;
        RECT 52.450 147.070 53.115 147.240 ;
        RECT 52.435 146.520 52.765 146.900 ;
        RECT 52.945 146.690 53.115 147.070 ;
        RECT 54.295 146.520 57.805 147.290 ;
        RECT 58.180 146.690 58.680 147.300 ;
        RECT 59.310 147.170 60.535 147.340 ;
        RECT 61.310 147.320 61.485 147.880 ;
        RECT 62.595 147.510 62.925 147.760 ;
        RECT 59.310 146.690 59.640 147.170 ;
        RECT 59.810 146.520 60.035 146.980 ;
        RECT 60.205 146.690 60.535 147.170 ;
        RECT 60.725 146.520 60.975 147.320 ;
        RECT 61.145 146.690 61.485 147.320 ;
        RECT 62.615 146.520 62.845 147.340 ;
        RECT 63.095 147.320 63.345 147.920 ;
        RECT 63.955 147.905 64.245 149.070 ;
        RECT 64.505 148.140 64.675 148.900 ;
        RECT 64.855 148.310 65.185 149.070 ;
        RECT 64.505 147.970 65.170 148.140 ;
        RECT 65.355 147.995 65.625 148.900 ;
        RECT 65.000 147.825 65.170 147.970 ;
        RECT 64.435 147.420 64.765 147.790 ;
        RECT 65.000 147.495 65.285 147.825 ;
        RECT 63.015 146.690 63.345 147.320 ;
        RECT 63.515 146.520 63.725 147.340 ;
        RECT 63.955 146.520 64.245 147.245 ;
        RECT 65.000 147.240 65.170 147.495 ;
        RECT 64.505 147.070 65.170 147.240 ;
        RECT 65.455 147.195 65.625 147.995 ;
        RECT 65.885 148.140 66.055 148.900 ;
        RECT 66.270 148.310 66.600 149.070 ;
        RECT 65.885 147.970 66.600 148.140 ;
        RECT 66.770 147.995 67.025 148.900 ;
        RECT 65.795 147.420 66.150 147.790 ;
        RECT 66.430 147.760 66.600 147.970 ;
        RECT 66.430 147.430 66.685 147.760 ;
        RECT 66.430 147.240 66.600 147.430 ;
        RECT 66.855 147.265 67.025 147.995 ;
        RECT 67.200 147.920 67.460 149.070 ;
        RECT 67.725 148.140 67.895 148.900 ;
        RECT 68.110 148.310 68.440 149.070 ;
        RECT 67.725 147.970 68.440 148.140 ;
        RECT 68.610 147.995 68.865 148.900 ;
        RECT 67.635 147.420 67.990 147.790 ;
        RECT 68.270 147.760 68.440 147.970 ;
        RECT 68.270 147.430 68.525 147.760 ;
        RECT 64.505 146.690 64.675 147.070 ;
        RECT 64.855 146.520 65.185 146.900 ;
        RECT 65.365 146.690 65.625 147.195 ;
        RECT 65.885 147.070 66.600 147.240 ;
        RECT 65.885 146.690 66.055 147.070 ;
        RECT 66.270 146.520 66.600 146.900 ;
        RECT 66.770 146.690 67.025 147.265 ;
        RECT 67.200 146.520 67.460 147.360 ;
        RECT 68.270 147.240 68.440 147.430 ;
        RECT 68.695 147.265 68.865 147.995 ;
        RECT 69.040 147.920 69.300 149.070 ;
        RECT 69.935 147.930 70.205 148.900 ;
        RECT 70.415 148.270 70.695 149.070 ;
        RECT 70.865 148.560 72.520 148.850 ;
        RECT 70.930 148.220 72.520 148.390 ;
        RECT 70.930 148.100 71.100 148.220 ;
        RECT 70.375 147.930 71.100 148.100 ;
        RECT 67.725 147.070 68.440 147.240 ;
        RECT 67.725 146.690 67.895 147.070 ;
        RECT 68.110 146.520 68.440 146.900 ;
        RECT 68.610 146.690 68.865 147.265 ;
        RECT 69.040 146.520 69.300 147.360 ;
        RECT 69.935 147.195 70.105 147.930 ;
        RECT 70.375 147.760 70.545 147.930 ;
        RECT 71.290 147.880 72.005 148.050 ;
        RECT 72.200 147.930 72.520 148.220 ;
        RECT 72.695 147.930 73.035 148.900 ;
        RECT 73.205 147.930 73.375 149.070 ;
        RECT 73.645 148.270 73.895 149.070 ;
        RECT 74.540 148.100 74.870 148.900 ;
        RECT 75.170 148.270 75.500 149.070 ;
        RECT 75.670 148.100 76.000 148.900 ;
        RECT 73.565 147.930 76.000 148.100 ;
        RECT 76.835 147.980 79.425 149.070 ;
        RECT 70.275 147.430 70.545 147.760 ;
        RECT 70.715 147.430 71.120 147.760 ;
        RECT 71.290 147.430 72.000 147.880 ;
        RECT 70.375 147.260 70.545 147.430 ;
        RECT 69.935 146.850 70.205 147.195 ;
        RECT 70.375 147.090 71.985 147.260 ;
        RECT 72.170 147.190 72.520 147.760 ;
        RECT 72.695 147.370 72.870 147.930 ;
        RECT 73.565 147.680 73.735 147.930 ;
        RECT 73.040 147.510 73.735 147.680 ;
        RECT 73.910 147.510 74.330 147.710 ;
        RECT 74.500 147.510 74.830 147.710 ;
        RECT 75.000 147.510 75.330 147.710 ;
        RECT 72.695 147.320 72.925 147.370 ;
        RECT 70.395 146.520 70.775 146.920 ;
        RECT 70.945 146.740 71.115 147.090 ;
        RECT 71.285 146.520 71.615 146.920 ;
        RECT 71.815 146.740 71.985 147.090 ;
        RECT 72.185 146.520 72.515 147.020 ;
        RECT 72.695 146.690 73.035 147.320 ;
        RECT 73.205 146.520 73.455 147.320 ;
        RECT 73.645 147.170 74.870 147.340 ;
        RECT 73.645 146.690 73.975 147.170 ;
        RECT 74.145 146.520 74.370 146.980 ;
        RECT 74.540 146.690 74.870 147.170 ;
        RECT 75.500 147.300 75.670 147.930 ;
        RECT 75.855 147.510 76.205 147.760 ;
        RECT 76.835 147.460 78.045 147.980 ;
        RECT 79.635 147.930 79.865 149.070 ;
        RECT 80.035 147.920 80.365 148.900 ;
        RECT 80.535 147.930 80.745 149.070 ;
        RECT 81.065 148.140 81.235 148.900 ;
        RECT 81.415 148.310 81.745 149.070 ;
        RECT 81.065 147.970 81.730 148.140 ;
        RECT 81.915 147.995 82.185 148.900 ;
        RECT 75.500 146.690 76.000 147.300 ;
        RECT 78.215 147.290 79.425 147.810 ;
        RECT 79.615 147.510 79.945 147.760 ;
        RECT 76.835 146.520 79.425 147.290 ;
        RECT 79.635 146.520 79.865 147.340 ;
        RECT 80.115 147.320 80.365 147.920 ;
        RECT 81.560 147.825 81.730 147.970 ;
        RECT 80.995 147.420 81.325 147.790 ;
        RECT 81.560 147.495 81.845 147.825 ;
        RECT 80.035 146.690 80.365 147.320 ;
        RECT 80.535 146.520 80.745 147.340 ;
        RECT 81.560 147.240 81.730 147.495 ;
        RECT 81.065 147.070 81.730 147.240 ;
        RECT 82.015 147.195 82.185 147.995 ;
        RECT 83.275 147.980 86.785 149.070 ;
        RECT 83.275 147.460 84.965 147.980 ;
        RECT 86.995 147.930 87.225 149.070 ;
        RECT 87.395 147.920 87.725 148.900 ;
        RECT 87.895 147.930 88.105 149.070 ;
        RECT 88.335 147.995 88.605 148.900 ;
        RECT 88.775 148.310 89.105 149.070 ;
        RECT 89.285 148.140 89.455 148.900 ;
        RECT 85.135 147.290 86.785 147.810 ;
        RECT 86.975 147.510 87.305 147.760 ;
        RECT 81.065 146.690 81.235 147.070 ;
        RECT 81.415 146.520 81.745 146.900 ;
        RECT 81.925 146.690 82.185 147.195 ;
        RECT 83.275 146.520 86.785 147.290 ;
        RECT 86.995 146.520 87.225 147.340 ;
        RECT 87.475 147.320 87.725 147.920 ;
        RECT 87.395 146.690 87.725 147.320 ;
        RECT 87.895 146.520 88.105 147.340 ;
        RECT 88.335 147.195 88.505 147.995 ;
        RECT 88.790 147.970 89.455 148.140 ;
        RECT 88.790 147.825 88.960 147.970 ;
        RECT 89.715 147.905 90.005 149.070 ;
        RECT 90.175 147.980 92.765 149.070 ;
        RECT 88.675 147.495 88.960 147.825 ;
        RECT 88.790 147.240 88.960 147.495 ;
        RECT 89.195 147.420 89.525 147.790 ;
        RECT 90.175 147.460 91.385 147.980 ;
        RECT 92.935 147.930 93.205 148.900 ;
        RECT 93.415 148.270 93.695 149.070 ;
        RECT 93.865 148.560 95.520 148.850 ;
        RECT 93.930 148.220 95.520 148.390 ;
        RECT 93.930 148.100 94.100 148.220 ;
        RECT 93.375 147.930 94.100 148.100 ;
        RECT 91.555 147.290 92.765 147.810 ;
        RECT 88.335 146.690 88.595 147.195 ;
        RECT 88.790 147.070 89.455 147.240 ;
        RECT 88.775 146.520 89.105 146.900 ;
        RECT 89.285 146.690 89.455 147.070 ;
        RECT 89.715 146.520 90.005 147.245 ;
        RECT 90.175 146.520 92.765 147.290 ;
        RECT 92.935 147.195 93.105 147.930 ;
        RECT 93.375 147.760 93.545 147.930 ;
        RECT 94.290 147.880 95.005 148.050 ;
        RECT 95.200 147.930 95.520 148.220 ;
        RECT 95.695 147.930 96.035 148.900 ;
        RECT 96.205 147.930 96.375 149.070 ;
        RECT 96.645 148.270 96.895 149.070 ;
        RECT 97.540 148.100 97.870 148.900 ;
        RECT 98.170 148.270 98.500 149.070 ;
        RECT 98.670 148.100 99.000 148.900 ;
        RECT 96.565 147.930 99.000 148.100 ;
        RECT 99.580 148.100 99.910 148.900 ;
        RECT 100.080 148.270 100.410 149.070 ;
        RECT 100.710 148.100 101.040 148.900 ;
        RECT 101.685 148.270 101.935 149.070 ;
        RECT 99.580 147.930 102.015 148.100 ;
        RECT 102.205 147.930 102.375 149.070 ;
        RECT 102.545 147.930 102.885 148.900 ;
        RECT 93.275 147.430 93.545 147.760 ;
        RECT 93.715 147.430 94.120 147.760 ;
        RECT 94.290 147.430 95.000 147.880 ;
        RECT 93.375 147.260 93.545 147.430 ;
        RECT 92.935 146.850 93.205 147.195 ;
        RECT 93.375 147.090 94.985 147.260 ;
        RECT 95.170 147.190 95.520 147.760 ;
        RECT 95.695 147.370 95.870 147.930 ;
        RECT 96.565 147.680 96.735 147.930 ;
        RECT 96.040 147.510 96.735 147.680 ;
        RECT 96.910 147.510 97.330 147.710 ;
        RECT 97.500 147.510 97.830 147.710 ;
        RECT 98.000 147.510 98.330 147.710 ;
        RECT 95.695 147.320 95.925 147.370 ;
        RECT 93.395 146.520 93.775 146.920 ;
        RECT 93.945 146.740 94.115 147.090 ;
        RECT 94.285 146.520 94.615 146.920 ;
        RECT 94.815 146.740 94.985 147.090 ;
        RECT 95.185 146.520 95.515 147.020 ;
        RECT 95.695 146.690 96.035 147.320 ;
        RECT 96.205 146.520 96.455 147.320 ;
        RECT 96.645 147.170 97.870 147.340 ;
        RECT 96.645 146.690 96.975 147.170 ;
        RECT 97.145 146.520 97.370 146.980 ;
        RECT 97.540 146.690 97.870 147.170 ;
        RECT 98.500 147.300 98.670 147.930 ;
        RECT 98.855 147.510 99.205 147.760 ;
        RECT 99.375 147.510 99.725 147.760 ;
        RECT 99.910 147.300 100.080 147.930 ;
        RECT 100.250 147.510 100.580 147.710 ;
        RECT 100.750 147.510 101.080 147.710 ;
        RECT 101.250 147.510 101.670 147.710 ;
        RECT 101.845 147.680 102.015 147.930 ;
        RECT 101.845 147.510 102.540 147.680 ;
        RECT 98.500 146.690 99.000 147.300 ;
        RECT 99.580 146.690 100.080 147.300 ;
        RECT 100.710 147.170 101.935 147.340 ;
        RECT 102.710 147.320 102.885 147.930 ;
        RECT 103.055 147.980 104.725 149.070 ;
        RECT 105.270 148.730 105.525 148.760 ;
        RECT 105.185 148.560 105.525 148.730 ;
        RECT 105.270 148.090 105.525 148.560 ;
        RECT 105.705 148.270 105.990 149.070 ;
        RECT 106.170 148.350 106.500 148.860 ;
        RECT 103.055 147.460 103.805 147.980 ;
        RECT 100.710 146.690 101.040 147.170 ;
        RECT 101.210 146.520 101.435 146.980 ;
        RECT 101.605 146.690 101.935 147.170 ;
        RECT 102.125 146.520 102.375 147.320 ;
        RECT 102.545 146.690 102.885 147.320 ;
        RECT 103.975 147.290 104.725 147.810 ;
        RECT 103.055 146.520 104.725 147.290 ;
        RECT 105.270 147.230 105.450 148.090 ;
        RECT 106.170 147.760 106.420 148.350 ;
        RECT 106.770 148.200 106.940 148.810 ;
        RECT 107.110 148.380 107.440 149.070 ;
        RECT 107.670 148.520 107.910 148.810 ;
        RECT 108.110 148.690 108.530 149.070 ;
        RECT 108.710 148.600 109.340 148.850 ;
        RECT 109.810 148.690 110.140 149.070 ;
        RECT 108.710 148.520 108.880 148.600 ;
        RECT 110.310 148.520 110.480 148.810 ;
        RECT 110.660 148.690 111.040 149.070 ;
        RECT 111.280 148.685 112.110 148.855 ;
        RECT 107.670 148.350 108.880 148.520 ;
        RECT 105.620 147.430 106.420 147.760 ;
        RECT 105.270 146.700 105.525 147.230 ;
        RECT 105.705 146.520 105.990 146.980 ;
        RECT 106.170 146.780 106.420 147.430 ;
        RECT 106.620 148.180 106.940 148.200 ;
        RECT 106.620 148.010 108.540 148.180 ;
        RECT 106.620 147.115 106.810 148.010 ;
        RECT 108.710 147.840 108.880 148.350 ;
        RECT 109.050 148.090 109.570 148.400 ;
        RECT 106.980 147.670 108.880 147.840 ;
        RECT 106.980 147.610 107.310 147.670 ;
        RECT 107.460 147.440 107.790 147.500 ;
        RECT 107.130 147.170 107.790 147.440 ;
        RECT 106.620 146.785 106.940 147.115 ;
        RECT 107.120 146.520 107.780 147.000 ;
        RECT 107.980 146.910 108.150 147.670 ;
        RECT 109.050 147.500 109.230 147.910 ;
        RECT 108.320 147.330 108.650 147.450 ;
        RECT 109.400 147.330 109.570 148.090 ;
        RECT 108.320 147.160 109.570 147.330 ;
        RECT 109.740 148.270 111.110 148.520 ;
        RECT 109.740 147.500 109.930 148.270 ;
        RECT 110.860 148.010 111.110 148.270 ;
        RECT 110.100 147.840 110.350 148.000 ;
        RECT 111.280 147.840 111.450 148.685 ;
        RECT 112.345 148.400 112.515 148.900 ;
        RECT 112.685 148.570 113.015 149.070 ;
        RECT 111.620 148.010 112.120 148.390 ;
        RECT 112.345 148.230 113.040 148.400 ;
        RECT 110.100 147.670 111.450 147.840 ;
        RECT 111.030 147.630 111.450 147.670 ;
        RECT 109.740 147.160 110.160 147.500 ;
        RECT 110.450 147.170 110.860 147.500 ;
        RECT 107.980 146.740 108.830 146.910 ;
        RECT 109.390 146.520 109.710 146.980 ;
        RECT 109.910 146.730 110.160 147.160 ;
        RECT 110.450 146.520 110.860 146.960 ;
        RECT 111.030 146.900 111.200 147.630 ;
        RECT 111.370 147.080 111.720 147.450 ;
        RECT 111.900 147.140 112.120 148.010 ;
        RECT 112.290 147.440 112.700 148.060 ;
        RECT 112.870 147.260 113.040 148.230 ;
        RECT 112.345 147.070 113.040 147.260 ;
        RECT 111.030 146.700 112.045 146.900 ;
        RECT 112.345 146.740 112.515 147.070 ;
        RECT 112.685 146.520 113.015 146.900 ;
        RECT 113.230 146.780 113.455 148.900 ;
        RECT 113.625 148.570 113.955 149.070 ;
        RECT 114.125 148.400 114.295 148.900 ;
        RECT 113.630 148.230 114.295 148.400 ;
        RECT 113.630 147.240 113.860 148.230 ;
        RECT 114.030 147.410 114.380 148.060 ;
        RECT 114.555 147.980 115.765 149.070 ;
        RECT 114.555 147.440 115.075 147.980 ;
        RECT 115.245 147.270 115.765 147.810 ;
        RECT 113.630 147.070 114.295 147.240 ;
        RECT 113.625 146.520 113.955 146.900 ;
        RECT 114.125 146.780 114.295 147.070 ;
        RECT 114.555 146.520 115.765 147.270 ;
        RECT 14.650 146.350 115.850 146.520 ;
        RECT 14.735 145.600 15.945 146.350 ;
        RECT 14.735 145.060 15.255 145.600 ;
        RECT 16.115 145.580 19.625 146.350 ;
        RECT 19.800 145.805 25.145 146.350 ;
        RECT 15.425 144.890 15.945 145.430 ;
        RECT 14.735 143.800 15.945 144.890 ;
        RECT 16.115 144.890 17.805 145.410 ;
        RECT 17.975 145.060 19.625 145.580 ;
        RECT 16.115 143.800 19.625 144.890 ;
        RECT 21.390 144.235 21.740 145.485 ;
        RECT 23.220 144.975 23.560 145.805 ;
        RECT 25.315 145.625 25.605 146.350 ;
        RECT 25.775 145.580 29.285 146.350 ;
        RECT 29.460 145.805 34.805 146.350 ;
        RECT 19.800 143.800 25.145 144.235 ;
        RECT 25.315 143.800 25.605 144.965 ;
        RECT 25.775 144.890 27.465 145.410 ;
        RECT 27.635 145.060 29.285 145.580 ;
        RECT 25.775 143.800 29.285 144.890 ;
        RECT 31.050 144.235 31.400 145.485 ;
        RECT 32.880 144.975 33.220 145.805 ;
        RECT 35.065 145.800 35.235 146.090 ;
        RECT 35.405 145.970 35.735 146.350 ;
        RECT 35.065 145.630 35.730 145.800 ;
        RECT 34.980 144.810 35.330 145.460 ;
        RECT 35.500 144.640 35.730 145.630 ;
        RECT 35.065 144.470 35.730 144.640 ;
        RECT 29.460 143.800 34.805 144.235 ;
        RECT 35.065 143.970 35.235 144.470 ;
        RECT 35.405 143.800 35.735 144.300 ;
        RECT 35.905 143.970 36.130 146.090 ;
        RECT 36.345 145.970 36.675 146.350 ;
        RECT 36.845 145.800 37.015 146.130 ;
        RECT 37.315 145.970 38.330 146.170 ;
        RECT 36.320 145.610 37.015 145.800 ;
        RECT 36.320 144.640 36.490 145.610 ;
        RECT 36.660 144.810 37.070 145.430 ;
        RECT 37.240 144.860 37.460 145.730 ;
        RECT 37.640 145.420 37.990 145.790 ;
        RECT 38.160 145.240 38.330 145.970 ;
        RECT 38.500 145.910 38.910 146.350 ;
        RECT 39.200 145.710 39.450 146.140 ;
        RECT 39.650 145.890 39.970 146.350 ;
        RECT 40.530 145.960 41.380 146.130 ;
        RECT 38.500 145.370 38.910 145.700 ;
        RECT 39.200 145.370 39.620 145.710 ;
        RECT 37.910 145.200 38.330 145.240 ;
        RECT 37.910 145.030 39.260 145.200 ;
        RECT 36.320 144.470 37.015 144.640 ;
        RECT 37.240 144.480 37.740 144.860 ;
        RECT 36.345 143.800 36.675 144.300 ;
        RECT 36.845 143.970 37.015 144.470 ;
        RECT 37.910 144.185 38.080 145.030 ;
        RECT 39.010 144.870 39.260 145.030 ;
        RECT 38.250 144.600 38.500 144.860 ;
        RECT 39.430 144.600 39.620 145.370 ;
        RECT 38.250 144.350 39.620 144.600 ;
        RECT 39.790 145.540 41.040 145.710 ;
        RECT 39.790 144.780 39.960 145.540 ;
        RECT 40.710 145.420 41.040 145.540 ;
        RECT 40.130 144.960 40.310 145.370 ;
        RECT 41.210 145.200 41.380 145.960 ;
        RECT 41.580 145.870 42.240 146.350 ;
        RECT 42.420 145.755 42.740 146.085 ;
        RECT 41.570 145.430 42.230 145.700 ;
        RECT 41.570 145.370 41.900 145.430 ;
        RECT 42.050 145.200 42.380 145.260 ;
        RECT 40.480 145.030 42.380 145.200 ;
        RECT 39.790 144.470 40.310 144.780 ;
        RECT 40.480 144.520 40.650 145.030 ;
        RECT 42.550 144.860 42.740 145.755 ;
        RECT 40.820 144.690 42.740 144.860 ;
        RECT 42.420 144.670 42.740 144.690 ;
        RECT 42.940 145.440 43.190 146.090 ;
        RECT 43.370 145.890 43.655 146.350 ;
        RECT 43.835 145.640 44.090 146.170 ;
        RECT 42.940 145.110 43.740 145.440 ;
        RECT 40.480 144.350 41.690 144.520 ;
        RECT 37.250 144.015 38.080 144.185 ;
        RECT 38.320 143.800 38.700 144.180 ;
        RECT 38.880 144.060 39.050 144.350 ;
        RECT 40.480 144.270 40.650 144.350 ;
        RECT 39.220 143.800 39.550 144.180 ;
        RECT 40.020 144.020 40.650 144.270 ;
        RECT 40.830 143.800 41.250 144.180 ;
        RECT 41.450 144.060 41.690 144.350 ;
        RECT 41.920 143.800 42.250 144.490 ;
        RECT 42.420 144.060 42.590 144.670 ;
        RECT 42.940 144.520 43.190 145.110 ;
        RECT 43.910 144.780 44.090 145.640 ;
        RECT 42.860 144.010 43.190 144.520 ;
        RECT 43.370 143.800 43.655 144.600 ;
        RECT 43.835 144.310 44.090 144.780 ;
        RECT 44.635 145.675 44.905 146.020 ;
        RECT 45.095 145.950 45.475 146.350 ;
        RECT 45.645 145.780 45.815 146.130 ;
        RECT 45.985 145.950 46.315 146.350 ;
        RECT 46.515 145.780 46.685 146.130 ;
        RECT 46.885 145.850 47.215 146.350 ;
        RECT 44.635 144.940 44.805 145.675 ;
        RECT 45.075 145.610 46.685 145.780 ;
        RECT 45.075 145.440 45.245 145.610 ;
        RECT 44.975 145.110 45.245 145.440 ;
        RECT 45.415 145.110 45.820 145.440 ;
        RECT 45.075 144.940 45.245 145.110 ;
        RECT 45.990 144.990 46.700 145.440 ;
        RECT 46.870 145.110 47.220 145.680 ;
        RECT 47.395 145.550 47.735 146.180 ;
        RECT 47.905 145.550 48.155 146.350 ;
        RECT 48.345 145.700 48.675 146.180 ;
        RECT 48.845 145.890 49.070 146.350 ;
        RECT 49.240 145.700 49.570 146.180 ;
        RECT 47.395 145.500 47.625 145.550 ;
        RECT 48.345 145.530 49.570 145.700 ;
        RECT 50.200 145.570 50.700 146.180 ;
        RECT 51.075 145.625 51.365 146.350 ;
        RECT 51.535 145.600 52.745 146.350 ;
        RECT 43.835 144.140 44.175 144.310 ;
        RECT 43.835 144.110 44.090 144.140 ;
        RECT 44.635 143.970 44.905 144.940 ;
        RECT 45.075 144.770 45.800 144.940 ;
        RECT 45.990 144.820 46.705 144.990 ;
        RECT 47.395 144.940 47.570 145.500 ;
        RECT 47.740 145.190 48.435 145.360 ;
        RECT 48.265 144.940 48.435 145.190 ;
        RECT 48.610 145.160 49.030 145.360 ;
        RECT 49.200 145.160 49.530 145.360 ;
        RECT 49.700 145.160 50.030 145.360 ;
        RECT 50.200 144.940 50.370 145.570 ;
        RECT 50.555 145.110 50.905 145.360 ;
        RECT 45.630 144.650 45.800 144.770 ;
        RECT 46.900 144.650 47.220 144.940 ;
        RECT 45.115 143.800 45.395 144.600 ;
        RECT 45.630 144.480 47.220 144.650 ;
        RECT 45.565 144.020 47.220 144.310 ;
        RECT 47.395 143.970 47.735 144.940 ;
        RECT 47.905 143.800 48.075 144.940 ;
        RECT 48.265 144.770 50.700 144.940 ;
        RECT 48.345 143.800 48.595 144.600 ;
        RECT 49.240 143.970 49.570 144.770 ;
        RECT 49.870 143.800 50.200 144.600 ;
        RECT 50.370 143.970 50.700 144.770 ;
        RECT 51.075 143.800 51.365 144.965 ;
        RECT 51.535 144.890 52.055 145.430 ;
        RECT 52.225 145.060 52.745 145.600 ;
        RECT 52.915 145.580 56.425 146.350 ;
        RECT 52.915 144.890 54.605 145.410 ;
        RECT 54.775 145.060 56.425 145.580 ;
        RECT 56.870 145.540 57.115 146.145 ;
        RECT 57.335 145.815 57.845 146.350 ;
        RECT 56.595 145.370 57.825 145.540 ;
        RECT 51.535 143.800 52.745 144.890 ;
        RECT 52.915 143.800 56.425 144.890 ;
        RECT 56.595 144.560 56.935 145.370 ;
        RECT 57.105 144.805 57.855 144.995 ;
        RECT 56.595 144.150 57.110 144.560 ;
        RECT 57.345 143.800 57.515 144.560 ;
        RECT 57.685 144.140 57.855 144.805 ;
        RECT 58.025 144.820 58.215 146.180 ;
        RECT 58.385 145.330 58.660 146.180 ;
        RECT 58.850 145.815 59.380 146.180 ;
        RECT 59.805 145.950 60.135 146.350 ;
        RECT 59.205 145.780 59.380 145.815 ;
        RECT 58.385 145.160 58.665 145.330 ;
        RECT 58.385 145.020 58.660 145.160 ;
        RECT 58.865 144.820 59.035 145.620 ;
        RECT 58.025 144.650 59.035 144.820 ;
        RECT 59.205 145.610 60.135 145.780 ;
        RECT 60.305 145.610 60.560 146.180 ;
        RECT 59.205 144.480 59.375 145.610 ;
        RECT 59.965 145.440 60.135 145.610 ;
        RECT 58.250 144.310 59.375 144.480 ;
        RECT 59.545 145.110 59.740 145.440 ;
        RECT 59.965 145.110 60.220 145.440 ;
        RECT 59.545 144.140 59.715 145.110 ;
        RECT 60.390 144.940 60.560 145.610 ;
        RECT 61.110 145.640 61.365 146.170 ;
        RECT 61.545 145.890 61.830 146.350 ;
        RECT 61.110 145.330 61.290 145.640 ;
        RECT 62.010 145.440 62.260 146.090 ;
        RECT 61.025 145.160 61.290 145.330 ;
        RECT 57.685 143.970 59.715 144.140 ;
        RECT 59.885 143.800 60.055 144.940 ;
        RECT 60.225 143.970 60.560 144.940 ;
        RECT 61.110 144.780 61.290 145.160 ;
        RECT 61.460 145.110 62.260 145.440 ;
        RECT 61.110 144.110 61.365 144.780 ;
        RECT 61.545 143.800 61.830 144.600 ;
        RECT 62.010 144.520 62.260 145.110 ;
        RECT 62.460 145.755 62.780 146.085 ;
        RECT 62.960 145.870 63.620 146.350 ;
        RECT 63.820 145.960 64.670 146.130 ;
        RECT 62.460 144.860 62.650 145.755 ;
        RECT 62.970 145.430 63.630 145.700 ;
        RECT 63.300 145.370 63.630 145.430 ;
        RECT 62.820 145.200 63.150 145.260 ;
        RECT 63.820 145.200 63.990 145.960 ;
        RECT 65.230 145.890 65.550 146.350 ;
        RECT 65.750 145.710 66.000 146.140 ;
        RECT 66.290 145.910 66.700 146.350 ;
        RECT 66.870 145.970 67.885 146.170 ;
        RECT 64.160 145.540 65.410 145.710 ;
        RECT 64.160 145.420 64.490 145.540 ;
        RECT 62.820 145.030 64.720 145.200 ;
        RECT 62.460 144.690 64.380 144.860 ;
        RECT 62.460 144.670 62.780 144.690 ;
        RECT 62.010 144.010 62.340 144.520 ;
        RECT 62.610 144.060 62.780 144.670 ;
        RECT 64.550 144.520 64.720 145.030 ;
        RECT 64.890 144.960 65.070 145.370 ;
        RECT 65.240 144.780 65.410 145.540 ;
        RECT 62.950 143.800 63.280 144.490 ;
        RECT 63.510 144.350 64.720 144.520 ;
        RECT 64.890 144.470 65.410 144.780 ;
        RECT 65.580 145.370 66.000 145.710 ;
        RECT 66.290 145.370 66.700 145.700 ;
        RECT 65.580 144.600 65.770 145.370 ;
        RECT 66.870 145.240 67.040 145.970 ;
        RECT 68.185 145.800 68.355 146.130 ;
        RECT 68.525 145.970 68.855 146.350 ;
        RECT 67.210 145.420 67.560 145.790 ;
        RECT 66.870 145.200 67.290 145.240 ;
        RECT 65.940 145.030 67.290 145.200 ;
        RECT 65.940 144.870 66.190 145.030 ;
        RECT 66.700 144.600 66.950 144.860 ;
        RECT 65.580 144.350 66.950 144.600 ;
        RECT 63.510 144.060 63.750 144.350 ;
        RECT 64.550 144.270 64.720 144.350 ;
        RECT 63.950 143.800 64.370 144.180 ;
        RECT 64.550 144.020 65.180 144.270 ;
        RECT 65.650 143.800 65.980 144.180 ;
        RECT 66.150 144.060 66.320 144.350 ;
        RECT 67.120 144.185 67.290 145.030 ;
        RECT 67.740 144.860 67.960 145.730 ;
        RECT 68.185 145.610 68.880 145.800 ;
        RECT 67.460 144.480 67.960 144.860 ;
        RECT 68.130 144.810 68.540 145.430 ;
        RECT 68.710 144.640 68.880 145.610 ;
        RECT 68.185 144.470 68.880 144.640 ;
        RECT 66.500 143.800 66.880 144.180 ;
        RECT 67.120 144.015 67.950 144.185 ;
        RECT 68.185 143.970 68.355 144.470 ;
        RECT 68.525 143.800 68.855 144.300 ;
        RECT 69.070 143.970 69.295 146.090 ;
        RECT 69.465 145.970 69.795 146.350 ;
        RECT 69.965 145.800 70.135 146.090 ;
        RECT 71.320 145.805 76.665 146.350 ;
        RECT 69.470 145.630 70.135 145.800 ;
        RECT 69.470 144.640 69.700 145.630 ;
        RECT 69.870 144.810 70.220 145.460 ;
        RECT 69.470 144.470 70.135 144.640 ;
        RECT 69.465 143.800 69.795 144.300 ;
        RECT 69.965 143.970 70.135 144.470 ;
        RECT 72.910 144.235 73.260 145.485 ;
        RECT 74.740 144.975 75.080 145.805 ;
        RECT 76.835 145.625 77.125 146.350 ;
        RECT 77.670 146.010 77.925 146.170 ;
        RECT 77.585 145.840 77.925 146.010 ;
        RECT 78.105 145.890 78.390 146.350 ;
        RECT 77.670 145.640 77.925 145.840 ;
        RECT 71.320 143.800 76.665 144.235 ;
        RECT 76.835 143.800 77.125 144.965 ;
        RECT 77.670 144.780 77.850 145.640 ;
        RECT 78.570 145.440 78.820 146.090 ;
        RECT 78.020 145.110 78.820 145.440 ;
        RECT 77.670 144.110 77.925 144.780 ;
        RECT 78.105 143.800 78.390 144.600 ;
        RECT 78.570 144.520 78.820 145.110 ;
        RECT 79.020 145.755 79.340 146.085 ;
        RECT 79.520 145.870 80.180 146.350 ;
        RECT 80.380 145.960 81.230 146.130 ;
        RECT 79.020 144.860 79.210 145.755 ;
        RECT 79.530 145.430 80.190 145.700 ;
        RECT 79.860 145.370 80.190 145.430 ;
        RECT 79.380 145.200 79.710 145.260 ;
        RECT 80.380 145.200 80.550 145.960 ;
        RECT 81.790 145.890 82.110 146.350 ;
        RECT 82.310 145.710 82.560 146.140 ;
        RECT 82.850 145.910 83.260 146.350 ;
        RECT 83.430 145.970 84.445 146.170 ;
        RECT 80.720 145.540 81.970 145.710 ;
        RECT 80.720 145.420 81.050 145.540 ;
        RECT 79.380 145.030 81.280 145.200 ;
        RECT 79.020 144.690 80.940 144.860 ;
        RECT 79.020 144.670 79.340 144.690 ;
        RECT 78.570 144.010 78.900 144.520 ;
        RECT 79.170 144.060 79.340 144.670 ;
        RECT 81.110 144.520 81.280 145.030 ;
        RECT 81.450 144.960 81.630 145.370 ;
        RECT 81.800 144.780 81.970 145.540 ;
        RECT 79.510 143.800 79.840 144.490 ;
        RECT 80.070 144.350 81.280 144.520 ;
        RECT 81.450 144.470 81.970 144.780 ;
        RECT 82.140 145.370 82.560 145.710 ;
        RECT 82.850 145.370 83.260 145.700 ;
        RECT 82.140 144.600 82.330 145.370 ;
        RECT 83.430 145.240 83.600 145.970 ;
        RECT 84.745 145.800 84.915 146.130 ;
        RECT 85.085 145.970 85.415 146.350 ;
        RECT 83.770 145.420 84.120 145.790 ;
        RECT 83.430 145.200 83.850 145.240 ;
        RECT 82.500 145.030 83.850 145.200 ;
        RECT 82.500 144.870 82.750 145.030 ;
        RECT 83.260 144.600 83.510 144.860 ;
        RECT 82.140 144.350 83.510 144.600 ;
        RECT 80.070 144.060 80.310 144.350 ;
        RECT 81.110 144.270 81.280 144.350 ;
        RECT 80.510 143.800 80.930 144.180 ;
        RECT 81.110 144.020 81.740 144.270 ;
        RECT 82.210 143.800 82.540 144.180 ;
        RECT 82.710 144.060 82.880 144.350 ;
        RECT 83.680 144.185 83.850 145.030 ;
        RECT 84.300 144.860 84.520 145.730 ;
        RECT 84.745 145.610 85.440 145.800 ;
        RECT 84.020 144.480 84.520 144.860 ;
        RECT 84.690 144.810 85.100 145.430 ;
        RECT 85.270 144.640 85.440 145.610 ;
        RECT 84.745 144.470 85.440 144.640 ;
        RECT 83.060 143.800 83.440 144.180 ;
        RECT 83.680 144.015 84.510 144.185 ;
        RECT 84.745 143.970 84.915 144.470 ;
        RECT 85.085 143.800 85.415 144.300 ;
        RECT 85.630 143.970 85.855 146.090 ;
        RECT 86.025 145.970 86.355 146.350 ;
        RECT 86.525 145.800 86.695 146.090 ;
        RECT 87.880 145.805 93.225 146.350 ;
        RECT 86.030 145.630 86.695 145.800 ;
        RECT 86.030 144.640 86.260 145.630 ;
        RECT 86.430 144.810 86.780 145.460 ;
        RECT 86.030 144.470 86.695 144.640 ;
        RECT 86.025 143.800 86.355 144.300 ;
        RECT 86.525 143.970 86.695 144.470 ;
        RECT 89.470 144.235 89.820 145.485 ;
        RECT 91.300 144.975 91.640 145.805 ;
        RECT 93.395 145.675 93.665 146.020 ;
        RECT 93.855 145.950 94.235 146.350 ;
        RECT 94.405 145.780 94.575 146.130 ;
        RECT 94.745 145.950 95.075 146.350 ;
        RECT 95.275 145.780 95.445 146.130 ;
        RECT 95.645 145.850 95.975 146.350 ;
        RECT 93.395 144.940 93.565 145.675 ;
        RECT 93.835 145.610 95.445 145.780 ;
        RECT 93.835 145.440 94.005 145.610 ;
        RECT 93.735 145.110 94.005 145.440 ;
        RECT 94.175 145.110 94.580 145.440 ;
        RECT 93.835 144.940 94.005 145.110 ;
        RECT 94.750 144.990 95.460 145.440 ;
        RECT 95.630 145.110 95.980 145.680 ;
        RECT 96.155 145.550 96.495 146.180 ;
        RECT 96.665 145.550 96.915 146.350 ;
        RECT 97.105 145.700 97.435 146.180 ;
        RECT 97.605 145.890 97.830 146.350 ;
        RECT 98.000 145.700 98.330 146.180 ;
        RECT 96.155 145.500 96.385 145.550 ;
        RECT 97.105 145.530 98.330 145.700 ;
        RECT 98.960 145.570 99.460 146.180 ;
        RECT 99.835 145.580 102.425 146.350 ;
        RECT 102.595 145.625 102.885 146.350 ;
        RECT 103.055 145.580 105.645 146.350 ;
        RECT 87.880 143.800 93.225 144.235 ;
        RECT 93.395 143.970 93.665 144.940 ;
        RECT 93.835 144.770 94.560 144.940 ;
        RECT 94.750 144.820 95.465 144.990 ;
        RECT 96.155 144.940 96.330 145.500 ;
        RECT 96.500 145.190 97.195 145.360 ;
        RECT 97.025 144.940 97.195 145.190 ;
        RECT 97.370 145.160 97.790 145.360 ;
        RECT 97.960 145.160 98.290 145.360 ;
        RECT 98.460 145.160 98.790 145.360 ;
        RECT 98.960 144.940 99.130 145.570 ;
        RECT 99.315 145.110 99.665 145.360 ;
        RECT 94.390 144.650 94.560 144.770 ;
        RECT 95.660 144.650 95.980 144.940 ;
        RECT 93.875 143.800 94.155 144.600 ;
        RECT 94.390 144.480 95.980 144.650 ;
        RECT 94.325 144.020 95.980 144.310 ;
        RECT 96.155 143.970 96.495 144.940 ;
        RECT 96.665 143.800 96.835 144.940 ;
        RECT 97.025 144.770 99.460 144.940 ;
        RECT 97.105 143.800 97.355 144.600 ;
        RECT 98.000 143.970 98.330 144.770 ;
        RECT 98.630 143.800 98.960 144.600 ;
        RECT 99.130 143.970 99.460 144.770 ;
        RECT 99.835 144.890 101.045 145.410 ;
        RECT 101.215 145.060 102.425 145.580 ;
        RECT 99.835 143.800 102.425 144.890 ;
        RECT 102.595 143.800 102.885 144.965 ;
        RECT 103.055 144.890 104.265 145.410 ;
        RECT 104.435 145.060 105.645 145.580 ;
        RECT 105.855 145.530 106.085 146.350 ;
        RECT 106.255 145.550 106.585 146.180 ;
        RECT 105.835 145.110 106.165 145.360 ;
        RECT 106.335 144.950 106.585 145.550 ;
        RECT 106.755 145.530 106.965 146.350 ;
        RECT 107.235 145.530 107.465 146.350 ;
        RECT 107.635 145.550 107.965 146.180 ;
        RECT 107.215 145.110 107.545 145.360 ;
        RECT 107.715 144.950 107.965 145.550 ;
        RECT 108.135 145.530 108.345 146.350 ;
        RECT 108.635 145.530 108.845 146.350 ;
        RECT 109.015 145.550 109.345 146.180 ;
        RECT 103.055 143.800 105.645 144.890 ;
        RECT 105.855 143.800 106.085 144.940 ;
        RECT 106.255 143.970 106.585 144.950 ;
        RECT 106.755 143.800 106.965 144.940 ;
        RECT 107.235 143.800 107.465 144.940 ;
        RECT 107.635 143.970 107.965 144.950 ;
        RECT 109.015 144.950 109.265 145.550 ;
        RECT 109.515 145.530 109.745 146.350 ;
        RECT 110.875 145.580 114.385 146.350 ;
        RECT 114.555 145.600 115.765 146.350 ;
        RECT 109.435 145.110 109.765 145.360 ;
        RECT 108.135 143.800 108.345 144.940 ;
        RECT 108.635 143.800 108.845 144.940 ;
        RECT 109.015 143.970 109.345 144.950 ;
        RECT 109.515 143.800 109.745 144.940 ;
        RECT 110.875 144.890 112.565 145.410 ;
        RECT 112.735 145.060 114.385 145.580 ;
        RECT 114.555 144.890 115.075 145.430 ;
        RECT 115.245 145.060 115.765 145.600 ;
        RECT 110.875 143.800 114.385 144.890 ;
        RECT 114.555 143.800 115.765 144.890 ;
        RECT 14.650 143.630 115.850 143.800 ;
        RECT 14.735 142.540 15.945 143.630 ;
        RECT 14.735 141.830 15.255 142.370 ;
        RECT 15.425 142.000 15.945 142.540 ;
        RECT 16.490 142.650 16.745 143.320 ;
        RECT 16.925 142.830 17.210 143.630 ;
        RECT 17.390 142.910 17.720 143.420 ;
        RECT 14.735 141.080 15.945 141.830 ;
        RECT 16.490 141.790 16.670 142.650 ;
        RECT 17.390 142.320 17.640 142.910 ;
        RECT 17.990 142.760 18.160 143.370 ;
        RECT 18.330 142.940 18.660 143.630 ;
        RECT 18.890 143.080 19.130 143.370 ;
        RECT 19.330 143.250 19.750 143.630 ;
        RECT 19.930 143.160 20.560 143.410 ;
        RECT 21.030 143.250 21.360 143.630 ;
        RECT 19.930 143.080 20.100 143.160 ;
        RECT 21.530 143.080 21.700 143.370 ;
        RECT 21.880 143.250 22.260 143.630 ;
        RECT 22.500 143.245 23.330 143.415 ;
        RECT 18.890 142.910 20.100 143.080 ;
        RECT 16.840 141.990 17.640 142.320 ;
        RECT 16.490 141.590 16.745 141.790 ;
        RECT 16.405 141.420 16.745 141.590 ;
        RECT 16.490 141.260 16.745 141.420 ;
        RECT 16.925 141.080 17.210 141.540 ;
        RECT 17.390 141.340 17.640 141.990 ;
        RECT 17.840 142.740 18.160 142.760 ;
        RECT 17.840 142.570 19.760 142.740 ;
        RECT 17.840 141.675 18.030 142.570 ;
        RECT 19.930 142.400 20.100 142.910 ;
        RECT 20.270 142.650 20.790 142.960 ;
        RECT 18.200 142.230 20.100 142.400 ;
        RECT 18.200 142.170 18.530 142.230 ;
        RECT 18.680 142.000 19.010 142.060 ;
        RECT 18.350 141.730 19.010 142.000 ;
        RECT 17.840 141.345 18.160 141.675 ;
        RECT 18.340 141.080 19.000 141.560 ;
        RECT 19.200 141.470 19.370 142.230 ;
        RECT 20.270 142.060 20.450 142.470 ;
        RECT 19.540 141.890 19.870 142.010 ;
        RECT 20.620 141.890 20.790 142.650 ;
        RECT 19.540 141.720 20.790 141.890 ;
        RECT 20.960 142.830 22.330 143.080 ;
        RECT 20.960 142.060 21.150 142.830 ;
        RECT 22.080 142.570 22.330 142.830 ;
        RECT 21.320 142.400 21.570 142.560 ;
        RECT 22.500 142.400 22.670 143.245 ;
        RECT 23.565 142.960 23.735 143.460 ;
        RECT 23.905 143.130 24.235 143.630 ;
        RECT 22.840 142.570 23.340 142.950 ;
        RECT 23.565 142.790 24.260 142.960 ;
        RECT 21.320 142.230 22.670 142.400 ;
        RECT 22.250 142.190 22.670 142.230 ;
        RECT 20.960 141.720 21.380 142.060 ;
        RECT 21.670 141.730 22.080 142.060 ;
        RECT 19.200 141.300 20.050 141.470 ;
        RECT 20.610 141.080 20.930 141.540 ;
        RECT 21.130 141.290 21.380 141.720 ;
        RECT 21.670 141.080 22.080 141.520 ;
        RECT 22.250 141.460 22.420 142.190 ;
        RECT 22.590 141.640 22.940 142.010 ;
        RECT 23.120 141.700 23.340 142.570 ;
        RECT 23.510 142.000 23.920 142.620 ;
        RECT 24.090 141.820 24.260 142.790 ;
        RECT 23.565 141.630 24.260 141.820 ;
        RECT 22.250 141.260 23.265 141.460 ;
        RECT 23.565 141.300 23.735 141.630 ;
        RECT 23.905 141.080 24.235 141.460 ;
        RECT 24.450 141.340 24.675 143.460 ;
        RECT 24.845 143.130 25.175 143.630 ;
        RECT 25.345 142.960 25.515 143.460 ;
        RECT 24.850 142.790 25.515 142.960 ;
        RECT 24.850 141.800 25.080 142.790 ;
        RECT 25.250 141.970 25.600 142.620 ;
        RECT 26.235 142.540 29.745 143.630 ;
        RECT 26.235 142.020 27.925 142.540 ;
        RECT 29.915 142.490 30.185 143.460 ;
        RECT 30.395 142.830 30.675 143.630 ;
        RECT 30.845 143.120 32.500 143.410 ;
        RECT 30.910 142.780 32.500 142.950 ;
        RECT 30.910 142.660 31.080 142.780 ;
        RECT 30.355 142.490 31.080 142.660 ;
        RECT 28.095 141.850 29.745 142.370 ;
        RECT 24.850 141.630 25.515 141.800 ;
        RECT 24.845 141.080 25.175 141.460 ;
        RECT 25.345 141.340 25.515 141.630 ;
        RECT 26.235 141.080 29.745 141.850 ;
        RECT 29.915 141.755 30.085 142.490 ;
        RECT 30.355 142.320 30.525 142.490 ;
        RECT 31.270 142.440 31.985 142.610 ;
        RECT 32.180 142.490 32.500 142.780 ;
        RECT 32.675 142.490 32.945 143.460 ;
        RECT 33.155 142.830 33.435 143.630 ;
        RECT 33.605 143.120 35.260 143.410 ;
        RECT 33.670 142.780 35.260 142.950 ;
        RECT 33.670 142.660 33.840 142.780 ;
        RECT 33.115 142.490 33.840 142.660 ;
        RECT 30.255 141.990 30.525 142.320 ;
        RECT 30.695 141.990 31.100 142.320 ;
        RECT 31.270 141.990 31.980 142.440 ;
        RECT 30.355 141.820 30.525 141.990 ;
        RECT 29.915 141.410 30.185 141.755 ;
        RECT 30.355 141.650 31.965 141.820 ;
        RECT 32.150 141.750 32.500 142.320 ;
        RECT 32.675 141.755 32.845 142.490 ;
        RECT 33.115 142.320 33.285 142.490 ;
        RECT 33.015 141.990 33.285 142.320 ;
        RECT 33.455 141.990 33.860 142.320 ;
        RECT 34.030 141.990 34.740 142.610 ;
        RECT 34.940 142.490 35.260 142.780 ;
        RECT 35.435 142.540 36.645 143.630 ;
        RECT 33.115 141.820 33.285 141.990 ;
        RECT 30.375 141.080 30.755 141.480 ;
        RECT 30.925 141.300 31.095 141.650 ;
        RECT 31.265 141.080 31.595 141.480 ;
        RECT 31.795 141.300 31.965 141.650 ;
        RECT 32.165 141.080 32.495 141.580 ;
        RECT 32.675 141.410 32.945 141.755 ;
        RECT 33.115 141.650 34.725 141.820 ;
        RECT 34.910 141.750 35.260 142.320 ;
        RECT 35.435 142.000 35.955 142.540 ;
        RECT 36.855 142.490 37.085 143.630 ;
        RECT 37.255 142.480 37.585 143.460 ;
        RECT 37.755 142.490 37.965 143.630 ;
        RECT 36.125 141.830 36.645 142.370 ;
        RECT 36.835 142.070 37.165 142.320 ;
        RECT 33.135 141.080 33.515 141.480 ;
        RECT 33.685 141.300 33.855 141.650 ;
        RECT 34.025 141.080 34.355 141.480 ;
        RECT 34.555 141.300 34.725 141.650 ;
        RECT 34.925 141.080 35.255 141.580 ;
        RECT 35.435 141.080 36.645 141.830 ;
        RECT 36.855 141.080 37.085 141.900 ;
        RECT 37.335 141.880 37.585 142.480 ;
        RECT 38.195 142.465 38.485 143.630 ;
        RECT 38.655 142.540 39.865 143.630 ;
        RECT 40.035 142.555 40.305 143.460 ;
        RECT 40.475 142.870 40.805 143.630 ;
        RECT 40.985 142.700 41.155 143.460 ;
        RECT 38.655 142.000 39.175 142.540 ;
        RECT 37.255 141.250 37.585 141.880 ;
        RECT 37.755 141.080 37.965 141.900 ;
        RECT 39.345 141.830 39.865 142.370 ;
        RECT 38.195 141.080 38.485 141.805 ;
        RECT 38.655 141.080 39.865 141.830 ;
        RECT 40.035 141.755 40.205 142.555 ;
        RECT 40.490 142.530 41.155 142.700 ;
        RECT 40.490 142.385 40.660 142.530 ;
        RECT 40.375 142.055 40.660 142.385 ;
        RECT 41.420 142.490 41.755 143.460 ;
        RECT 41.925 142.490 42.095 143.630 ;
        RECT 42.265 143.290 44.295 143.460 ;
        RECT 40.490 141.800 40.660 142.055 ;
        RECT 40.895 141.980 41.225 142.350 ;
        RECT 41.420 141.820 41.590 142.490 ;
        RECT 42.265 142.320 42.435 143.290 ;
        RECT 41.760 141.990 42.015 142.320 ;
        RECT 42.240 141.990 42.435 142.320 ;
        RECT 42.605 142.950 43.730 143.120 ;
        RECT 41.845 141.820 42.015 141.990 ;
        RECT 42.605 141.820 42.775 142.950 ;
        RECT 40.035 141.250 40.295 141.755 ;
        RECT 40.490 141.630 41.155 141.800 ;
        RECT 40.475 141.080 40.805 141.460 ;
        RECT 40.985 141.250 41.155 141.630 ;
        RECT 41.420 141.250 41.675 141.820 ;
        RECT 41.845 141.650 42.775 141.820 ;
        RECT 42.945 142.610 43.955 142.780 ;
        RECT 42.945 141.810 43.115 142.610 ;
        RECT 43.320 142.270 43.595 142.410 ;
        RECT 43.315 142.100 43.595 142.270 ;
        RECT 42.600 141.615 42.775 141.650 ;
        RECT 41.845 141.080 42.175 141.480 ;
        RECT 42.600 141.250 43.130 141.615 ;
        RECT 43.320 141.250 43.595 142.100 ;
        RECT 43.765 141.250 43.955 142.610 ;
        RECT 44.125 142.625 44.295 143.290 ;
        RECT 44.465 142.870 44.635 143.630 ;
        RECT 44.870 142.870 45.385 143.280 ;
        RECT 44.125 142.435 44.875 142.625 ;
        RECT 45.045 142.060 45.385 142.870 ;
        RECT 44.155 141.890 45.385 142.060 ;
        RECT 46.015 142.540 47.685 143.630 ;
        RECT 48.230 142.650 48.485 143.320 ;
        RECT 48.665 142.830 48.950 143.630 ;
        RECT 49.130 142.910 49.460 143.420 ;
        RECT 46.015 142.020 46.765 142.540 ;
        RECT 44.135 141.080 44.645 141.615 ;
        RECT 44.865 141.285 45.110 141.890 ;
        RECT 46.935 141.850 47.685 142.370 ;
        RECT 46.015 141.080 47.685 141.850 ;
        RECT 48.230 141.790 48.410 142.650 ;
        RECT 49.130 142.320 49.380 142.910 ;
        RECT 49.730 142.760 49.900 143.370 ;
        RECT 50.070 142.940 50.400 143.630 ;
        RECT 50.630 143.080 50.870 143.370 ;
        RECT 51.070 143.250 51.490 143.630 ;
        RECT 51.670 143.160 52.300 143.410 ;
        RECT 52.770 143.250 53.100 143.630 ;
        RECT 51.670 143.080 51.840 143.160 ;
        RECT 53.270 143.080 53.440 143.370 ;
        RECT 53.620 143.250 54.000 143.630 ;
        RECT 54.240 143.245 55.070 143.415 ;
        RECT 50.630 142.910 51.840 143.080 ;
        RECT 48.580 141.990 49.380 142.320 ;
        RECT 48.230 141.590 48.485 141.790 ;
        RECT 48.145 141.420 48.485 141.590 ;
        RECT 48.230 141.260 48.485 141.420 ;
        RECT 48.665 141.080 48.950 141.540 ;
        RECT 49.130 141.340 49.380 141.990 ;
        RECT 49.580 142.740 49.900 142.760 ;
        RECT 49.580 142.570 51.500 142.740 ;
        RECT 49.580 141.675 49.770 142.570 ;
        RECT 51.670 142.400 51.840 142.910 ;
        RECT 52.010 142.650 52.530 142.960 ;
        RECT 49.940 142.230 51.840 142.400 ;
        RECT 49.940 142.170 50.270 142.230 ;
        RECT 50.420 142.000 50.750 142.060 ;
        RECT 50.090 141.730 50.750 142.000 ;
        RECT 49.580 141.345 49.900 141.675 ;
        RECT 50.080 141.080 50.740 141.560 ;
        RECT 50.940 141.470 51.110 142.230 ;
        RECT 52.010 142.060 52.190 142.470 ;
        RECT 51.280 141.890 51.610 142.010 ;
        RECT 52.360 141.890 52.530 142.650 ;
        RECT 51.280 141.720 52.530 141.890 ;
        RECT 52.700 142.830 54.070 143.080 ;
        RECT 52.700 142.060 52.890 142.830 ;
        RECT 53.820 142.570 54.070 142.830 ;
        RECT 53.060 142.400 53.310 142.560 ;
        RECT 54.240 142.400 54.410 143.245 ;
        RECT 55.305 142.960 55.475 143.460 ;
        RECT 55.645 143.130 55.975 143.630 ;
        RECT 54.580 142.570 55.080 142.950 ;
        RECT 55.305 142.790 56.000 142.960 ;
        RECT 53.060 142.230 54.410 142.400 ;
        RECT 53.990 142.190 54.410 142.230 ;
        RECT 52.700 141.720 53.120 142.060 ;
        RECT 53.410 141.730 53.820 142.060 ;
        RECT 50.940 141.300 51.790 141.470 ;
        RECT 52.350 141.080 52.670 141.540 ;
        RECT 52.870 141.290 53.120 141.720 ;
        RECT 53.410 141.080 53.820 141.520 ;
        RECT 53.990 141.460 54.160 142.190 ;
        RECT 54.330 141.640 54.680 142.010 ;
        RECT 54.860 141.700 55.080 142.570 ;
        RECT 55.250 142.000 55.660 142.620 ;
        RECT 55.830 141.820 56.000 142.790 ;
        RECT 55.305 141.630 56.000 141.820 ;
        RECT 53.990 141.260 55.005 141.460 ;
        RECT 55.305 141.300 55.475 141.630 ;
        RECT 55.645 141.080 55.975 141.460 ;
        RECT 56.190 141.340 56.415 143.460 ;
        RECT 56.585 143.130 56.915 143.630 ;
        RECT 57.085 142.960 57.255 143.460 ;
        RECT 56.590 142.790 57.255 142.960 ;
        RECT 56.590 141.800 56.820 142.790 ;
        RECT 56.990 141.970 57.340 142.620 ;
        RECT 57.515 142.490 57.855 143.460 ;
        RECT 58.025 142.490 58.195 143.630 ;
        RECT 58.465 142.830 58.715 143.630 ;
        RECT 59.360 142.660 59.690 143.460 ;
        RECT 59.990 142.830 60.320 143.630 ;
        RECT 60.490 142.660 60.820 143.460 ;
        RECT 58.385 142.490 60.820 142.660 ;
        RECT 61.195 142.540 63.785 143.630 ;
        RECT 57.515 141.880 57.690 142.490 ;
        RECT 58.385 142.240 58.555 142.490 ;
        RECT 57.860 142.070 58.555 142.240 ;
        RECT 58.730 142.070 59.150 142.270 ;
        RECT 59.320 142.070 59.650 142.270 ;
        RECT 59.820 142.070 60.150 142.270 ;
        RECT 56.590 141.630 57.255 141.800 ;
        RECT 56.585 141.080 56.915 141.460 ;
        RECT 57.085 141.340 57.255 141.630 ;
        RECT 57.515 141.250 57.855 141.880 ;
        RECT 58.025 141.080 58.275 141.880 ;
        RECT 58.465 141.730 59.690 141.900 ;
        RECT 58.465 141.250 58.795 141.730 ;
        RECT 58.965 141.080 59.190 141.540 ;
        RECT 59.360 141.250 59.690 141.730 ;
        RECT 60.320 141.860 60.490 142.490 ;
        RECT 60.675 142.070 61.025 142.320 ;
        RECT 61.195 142.020 62.405 142.540 ;
        RECT 63.955 142.465 64.245 143.630 ;
        RECT 64.475 142.490 64.685 143.630 ;
        RECT 64.855 142.480 65.185 143.460 ;
        RECT 65.355 142.490 65.585 143.630 ;
        RECT 65.885 142.700 66.055 143.460 ;
        RECT 66.235 142.870 66.565 143.630 ;
        RECT 65.885 142.530 66.550 142.700 ;
        RECT 66.735 142.555 67.005 143.460 ;
        RECT 60.320 141.250 60.820 141.860 ;
        RECT 62.575 141.850 63.785 142.370 ;
        RECT 61.195 141.080 63.785 141.850 ;
        RECT 63.955 141.080 64.245 141.805 ;
        RECT 64.475 141.080 64.685 141.900 ;
        RECT 64.855 141.880 65.105 142.480 ;
        RECT 66.380 142.385 66.550 142.530 ;
        RECT 65.275 142.070 65.605 142.320 ;
        RECT 65.815 141.980 66.145 142.350 ;
        RECT 66.380 142.055 66.665 142.385 ;
        RECT 64.855 141.250 65.185 141.880 ;
        RECT 65.355 141.080 65.585 141.900 ;
        RECT 66.380 141.800 66.550 142.055 ;
        RECT 65.885 141.630 66.550 141.800 ;
        RECT 66.835 141.755 67.005 142.555 ;
        RECT 67.175 142.540 70.685 143.630 ;
        RECT 70.860 143.195 76.205 143.630 ;
        RECT 67.175 142.020 68.865 142.540 ;
        RECT 69.035 141.850 70.685 142.370 ;
        RECT 72.450 141.945 72.800 143.195 ;
        RECT 76.375 142.870 76.890 143.280 ;
        RECT 77.125 142.870 77.295 143.630 ;
        RECT 77.465 143.290 79.495 143.460 ;
        RECT 65.885 141.250 66.055 141.630 ;
        RECT 66.235 141.080 66.565 141.460 ;
        RECT 66.745 141.250 67.005 141.755 ;
        RECT 67.175 141.080 70.685 141.850 ;
        RECT 74.280 141.625 74.620 142.455 ;
        RECT 76.375 142.060 76.715 142.870 ;
        RECT 77.465 142.625 77.635 143.290 ;
        RECT 78.030 142.950 79.155 143.120 ;
        RECT 76.885 142.435 77.635 142.625 ;
        RECT 77.805 142.610 78.815 142.780 ;
        RECT 76.375 141.890 77.605 142.060 ;
        RECT 70.860 141.080 76.205 141.625 ;
        RECT 76.650 141.285 76.895 141.890 ;
        RECT 77.115 141.080 77.625 141.615 ;
        RECT 77.805 141.250 77.995 142.610 ;
        RECT 78.165 141.590 78.440 142.410 ;
        RECT 78.645 141.810 78.815 142.610 ;
        RECT 78.985 141.820 79.155 142.950 ;
        RECT 79.325 142.320 79.495 143.290 ;
        RECT 79.665 142.490 79.835 143.630 ;
        RECT 80.005 142.490 80.340 143.460 ;
        RECT 81.440 143.195 86.785 143.630 ;
        RECT 79.325 141.990 79.520 142.320 ;
        RECT 79.745 141.990 80.000 142.320 ;
        RECT 79.745 141.820 79.915 141.990 ;
        RECT 80.170 141.820 80.340 142.490 ;
        RECT 83.030 141.945 83.380 143.195 ;
        RECT 86.955 142.490 87.225 143.460 ;
        RECT 87.435 142.830 87.715 143.630 ;
        RECT 87.885 143.120 89.540 143.410 ;
        RECT 87.950 142.780 89.540 142.950 ;
        RECT 87.950 142.660 88.120 142.780 ;
        RECT 87.395 142.490 88.120 142.660 ;
        RECT 78.985 141.650 79.915 141.820 ;
        RECT 78.985 141.615 79.160 141.650 ;
        RECT 78.165 141.420 78.445 141.590 ;
        RECT 78.165 141.250 78.440 141.420 ;
        RECT 78.630 141.250 79.160 141.615 ;
        RECT 79.585 141.080 79.915 141.480 ;
        RECT 80.085 141.250 80.340 141.820 ;
        RECT 84.860 141.625 85.200 142.455 ;
        RECT 86.955 141.755 87.125 142.490 ;
        RECT 87.395 142.320 87.565 142.490 ;
        RECT 88.310 142.440 89.025 142.610 ;
        RECT 89.220 142.490 89.540 142.780 ;
        RECT 89.715 142.465 90.005 143.630 ;
        RECT 90.175 142.490 90.515 143.460 ;
        RECT 90.685 142.490 90.855 143.630 ;
        RECT 91.125 142.830 91.375 143.630 ;
        RECT 92.020 142.660 92.350 143.460 ;
        RECT 92.650 142.830 92.980 143.630 ;
        RECT 93.150 142.660 93.480 143.460 ;
        RECT 91.045 142.490 93.480 142.660 ;
        RECT 93.860 142.490 94.195 143.460 ;
        RECT 94.365 142.490 94.535 143.630 ;
        RECT 94.705 143.290 96.735 143.460 ;
        RECT 87.295 141.990 87.565 142.320 ;
        RECT 87.735 141.990 88.140 142.320 ;
        RECT 88.310 141.990 89.020 142.440 ;
        RECT 87.395 141.820 87.565 141.990 ;
        RECT 81.440 141.080 86.785 141.625 ;
        RECT 86.955 141.410 87.225 141.755 ;
        RECT 87.395 141.650 89.005 141.820 ;
        RECT 89.190 141.750 89.540 142.320 ;
        RECT 90.175 141.930 90.350 142.490 ;
        RECT 91.045 142.240 91.215 142.490 ;
        RECT 90.520 142.070 91.215 142.240 ;
        RECT 91.390 142.070 91.810 142.270 ;
        RECT 91.980 142.070 92.310 142.270 ;
        RECT 92.480 142.070 92.810 142.270 ;
        RECT 90.175 141.880 90.405 141.930 ;
        RECT 87.415 141.080 87.795 141.480 ;
        RECT 87.965 141.300 88.135 141.650 ;
        RECT 88.305 141.080 88.635 141.480 ;
        RECT 88.835 141.300 89.005 141.650 ;
        RECT 89.205 141.080 89.535 141.580 ;
        RECT 89.715 141.080 90.005 141.805 ;
        RECT 90.175 141.250 90.515 141.880 ;
        RECT 90.685 141.080 90.935 141.880 ;
        RECT 91.125 141.730 92.350 141.900 ;
        RECT 91.125 141.250 91.455 141.730 ;
        RECT 91.625 141.080 91.850 141.540 ;
        RECT 92.020 141.250 92.350 141.730 ;
        RECT 92.980 141.860 93.150 142.490 ;
        RECT 93.335 142.070 93.685 142.320 ;
        RECT 92.980 141.250 93.480 141.860 ;
        RECT 93.860 141.820 94.030 142.490 ;
        RECT 94.705 142.320 94.875 143.290 ;
        RECT 94.200 141.990 94.455 142.320 ;
        RECT 94.680 141.990 94.875 142.320 ;
        RECT 95.045 142.950 96.170 143.120 ;
        RECT 94.285 141.820 94.455 141.990 ;
        RECT 95.045 141.820 95.215 142.950 ;
        RECT 93.860 141.250 94.115 141.820 ;
        RECT 94.285 141.650 95.215 141.820 ;
        RECT 95.385 142.610 96.395 142.780 ;
        RECT 95.385 141.810 95.555 142.610 ;
        RECT 95.040 141.615 95.215 141.650 ;
        RECT 94.285 141.080 94.615 141.480 ;
        RECT 95.040 141.250 95.570 141.615 ;
        RECT 95.760 141.590 96.035 142.410 ;
        RECT 95.755 141.420 96.035 141.590 ;
        RECT 95.760 141.250 96.035 141.420 ;
        RECT 96.205 141.250 96.395 142.610 ;
        RECT 96.565 142.625 96.735 143.290 ;
        RECT 96.905 142.870 97.075 143.630 ;
        RECT 97.310 142.870 97.825 143.280 ;
        RECT 96.565 142.435 97.315 142.625 ;
        RECT 97.485 142.060 97.825 142.870 ;
        RECT 96.595 141.890 97.825 142.060 ;
        RECT 97.995 142.540 100.585 143.630 ;
        RECT 100.755 142.870 101.270 143.280 ;
        RECT 101.505 142.870 101.675 143.630 ;
        RECT 101.845 143.290 103.875 143.460 ;
        RECT 97.995 142.020 99.205 142.540 ;
        RECT 96.575 141.080 97.085 141.615 ;
        RECT 97.305 141.285 97.550 141.890 ;
        RECT 99.375 141.850 100.585 142.370 ;
        RECT 100.755 142.060 101.095 142.870 ;
        RECT 101.845 142.625 102.015 143.290 ;
        RECT 102.410 142.950 103.535 143.120 ;
        RECT 101.265 142.435 102.015 142.625 ;
        RECT 102.185 142.610 103.195 142.780 ;
        RECT 100.755 141.890 101.985 142.060 ;
        RECT 97.995 141.080 100.585 141.850 ;
        RECT 101.030 141.285 101.275 141.890 ;
        RECT 101.495 141.080 102.005 141.615 ;
        RECT 102.185 141.250 102.375 142.610 ;
        RECT 102.545 142.270 102.820 142.410 ;
        RECT 102.545 142.100 102.825 142.270 ;
        RECT 102.545 141.250 102.820 142.100 ;
        RECT 103.025 141.810 103.195 142.610 ;
        RECT 103.365 141.820 103.535 142.950 ;
        RECT 103.705 142.320 103.875 143.290 ;
        RECT 104.045 142.490 104.215 143.630 ;
        RECT 104.385 142.490 104.720 143.460 ;
        RECT 103.705 141.990 103.900 142.320 ;
        RECT 104.125 141.990 104.380 142.320 ;
        RECT 104.125 141.820 104.295 141.990 ;
        RECT 104.550 141.820 104.720 142.490 ;
        RECT 105.270 142.650 105.525 143.320 ;
        RECT 105.705 142.830 105.990 143.630 ;
        RECT 106.170 142.910 106.500 143.420 ;
        RECT 105.270 141.930 105.450 142.650 ;
        RECT 106.170 142.320 106.420 142.910 ;
        RECT 106.770 142.760 106.940 143.370 ;
        RECT 107.110 142.940 107.440 143.630 ;
        RECT 107.670 143.080 107.910 143.370 ;
        RECT 108.110 143.250 108.530 143.630 ;
        RECT 108.710 143.160 109.340 143.410 ;
        RECT 109.810 143.250 110.140 143.630 ;
        RECT 108.710 143.080 108.880 143.160 ;
        RECT 110.310 143.080 110.480 143.370 ;
        RECT 110.660 143.250 111.040 143.630 ;
        RECT 111.280 143.245 112.110 143.415 ;
        RECT 107.670 142.910 108.880 143.080 ;
        RECT 105.620 141.990 106.420 142.320 ;
        RECT 103.365 141.650 104.295 141.820 ;
        RECT 103.365 141.615 103.540 141.650 ;
        RECT 103.010 141.250 103.540 141.615 ;
        RECT 103.965 141.080 104.295 141.480 ;
        RECT 104.465 141.250 104.720 141.820 ;
        RECT 105.185 141.790 105.450 141.930 ;
        RECT 105.185 141.760 105.525 141.790 ;
        RECT 105.270 141.260 105.525 141.760 ;
        RECT 105.705 141.080 105.990 141.540 ;
        RECT 106.170 141.340 106.420 141.990 ;
        RECT 106.620 142.740 106.940 142.760 ;
        RECT 106.620 142.570 108.540 142.740 ;
        RECT 106.620 141.675 106.810 142.570 ;
        RECT 108.710 142.400 108.880 142.910 ;
        RECT 109.050 142.650 109.570 142.960 ;
        RECT 106.980 142.230 108.880 142.400 ;
        RECT 106.980 142.170 107.310 142.230 ;
        RECT 107.460 142.000 107.790 142.060 ;
        RECT 107.130 141.730 107.790 142.000 ;
        RECT 106.620 141.345 106.940 141.675 ;
        RECT 107.120 141.080 107.780 141.560 ;
        RECT 107.980 141.470 108.150 142.230 ;
        RECT 109.050 142.060 109.230 142.470 ;
        RECT 108.320 141.890 108.650 142.010 ;
        RECT 109.400 141.890 109.570 142.650 ;
        RECT 108.320 141.720 109.570 141.890 ;
        RECT 109.740 142.830 111.110 143.080 ;
        RECT 109.740 142.060 109.930 142.830 ;
        RECT 110.860 142.570 111.110 142.830 ;
        RECT 110.100 142.400 110.350 142.560 ;
        RECT 111.280 142.400 111.450 143.245 ;
        RECT 112.345 142.960 112.515 143.460 ;
        RECT 112.685 143.130 113.015 143.630 ;
        RECT 111.620 142.570 112.120 142.950 ;
        RECT 112.345 142.790 113.040 142.960 ;
        RECT 110.100 142.230 111.450 142.400 ;
        RECT 111.030 142.190 111.450 142.230 ;
        RECT 109.740 141.720 110.160 142.060 ;
        RECT 110.450 141.730 110.860 142.060 ;
        RECT 107.980 141.300 108.830 141.470 ;
        RECT 109.390 141.080 109.710 141.540 ;
        RECT 109.910 141.290 110.160 141.720 ;
        RECT 110.450 141.080 110.860 141.520 ;
        RECT 111.030 141.460 111.200 142.190 ;
        RECT 111.370 141.640 111.720 142.010 ;
        RECT 111.900 141.700 112.120 142.570 ;
        RECT 112.290 142.000 112.700 142.620 ;
        RECT 112.870 141.820 113.040 142.790 ;
        RECT 112.345 141.630 113.040 141.820 ;
        RECT 111.030 141.260 112.045 141.460 ;
        RECT 112.345 141.300 112.515 141.630 ;
        RECT 112.685 141.080 113.015 141.460 ;
        RECT 113.230 141.340 113.455 143.460 ;
        RECT 113.625 143.130 113.955 143.630 ;
        RECT 114.125 142.960 114.295 143.460 ;
        RECT 113.630 142.790 114.295 142.960 ;
        RECT 113.630 141.800 113.860 142.790 ;
        RECT 114.030 141.970 114.380 142.620 ;
        RECT 114.555 142.540 115.765 143.630 ;
        RECT 114.555 142.000 115.075 142.540 ;
        RECT 115.245 141.830 115.765 142.370 ;
        RECT 113.630 141.630 114.295 141.800 ;
        RECT 113.625 141.080 113.955 141.460 ;
        RECT 114.125 141.340 114.295 141.630 ;
        RECT 114.555 141.080 115.765 141.830 ;
        RECT 14.650 140.910 115.850 141.080 ;
        RECT 14.735 140.160 15.945 140.910 ;
        RECT 16.115 140.160 17.325 140.910 ;
        RECT 14.735 139.620 15.255 140.160 ;
        RECT 15.425 139.450 15.945 139.990 ;
        RECT 14.735 138.360 15.945 139.450 ;
        RECT 16.115 139.450 16.635 139.990 ;
        RECT 16.805 139.620 17.325 140.160 ;
        RECT 17.495 140.140 21.005 140.910 ;
        RECT 17.495 139.450 19.185 139.970 ;
        RECT 19.355 139.620 21.005 140.140 ;
        RECT 21.215 140.090 21.445 140.910 ;
        RECT 21.615 140.110 21.945 140.740 ;
        RECT 21.195 139.670 21.525 139.920 ;
        RECT 21.695 139.510 21.945 140.110 ;
        RECT 22.115 140.090 22.325 140.910 ;
        RECT 22.645 140.360 22.815 140.740 ;
        RECT 22.995 140.530 23.325 140.910 ;
        RECT 22.645 140.190 23.310 140.360 ;
        RECT 23.505 140.235 23.765 140.740 ;
        RECT 22.575 139.640 22.905 140.010 ;
        RECT 23.140 139.935 23.310 140.190 ;
        RECT 16.115 138.360 17.325 139.450 ;
        RECT 17.495 138.360 21.005 139.450 ;
        RECT 21.215 138.360 21.445 139.500 ;
        RECT 21.615 138.530 21.945 139.510 ;
        RECT 23.140 139.605 23.425 139.935 ;
        RECT 22.115 138.360 22.325 139.500 ;
        RECT 23.140 139.460 23.310 139.605 ;
        RECT 22.645 139.290 23.310 139.460 ;
        RECT 23.595 139.435 23.765 140.235 ;
        RECT 23.935 140.160 25.145 140.910 ;
        RECT 25.315 140.185 25.605 140.910 ;
        RECT 25.775 140.160 26.985 140.910 ;
        RECT 22.645 138.530 22.815 139.290 ;
        RECT 22.995 138.360 23.325 139.120 ;
        RECT 23.495 138.530 23.765 139.435 ;
        RECT 23.935 139.450 24.455 139.990 ;
        RECT 24.625 139.620 25.145 140.160 ;
        RECT 23.935 138.360 25.145 139.450 ;
        RECT 25.315 138.360 25.605 139.525 ;
        RECT 25.775 139.450 26.295 139.990 ;
        RECT 26.465 139.620 26.985 140.160 ;
        RECT 27.155 140.235 27.415 140.740 ;
        RECT 27.595 140.530 27.925 140.910 ;
        RECT 28.105 140.360 28.275 140.740 ;
        RECT 25.775 138.360 26.985 139.450 ;
        RECT 27.155 139.435 27.325 140.235 ;
        RECT 27.610 140.190 28.275 140.360 ;
        RECT 27.610 139.935 27.780 140.190 ;
        RECT 28.535 140.160 29.745 140.910 ;
        RECT 27.495 139.605 27.780 139.935 ;
        RECT 28.015 139.640 28.345 140.010 ;
        RECT 27.610 139.460 27.780 139.605 ;
        RECT 27.155 138.530 27.425 139.435 ;
        RECT 27.610 139.290 28.275 139.460 ;
        RECT 27.595 138.360 27.925 139.120 ;
        RECT 28.105 138.530 28.275 139.290 ;
        RECT 28.535 139.450 29.055 139.990 ;
        RECT 29.225 139.620 29.745 140.160 ;
        RECT 30.115 140.280 30.445 140.640 ;
        RECT 31.065 140.450 31.315 140.910 ;
        RECT 31.485 140.450 32.045 140.740 ;
        RECT 30.115 140.090 31.505 140.280 ;
        RECT 31.335 140.000 31.505 140.090 ;
        RECT 29.930 139.670 30.605 139.920 ;
        RECT 30.825 139.670 31.165 139.920 ;
        RECT 31.335 139.670 31.625 140.000 ;
        RECT 28.535 138.360 29.745 139.450 ;
        RECT 29.930 139.310 30.195 139.670 ;
        RECT 31.335 139.420 31.505 139.670 ;
        RECT 30.565 139.250 31.505 139.420 ;
        RECT 30.115 138.360 30.395 139.030 ;
        RECT 30.565 138.700 30.865 139.250 ;
        RECT 31.795 139.080 32.045 140.450 ;
        RECT 32.215 140.140 35.725 140.910 ;
        RECT 35.900 140.365 41.245 140.910 ;
        RECT 41.420 140.365 46.765 140.910 ;
        RECT 31.065 138.360 31.395 139.080 ;
        RECT 31.585 138.530 32.045 139.080 ;
        RECT 32.215 139.450 33.905 139.970 ;
        RECT 34.075 139.620 35.725 140.140 ;
        RECT 32.215 138.360 35.725 139.450 ;
        RECT 37.490 138.795 37.840 140.045 ;
        RECT 39.320 139.535 39.660 140.365 ;
        RECT 43.010 138.795 43.360 140.045 ;
        RECT 44.840 139.535 45.180 140.365 ;
        RECT 47.210 140.100 47.455 140.705 ;
        RECT 47.675 140.375 48.185 140.910 ;
        RECT 46.935 139.930 48.165 140.100 ;
        RECT 46.935 139.120 47.275 139.930 ;
        RECT 47.445 139.365 48.195 139.555 ;
        RECT 35.900 138.360 41.245 138.795 ;
        RECT 41.420 138.360 46.765 138.795 ;
        RECT 46.935 138.710 47.450 139.120 ;
        RECT 47.685 138.360 47.855 139.120 ;
        RECT 48.025 138.700 48.195 139.365 ;
        RECT 48.365 139.380 48.555 140.740 ;
        RECT 48.725 140.570 49.000 140.740 ;
        RECT 48.725 140.400 49.005 140.570 ;
        RECT 48.725 139.580 49.000 140.400 ;
        RECT 49.190 140.375 49.720 140.740 ;
        RECT 50.145 140.510 50.475 140.910 ;
        RECT 49.545 140.340 49.720 140.375 ;
        RECT 49.205 139.380 49.375 140.180 ;
        RECT 48.365 139.210 49.375 139.380 ;
        RECT 49.545 140.170 50.475 140.340 ;
        RECT 50.645 140.170 50.900 140.740 ;
        RECT 51.075 140.185 51.365 140.910 ;
        RECT 49.545 139.040 49.715 140.170 ;
        RECT 50.305 140.000 50.475 140.170 ;
        RECT 48.590 138.870 49.715 139.040 ;
        RECT 49.885 139.670 50.080 140.000 ;
        RECT 50.305 139.670 50.560 140.000 ;
        RECT 49.885 138.700 50.055 139.670 ;
        RECT 50.730 139.500 50.900 140.170 ;
        RECT 51.595 140.090 51.805 140.910 ;
        RECT 51.975 140.110 52.305 140.740 ;
        RECT 48.025 138.530 50.055 138.700 ;
        RECT 50.225 138.360 50.395 139.500 ;
        RECT 50.565 138.530 50.900 139.500 ;
        RECT 51.075 138.360 51.365 139.525 ;
        RECT 51.975 139.510 52.225 140.110 ;
        RECT 52.475 140.090 52.705 140.910 ;
        RECT 53.465 140.360 53.635 140.740 ;
        RECT 53.815 140.530 54.145 140.910 ;
        RECT 53.465 140.190 54.130 140.360 ;
        RECT 54.325 140.235 54.585 140.740 ;
        RECT 52.395 139.670 52.725 139.920 ;
        RECT 53.395 139.640 53.725 140.010 ;
        RECT 53.960 139.935 54.130 140.190 ;
        RECT 53.960 139.605 54.245 139.935 ;
        RECT 51.595 138.360 51.805 139.500 ;
        RECT 51.975 138.530 52.305 139.510 ;
        RECT 52.475 138.360 52.705 139.500 ;
        RECT 53.960 139.460 54.130 139.605 ;
        RECT 53.465 139.290 54.130 139.460 ;
        RECT 54.415 139.435 54.585 140.235 ;
        RECT 54.755 140.140 56.425 140.910 ;
        RECT 53.465 138.530 53.635 139.290 ;
        RECT 53.815 138.360 54.145 139.120 ;
        RECT 54.315 138.530 54.585 139.435 ;
        RECT 54.755 139.450 55.505 139.970 ;
        RECT 55.675 139.620 56.425 140.140 ;
        RECT 56.595 140.110 56.935 140.740 ;
        RECT 57.105 140.110 57.355 140.910 ;
        RECT 57.545 140.260 57.875 140.740 ;
        RECT 58.045 140.450 58.270 140.910 ;
        RECT 58.440 140.260 58.770 140.740 ;
        RECT 56.595 140.060 56.825 140.110 ;
        RECT 57.545 140.090 58.770 140.260 ;
        RECT 59.400 140.130 59.900 140.740 ;
        RECT 56.595 139.500 56.770 140.060 ;
        RECT 56.940 139.750 57.635 139.920 ;
        RECT 57.465 139.500 57.635 139.750 ;
        RECT 57.810 139.720 58.230 139.920 ;
        RECT 58.400 139.720 58.730 139.920 ;
        RECT 58.900 139.720 59.230 139.920 ;
        RECT 59.400 139.500 59.570 140.130 ;
        RECT 61.010 140.100 61.255 140.705 ;
        RECT 61.475 140.375 61.985 140.910 ;
        RECT 60.735 139.930 61.965 140.100 ;
        RECT 59.755 139.670 60.105 139.920 ;
        RECT 54.755 138.360 56.425 139.450 ;
        RECT 56.595 138.530 56.935 139.500 ;
        RECT 57.105 138.360 57.275 139.500 ;
        RECT 57.465 139.330 59.900 139.500 ;
        RECT 57.545 138.360 57.795 139.160 ;
        RECT 58.440 138.530 58.770 139.330 ;
        RECT 59.070 138.360 59.400 139.160 ;
        RECT 59.570 138.530 59.900 139.330 ;
        RECT 60.735 139.120 61.075 139.930 ;
        RECT 61.245 139.365 61.995 139.555 ;
        RECT 60.735 138.710 61.250 139.120 ;
        RECT 61.485 138.360 61.655 139.120 ;
        RECT 61.825 138.700 61.995 139.365 ;
        RECT 62.165 139.380 62.355 140.740 ;
        RECT 62.525 139.890 62.800 140.740 ;
        RECT 62.990 140.375 63.520 140.740 ;
        RECT 63.945 140.510 64.275 140.910 ;
        RECT 63.345 140.340 63.520 140.375 ;
        RECT 62.525 139.720 62.805 139.890 ;
        RECT 62.525 139.580 62.800 139.720 ;
        RECT 63.005 139.380 63.175 140.180 ;
        RECT 62.165 139.210 63.175 139.380 ;
        RECT 63.345 140.170 64.275 140.340 ;
        RECT 64.445 140.170 64.700 140.740 ;
        RECT 63.345 139.040 63.515 140.170 ;
        RECT 64.105 140.000 64.275 140.170 ;
        RECT 62.390 138.870 63.515 139.040 ;
        RECT 63.685 139.670 63.880 140.000 ;
        RECT 64.105 139.670 64.360 140.000 ;
        RECT 63.685 138.700 63.855 139.670 ;
        RECT 64.530 139.500 64.700 140.170 ;
        RECT 64.875 140.140 67.465 140.910 ;
        RECT 67.640 140.365 72.985 140.910 ;
        RECT 61.825 138.530 63.855 138.700 ;
        RECT 64.025 138.360 64.195 139.500 ;
        RECT 64.365 138.530 64.700 139.500 ;
        RECT 64.875 139.450 66.085 139.970 ;
        RECT 66.255 139.620 67.465 140.140 ;
        RECT 64.875 138.360 67.465 139.450 ;
        RECT 69.230 138.795 69.580 140.045 ;
        RECT 71.060 139.535 71.400 140.365 ;
        RECT 73.360 140.130 73.860 140.740 ;
        RECT 73.155 139.670 73.505 139.920 ;
        RECT 73.690 139.500 73.860 140.130 ;
        RECT 74.490 140.260 74.820 140.740 ;
        RECT 74.990 140.450 75.215 140.910 ;
        RECT 75.385 140.260 75.715 140.740 ;
        RECT 74.490 140.090 75.715 140.260 ;
        RECT 75.905 140.110 76.155 140.910 ;
        RECT 76.325 140.110 76.665 140.740 ;
        RECT 76.835 140.185 77.125 140.910 ;
        RECT 77.385 140.360 77.555 140.740 ;
        RECT 77.735 140.530 78.065 140.910 ;
        RECT 77.385 140.190 78.050 140.360 ;
        RECT 78.245 140.235 78.505 140.740 ;
        RECT 74.030 139.720 74.360 139.920 ;
        RECT 74.530 139.720 74.860 139.920 ;
        RECT 75.030 139.720 75.450 139.920 ;
        RECT 75.625 139.750 76.320 139.920 ;
        RECT 75.625 139.500 75.795 139.750 ;
        RECT 76.490 139.500 76.665 140.110 ;
        RECT 77.315 139.640 77.645 140.010 ;
        RECT 77.880 139.935 78.050 140.190 ;
        RECT 77.880 139.605 78.165 139.935 ;
        RECT 73.360 139.330 75.795 139.500 ;
        RECT 67.640 138.360 72.985 138.795 ;
        RECT 73.360 138.530 73.690 139.330 ;
        RECT 73.860 138.360 74.190 139.160 ;
        RECT 74.490 138.530 74.820 139.330 ;
        RECT 75.465 138.360 75.715 139.160 ;
        RECT 75.985 138.360 76.155 139.500 ;
        RECT 76.325 138.530 76.665 139.500 ;
        RECT 76.835 138.360 77.125 139.525 ;
        RECT 77.880 139.460 78.050 139.605 ;
        RECT 77.385 139.290 78.050 139.460 ;
        RECT 78.335 139.435 78.505 140.235 ;
        RECT 78.735 140.090 78.945 140.910 ;
        RECT 79.115 140.110 79.445 140.740 ;
        RECT 79.115 139.510 79.365 140.110 ;
        RECT 79.615 140.090 79.845 140.910 ;
        RECT 80.430 140.200 80.685 140.730 ;
        RECT 80.865 140.450 81.150 140.910 ;
        RECT 79.535 139.670 79.865 139.920 ;
        RECT 77.385 138.530 77.555 139.290 ;
        RECT 77.735 138.360 78.065 139.120 ;
        RECT 78.235 138.530 78.505 139.435 ;
        RECT 78.735 138.360 78.945 139.500 ;
        RECT 79.115 138.530 79.445 139.510 ;
        RECT 79.615 138.360 79.845 139.500 ;
        RECT 80.430 139.340 80.610 140.200 ;
        RECT 81.330 140.000 81.580 140.650 ;
        RECT 80.780 139.670 81.580 140.000 ;
        RECT 80.430 138.870 80.685 139.340 ;
        RECT 80.345 138.700 80.685 138.870 ;
        RECT 80.430 138.670 80.685 138.700 ;
        RECT 80.865 138.360 81.150 139.160 ;
        RECT 81.330 139.080 81.580 139.670 ;
        RECT 81.780 140.315 82.100 140.645 ;
        RECT 82.280 140.430 82.940 140.910 ;
        RECT 83.140 140.520 83.990 140.690 ;
        RECT 81.780 139.420 81.970 140.315 ;
        RECT 82.290 139.990 82.950 140.260 ;
        RECT 82.620 139.930 82.950 139.990 ;
        RECT 82.140 139.760 82.470 139.820 ;
        RECT 83.140 139.760 83.310 140.520 ;
        RECT 84.550 140.450 84.870 140.910 ;
        RECT 85.070 140.270 85.320 140.700 ;
        RECT 85.610 140.470 86.020 140.910 ;
        RECT 86.190 140.530 87.205 140.730 ;
        RECT 83.480 140.100 84.730 140.270 ;
        RECT 83.480 139.980 83.810 140.100 ;
        RECT 82.140 139.590 84.040 139.760 ;
        RECT 81.780 139.250 83.700 139.420 ;
        RECT 81.780 139.230 82.100 139.250 ;
        RECT 81.330 138.570 81.660 139.080 ;
        RECT 81.930 138.620 82.100 139.230 ;
        RECT 83.870 139.080 84.040 139.590 ;
        RECT 84.210 139.520 84.390 139.930 ;
        RECT 84.560 139.340 84.730 140.100 ;
        RECT 82.270 138.360 82.600 139.050 ;
        RECT 82.830 138.910 84.040 139.080 ;
        RECT 84.210 139.030 84.730 139.340 ;
        RECT 84.900 139.930 85.320 140.270 ;
        RECT 85.610 139.930 86.020 140.260 ;
        RECT 84.900 139.160 85.090 139.930 ;
        RECT 86.190 139.800 86.360 140.530 ;
        RECT 87.505 140.360 87.675 140.690 ;
        RECT 87.845 140.530 88.175 140.910 ;
        RECT 86.530 139.980 86.880 140.350 ;
        RECT 86.190 139.760 86.610 139.800 ;
        RECT 85.260 139.590 86.610 139.760 ;
        RECT 85.260 139.430 85.510 139.590 ;
        RECT 86.020 139.160 86.270 139.420 ;
        RECT 84.900 138.910 86.270 139.160 ;
        RECT 82.830 138.620 83.070 138.910 ;
        RECT 83.870 138.830 84.040 138.910 ;
        RECT 83.270 138.360 83.690 138.740 ;
        RECT 83.870 138.580 84.500 138.830 ;
        RECT 84.970 138.360 85.300 138.740 ;
        RECT 85.470 138.620 85.640 138.910 ;
        RECT 86.440 138.745 86.610 139.590 ;
        RECT 87.060 139.420 87.280 140.290 ;
        RECT 87.505 140.170 88.200 140.360 ;
        RECT 86.780 139.040 87.280 139.420 ;
        RECT 87.450 139.370 87.860 139.990 ;
        RECT 88.030 139.200 88.200 140.170 ;
        RECT 87.505 139.030 88.200 139.200 ;
        RECT 85.820 138.360 86.200 138.740 ;
        RECT 86.440 138.575 87.270 138.745 ;
        RECT 87.505 138.530 87.675 139.030 ;
        RECT 87.845 138.360 88.175 138.860 ;
        RECT 88.390 138.530 88.615 140.650 ;
        RECT 88.785 140.530 89.115 140.910 ;
        RECT 89.285 140.360 89.455 140.650 ;
        RECT 90.090 140.570 90.345 140.730 ;
        RECT 90.005 140.400 90.345 140.570 ;
        RECT 90.525 140.450 90.810 140.910 ;
        RECT 88.790 140.190 89.455 140.360 ;
        RECT 90.090 140.200 90.345 140.400 ;
        RECT 88.790 139.200 89.020 140.190 ;
        RECT 89.190 139.370 89.540 140.020 ;
        RECT 90.090 139.340 90.270 140.200 ;
        RECT 90.990 140.000 91.240 140.650 ;
        RECT 90.440 139.670 91.240 140.000 ;
        RECT 88.790 139.030 89.455 139.200 ;
        RECT 88.785 138.360 89.115 138.860 ;
        RECT 89.285 138.530 89.455 139.030 ;
        RECT 90.090 138.670 90.345 139.340 ;
        RECT 90.525 138.360 90.810 139.160 ;
        RECT 90.990 139.080 91.240 139.670 ;
        RECT 91.440 140.315 91.760 140.645 ;
        RECT 91.940 140.430 92.600 140.910 ;
        RECT 92.800 140.520 93.650 140.690 ;
        RECT 91.440 139.420 91.630 140.315 ;
        RECT 91.950 139.990 92.610 140.260 ;
        RECT 92.280 139.930 92.610 139.990 ;
        RECT 91.800 139.760 92.130 139.820 ;
        RECT 92.800 139.760 92.970 140.520 ;
        RECT 94.210 140.450 94.530 140.910 ;
        RECT 94.730 140.270 94.980 140.700 ;
        RECT 95.270 140.470 95.680 140.910 ;
        RECT 95.850 140.530 96.865 140.730 ;
        RECT 93.140 140.100 94.390 140.270 ;
        RECT 93.140 139.980 93.470 140.100 ;
        RECT 91.800 139.590 93.700 139.760 ;
        RECT 91.440 139.250 93.360 139.420 ;
        RECT 91.440 139.230 91.760 139.250 ;
        RECT 90.990 138.570 91.320 139.080 ;
        RECT 91.590 138.620 91.760 139.230 ;
        RECT 93.530 139.080 93.700 139.590 ;
        RECT 93.870 139.520 94.050 139.930 ;
        RECT 94.220 139.340 94.390 140.100 ;
        RECT 91.930 138.360 92.260 139.050 ;
        RECT 92.490 138.910 93.700 139.080 ;
        RECT 93.870 139.030 94.390 139.340 ;
        RECT 94.560 139.930 94.980 140.270 ;
        RECT 95.270 139.930 95.680 140.260 ;
        RECT 94.560 139.160 94.750 139.930 ;
        RECT 95.850 139.800 96.020 140.530 ;
        RECT 97.165 140.360 97.335 140.690 ;
        RECT 97.505 140.530 97.835 140.910 ;
        RECT 96.190 139.980 96.540 140.350 ;
        RECT 95.850 139.760 96.270 139.800 ;
        RECT 94.920 139.590 96.270 139.760 ;
        RECT 94.920 139.430 95.170 139.590 ;
        RECT 95.680 139.160 95.930 139.420 ;
        RECT 94.560 138.910 95.930 139.160 ;
        RECT 92.490 138.620 92.730 138.910 ;
        RECT 93.530 138.830 93.700 138.910 ;
        RECT 92.930 138.360 93.350 138.740 ;
        RECT 93.530 138.580 94.160 138.830 ;
        RECT 94.630 138.360 94.960 138.740 ;
        RECT 95.130 138.620 95.300 138.910 ;
        RECT 96.100 138.745 96.270 139.590 ;
        RECT 96.720 139.420 96.940 140.290 ;
        RECT 97.165 140.170 97.860 140.360 ;
        RECT 96.440 139.040 96.940 139.420 ;
        RECT 97.110 139.370 97.520 139.990 ;
        RECT 97.690 139.200 97.860 140.170 ;
        RECT 97.165 139.030 97.860 139.200 ;
        RECT 95.480 138.360 95.860 138.740 ;
        RECT 96.100 138.575 96.930 138.745 ;
        RECT 97.165 138.530 97.335 139.030 ;
        RECT 97.505 138.360 97.835 138.860 ;
        RECT 98.050 138.530 98.275 140.650 ;
        RECT 98.445 140.530 98.775 140.910 ;
        RECT 98.945 140.360 99.115 140.650 ;
        RECT 98.450 140.190 99.115 140.360 ;
        RECT 99.375 140.235 99.645 140.580 ;
        RECT 99.835 140.510 100.215 140.910 ;
        RECT 100.385 140.340 100.555 140.690 ;
        RECT 100.725 140.510 101.055 140.910 ;
        RECT 101.255 140.340 101.425 140.690 ;
        RECT 101.625 140.410 101.955 140.910 ;
        RECT 98.450 139.200 98.680 140.190 ;
        RECT 98.850 139.370 99.200 140.020 ;
        RECT 99.375 139.500 99.545 140.235 ;
        RECT 99.815 140.170 101.425 140.340 ;
        RECT 99.815 140.000 99.985 140.170 ;
        RECT 99.715 139.670 99.985 140.000 ;
        RECT 100.155 139.670 100.560 140.000 ;
        RECT 99.815 139.500 99.985 139.670 ;
        RECT 100.730 139.550 101.440 140.000 ;
        RECT 101.610 139.670 101.960 140.240 ;
        RECT 102.595 140.185 102.885 140.910 ;
        RECT 103.430 140.200 103.685 140.730 ;
        RECT 103.865 140.450 104.150 140.910 ;
        RECT 98.450 139.030 99.115 139.200 ;
        RECT 98.445 138.360 98.775 138.860 ;
        RECT 98.945 138.530 99.115 139.030 ;
        RECT 99.375 138.530 99.645 139.500 ;
        RECT 99.815 139.330 100.540 139.500 ;
        RECT 100.730 139.380 101.445 139.550 ;
        RECT 100.370 139.210 100.540 139.330 ;
        RECT 101.640 139.210 101.960 139.500 ;
        RECT 99.855 138.360 100.135 139.160 ;
        RECT 100.370 139.040 101.960 139.210 ;
        RECT 100.305 138.580 101.960 138.870 ;
        RECT 102.595 138.360 102.885 139.525 ;
        RECT 103.430 139.340 103.610 140.200 ;
        RECT 104.330 140.000 104.580 140.650 ;
        RECT 103.780 139.670 104.580 140.000 ;
        RECT 103.430 138.870 103.685 139.340 ;
        RECT 103.345 138.700 103.685 138.870 ;
        RECT 103.430 138.670 103.685 138.700 ;
        RECT 103.865 138.360 104.150 139.160 ;
        RECT 104.330 139.080 104.580 139.670 ;
        RECT 104.780 140.315 105.100 140.645 ;
        RECT 105.280 140.430 105.940 140.910 ;
        RECT 106.140 140.520 106.990 140.690 ;
        RECT 104.780 139.420 104.970 140.315 ;
        RECT 105.290 139.990 105.950 140.260 ;
        RECT 105.620 139.930 105.950 139.990 ;
        RECT 105.140 139.760 105.470 139.820 ;
        RECT 106.140 139.760 106.310 140.520 ;
        RECT 107.550 140.450 107.870 140.910 ;
        RECT 108.070 140.270 108.320 140.700 ;
        RECT 108.610 140.470 109.020 140.910 ;
        RECT 109.190 140.530 110.205 140.730 ;
        RECT 106.480 140.100 107.730 140.270 ;
        RECT 106.480 139.980 106.810 140.100 ;
        RECT 105.140 139.590 107.040 139.760 ;
        RECT 104.780 139.250 106.700 139.420 ;
        RECT 104.780 139.230 105.100 139.250 ;
        RECT 104.330 138.570 104.660 139.080 ;
        RECT 104.930 138.620 105.100 139.230 ;
        RECT 106.870 139.080 107.040 139.590 ;
        RECT 107.210 139.520 107.390 139.930 ;
        RECT 107.560 139.340 107.730 140.100 ;
        RECT 105.270 138.360 105.600 139.050 ;
        RECT 105.830 138.910 107.040 139.080 ;
        RECT 107.210 139.030 107.730 139.340 ;
        RECT 107.900 139.930 108.320 140.270 ;
        RECT 108.610 139.930 109.020 140.260 ;
        RECT 107.900 139.160 108.090 139.930 ;
        RECT 109.190 139.800 109.360 140.530 ;
        RECT 110.505 140.360 110.675 140.690 ;
        RECT 110.845 140.530 111.175 140.910 ;
        RECT 109.530 139.980 109.880 140.350 ;
        RECT 109.190 139.760 109.610 139.800 ;
        RECT 108.260 139.590 109.610 139.760 ;
        RECT 108.260 139.430 108.510 139.590 ;
        RECT 109.020 139.160 109.270 139.420 ;
        RECT 107.900 138.910 109.270 139.160 ;
        RECT 105.830 138.620 106.070 138.910 ;
        RECT 106.870 138.830 107.040 138.910 ;
        RECT 106.270 138.360 106.690 138.740 ;
        RECT 106.870 138.580 107.500 138.830 ;
        RECT 107.970 138.360 108.300 138.740 ;
        RECT 108.470 138.620 108.640 138.910 ;
        RECT 109.440 138.745 109.610 139.590 ;
        RECT 110.060 139.420 110.280 140.290 ;
        RECT 110.505 140.170 111.200 140.360 ;
        RECT 109.780 139.040 110.280 139.420 ;
        RECT 110.450 139.370 110.860 139.990 ;
        RECT 111.030 139.200 111.200 140.170 ;
        RECT 110.505 139.030 111.200 139.200 ;
        RECT 108.820 138.360 109.200 138.740 ;
        RECT 109.440 138.575 110.270 138.745 ;
        RECT 110.505 138.530 110.675 139.030 ;
        RECT 110.845 138.360 111.175 138.860 ;
        RECT 111.390 138.530 111.615 140.650 ;
        RECT 111.785 140.530 112.115 140.910 ;
        RECT 112.285 140.360 112.455 140.650 ;
        RECT 111.790 140.190 112.455 140.360 ;
        RECT 112.715 140.235 112.975 140.740 ;
        RECT 113.155 140.530 113.485 140.910 ;
        RECT 113.665 140.360 113.835 140.740 ;
        RECT 111.790 139.200 112.020 140.190 ;
        RECT 112.190 139.370 112.540 140.020 ;
        RECT 112.715 139.435 112.885 140.235 ;
        RECT 113.170 140.190 113.835 140.360 ;
        RECT 113.170 139.935 113.340 140.190 ;
        RECT 114.555 140.160 115.765 140.910 ;
        RECT 113.055 139.605 113.340 139.935 ;
        RECT 113.575 139.640 113.905 140.010 ;
        RECT 113.170 139.460 113.340 139.605 ;
        RECT 111.790 139.030 112.455 139.200 ;
        RECT 111.785 138.360 112.115 138.860 ;
        RECT 112.285 138.530 112.455 139.030 ;
        RECT 112.715 138.530 112.985 139.435 ;
        RECT 113.170 139.290 113.835 139.460 ;
        RECT 113.155 138.360 113.485 139.120 ;
        RECT 113.665 138.530 113.835 139.290 ;
        RECT 114.555 139.450 115.075 139.990 ;
        RECT 115.245 139.620 115.765 140.160 ;
        RECT 114.555 138.360 115.765 139.450 ;
        RECT 14.650 138.190 115.850 138.360 ;
        RECT 14.735 137.100 15.945 138.190 ;
        RECT 14.735 136.390 15.255 136.930 ;
        RECT 15.425 136.560 15.945 137.100 ;
        RECT 16.115 137.100 17.325 138.190 ;
        RECT 16.115 136.560 16.635 137.100 ;
        RECT 17.535 137.050 17.765 138.190 ;
        RECT 17.935 137.040 18.265 138.020 ;
        RECT 18.435 137.050 18.645 138.190 ;
        RECT 19.250 137.210 19.505 137.880 ;
        RECT 19.685 137.390 19.970 138.190 ;
        RECT 20.150 137.470 20.480 137.980 ;
        RECT 16.805 136.390 17.325 136.930 ;
        RECT 17.515 136.630 17.845 136.880 ;
        RECT 14.735 135.640 15.945 136.390 ;
        RECT 16.115 135.640 17.325 136.390 ;
        RECT 17.535 135.640 17.765 136.460 ;
        RECT 18.015 136.440 18.265 137.040 ;
        RECT 17.935 135.810 18.265 136.440 ;
        RECT 18.435 135.640 18.645 136.460 ;
        RECT 19.250 136.350 19.430 137.210 ;
        RECT 20.150 136.880 20.400 137.470 ;
        RECT 20.750 137.320 20.920 137.930 ;
        RECT 21.090 137.500 21.420 138.190 ;
        RECT 21.650 137.640 21.890 137.930 ;
        RECT 22.090 137.810 22.510 138.190 ;
        RECT 22.690 137.720 23.320 137.970 ;
        RECT 23.790 137.810 24.120 138.190 ;
        RECT 22.690 137.640 22.860 137.720 ;
        RECT 24.290 137.640 24.460 137.930 ;
        RECT 24.640 137.810 25.020 138.190 ;
        RECT 25.260 137.805 26.090 137.975 ;
        RECT 21.650 137.470 22.860 137.640 ;
        RECT 19.600 136.550 20.400 136.880 ;
        RECT 19.250 136.150 19.505 136.350 ;
        RECT 19.165 135.980 19.505 136.150 ;
        RECT 19.250 135.820 19.505 135.980 ;
        RECT 19.685 135.640 19.970 136.100 ;
        RECT 20.150 135.900 20.400 136.550 ;
        RECT 20.600 137.300 20.920 137.320 ;
        RECT 20.600 137.130 22.520 137.300 ;
        RECT 20.600 136.235 20.790 137.130 ;
        RECT 22.690 136.960 22.860 137.470 ;
        RECT 23.030 137.210 23.550 137.520 ;
        RECT 20.960 136.790 22.860 136.960 ;
        RECT 20.960 136.730 21.290 136.790 ;
        RECT 21.440 136.560 21.770 136.620 ;
        RECT 21.110 136.290 21.770 136.560 ;
        RECT 20.600 135.905 20.920 136.235 ;
        RECT 21.100 135.640 21.760 136.120 ;
        RECT 21.960 136.030 22.130 136.790 ;
        RECT 23.030 136.620 23.210 137.030 ;
        RECT 22.300 136.450 22.630 136.570 ;
        RECT 23.380 136.450 23.550 137.210 ;
        RECT 22.300 136.280 23.550 136.450 ;
        RECT 23.720 137.390 25.090 137.640 ;
        RECT 23.720 136.620 23.910 137.390 ;
        RECT 24.840 137.130 25.090 137.390 ;
        RECT 24.080 136.960 24.330 137.120 ;
        RECT 25.260 136.960 25.430 137.805 ;
        RECT 26.325 137.520 26.495 138.020 ;
        RECT 26.665 137.690 26.995 138.190 ;
        RECT 25.600 137.130 26.100 137.510 ;
        RECT 26.325 137.350 27.020 137.520 ;
        RECT 24.080 136.790 25.430 136.960 ;
        RECT 25.010 136.750 25.430 136.790 ;
        RECT 23.720 136.280 24.140 136.620 ;
        RECT 24.430 136.290 24.840 136.620 ;
        RECT 21.960 135.860 22.810 136.030 ;
        RECT 23.370 135.640 23.690 136.100 ;
        RECT 23.890 135.850 24.140 136.280 ;
        RECT 24.430 135.640 24.840 136.080 ;
        RECT 25.010 136.020 25.180 136.750 ;
        RECT 25.350 136.200 25.700 136.570 ;
        RECT 25.880 136.260 26.100 137.130 ;
        RECT 26.270 136.560 26.680 137.180 ;
        RECT 26.850 136.380 27.020 137.350 ;
        RECT 26.325 136.190 27.020 136.380 ;
        RECT 25.010 135.820 26.025 136.020 ;
        RECT 26.325 135.860 26.495 136.190 ;
        RECT 26.665 135.640 26.995 136.020 ;
        RECT 27.210 135.900 27.435 138.020 ;
        RECT 27.605 137.690 27.935 138.190 ;
        RECT 28.105 137.520 28.275 138.020 ;
        RECT 28.735 137.520 29.015 138.190 ;
        RECT 27.610 137.350 28.275 137.520 ;
        RECT 27.610 136.360 27.840 137.350 ;
        RECT 29.185 137.300 29.485 137.850 ;
        RECT 29.685 137.470 30.015 138.190 ;
        RECT 30.205 137.470 30.665 138.020 ;
        RECT 31.035 137.520 31.315 138.190 ;
        RECT 28.010 136.530 28.360 137.180 ;
        RECT 28.550 136.880 28.815 137.240 ;
        RECT 29.185 137.130 30.125 137.300 ;
        RECT 29.955 136.880 30.125 137.130 ;
        RECT 28.550 136.630 29.225 136.880 ;
        RECT 29.445 136.630 29.785 136.880 ;
        RECT 29.955 136.550 30.245 136.880 ;
        RECT 29.955 136.460 30.125 136.550 ;
        RECT 27.610 136.190 28.275 136.360 ;
        RECT 27.605 135.640 27.935 136.020 ;
        RECT 28.105 135.900 28.275 136.190 ;
        RECT 28.735 136.270 30.125 136.460 ;
        RECT 28.735 135.910 29.065 136.270 ;
        RECT 30.415 136.100 30.665 137.470 ;
        RECT 31.485 137.300 31.785 137.850 ;
        RECT 31.985 137.470 32.315 138.190 ;
        RECT 32.505 137.470 32.965 138.020 ;
        RECT 33.335 137.520 33.615 138.190 ;
        RECT 30.850 136.880 31.115 137.240 ;
        RECT 31.485 137.130 32.425 137.300 ;
        RECT 32.255 136.880 32.425 137.130 ;
        RECT 30.850 136.630 31.525 136.880 ;
        RECT 31.745 136.630 32.085 136.880 ;
        RECT 32.255 136.550 32.545 136.880 ;
        RECT 32.255 136.460 32.425 136.550 ;
        RECT 29.685 135.640 29.935 136.100 ;
        RECT 30.105 135.810 30.665 136.100 ;
        RECT 31.035 136.270 32.425 136.460 ;
        RECT 31.035 135.910 31.365 136.270 ;
        RECT 32.715 136.100 32.965 137.470 ;
        RECT 33.785 137.300 34.085 137.850 ;
        RECT 34.285 137.470 34.615 138.190 ;
        RECT 34.805 137.470 35.265 138.020 ;
        RECT 36.095 137.520 36.375 138.190 ;
        RECT 33.150 136.880 33.415 137.240 ;
        RECT 33.785 137.130 34.725 137.300 ;
        RECT 34.555 136.880 34.725 137.130 ;
        RECT 33.150 136.630 33.825 136.880 ;
        RECT 34.045 136.630 34.385 136.880 ;
        RECT 34.555 136.550 34.845 136.880 ;
        RECT 34.555 136.460 34.725 136.550 ;
        RECT 31.985 135.640 32.235 136.100 ;
        RECT 32.405 135.810 32.965 136.100 ;
        RECT 33.335 136.270 34.725 136.460 ;
        RECT 33.335 135.910 33.665 136.270 ;
        RECT 35.015 136.100 35.265 137.470 ;
        RECT 36.545 137.300 36.845 137.850 ;
        RECT 37.045 137.470 37.375 138.190 ;
        RECT 37.565 137.470 38.025 138.020 ;
        RECT 35.910 136.880 36.175 137.240 ;
        RECT 36.545 137.130 37.485 137.300 ;
        RECT 37.315 136.880 37.485 137.130 ;
        RECT 35.910 136.630 36.585 136.880 ;
        RECT 36.805 136.630 37.145 136.880 ;
        RECT 37.315 136.550 37.605 136.880 ;
        RECT 37.315 136.460 37.485 136.550 ;
        RECT 34.285 135.640 34.535 136.100 ;
        RECT 34.705 135.810 35.265 136.100 ;
        RECT 36.095 136.270 37.485 136.460 ;
        RECT 36.095 135.910 36.425 136.270 ;
        RECT 37.775 136.100 38.025 137.470 ;
        RECT 38.195 137.025 38.485 138.190 ;
        RECT 38.655 137.050 38.925 138.020 ;
        RECT 39.135 137.390 39.415 138.190 ;
        RECT 39.585 137.680 41.240 137.970 ;
        RECT 41.420 137.755 46.765 138.190 ;
        RECT 39.650 137.340 41.240 137.510 ;
        RECT 39.650 137.220 39.820 137.340 ;
        RECT 39.095 137.050 39.820 137.220 ;
        RECT 37.045 135.640 37.295 136.100 ;
        RECT 37.465 135.810 38.025 136.100 ;
        RECT 38.195 135.640 38.485 136.365 ;
        RECT 38.655 136.315 38.825 137.050 ;
        RECT 39.095 136.880 39.265 137.050 ;
        RECT 38.995 136.550 39.265 136.880 ;
        RECT 39.435 136.550 39.840 136.880 ;
        RECT 40.010 136.550 40.720 137.170 ;
        RECT 40.920 137.050 41.240 137.340 ;
        RECT 39.095 136.380 39.265 136.550 ;
        RECT 38.655 135.970 38.925 136.315 ;
        RECT 39.095 136.210 40.705 136.380 ;
        RECT 40.890 136.310 41.240 136.880 ;
        RECT 43.010 136.505 43.360 137.755 ;
        RECT 46.935 137.050 47.275 138.020 ;
        RECT 47.445 137.050 47.615 138.190 ;
        RECT 47.885 137.390 48.135 138.190 ;
        RECT 48.780 137.220 49.110 138.020 ;
        RECT 49.410 137.390 49.740 138.190 ;
        RECT 49.910 137.220 50.240 138.020 ;
        RECT 47.805 137.050 50.240 137.220 ;
        RECT 51.575 137.050 51.805 138.190 ;
        RECT 39.115 135.640 39.495 136.040 ;
        RECT 39.665 135.860 39.835 136.210 ;
        RECT 40.005 135.640 40.335 136.040 ;
        RECT 40.535 135.860 40.705 136.210 ;
        RECT 44.840 136.185 45.180 137.015 ;
        RECT 46.935 136.490 47.110 137.050 ;
        RECT 47.805 136.800 47.975 137.050 ;
        RECT 47.280 136.630 47.975 136.800 ;
        RECT 48.150 136.630 48.570 136.830 ;
        RECT 48.740 136.630 49.070 136.830 ;
        RECT 49.240 136.630 49.570 136.830 ;
        RECT 46.935 136.440 47.165 136.490 ;
        RECT 40.905 135.640 41.235 136.140 ;
        RECT 41.420 135.640 46.765 136.185 ;
        RECT 46.935 135.810 47.275 136.440 ;
        RECT 47.445 135.640 47.695 136.440 ;
        RECT 47.885 136.290 49.110 136.460 ;
        RECT 47.885 135.810 48.215 136.290 ;
        RECT 48.385 135.640 48.610 136.100 ;
        RECT 48.780 135.810 49.110 136.290 ;
        RECT 49.740 136.420 49.910 137.050 ;
        RECT 51.975 137.040 52.305 138.020 ;
        RECT 52.475 137.050 52.685 138.190 ;
        RECT 53.375 137.100 56.885 138.190 ;
        RECT 57.060 137.755 62.405 138.190 ;
        RECT 50.095 136.630 50.445 136.880 ;
        RECT 51.555 136.630 51.885 136.880 ;
        RECT 49.740 135.810 50.240 136.420 ;
        RECT 51.575 135.640 51.805 136.460 ;
        RECT 52.055 136.440 52.305 137.040 ;
        RECT 53.375 136.580 55.065 137.100 ;
        RECT 51.975 135.810 52.305 136.440 ;
        RECT 52.475 135.640 52.685 136.460 ;
        RECT 55.235 136.410 56.885 136.930 ;
        RECT 58.650 136.505 59.000 137.755 ;
        RECT 62.635 137.050 62.845 138.190 ;
        RECT 63.015 137.040 63.345 138.020 ;
        RECT 63.515 137.050 63.745 138.190 ;
        RECT 53.375 135.640 56.885 136.410 ;
        RECT 60.480 136.185 60.820 137.015 ;
        RECT 57.060 135.640 62.405 136.185 ;
        RECT 62.635 135.640 62.845 136.460 ;
        RECT 63.015 136.440 63.265 137.040 ;
        RECT 63.955 137.025 64.245 138.190 ;
        RECT 64.415 137.100 65.625 138.190 ;
        RECT 65.800 137.765 66.135 138.190 ;
        RECT 66.305 137.585 66.490 137.990 ;
        RECT 65.825 137.410 66.490 137.585 ;
        RECT 66.695 137.410 67.025 138.190 ;
        RECT 63.435 136.630 63.765 136.880 ;
        RECT 64.415 136.560 64.935 137.100 ;
        RECT 63.015 135.810 63.345 136.440 ;
        RECT 63.515 135.640 63.745 136.460 ;
        RECT 65.105 136.390 65.625 136.930 ;
        RECT 63.955 135.640 64.245 136.365 ;
        RECT 64.415 135.640 65.625 136.390 ;
        RECT 65.825 136.380 66.165 137.410 ;
        RECT 67.195 137.220 67.465 137.990 ;
        RECT 66.335 137.050 67.465 137.220 ;
        RECT 66.335 136.550 66.585 137.050 ;
        RECT 65.825 136.210 66.510 136.380 ;
        RECT 66.765 136.300 67.125 136.880 ;
        RECT 65.800 135.640 66.135 136.040 ;
        RECT 66.305 135.810 66.510 136.210 ;
        RECT 67.295 136.140 67.465 137.050 ;
        RECT 66.720 135.640 66.995 136.120 ;
        RECT 67.205 135.810 67.465 136.140 ;
        RECT 68.555 137.050 68.825 138.020 ;
        RECT 69.035 137.390 69.315 138.190 ;
        RECT 69.485 137.680 71.140 137.970 ;
        RECT 69.550 137.340 71.140 137.510 ;
        RECT 69.550 137.220 69.720 137.340 ;
        RECT 68.995 137.050 69.720 137.220 ;
        RECT 68.555 136.315 68.725 137.050 ;
        RECT 68.995 136.880 69.165 137.050 ;
        RECT 69.910 137.000 70.625 137.170 ;
        RECT 70.820 137.050 71.140 137.340 ;
        RECT 71.315 137.050 71.655 138.020 ;
        RECT 71.825 137.050 71.995 138.190 ;
        RECT 72.265 137.390 72.515 138.190 ;
        RECT 73.160 137.220 73.490 138.020 ;
        RECT 73.790 137.390 74.120 138.190 ;
        RECT 74.290 137.220 74.620 138.020 ;
        RECT 72.185 137.050 74.620 137.220 ;
        RECT 75.370 137.210 75.625 137.880 ;
        RECT 75.805 137.390 76.090 138.190 ;
        RECT 76.270 137.470 76.600 137.980 ;
        RECT 68.895 136.550 69.165 136.880 ;
        RECT 69.335 136.550 69.740 136.880 ;
        RECT 69.910 136.550 70.620 137.000 ;
        RECT 68.995 136.380 69.165 136.550 ;
        RECT 68.555 135.970 68.825 136.315 ;
        RECT 68.995 136.210 70.605 136.380 ;
        RECT 70.790 136.310 71.140 136.880 ;
        RECT 71.315 136.490 71.490 137.050 ;
        RECT 72.185 136.800 72.355 137.050 ;
        RECT 71.660 136.630 72.355 136.800 ;
        RECT 72.530 136.630 72.950 136.830 ;
        RECT 73.120 136.630 73.450 136.830 ;
        RECT 73.620 136.630 73.950 136.830 ;
        RECT 71.315 136.440 71.545 136.490 ;
        RECT 69.015 135.640 69.395 136.040 ;
        RECT 69.565 135.860 69.735 136.210 ;
        RECT 69.905 135.640 70.235 136.040 ;
        RECT 70.435 135.860 70.605 136.210 ;
        RECT 70.805 135.640 71.135 136.140 ;
        RECT 71.315 135.810 71.655 136.440 ;
        RECT 71.825 135.640 72.075 136.440 ;
        RECT 72.265 136.290 73.490 136.460 ;
        RECT 72.265 135.810 72.595 136.290 ;
        RECT 72.765 135.640 72.990 136.100 ;
        RECT 73.160 135.810 73.490 136.290 ;
        RECT 74.120 136.420 74.290 137.050 ;
        RECT 74.475 136.630 74.825 136.880 ;
        RECT 74.120 135.810 74.620 136.420 ;
        RECT 75.370 136.350 75.550 137.210 ;
        RECT 76.270 136.880 76.520 137.470 ;
        RECT 76.870 137.320 77.040 137.930 ;
        RECT 77.210 137.500 77.540 138.190 ;
        RECT 77.770 137.640 78.010 137.930 ;
        RECT 78.210 137.810 78.630 138.190 ;
        RECT 78.810 137.720 79.440 137.970 ;
        RECT 79.910 137.810 80.240 138.190 ;
        RECT 78.810 137.640 78.980 137.720 ;
        RECT 80.410 137.640 80.580 137.930 ;
        RECT 80.760 137.810 81.140 138.190 ;
        RECT 81.380 137.805 82.210 137.975 ;
        RECT 77.770 137.470 78.980 137.640 ;
        RECT 75.720 136.550 76.520 136.880 ;
        RECT 75.370 136.150 75.625 136.350 ;
        RECT 75.285 135.980 75.625 136.150 ;
        RECT 75.370 135.820 75.625 135.980 ;
        RECT 75.805 135.640 76.090 136.100 ;
        RECT 76.270 135.900 76.520 136.550 ;
        RECT 76.720 137.300 77.040 137.320 ;
        RECT 76.720 137.130 78.640 137.300 ;
        RECT 76.720 136.235 76.910 137.130 ;
        RECT 78.810 136.960 78.980 137.470 ;
        RECT 79.150 137.210 79.670 137.520 ;
        RECT 77.080 136.790 78.980 136.960 ;
        RECT 77.080 136.730 77.410 136.790 ;
        RECT 77.560 136.560 77.890 136.620 ;
        RECT 77.230 136.290 77.890 136.560 ;
        RECT 76.720 135.905 77.040 136.235 ;
        RECT 77.220 135.640 77.880 136.120 ;
        RECT 78.080 136.030 78.250 136.790 ;
        RECT 79.150 136.620 79.330 137.030 ;
        RECT 78.420 136.450 78.750 136.570 ;
        RECT 79.500 136.450 79.670 137.210 ;
        RECT 78.420 136.280 79.670 136.450 ;
        RECT 79.840 137.390 81.210 137.640 ;
        RECT 79.840 136.620 80.030 137.390 ;
        RECT 80.960 137.130 81.210 137.390 ;
        RECT 80.200 136.960 80.450 137.120 ;
        RECT 81.380 136.960 81.550 137.805 ;
        RECT 82.445 137.520 82.615 138.020 ;
        RECT 82.785 137.690 83.115 138.190 ;
        RECT 81.720 137.130 82.220 137.510 ;
        RECT 82.445 137.350 83.140 137.520 ;
        RECT 80.200 136.790 81.550 136.960 ;
        RECT 81.130 136.750 81.550 136.790 ;
        RECT 79.840 136.280 80.260 136.620 ;
        RECT 80.550 136.290 80.960 136.620 ;
        RECT 78.080 135.860 78.930 136.030 ;
        RECT 79.490 135.640 79.810 136.100 ;
        RECT 80.010 135.850 80.260 136.280 ;
        RECT 80.550 135.640 80.960 136.080 ;
        RECT 81.130 136.020 81.300 136.750 ;
        RECT 81.470 136.200 81.820 136.570 ;
        RECT 82.000 136.260 82.220 137.130 ;
        RECT 82.390 136.560 82.800 137.180 ;
        RECT 82.970 136.380 83.140 137.350 ;
        RECT 82.445 136.190 83.140 136.380 ;
        RECT 81.130 135.820 82.145 136.020 ;
        RECT 82.445 135.860 82.615 136.190 ;
        RECT 82.785 135.640 83.115 136.020 ;
        RECT 83.330 135.900 83.555 138.020 ;
        RECT 83.725 137.690 84.055 138.190 ;
        RECT 84.225 137.520 84.395 138.020 ;
        RECT 83.730 137.350 84.395 137.520 ;
        RECT 84.655 137.430 85.170 137.840 ;
        RECT 85.405 137.430 85.575 138.190 ;
        RECT 85.745 137.850 87.775 138.020 ;
        RECT 83.730 136.360 83.960 137.350 ;
        RECT 84.130 136.530 84.480 137.180 ;
        RECT 84.655 136.620 84.995 137.430 ;
        RECT 85.745 137.185 85.915 137.850 ;
        RECT 86.310 137.510 87.435 137.680 ;
        RECT 85.165 136.995 85.915 137.185 ;
        RECT 86.085 137.170 87.095 137.340 ;
        RECT 84.655 136.450 85.885 136.620 ;
        RECT 83.730 136.190 84.395 136.360 ;
        RECT 83.725 135.640 84.055 136.020 ;
        RECT 84.225 135.900 84.395 136.190 ;
        RECT 84.930 135.845 85.175 136.450 ;
        RECT 85.395 135.640 85.905 136.175 ;
        RECT 86.085 135.810 86.275 137.170 ;
        RECT 86.445 136.490 86.720 136.970 ;
        RECT 86.445 136.320 86.725 136.490 ;
        RECT 86.925 136.370 87.095 137.170 ;
        RECT 87.265 136.380 87.435 137.510 ;
        RECT 87.605 136.880 87.775 137.850 ;
        RECT 87.945 137.050 88.115 138.190 ;
        RECT 88.285 137.050 88.620 138.020 ;
        RECT 87.605 136.550 87.800 136.880 ;
        RECT 88.025 136.550 88.280 136.880 ;
        RECT 88.025 136.380 88.195 136.550 ;
        RECT 88.450 136.380 88.620 137.050 ;
        RECT 89.715 137.025 90.005 138.190 ;
        RECT 90.175 137.100 91.385 138.190 ;
        RECT 90.175 136.560 90.695 137.100 ;
        RECT 91.595 137.050 91.825 138.190 ;
        RECT 91.995 137.040 92.325 138.020 ;
        RECT 92.495 137.050 92.705 138.190 ;
        RECT 92.935 137.100 94.145 138.190 ;
        RECT 94.405 137.260 94.575 138.020 ;
        RECT 94.755 137.430 95.085 138.190 ;
        RECT 90.865 136.390 91.385 136.930 ;
        RECT 91.575 136.630 91.905 136.880 ;
        RECT 86.445 135.810 86.720 136.320 ;
        RECT 87.265 136.210 88.195 136.380 ;
        RECT 87.265 136.175 87.440 136.210 ;
        RECT 86.910 135.810 87.440 136.175 ;
        RECT 87.865 135.640 88.195 136.040 ;
        RECT 88.365 135.810 88.620 136.380 ;
        RECT 89.715 135.640 90.005 136.365 ;
        RECT 90.175 135.640 91.385 136.390 ;
        RECT 91.595 135.640 91.825 136.460 ;
        RECT 92.075 136.440 92.325 137.040 ;
        RECT 92.935 136.560 93.455 137.100 ;
        RECT 94.405 137.090 95.070 137.260 ;
        RECT 95.255 137.115 95.525 138.020 ;
        RECT 94.900 136.945 95.070 137.090 ;
        RECT 91.995 135.810 92.325 136.440 ;
        RECT 92.495 135.640 92.705 136.460 ;
        RECT 93.625 136.390 94.145 136.930 ;
        RECT 94.335 136.540 94.665 136.910 ;
        RECT 94.900 136.615 95.185 136.945 ;
        RECT 92.935 135.640 94.145 136.390 ;
        RECT 94.900 136.360 95.070 136.615 ;
        RECT 94.405 136.190 95.070 136.360 ;
        RECT 95.355 136.315 95.525 137.115 ;
        RECT 94.405 135.810 94.575 136.190 ;
        RECT 94.755 135.640 95.085 136.020 ;
        RECT 95.265 135.810 95.525 136.315 ;
        RECT 95.695 137.470 96.155 138.020 ;
        RECT 96.345 137.470 96.675 138.190 ;
        RECT 95.695 136.100 95.945 137.470 ;
        RECT 96.875 137.300 97.175 137.850 ;
        RECT 97.345 137.520 97.625 138.190 ;
        RECT 96.235 137.130 97.175 137.300 ;
        RECT 96.235 136.880 96.405 137.130 ;
        RECT 97.545 136.880 97.810 137.240 ;
        RECT 96.115 136.550 96.405 136.880 ;
        RECT 96.575 136.630 96.915 136.880 ;
        RECT 97.135 136.630 97.810 136.880 ;
        RECT 97.995 137.100 99.205 138.190 ;
        RECT 99.375 137.100 102.885 138.190 ;
        RECT 103.055 137.430 103.570 137.840 ;
        RECT 103.805 137.430 103.975 138.190 ;
        RECT 104.145 137.850 106.175 138.020 ;
        RECT 97.995 136.560 98.515 137.100 ;
        RECT 96.235 136.460 96.405 136.550 ;
        RECT 96.235 136.270 97.625 136.460 ;
        RECT 98.685 136.390 99.205 136.930 ;
        RECT 99.375 136.580 101.065 137.100 ;
        RECT 101.235 136.410 102.885 136.930 ;
        RECT 103.055 136.620 103.395 137.430 ;
        RECT 104.145 137.185 104.315 137.850 ;
        RECT 104.710 137.510 105.835 137.680 ;
        RECT 103.565 136.995 104.315 137.185 ;
        RECT 104.485 137.170 105.495 137.340 ;
        RECT 103.055 136.450 104.285 136.620 ;
        RECT 95.695 135.810 96.255 136.100 ;
        RECT 96.425 135.640 96.675 136.100 ;
        RECT 97.295 135.910 97.625 136.270 ;
        RECT 97.995 135.640 99.205 136.390 ;
        RECT 99.375 135.640 102.885 136.410 ;
        RECT 103.330 135.845 103.575 136.450 ;
        RECT 103.795 135.640 104.305 136.175 ;
        RECT 104.485 135.810 104.675 137.170 ;
        RECT 104.845 136.830 105.120 136.970 ;
        RECT 104.845 136.660 105.125 136.830 ;
        RECT 104.845 135.810 105.120 136.660 ;
        RECT 105.325 136.370 105.495 137.170 ;
        RECT 105.665 136.380 105.835 137.510 ;
        RECT 106.005 136.880 106.175 137.850 ;
        RECT 106.345 137.050 106.515 138.190 ;
        RECT 106.685 137.050 107.020 138.020 ;
        RECT 107.745 137.260 107.915 138.020 ;
        RECT 108.095 137.430 108.425 138.190 ;
        RECT 107.745 137.090 108.410 137.260 ;
        RECT 108.595 137.115 108.865 138.020 ;
        RECT 109.040 137.755 114.385 138.190 ;
        RECT 106.005 136.550 106.200 136.880 ;
        RECT 106.425 136.550 106.680 136.880 ;
        RECT 106.425 136.380 106.595 136.550 ;
        RECT 106.850 136.380 107.020 137.050 ;
        RECT 108.240 136.945 108.410 137.090 ;
        RECT 107.675 136.540 108.005 136.910 ;
        RECT 108.240 136.615 108.525 136.945 ;
        RECT 105.665 136.210 106.595 136.380 ;
        RECT 105.665 136.175 105.840 136.210 ;
        RECT 105.310 135.810 105.840 136.175 ;
        RECT 106.265 135.640 106.595 136.040 ;
        RECT 106.765 135.810 107.020 136.380 ;
        RECT 108.240 136.360 108.410 136.615 ;
        RECT 107.745 136.190 108.410 136.360 ;
        RECT 108.695 136.315 108.865 137.115 ;
        RECT 110.630 136.505 110.980 137.755 ;
        RECT 114.555 137.100 115.765 138.190 ;
        RECT 107.745 135.810 107.915 136.190 ;
        RECT 108.095 135.640 108.425 136.020 ;
        RECT 108.605 135.810 108.865 136.315 ;
        RECT 112.460 136.185 112.800 137.015 ;
        RECT 114.555 136.560 115.075 137.100 ;
        RECT 115.245 136.390 115.765 136.930 ;
        RECT 109.040 135.640 114.385 136.185 ;
        RECT 114.555 135.640 115.765 136.390 ;
        RECT 14.650 135.470 115.850 135.640 ;
        RECT 14.735 134.720 15.945 135.470 ;
        RECT 14.735 134.180 15.255 134.720 ;
        RECT 16.575 134.700 20.085 135.470 ;
        RECT 15.425 134.010 15.945 134.550 ;
        RECT 14.735 132.920 15.945 134.010 ;
        RECT 16.575 134.010 18.265 134.530 ;
        RECT 18.435 134.180 20.085 134.700 ;
        RECT 20.530 134.660 20.775 135.265 ;
        RECT 20.995 134.935 21.505 135.470 ;
        RECT 20.255 134.490 21.485 134.660 ;
        RECT 16.575 132.920 20.085 134.010 ;
        RECT 20.255 133.680 20.595 134.490 ;
        RECT 20.765 133.925 21.515 134.115 ;
        RECT 20.255 133.270 20.770 133.680 ;
        RECT 21.005 132.920 21.175 133.680 ;
        RECT 21.345 133.260 21.515 133.925 ;
        RECT 21.685 133.940 21.875 135.300 ;
        RECT 22.045 135.130 22.320 135.300 ;
        RECT 22.045 134.960 22.325 135.130 ;
        RECT 22.045 134.140 22.320 134.960 ;
        RECT 22.510 134.935 23.040 135.300 ;
        RECT 23.465 135.070 23.795 135.470 ;
        RECT 22.865 134.900 23.040 134.935 ;
        RECT 22.525 133.940 22.695 134.740 ;
        RECT 21.685 133.770 22.695 133.940 ;
        RECT 22.865 134.730 23.795 134.900 ;
        RECT 23.965 134.730 24.220 135.300 ;
        RECT 25.315 134.745 25.605 135.470 ;
        RECT 22.865 133.600 23.035 134.730 ;
        RECT 23.625 134.560 23.795 134.730 ;
        RECT 21.910 133.430 23.035 133.600 ;
        RECT 23.205 134.230 23.400 134.560 ;
        RECT 23.625 134.230 23.880 134.560 ;
        RECT 23.205 133.260 23.375 134.230 ;
        RECT 24.050 134.060 24.220 134.730 ;
        RECT 26.240 134.730 26.495 135.300 ;
        RECT 26.665 135.070 26.995 135.470 ;
        RECT 27.420 134.935 27.950 135.300 ;
        RECT 28.140 135.130 28.415 135.300 ;
        RECT 28.135 134.960 28.415 135.130 ;
        RECT 27.420 134.900 27.595 134.935 ;
        RECT 26.665 134.730 27.595 134.900 ;
        RECT 21.345 133.090 23.375 133.260 ;
        RECT 23.545 132.920 23.715 134.060 ;
        RECT 23.885 133.090 24.220 134.060 ;
        RECT 25.315 132.920 25.605 134.085 ;
        RECT 26.240 134.060 26.410 134.730 ;
        RECT 26.665 134.560 26.835 134.730 ;
        RECT 26.580 134.230 26.835 134.560 ;
        RECT 27.060 134.230 27.255 134.560 ;
        RECT 26.240 133.090 26.575 134.060 ;
        RECT 26.745 132.920 26.915 134.060 ;
        RECT 27.085 133.260 27.255 134.230 ;
        RECT 27.425 133.600 27.595 134.730 ;
        RECT 27.765 133.940 27.935 134.740 ;
        RECT 28.140 134.140 28.415 134.960 ;
        RECT 28.585 133.940 28.775 135.300 ;
        RECT 28.955 134.935 29.465 135.470 ;
        RECT 29.685 134.660 29.930 135.265 ;
        RECT 28.975 134.490 30.205 134.660 ;
        RECT 30.415 134.650 30.645 135.470 ;
        RECT 30.815 134.670 31.145 135.300 ;
        RECT 27.765 133.770 28.775 133.940 ;
        RECT 28.945 133.925 29.695 134.115 ;
        RECT 27.425 133.430 28.550 133.600 ;
        RECT 28.945 133.260 29.115 133.925 ;
        RECT 29.865 133.680 30.205 134.490 ;
        RECT 30.395 134.230 30.725 134.480 ;
        RECT 30.895 134.070 31.145 134.670 ;
        RECT 31.315 134.650 31.525 135.470 ;
        RECT 32.030 134.660 32.275 135.265 ;
        RECT 32.495 134.935 33.005 135.470 ;
        RECT 27.085 133.090 29.115 133.260 ;
        RECT 29.285 132.920 29.455 133.680 ;
        RECT 29.690 133.270 30.205 133.680 ;
        RECT 30.415 132.920 30.645 134.060 ;
        RECT 30.815 133.090 31.145 134.070 ;
        RECT 31.755 134.490 32.985 134.660 ;
        RECT 31.315 132.920 31.525 134.060 ;
        RECT 31.755 133.680 32.095 134.490 ;
        RECT 32.265 133.925 33.015 134.115 ;
        RECT 31.755 133.270 32.270 133.680 ;
        RECT 32.505 132.920 32.675 133.680 ;
        RECT 32.845 133.260 33.015 133.925 ;
        RECT 33.185 133.940 33.375 135.300 ;
        RECT 33.545 134.790 33.820 135.300 ;
        RECT 34.010 134.935 34.540 135.300 ;
        RECT 34.965 135.070 35.295 135.470 ;
        RECT 34.365 134.900 34.540 134.935 ;
        RECT 33.545 134.620 33.825 134.790 ;
        RECT 33.545 134.140 33.820 134.620 ;
        RECT 34.025 133.940 34.195 134.740 ;
        RECT 33.185 133.770 34.195 133.940 ;
        RECT 34.365 134.730 35.295 134.900 ;
        RECT 35.465 134.730 35.720 135.300 ;
        RECT 34.365 133.600 34.535 134.730 ;
        RECT 35.125 134.560 35.295 134.730 ;
        RECT 33.410 133.430 34.535 133.600 ;
        RECT 34.705 134.230 34.900 134.560 ;
        RECT 35.125 134.230 35.380 134.560 ;
        RECT 34.705 133.260 34.875 134.230 ;
        RECT 35.550 134.060 35.720 134.730 ;
        RECT 35.895 134.700 37.565 135.470 ;
        RECT 32.845 133.090 34.875 133.260 ;
        RECT 35.045 132.920 35.215 134.060 ;
        RECT 35.385 133.090 35.720 134.060 ;
        RECT 35.895 134.010 36.645 134.530 ;
        RECT 36.815 134.180 37.565 134.700 ;
        RECT 37.735 134.795 38.005 135.140 ;
        RECT 38.195 135.070 38.575 135.470 ;
        RECT 38.745 134.900 38.915 135.250 ;
        RECT 39.085 135.070 39.415 135.470 ;
        RECT 39.615 134.900 39.785 135.250 ;
        RECT 39.985 134.970 40.315 135.470 ;
        RECT 37.735 134.060 37.905 134.795 ;
        RECT 38.175 134.730 39.785 134.900 ;
        RECT 38.175 134.560 38.345 134.730 ;
        RECT 38.075 134.230 38.345 134.560 ;
        RECT 38.515 134.230 38.920 134.560 ;
        RECT 38.175 134.060 38.345 134.230 ;
        RECT 39.090 134.110 39.800 134.560 ;
        RECT 39.970 134.230 40.320 134.800 ;
        RECT 40.495 134.795 40.765 135.140 ;
        RECT 40.955 135.070 41.335 135.470 ;
        RECT 41.505 134.900 41.675 135.250 ;
        RECT 41.845 135.070 42.175 135.470 ;
        RECT 42.375 134.900 42.545 135.250 ;
        RECT 42.745 134.970 43.075 135.470 ;
        RECT 35.895 132.920 37.565 134.010 ;
        RECT 37.735 133.090 38.005 134.060 ;
        RECT 38.175 133.890 38.900 134.060 ;
        RECT 39.090 133.940 39.805 134.110 ;
        RECT 40.495 134.060 40.665 134.795 ;
        RECT 40.935 134.730 42.545 134.900 ;
        RECT 40.935 134.560 41.105 134.730 ;
        RECT 40.835 134.230 41.105 134.560 ;
        RECT 41.275 134.230 41.680 134.560 ;
        RECT 40.935 134.060 41.105 134.230 ;
        RECT 41.850 134.110 42.560 134.560 ;
        RECT 42.730 134.230 43.080 134.800 ;
        RECT 43.255 134.670 43.595 135.300 ;
        RECT 43.765 134.670 44.015 135.470 ;
        RECT 44.205 134.820 44.535 135.300 ;
        RECT 44.705 135.010 44.930 135.470 ;
        RECT 45.100 134.820 45.430 135.300 ;
        RECT 43.255 134.620 43.485 134.670 ;
        RECT 44.205 134.650 45.430 134.820 ;
        RECT 46.060 134.690 46.560 135.300 ;
        RECT 38.730 133.770 38.900 133.890 ;
        RECT 40.000 133.770 40.320 134.060 ;
        RECT 38.215 132.920 38.495 133.720 ;
        RECT 38.730 133.600 40.320 133.770 ;
        RECT 38.665 133.140 40.320 133.430 ;
        RECT 40.495 133.090 40.765 134.060 ;
        RECT 40.935 133.890 41.660 134.060 ;
        RECT 41.850 133.940 42.565 134.110 ;
        RECT 43.255 134.060 43.430 134.620 ;
        RECT 43.600 134.310 44.295 134.480 ;
        RECT 44.125 134.060 44.295 134.310 ;
        RECT 44.470 134.280 44.890 134.480 ;
        RECT 45.060 134.280 45.390 134.480 ;
        RECT 45.560 134.280 45.890 134.480 ;
        RECT 46.060 134.060 46.230 134.690 ;
        RECT 47.210 134.660 47.455 135.265 ;
        RECT 47.675 134.935 48.185 135.470 ;
        RECT 46.935 134.490 48.165 134.660 ;
        RECT 46.415 134.230 46.765 134.480 ;
        RECT 41.490 133.770 41.660 133.890 ;
        RECT 42.760 133.770 43.080 134.060 ;
        RECT 40.975 132.920 41.255 133.720 ;
        RECT 41.490 133.600 43.080 133.770 ;
        RECT 41.425 133.140 43.080 133.430 ;
        RECT 43.255 133.090 43.595 134.060 ;
        RECT 43.765 132.920 43.935 134.060 ;
        RECT 44.125 133.890 46.560 134.060 ;
        RECT 44.205 132.920 44.455 133.720 ;
        RECT 45.100 133.090 45.430 133.890 ;
        RECT 45.730 132.920 46.060 133.720 ;
        RECT 46.230 133.090 46.560 133.890 ;
        RECT 46.935 133.680 47.275 134.490 ;
        RECT 47.445 133.925 48.195 134.115 ;
        RECT 46.935 133.270 47.450 133.680 ;
        RECT 47.685 132.920 47.855 133.680 ;
        RECT 48.025 133.260 48.195 133.925 ;
        RECT 48.365 133.940 48.555 135.300 ;
        RECT 48.725 134.790 49.000 135.300 ;
        RECT 49.190 134.935 49.720 135.300 ;
        RECT 50.145 135.070 50.475 135.470 ;
        RECT 49.545 134.900 49.720 134.935 ;
        RECT 48.725 134.620 49.005 134.790 ;
        RECT 48.725 134.140 49.000 134.620 ;
        RECT 49.205 133.940 49.375 134.740 ;
        RECT 48.365 133.770 49.375 133.940 ;
        RECT 49.545 134.730 50.475 134.900 ;
        RECT 50.645 134.730 50.900 135.300 ;
        RECT 51.075 134.745 51.365 135.470 ;
        RECT 52.085 134.920 52.255 135.300 ;
        RECT 52.435 135.090 52.765 135.470 ;
        RECT 52.085 134.750 52.750 134.920 ;
        RECT 52.945 134.795 53.205 135.300 ;
        RECT 49.545 133.600 49.715 134.730 ;
        RECT 50.305 134.560 50.475 134.730 ;
        RECT 48.590 133.430 49.715 133.600 ;
        RECT 49.885 134.230 50.080 134.560 ;
        RECT 50.305 134.230 50.560 134.560 ;
        RECT 49.885 133.260 50.055 134.230 ;
        RECT 50.730 134.060 50.900 134.730 ;
        RECT 52.015 134.200 52.345 134.570 ;
        RECT 52.580 134.495 52.750 134.750 ;
        RECT 52.580 134.165 52.865 134.495 ;
        RECT 48.025 133.090 50.055 133.260 ;
        RECT 50.225 132.920 50.395 134.060 ;
        RECT 50.565 133.090 50.900 134.060 ;
        RECT 51.075 132.920 51.365 134.085 ;
        RECT 52.580 134.020 52.750 134.165 ;
        RECT 52.085 133.850 52.750 134.020 ;
        RECT 53.035 133.995 53.205 134.795 ;
        RECT 53.650 134.660 53.895 135.265 ;
        RECT 54.115 134.935 54.625 135.470 ;
        RECT 52.085 133.090 52.255 133.850 ;
        RECT 52.435 132.920 52.765 133.680 ;
        RECT 52.935 133.090 53.205 133.995 ;
        RECT 53.375 134.490 54.605 134.660 ;
        RECT 53.375 133.680 53.715 134.490 ;
        RECT 53.885 133.925 54.635 134.115 ;
        RECT 53.375 133.270 53.890 133.680 ;
        RECT 54.125 132.920 54.295 133.680 ;
        RECT 54.465 133.260 54.635 133.925 ;
        RECT 54.805 133.940 54.995 135.300 ;
        RECT 55.165 134.450 55.440 135.300 ;
        RECT 55.630 134.935 56.160 135.300 ;
        RECT 56.585 135.070 56.915 135.470 ;
        RECT 55.985 134.900 56.160 134.935 ;
        RECT 55.165 134.280 55.445 134.450 ;
        RECT 55.165 134.140 55.440 134.280 ;
        RECT 55.645 133.940 55.815 134.740 ;
        RECT 54.805 133.770 55.815 133.940 ;
        RECT 55.985 134.730 56.915 134.900 ;
        RECT 57.085 134.730 57.340 135.300 ;
        RECT 55.985 133.600 56.155 134.730 ;
        RECT 56.745 134.560 56.915 134.730 ;
        RECT 55.030 133.430 56.155 133.600 ;
        RECT 56.325 134.230 56.520 134.560 ;
        RECT 56.745 134.230 57.000 134.560 ;
        RECT 56.325 133.260 56.495 134.230 ;
        RECT 57.170 134.060 57.340 134.730 ;
        RECT 57.515 134.720 58.725 135.470 ;
        RECT 54.465 133.090 56.495 133.260 ;
        RECT 56.665 132.920 56.835 134.060 ;
        RECT 57.005 133.090 57.340 134.060 ;
        RECT 57.515 134.010 58.035 134.550 ;
        RECT 58.205 134.180 58.725 134.720 ;
        RECT 59.270 134.760 59.525 135.290 ;
        RECT 59.705 135.010 59.990 135.470 ;
        RECT 57.515 132.920 58.725 134.010 ;
        RECT 59.270 133.900 59.450 134.760 ;
        RECT 60.170 134.560 60.420 135.210 ;
        RECT 59.620 134.230 60.420 134.560 ;
        RECT 59.270 133.430 59.525 133.900 ;
        RECT 59.185 133.260 59.525 133.430 ;
        RECT 59.270 133.230 59.525 133.260 ;
        RECT 59.705 132.920 59.990 133.720 ;
        RECT 60.170 133.640 60.420 134.230 ;
        RECT 60.620 134.875 60.940 135.205 ;
        RECT 61.120 134.990 61.780 135.470 ;
        RECT 61.980 135.080 62.830 135.250 ;
        RECT 60.620 133.980 60.810 134.875 ;
        RECT 61.130 134.550 61.790 134.820 ;
        RECT 61.460 134.490 61.790 134.550 ;
        RECT 60.980 134.320 61.310 134.380 ;
        RECT 61.980 134.320 62.150 135.080 ;
        RECT 63.390 135.010 63.710 135.470 ;
        RECT 63.910 134.830 64.160 135.260 ;
        RECT 64.450 135.030 64.860 135.470 ;
        RECT 65.030 135.090 66.045 135.290 ;
        RECT 62.320 134.660 63.570 134.830 ;
        RECT 62.320 134.540 62.650 134.660 ;
        RECT 60.980 134.150 62.880 134.320 ;
        RECT 60.620 133.810 62.540 133.980 ;
        RECT 60.620 133.790 60.940 133.810 ;
        RECT 60.170 133.130 60.500 133.640 ;
        RECT 60.770 133.180 60.940 133.790 ;
        RECT 62.710 133.640 62.880 134.150 ;
        RECT 63.050 134.080 63.230 134.490 ;
        RECT 63.400 133.900 63.570 134.660 ;
        RECT 61.110 132.920 61.440 133.610 ;
        RECT 61.670 133.470 62.880 133.640 ;
        RECT 63.050 133.590 63.570 133.900 ;
        RECT 63.740 134.490 64.160 134.830 ;
        RECT 64.450 134.490 64.860 134.820 ;
        RECT 63.740 133.720 63.930 134.490 ;
        RECT 65.030 134.360 65.200 135.090 ;
        RECT 66.345 134.920 66.515 135.250 ;
        RECT 66.685 135.090 67.015 135.470 ;
        RECT 65.370 134.540 65.720 134.910 ;
        RECT 65.030 134.320 65.450 134.360 ;
        RECT 64.100 134.150 65.450 134.320 ;
        RECT 64.100 133.990 64.350 134.150 ;
        RECT 64.860 133.720 65.110 133.980 ;
        RECT 63.740 133.470 65.110 133.720 ;
        RECT 61.670 133.180 61.910 133.470 ;
        RECT 62.710 133.390 62.880 133.470 ;
        RECT 62.110 132.920 62.530 133.300 ;
        RECT 62.710 133.140 63.340 133.390 ;
        RECT 63.810 132.920 64.140 133.300 ;
        RECT 64.310 133.180 64.480 133.470 ;
        RECT 65.280 133.305 65.450 134.150 ;
        RECT 65.900 133.980 66.120 134.850 ;
        RECT 66.345 134.730 67.040 134.920 ;
        RECT 65.620 133.600 66.120 133.980 ;
        RECT 66.290 133.930 66.700 134.550 ;
        RECT 66.870 133.760 67.040 134.730 ;
        RECT 66.345 133.590 67.040 133.760 ;
        RECT 64.660 132.920 65.040 133.300 ;
        RECT 65.280 133.135 66.110 133.305 ;
        RECT 66.345 133.090 66.515 133.590 ;
        RECT 66.685 132.920 67.015 133.420 ;
        RECT 67.230 133.090 67.455 135.210 ;
        RECT 67.625 135.090 67.955 135.470 ;
        RECT 68.125 134.920 68.295 135.210 ;
        RECT 67.630 134.750 68.295 134.920 ;
        RECT 67.630 133.760 67.860 134.750 ;
        RECT 68.555 134.700 72.065 135.470 ;
        RECT 68.030 133.930 68.380 134.580 ;
        RECT 68.555 134.010 70.245 134.530 ;
        RECT 70.415 134.180 72.065 134.700 ;
        RECT 72.235 134.795 72.505 135.140 ;
        RECT 72.695 135.070 73.075 135.470 ;
        RECT 73.245 134.900 73.415 135.250 ;
        RECT 73.585 135.070 73.915 135.470 ;
        RECT 74.115 134.900 74.285 135.250 ;
        RECT 74.485 134.970 74.815 135.470 ;
        RECT 72.235 134.060 72.405 134.795 ;
        RECT 72.675 134.730 74.285 134.900 ;
        RECT 72.675 134.560 72.845 134.730 ;
        RECT 72.575 134.230 72.845 134.560 ;
        RECT 73.015 134.230 73.420 134.560 ;
        RECT 72.675 134.060 72.845 134.230 ;
        RECT 73.590 134.110 74.300 134.560 ;
        RECT 74.470 134.230 74.820 134.800 ;
        RECT 74.995 134.700 76.665 135.470 ;
        RECT 76.835 134.745 77.125 135.470 ;
        RECT 67.630 133.590 68.295 133.760 ;
        RECT 67.625 132.920 67.955 133.420 ;
        RECT 68.125 133.090 68.295 133.590 ;
        RECT 68.555 132.920 72.065 134.010 ;
        RECT 72.235 133.090 72.505 134.060 ;
        RECT 72.675 133.890 73.400 134.060 ;
        RECT 73.590 133.940 74.305 134.110 ;
        RECT 73.230 133.770 73.400 133.890 ;
        RECT 74.500 133.770 74.820 134.060 ;
        RECT 72.715 132.920 72.995 133.720 ;
        RECT 73.230 133.600 74.820 133.770 ;
        RECT 74.995 134.010 75.745 134.530 ;
        RECT 75.915 134.180 76.665 134.700 ;
        RECT 77.300 134.730 77.555 135.300 ;
        RECT 77.725 135.070 78.055 135.470 ;
        RECT 78.480 134.935 79.010 135.300 ;
        RECT 78.480 134.900 78.655 134.935 ;
        RECT 77.725 134.730 78.655 134.900 ;
        RECT 79.200 134.790 79.475 135.300 ;
        RECT 73.165 133.140 74.820 133.430 ;
        RECT 74.995 132.920 76.665 134.010 ;
        RECT 76.835 132.920 77.125 134.085 ;
        RECT 77.300 134.060 77.470 134.730 ;
        RECT 77.725 134.560 77.895 134.730 ;
        RECT 77.640 134.230 77.895 134.560 ;
        RECT 78.120 134.230 78.315 134.560 ;
        RECT 77.300 133.090 77.635 134.060 ;
        RECT 77.805 132.920 77.975 134.060 ;
        RECT 78.145 133.260 78.315 134.230 ;
        RECT 78.485 133.600 78.655 134.730 ;
        RECT 78.825 133.940 78.995 134.740 ;
        RECT 79.195 134.620 79.475 134.790 ;
        RECT 79.200 134.140 79.475 134.620 ;
        RECT 79.645 133.940 79.835 135.300 ;
        RECT 80.015 134.935 80.525 135.470 ;
        RECT 80.745 134.660 80.990 135.265 ;
        RECT 81.895 134.700 83.565 135.470 ;
        RECT 80.035 134.490 81.265 134.660 ;
        RECT 78.825 133.770 79.835 133.940 ;
        RECT 80.005 133.925 80.755 134.115 ;
        RECT 78.485 133.430 79.610 133.600 ;
        RECT 80.005 133.260 80.175 133.925 ;
        RECT 80.925 133.680 81.265 134.490 ;
        RECT 78.145 133.090 80.175 133.260 ;
        RECT 80.345 132.920 80.515 133.680 ;
        RECT 80.750 133.270 81.265 133.680 ;
        RECT 81.895 134.010 82.645 134.530 ;
        RECT 82.815 134.180 83.565 134.700 ;
        RECT 83.795 134.650 84.005 135.470 ;
        RECT 84.175 134.670 84.505 135.300 ;
        RECT 84.175 134.070 84.425 134.670 ;
        RECT 84.675 134.650 84.905 135.470 ;
        RECT 86.035 134.795 86.295 135.300 ;
        RECT 86.475 135.090 86.805 135.470 ;
        RECT 86.985 134.920 87.155 135.300 ;
        RECT 84.595 134.230 84.925 134.480 ;
        RECT 81.895 132.920 83.565 134.010 ;
        RECT 83.795 132.920 84.005 134.060 ;
        RECT 84.175 133.090 84.505 134.070 ;
        RECT 84.675 132.920 84.905 134.060 ;
        RECT 86.035 133.995 86.205 134.795 ;
        RECT 86.490 134.750 87.155 134.920 ;
        RECT 87.415 134.795 87.675 135.300 ;
        RECT 87.855 135.090 88.185 135.470 ;
        RECT 88.365 134.920 88.535 135.300 ;
        RECT 86.490 134.495 86.660 134.750 ;
        RECT 86.375 134.165 86.660 134.495 ;
        RECT 86.895 134.200 87.225 134.570 ;
        RECT 86.490 134.020 86.660 134.165 ;
        RECT 86.035 133.090 86.305 133.995 ;
        RECT 86.490 133.850 87.155 134.020 ;
        RECT 86.475 132.920 86.805 133.680 ;
        RECT 86.985 133.090 87.155 133.850 ;
        RECT 87.415 133.995 87.585 134.795 ;
        RECT 87.870 134.750 88.535 134.920 ;
        RECT 87.870 134.495 88.040 134.750 ;
        RECT 88.795 134.720 90.005 135.470 ;
        RECT 87.755 134.165 88.040 134.495 ;
        RECT 88.275 134.200 88.605 134.570 ;
        RECT 87.870 134.020 88.040 134.165 ;
        RECT 87.415 133.090 87.685 133.995 ;
        RECT 87.870 133.850 88.535 134.020 ;
        RECT 87.855 132.920 88.185 133.680 ;
        RECT 88.365 133.090 88.535 133.850 ;
        RECT 88.795 134.010 89.315 134.550 ;
        RECT 89.485 134.180 90.005 134.720 ;
        RECT 90.175 135.010 90.735 135.300 ;
        RECT 90.905 135.010 91.155 135.470 ;
        RECT 88.795 132.920 90.005 134.010 ;
        RECT 90.175 133.640 90.425 135.010 ;
        RECT 91.775 134.840 92.105 135.200 ;
        RECT 90.715 134.650 92.105 134.840 ;
        RECT 92.475 135.010 93.035 135.300 ;
        RECT 93.205 135.010 93.455 135.470 ;
        RECT 90.715 134.560 90.885 134.650 ;
        RECT 90.595 134.230 90.885 134.560 ;
        RECT 91.055 134.230 91.395 134.480 ;
        RECT 91.615 134.230 92.290 134.480 ;
        RECT 90.715 133.980 90.885 134.230 ;
        RECT 90.715 133.810 91.655 133.980 ;
        RECT 92.025 133.870 92.290 134.230 ;
        RECT 90.175 133.090 90.635 133.640 ;
        RECT 90.825 132.920 91.155 133.640 ;
        RECT 91.355 133.260 91.655 133.810 ;
        RECT 92.475 133.640 92.725 135.010 ;
        RECT 94.075 134.840 94.405 135.200 ;
        RECT 95.755 134.990 96.035 135.470 ;
        RECT 93.015 134.650 94.405 134.840 ;
        RECT 96.205 134.820 96.465 135.210 ;
        RECT 96.640 134.990 96.895 135.470 ;
        RECT 97.065 134.820 97.360 135.210 ;
        RECT 97.540 134.990 97.815 135.470 ;
        RECT 97.985 134.970 98.285 135.300 ;
        RECT 95.710 134.650 97.360 134.820 ;
        RECT 93.015 134.560 93.185 134.650 ;
        RECT 92.895 134.230 93.185 134.560 ;
        RECT 93.355 134.230 93.695 134.480 ;
        RECT 93.915 134.230 94.590 134.480 ;
        RECT 93.015 133.980 93.185 134.230 ;
        RECT 93.015 133.810 93.955 133.980 ;
        RECT 94.325 133.870 94.590 134.230 ;
        RECT 95.710 134.140 96.115 134.650 ;
        RECT 96.285 134.310 97.425 134.480 ;
        RECT 95.710 133.970 96.465 134.140 ;
        RECT 91.825 132.920 92.105 133.590 ;
        RECT 92.475 133.090 92.935 133.640 ;
        RECT 93.125 132.920 93.455 133.640 ;
        RECT 93.655 133.260 93.955 133.810 ;
        RECT 94.125 132.920 94.405 133.590 ;
        RECT 95.750 132.920 96.035 133.790 ;
        RECT 96.205 133.720 96.465 133.970 ;
        RECT 97.255 134.060 97.425 134.310 ;
        RECT 97.595 134.230 97.945 134.800 ;
        RECT 98.115 134.060 98.285 134.970 ;
        RECT 98.655 134.840 98.985 135.200 ;
        RECT 99.605 135.010 99.855 135.470 ;
        RECT 100.025 135.010 100.585 135.300 ;
        RECT 98.655 134.650 100.045 134.840 ;
        RECT 99.875 134.560 100.045 134.650 ;
        RECT 97.255 133.890 98.285 134.060 ;
        RECT 96.205 133.550 97.325 133.720 ;
        RECT 96.205 133.090 96.465 133.550 ;
        RECT 96.640 132.920 96.895 133.380 ;
        RECT 97.065 133.090 97.325 133.550 ;
        RECT 97.495 132.920 97.805 133.720 ;
        RECT 97.975 133.090 98.285 133.890 ;
        RECT 98.470 134.230 99.145 134.480 ;
        RECT 99.365 134.230 99.705 134.480 ;
        RECT 99.875 134.230 100.165 134.560 ;
        RECT 98.470 133.870 98.735 134.230 ;
        RECT 99.875 133.980 100.045 134.230 ;
        RECT 99.105 133.810 100.045 133.980 ;
        RECT 98.655 132.920 98.935 133.590 ;
        RECT 99.105 133.260 99.405 133.810 ;
        RECT 100.335 133.640 100.585 135.010 ;
        RECT 100.755 134.700 102.425 135.470 ;
        RECT 102.595 134.745 102.885 135.470 ;
        RECT 103.520 134.925 108.865 135.470 ;
        RECT 109.040 134.925 114.385 135.470 ;
        RECT 99.605 132.920 99.935 133.640 ;
        RECT 100.125 133.090 100.585 133.640 ;
        RECT 100.755 134.010 101.505 134.530 ;
        RECT 101.675 134.180 102.425 134.700 ;
        RECT 100.755 132.920 102.425 134.010 ;
        RECT 102.595 132.920 102.885 134.085 ;
        RECT 105.110 133.355 105.460 134.605 ;
        RECT 106.940 134.095 107.280 134.925 ;
        RECT 110.630 133.355 110.980 134.605 ;
        RECT 112.460 134.095 112.800 134.925 ;
        RECT 114.555 134.720 115.765 135.470 ;
        RECT 114.555 134.010 115.075 134.550 ;
        RECT 115.245 134.180 115.765 134.720 ;
        RECT 103.520 132.920 108.865 133.355 ;
        RECT 109.040 132.920 114.385 133.355 ;
        RECT 114.555 132.920 115.765 134.010 ;
        RECT 14.650 132.750 115.850 132.920 ;
        RECT 14.735 131.660 15.945 132.750 ;
        RECT 16.950 132.410 17.205 132.440 ;
        RECT 16.865 132.240 17.205 132.410 ;
        RECT 14.735 130.950 15.255 131.490 ;
        RECT 15.425 131.120 15.945 131.660 ;
        RECT 16.950 131.770 17.205 132.240 ;
        RECT 17.385 131.950 17.670 132.750 ;
        RECT 17.850 132.030 18.180 132.540 ;
        RECT 14.735 130.200 15.945 130.950 ;
        RECT 16.950 130.910 17.130 131.770 ;
        RECT 17.850 131.440 18.100 132.030 ;
        RECT 18.450 131.880 18.620 132.490 ;
        RECT 18.790 132.060 19.120 132.750 ;
        RECT 19.350 132.200 19.590 132.490 ;
        RECT 19.790 132.370 20.210 132.750 ;
        RECT 20.390 132.280 21.020 132.530 ;
        RECT 21.490 132.370 21.820 132.750 ;
        RECT 20.390 132.200 20.560 132.280 ;
        RECT 21.990 132.200 22.160 132.490 ;
        RECT 22.340 132.370 22.720 132.750 ;
        RECT 22.960 132.365 23.790 132.535 ;
        RECT 19.350 132.030 20.560 132.200 ;
        RECT 17.300 131.110 18.100 131.440 ;
        RECT 16.950 130.380 17.205 130.910 ;
        RECT 17.385 130.200 17.670 130.660 ;
        RECT 17.850 130.460 18.100 131.110 ;
        RECT 18.300 131.860 18.620 131.880 ;
        RECT 18.300 131.690 20.220 131.860 ;
        RECT 18.300 130.795 18.490 131.690 ;
        RECT 20.390 131.520 20.560 132.030 ;
        RECT 20.730 131.770 21.250 132.080 ;
        RECT 18.660 131.350 20.560 131.520 ;
        RECT 18.660 131.290 18.990 131.350 ;
        RECT 19.140 131.120 19.470 131.180 ;
        RECT 18.810 130.850 19.470 131.120 ;
        RECT 18.300 130.465 18.620 130.795 ;
        RECT 18.800 130.200 19.460 130.680 ;
        RECT 19.660 130.590 19.830 131.350 ;
        RECT 20.730 131.180 20.910 131.590 ;
        RECT 20.000 131.010 20.330 131.130 ;
        RECT 21.080 131.010 21.250 131.770 ;
        RECT 20.000 130.840 21.250 131.010 ;
        RECT 21.420 131.950 22.790 132.200 ;
        RECT 21.420 131.180 21.610 131.950 ;
        RECT 22.540 131.690 22.790 131.950 ;
        RECT 21.780 131.520 22.030 131.680 ;
        RECT 22.960 131.520 23.130 132.365 ;
        RECT 24.025 132.080 24.195 132.580 ;
        RECT 24.365 132.250 24.695 132.750 ;
        RECT 23.300 131.690 23.800 132.070 ;
        RECT 24.025 131.910 24.720 132.080 ;
        RECT 21.780 131.350 23.130 131.520 ;
        RECT 22.710 131.310 23.130 131.350 ;
        RECT 21.420 130.840 21.840 131.180 ;
        RECT 22.130 130.850 22.540 131.180 ;
        RECT 19.660 130.420 20.510 130.590 ;
        RECT 21.070 130.200 21.390 130.660 ;
        RECT 21.590 130.410 21.840 130.840 ;
        RECT 22.130 130.200 22.540 130.640 ;
        RECT 22.710 130.580 22.880 131.310 ;
        RECT 23.050 130.760 23.400 131.130 ;
        RECT 23.580 130.820 23.800 131.690 ;
        RECT 23.970 131.120 24.380 131.740 ;
        RECT 24.550 130.940 24.720 131.910 ;
        RECT 24.025 130.750 24.720 130.940 ;
        RECT 22.710 130.380 23.725 130.580 ;
        RECT 24.025 130.420 24.195 130.750 ;
        RECT 24.365 130.200 24.695 130.580 ;
        RECT 24.910 130.460 25.135 132.580 ;
        RECT 25.305 132.250 25.635 132.750 ;
        RECT 25.805 132.080 25.975 132.580 ;
        RECT 25.310 131.910 25.975 132.080 ;
        RECT 25.310 130.920 25.540 131.910 ;
        RECT 25.710 131.090 26.060 131.740 ;
        RECT 26.275 131.610 26.505 132.750 ;
        RECT 26.675 131.600 27.005 132.580 ;
        RECT 27.175 131.610 27.385 132.750 ;
        RECT 27.990 132.410 28.245 132.440 ;
        RECT 27.905 132.240 28.245 132.410 ;
        RECT 27.990 131.770 28.245 132.240 ;
        RECT 28.425 131.950 28.710 132.750 ;
        RECT 28.890 132.030 29.220 132.540 ;
        RECT 26.255 131.190 26.585 131.440 ;
        RECT 25.310 130.750 25.975 130.920 ;
        RECT 25.305 130.200 25.635 130.580 ;
        RECT 25.805 130.460 25.975 130.750 ;
        RECT 26.275 130.200 26.505 131.020 ;
        RECT 26.755 131.000 27.005 131.600 ;
        RECT 26.675 130.370 27.005 131.000 ;
        RECT 27.175 130.200 27.385 131.020 ;
        RECT 27.990 130.910 28.170 131.770 ;
        RECT 28.890 131.440 29.140 132.030 ;
        RECT 29.490 131.880 29.660 132.490 ;
        RECT 29.830 132.060 30.160 132.750 ;
        RECT 30.390 132.200 30.630 132.490 ;
        RECT 30.830 132.370 31.250 132.750 ;
        RECT 31.430 132.280 32.060 132.530 ;
        RECT 32.530 132.370 32.860 132.750 ;
        RECT 31.430 132.200 31.600 132.280 ;
        RECT 33.030 132.200 33.200 132.490 ;
        RECT 33.380 132.370 33.760 132.750 ;
        RECT 34.000 132.365 34.830 132.535 ;
        RECT 30.390 132.030 31.600 132.200 ;
        RECT 28.340 131.110 29.140 131.440 ;
        RECT 27.990 130.380 28.245 130.910 ;
        RECT 28.425 130.200 28.710 130.660 ;
        RECT 28.890 130.460 29.140 131.110 ;
        RECT 29.340 131.860 29.660 131.880 ;
        RECT 29.340 131.690 31.260 131.860 ;
        RECT 29.340 130.795 29.530 131.690 ;
        RECT 31.430 131.520 31.600 132.030 ;
        RECT 31.770 131.770 32.290 132.080 ;
        RECT 29.700 131.350 31.600 131.520 ;
        RECT 29.700 131.290 30.030 131.350 ;
        RECT 30.180 131.120 30.510 131.180 ;
        RECT 29.850 130.850 30.510 131.120 ;
        RECT 29.340 130.465 29.660 130.795 ;
        RECT 29.840 130.200 30.500 130.680 ;
        RECT 30.700 130.590 30.870 131.350 ;
        RECT 31.770 131.180 31.950 131.590 ;
        RECT 31.040 131.010 31.370 131.130 ;
        RECT 32.120 131.010 32.290 131.770 ;
        RECT 31.040 130.840 32.290 131.010 ;
        RECT 32.460 131.950 33.830 132.200 ;
        RECT 32.460 131.180 32.650 131.950 ;
        RECT 33.580 131.690 33.830 131.950 ;
        RECT 32.820 131.520 33.070 131.680 ;
        RECT 34.000 131.520 34.170 132.365 ;
        RECT 35.065 132.080 35.235 132.580 ;
        RECT 35.405 132.250 35.735 132.750 ;
        RECT 34.340 131.690 34.840 132.070 ;
        RECT 35.065 131.910 35.760 132.080 ;
        RECT 32.820 131.350 34.170 131.520 ;
        RECT 33.750 131.310 34.170 131.350 ;
        RECT 32.460 130.840 32.880 131.180 ;
        RECT 33.170 130.850 33.580 131.180 ;
        RECT 30.700 130.420 31.550 130.590 ;
        RECT 32.110 130.200 32.430 130.660 ;
        RECT 32.630 130.410 32.880 130.840 ;
        RECT 33.170 130.200 33.580 130.640 ;
        RECT 33.750 130.580 33.920 131.310 ;
        RECT 34.090 130.760 34.440 131.130 ;
        RECT 34.620 130.820 34.840 131.690 ;
        RECT 35.010 131.120 35.420 131.740 ;
        RECT 35.590 130.940 35.760 131.910 ;
        RECT 35.065 130.750 35.760 130.940 ;
        RECT 33.750 130.380 34.765 130.580 ;
        RECT 35.065 130.420 35.235 130.750 ;
        RECT 35.405 130.200 35.735 130.580 ;
        RECT 35.950 130.460 36.175 132.580 ;
        RECT 36.345 132.250 36.675 132.750 ;
        RECT 36.845 132.080 37.015 132.580 ;
        RECT 36.350 131.910 37.015 132.080 ;
        RECT 36.350 130.920 36.580 131.910 ;
        RECT 36.750 131.090 37.100 131.740 ;
        RECT 38.195 131.585 38.485 132.750 ;
        RECT 38.855 132.080 39.135 132.750 ;
        RECT 39.305 131.860 39.605 132.410 ;
        RECT 39.805 132.030 40.135 132.750 ;
        RECT 40.325 132.030 40.785 132.580 ;
        RECT 38.670 131.440 38.935 131.800 ;
        RECT 39.305 131.690 40.245 131.860 ;
        RECT 40.075 131.440 40.245 131.690 ;
        RECT 38.670 131.190 39.345 131.440 ;
        RECT 39.565 131.190 39.905 131.440 ;
        RECT 40.075 131.110 40.365 131.440 ;
        RECT 40.075 131.020 40.245 131.110 ;
        RECT 36.350 130.750 37.015 130.920 ;
        RECT 36.345 130.200 36.675 130.580 ;
        RECT 36.845 130.460 37.015 130.750 ;
        RECT 38.195 130.200 38.485 130.925 ;
        RECT 38.855 130.830 40.245 131.020 ;
        RECT 38.855 130.470 39.185 130.830 ;
        RECT 40.535 130.660 40.785 132.030 ;
        RECT 40.955 131.660 42.165 132.750 ;
        RECT 42.335 132.030 42.795 132.580 ;
        RECT 42.985 132.030 43.315 132.750 ;
        RECT 40.955 131.120 41.475 131.660 ;
        RECT 41.645 130.950 42.165 131.490 ;
        RECT 39.805 130.200 40.055 130.660 ;
        RECT 40.225 130.370 40.785 130.660 ;
        RECT 40.955 130.200 42.165 130.950 ;
        RECT 42.335 130.660 42.585 132.030 ;
        RECT 43.515 131.860 43.815 132.410 ;
        RECT 43.985 132.080 44.265 132.750 ;
        RECT 42.875 131.690 43.815 131.860 ;
        RECT 42.875 131.440 43.045 131.690 ;
        RECT 44.185 131.440 44.450 131.800 ;
        RECT 42.755 131.110 43.045 131.440 ;
        RECT 43.215 131.190 43.555 131.440 ;
        RECT 43.775 131.190 44.450 131.440 ;
        RECT 44.635 131.610 44.975 132.580 ;
        RECT 45.145 131.610 45.315 132.750 ;
        RECT 45.585 131.950 45.835 132.750 ;
        RECT 46.480 131.780 46.810 132.580 ;
        RECT 47.110 131.950 47.440 132.750 ;
        RECT 47.610 131.780 47.940 132.580 ;
        RECT 45.505 131.610 47.940 131.780 ;
        RECT 48.690 131.770 48.945 132.440 ;
        RECT 49.125 131.950 49.410 132.750 ;
        RECT 49.590 132.030 49.920 132.540 ;
        RECT 48.690 131.730 48.870 131.770 ;
        RECT 42.875 131.020 43.045 131.110 ;
        RECT 42.875 130.830 44.265 131.020 ;
        RECT 42.335 130.370 42.895 130.660 ;
        RECT 43.065 130.200 43.315 130.660 ;
        RECT 43.935 130.470 44.265 130.830 ;
        RECT 44.635 131.000 44.810 131.610 ;
        RECT 45.505 131.360 45.675 131.610 ;
        RECT 44.980 131.190 45.675 131.360 ;
        RECT 45.850 131.190 46.270 131.390 ;
        RECT 46.440 131.190 46.770 131.390 ;
        RECT 46.940 131.190 47.270 131.390 ;
        RECT 44.635 130.370 44.975 131.000 ;
        RECT 45.145 130.200 45.395 131.000 ;
        RECT 45.585 130.850 46.810 131.020 ;
        RECT 45.585 130.370 45.915 130.850 ;
        RECT 46.085 130.200 46.310 130.660 ;
        RECT 46.480 130.370 46.810 130.850 ;
        RECT 47.440 130.980 47.610 131.610 ;
        RECT 48.605 131.560 48.870 131.730 ;
        RECT 47.795 131.190 48.145 131.440 ;
        RECT 47.440 130.370 47.940 130.980 ;
        RECT 48.690 130.910 48.870 131.560 ;
        RECT 49.590 131.440 49.840 132.030 ;
        RECT 50.190 131.880 50.360 132.490 ;
        RECT 50.530 132.060 50.860 132.750 ;
        RECT 51.090 132.200 51.330 132.490 ;
        RECT 51.530 132.370 51.950 132.750 ;
        RECT 52.130 132.280 52.760 132.530 ;
        RECT 53.230 132.370 53.560 132.750 ;
        RECT 52.130 132.200 52.300 132.280 ;
        RECT 53.730 132.200 53.900 132.490 ;
        RECT 54.080 132.370 54.460 132.750 ;
        RECT 54.700 132.365 55.530 132.535 ;
        RECT 51.090 132.030 52.300 132.200 ;
        RECT 49.040 131.110 49.840 131.440 ;
        RECT 48.690 130.380 48.945 130.910 ;
        RECT 49.125 130.200 49.410 130.660 ;
        RECT 49.590 130.460 49.840 131.110 ;
        RECT 50.040 131.860 50.360 131.880 ;
        RECT 50.040 131.690 51.960 131.860 ;
        RECT 50.040 130.795 50.230 131.690 ;
        RECT 52.130 131.520 52.300 132.030 ;
        RECT 52.470 131.770 52.990 132.080 ;
        RECT 50.400 131.350 52.300 131.520 ;
        RECT 50.400 131.290 50.730 131.350 ;
        RECT 50.880 131.120 51.210 131.180 ;
        RECT 50.550 130.850 51.210 131.120 ;
        RECT 50.040 130.465 50.360 130.795 ;
        RECT 50.540 130.200 51.200 130.680 ;
        RECT 51.400 130.590 51.570 131.350 ;
        RECT 52.470 131.180 52.650 131.590 ;
        RECT 51.740 131.010 52.070 131.130 ;
        RECT 52.820 131.010 52.990 131.770 ;
        RECT 51.740 130.840 52.990 131.010 ;
        RECT 53.160 131.950 54.530 132.200 ;
        RECT 53.160 131.180 53.350 131.950 ;
        RECT 54.280 131.690 54.530 131.950 ;
        RECT 53.520 131.520 53.770 131.680 ;
        RECT 54.700 131.520 54.870 132.365 ;
        RECT 55.765 132.080 55.935 132.580 ;
        RECT 56.105 132.250 56.435 132.750 ;
        RECT 55.040 131.690 55.540 132.070 ;
        RECT 55.765 131.910 56.460 132.080 ;
        RECT 53.520 131.350 54.870 131.520 ;
        RECT 54.450 131.310 54.870 131.350 ;
        RECT 53.160 130.840 53.580 131.180 ;
        RECT 53.870 130.850 54.280 131.180 ;
        RECT 51.400 130.420 52.250 130.590 ;
        RECT 52.810 130.200 53.130 130.660 ;
        RECT 53.330 130.410 53.580 130.840 ;
        RECT 53.870 130.200 54.280 130.640 ;
        RECT 54.450 130.580 54.620 131.310 ;
        RECT 54.790 130.760 55.140 131.130 ;
        RECT 55.320 130.820 55.540 131.690 ;
        RECT 55.710 131.120 56.120 131.740 ;
        RECT 56.290 130.940 56.460 131.910 ;
        RECT 55.765 130.750 56.460 130.940 ;
        RECT 54.450 130.380 55.465 130.580 ;
        RECT 55.765 130.420 55.935 130.750 ;
        RECT 56.105 130.200 56.435 130.580 ;
        RECT 56.650 130.460 56.875 132.580 ;
        RECT 57.045 132.250 57.375 132.750 ;
        RECT 57.545 132.080 57.715 132.580 ;
        RECT 57.050 131.910 57.715 132.080 ;
        RECT 58.895 131.990 59.410 132.400 ;
        RECT 59.645 131.990 59.815 132.750 ;
        RECT 59.985 132.410 62.015 132.580 ;
        RECT 57.050 130.920 57.280 131.910 ;
        RECT 57.450 131.090 57.800 131.740 ;
        RECT 58.895 131.180 59.235 131.990 ;
        RECT 59.985 131.745 60.155 132.410 ;
        RECT 60.550 132.070 61.675 132.240 ;
        RECT 59.405 131.555 60.155 131.745 ;
        RECT 60.325 131.730 61.335 131.900 ;
        RECT 58.895 131.010 60.125 131.180 ;
        RECT 57.050 130.750 57.715 130.920 ;
        RECT 57.045 130.200 57.375 130.580 ;
        RECT 57.545 130.460 57.715 130.750 ;
        RECT 59.170 130.405 59.415 131.010 ;
        RECT 59.635 130.200 60.145 130.735 ;
        RECT 60.325 130.370 60.515 131.730 ;
        RECT 60.685 130.710 60.960 131.530 ;
        RECT 61.165 130.930 61.335 131.730 ;
        RECT 61.505 130.940 61.675 132.070 ;
        RECT 61.845 131.440 62.015 132.410 ;
        RECT 62.185 131.610 62.355 132.750 ;
        RECT 62.525 131.610 62.860 132.580 ;
        RECT 61.845 131.110 62.040 131.440 ;
        RECT 62.265 131.110 62.520 131.440 ;
        RECT 62.265 130.940 62.435 131.110 ;
        RECT 62.690 130.940 62.860 131.610 ;
        RECT 63.955 131.585 64.245 132.750 ;
        RECT 65.335 132.030 65.795 132.580 ;
        RECT 65.985 132.030 66.315 132.750 ;
        RECT 61.505 130.770 62.435 130.940 ;
        RECT 61.505 130.735 61.680 130.770 ;
        RECT 60.685 130.540 60.965 130.710 ;
        RECT 60.685 130.370 60.960 130.540 ;
        RECT 61.150 130.370 61.680 130.735 ;
        RECT 62.105 130.200 62.435 130.600 ;
        RECT 62.605 130.370 62.860 130.940 ;
        RECT 63.955 130.200 64.245 130.925 ;
        RECT 65.335 130.660 65.585 132.030 ;
        RECT 66.515 131.860 66.815 132.410 ;
        RECT 66.985 132.080 67.265 132.750 ;
        RECT 65.875 131.690 66.815 131.860 ;
        RECT 65.875 131.440 66.045 131.690 ;
        RECT 67.185 131.440 67.450 131.800 ;
        RECT 65.755 131.110 66.045 131.440 ;
        RECT 66.215 131.190 66.555 131.440 ;
        RECT 66.775 131.190 67.450 131.440 ;
        RECT 67.635 131.780 67.905 132.550 ;
        RECT 68.075 131.970 68.405 132.750 ;
        RECT 68.610 132.145 68.795 132.550 ;
        RECT 68.965 132.325 69.300 132.750 ;
        RECT 68.610 131.970 69.275 132.145 ;
        RECT 67.635 131.610 68.765 131.780 ;
        RECT 65.875 131.020 66.045 131.110 ;
        RECT 65.875 130.830 67.265 131.020 ;
        RECT 65.335 130.370 65.895 130.660 ;
        RECT 66.065 130.200 66.315 130.660 ;
        RECT 66.935 130.470 67.265 130.830 ;
        RECT 67.635 130.700 67.805 131.610 ;
        RECT 67.975 130.860 68.335 131.440 ;
        RECT 68.515 131.110 68.765 131.610 ;
        RECT 68.935 130.940 69.275 131.970 ;
        RECT 68.590 130.770 69.275 130.940 ;
        RECT 69.475 131.675 69.745 132.580 ;
        RECT 69.915 131.990 70.245 132.750 ;
        RECT 70.425 131.820 70.595 132.580 ;
        RECT 69.475 130.875 69.645 131.675 ;
        RECT 69.930 131.650 70.595 131.820 ;
        RECT 70.855 131.660 72.065 132.750 ;
        RECT 72.235 132.030 72.695 132.580 ;
        RECT 72.885 132.030 73.215 132.750 ;
        RECT 69.930 131.505 70.100 131.650 ;
        RECT 69.815 131.175 70.100 131.505 ;
        RECT 69.930 130.920 70.100 131.175 ;
        RECT 70.335 131.100 70.665 131.470 ;
        RECT 70.855 131.120 71.375 131.660 ;
        RECT 71.545 130.950 72.065 131.490 ;
        RECT 67.635 130.370 67.895 130.700 ;
        RECT 68.105 130.200 68.380 130.680 ;
        RECT 68.590 130.370 68.795 130.770 ;
        RECT 68.965 130.200 69.300 130.600 ;
        RECT 69.475 130.370 69.735 130.875 ;
        RECT 69.930 130.750 70.595 130.920 ;
        RECT 69.915 130.200 70.245 130.580 ;
        RECT 70.425 130.370 70.595 130.750 ;
        RECT 70.855 130.200 72.065 130.950 ;
        RECT 72.235 130.660 72.485 132.030 ;
        RECT 73.415 131.860 73.715 132.410 ;
        RECT 73.885 132.080 74.165 132.750 ;
        RECT 72.775 131.690 73.715 131.860 ;
        RECT 72.775 131.440 72.945 131.690 ;
        RECT 74.085 131.440 74.350 131.800 ;
        RECT 72.655 131.110 72.945 131.440 ;
        RECT 73.115 131.190 73.455 131.440 ;
        RECT 73.675 131.190 74.350 131.440 ;
        RECT 74.535 131.660 75.745 132.750 ;
        RECT 76.005 132.005 76.275 132.750 ;
        RECT 76.905 132.745 83.180 132.750 ;
        RECT 76.445 131.835 76.735 132.575 ;
        RECT 76.905 132.020 77.160 132.745 ;
        RECT 77.345 131.850 77.605 132.575 ;
        RECT 77.775 132.020 78.020 132.745 ;
        RECT 78.205 131.850 78.465 132.575 ;
        RECT 78.635 132.020 78.880 132.745 ;
        RECT 79.065 131.850 79.325 132.575 ;
        RECT 79.495 132.020 79.740 132.745 ;
        RECT 79.910 131.850 80.170 132.575 ;
        RECT 80.340 132.020 80.600 132.745 ;
        RECT 80.770 131.850 81.030 132.575 ;
        RECT 81.200 132.020 81.460 132.745 ;
        RECT 81.630 131.850 81.890 132.575 ;
        RECT 82.060 132.020 82.320 132.745 ;
        RECT 82.490 131.850 82.750 132.575 ;
        RECT 82.920 131.950 83.180 132.745 ;
        RECT 77.345 131.835 82.750 131.850 ;
        RECT 74.535 131.120 75.055 131.660 ;
        RECT 76.005 131.610 82.750 131.835 ;
        RECT 72.775 131.020 72.945 131.110 ;
        RECT 72.775 130.830 74.165 131.020 ;
        RECT 75.225 130.950 75.745 131.490 ;
        RECT 72.235 130.370 72.795 130.660 ;
        RECT 72.965 130.200 73.215 130.660 ;
        RECT 73.835 130.470 74.165 130.830 ;
        RECT 74.535 130.200 75.745 130.950 ;
        RECT 76.005 131.020 77.170 131.610 ;
        RECT 83.350 131.440 83.600 132.575 ;
        RECT 83.780 131.940 84.040 132.750 ;
        RECT 84.215 131.440 84.460 132.580 ;
        RECT 84.640 131.940 84.935 132.750 ;
        RECT 85.120 131.610 85.455 132.580 ;
        RECT 85.625 131.610 85.795 132.750 ;
        RECT 85.965 132.410 87.995 132.580 ;
        RECT 77.340 131.190 84.460 131.440 ;
        RECT 76.005 130.850 82.750 131.020 ;
        RECT 76.005 130.200 76.305 130.680 ;
        RECT 76.475 130.395 76.735 130.850 ;
        RECT 76.905 130.200 77.165 130.680 ;
        RECT 77.345 130.395 77.605 130.850 ;
        RECT 77.775 130.200 78.025 130.680 ;
        RECT 78.205 130.395 78.465 130.850 ;
        RECT 78.635 130.200 78.885 130.680 ;
        RECT 79.065 130.395 79.325 130.850 ;
        RECT 79.495 130.200 79.740 130.680 ;
        RECT 79.910 130.395 80.185 130.850 ;
        RECT 80.355 130.200 80.600 130.680 ;
        RECT 80.770 130.395 81.030 130.850 ;
        RECT 81.200 130.200 81.460 130.680 ;
        RECT 81.630 130.395 81.890 130.850 ;
        RECT 82.060 130.200 82.320 130.680 ;
        RECT 82.490 130.395 82.750 130.850 ;
        RECT 82.920 130.200 83.180 130.760 ;
        RECT 83.350 130.380 83.600 131.190 ;
        RECT 83.780 130.200 84.040 130.725 ;
        RECT 84.210 130.380 84.460 131.190 ;
        RECT 84.630 130.880 84.945 131.440 ;
        RECT 85.120 130.940 85.290 131.610 ;
        RECT 85.965 131.440 86.135 132.410 ;
        RECT 85.460 131.110 85.715 131.440 ;
        RECT 85.940 131.110 86.135 131.440 ;
        RECT 86.305 132.070 87.430 132.240 ;
        RECT 85.545 130.940 85.715 131.110 ;
        RECT 86.305 130.940 86.475 132.070 ;
        RECT 84.640 130.200 84.945 130.710 ;
        RECT 85.120 130.370 85.375 130.940 ;
        RECT 85.545 130.770 86.475 130.940 ;
        RECT 86.645 131.730 87.655 131.900 ;
        RECT 86.645 130.930 86.815 131.730 ;
        RECT 87.020 131.390 87.295 131.530 ;
        RECT 87.015 131.220 87.295 131.390 ;
        RECT 86.300 130.735 86.475 130.770 ;
        RECT 85.545 130.200 85.875 130.600 ;
        RECT 86.300 130.370 86.830 130.735 ;
        RECT 87.020 130.370 87.295 131.220 ;
        RECT 87.465 130.370 87.655 131.730 ;
        RECT 87.825 131.745 87.995 132.410 ;
        RECT 88.165 131.990 88.335 132.750 ;
        RECT 88.570 131.990 89.085 132.400 ;
        RECT 87.825 131.555 88.575 131.745 ;
        RECT 88.745 131.180 89.085 131.990 ;
        RECT 89.715 131.585 90.005 132.750 ;
        RECT 90.265 132.005 90.535 132.750 ;
        RECT 91.165 132.745 97.440 132.750 ;
        RECT 90.705 131.835 90.995 132.575 ;
        RECT 91.165 132.020 91.420 132.745 ;
        RECT 91.605 131.850 91.865 132.575 ;
        RECT 92.035 132.020 92.280 132.745 ;
        RECT 92.465 131.850 92.725 132.575 ;
        RECT 92.895 132.020 93.140 132.745 ;
        RECT 93.325 131.850 93.585 132.575 ;
        RECT 93.755 132.020 94.000 132.745 ;
        RECT 94.170 131.850 94.430 132.575 ;
        RECT 94.600 132.020 94.860 132.745 ;
        RECT 95.030 131.850 95.290 132.575 ;
        RECT 95.460 132.020 95.720 132.745 ;
        RECT 95.890 131.850 96.150 132.575 ;
        RECT 96.320 132.020 96.580 132.745 ;
        RECT 96.750 131.850 97.010 132.575 ;
        RECT 97.180 131.950 97.440 132.745 ;
        RECT 91.605 131.835 97.010 131.850 ;
        RECT 90.265 131.610 97.010 131.835 ;
        RECT 87.855 131.010 89.085 131.180 ;
        RECT 90.265 131.020 91.430 131.610 ;
        RECT 97.610 131.440 97.860 132.575 ;
        RECT 98.040 131.940 98.300 132.750 ;
        RECT 98.475 131.440 98.720 132.580 ;
        RECT 98.900 131.940 99.195 132.750 ;
        RECT 99.575 132.080 99.855 132.750 ;
        RECT 100.025 131.860 100.325 132.410 ;
        RECT 100.525 132.030 100.855 132.750 ;
        RECT 101.045 132.030 101.505 132.580 ;
        RECT 99.390 131.440 99.655 131.800 ;
        RECT 100.025 131.690 100.965 131.860 ;
        RECT 100.795 131.440 100.965 131.690 ;
        RECT 91.600 131.190 98.720 131.440 ;
        RECT 87.835 130.200 88.345 130.735 ;
        RECT 88.565 130.405 88.810 131.010 ;
        RECT 89.715 130.200 90.005 130.925 ;
        RECT 90.265 130.850 97.010 131.020 ;
        RECT 90.265 130.200 90.565 130.680 ;
        RECT 90.735 130.395 90.995 130.850 ;
        RECT 91.165 130.200 91.425 130.680 ;
        RECT 91.605 130.395 91.865 130.850 ;
        RECT 92.035 130.200 92.285 130.680 ;
        RECT 92.465 130.395 92.725 130.850 ;
        RECT 92.895 130.200 93.145 130.680 ;
        RECT 93.325 130.395 93.585 130.850 ;
        RECT 93.755 130.200 94.000 130.680 ;
        RECT 94.170 130.395 94.445 130.850 ;
        RECT 94.615 130.200 94.860 130.680 ;
        RECT 95.030 130.395 95.290 130.850 ;
        RECT 95.460 130.200 95.720 130.680 ;
        RECT 95.890 130.395 96.150 130.850 ;
        RECT 96.320 130.200 96.580 130.680 ;
        RECT 96.750 130.395 97.010 130.850 ;
        RECT 97.180 130.200 97.440 130.760 ;
        RECT 97.610 130.380 97.860 131.190 ;
        RECT 98.040 130.200 98.300 130.725 ;
        RECT 98.470 130.380 98.720 131.190 ;
        RECT 98.890 130.880 99.205 131.440 ;
        RECT 99.390 131.190 100.065 131.440 ;
        RECT 100.285 131.190 100.625 131.440 ;
        RECT 100.795 131.110 101.085 131.440 ;
        RECT 100.795 131.020 100.965 131.110 ;
        RECT 99.575 130.830 100.965 131.020 ;
        RECT 98.900 130.200 99.205 130.710 ;
        RECT 99.575 130.470 99.905 130.830 ;
        RECT 101.255 130.660 101.505 132.030 ;
        RECT 101.675 131.990 102.190 132.400 ;
        RECT 102.425 131.990 102.595 132.750 ;
        RECT 102.765 132.410 104.795 132.580 ;
        RECT 101.675 131.180 102.015 131.990 ;
        RECT 102.765 131.745 102.935 132.410 ;
        RECT 103.330 132.070 104.455 132.240 ;
        RECT 102.185 131.555 102.935 131.745 ;
        RECT 103.105 131.730 104.115 131.900 ;
        RECT 101.675 131.010 102.905 131.180 ;
        RECT 100.525 130.200 100.775 130.660 ;
        RECT 100.945 130.370 101.505 130.660 ;
        RECT 101.950 130.405 102.195 131.010 ;
        RECT 102.415 130.200 102.925 130.735 ;
        RECT 103.105 130.370 103.295 131.730 ;
        RECT 103.465 130.710 103.740 131.530 ;
        RECT 103.945 130.930 104.115 131.730 ;
        RECT 104.285 130.940 104.455 132.070 ;
        RECT 104.625 131.440 104.795 132.410 ;
        RECT 104.965 131.610 105.135 132.750 ;
        RECT 105.305 131.610 105.640 132.580 ;
        RECT 104.625 131.110 104.820 131.440 ;
        RECT 105.045 131.110 105.300 131.440 ;
        RECT 105.045 130.940 105.215 131.110 ;
        RECT 105.470 130.940 105.640 131.610 ;
        RECT 105.815 131.660 107.485 132.750 ;
        RECT 105.815 131.140 106.565 131.660 ;
        RECT 107.695 131.610 107.925 132.750 ;
        RECT 108.095 131.600 108.425 132.580 ;
        RECT 108.595 131.610 108.805 132.750 ;
        RECT 109.585 131.820 109.755 132.580 ;
        RECT 109.935 131.990 110.265 132.750 ;
        RECT 109.585 131.650 110.250 131.820 ;
        RECT 110.435 131.675 110.705 132.580 ;
        RECT 106.735 130.970 107.485 131.490 ;
        RECT 107.675 131.190 108.005 131.440 ;
        RECT 104.285 130.770 105.215 130.940 ;
        RECT 104.285 130.735 104.460 130.770 ;
        RECT 103.465 130.540 103.745 130.710 ;
        RECT 103.465 130.370 103.740 130.540 ;
        RECT 103.930 130.370 104.460 130.735 ;
        RECT 104.885 130.200 105.215 130.600 ;
        RECT 105.385 130.370 105.640 130.940 ;
        RECT 105.815 130.200 107.485 130.970 ;
        RECT 107.695 130.200 107.925 131.020 ;
        RECT 108.175 131.000 108.425 131.600 ;
        RECT 110.080 131.505 110.250 131.650 ;
        RECT 109.515 131.100 109.845 131.470 ;
        RECT 110.080 131.175 110.365 131.505 ;
        RECT 108.095 130.370 108.425 131.000 ;
        RECT 108.595 130.200 108.805 131.020 ;
        RECT 110.080 130.920 110.250 131.175 ;
        RECT 109.585 130.750 110.250 130.920 ;
        RECT 110.535 130.875 110.705 131.675 ;
        RECT 110.875 131.660 114.385 132.750 ;
        RECT 114.555 131.660 115.765 132.750 ;
        RECT 110.875 131.140 112.565 131.660 ;
        RECT 112.735 130.970 114.385 131.490 ;
        RECT 114.555 131.120 115.075 131.660 ;
        RECT 109.585 130.370 109.755 130.750 ;
        RECT 109.935 130.200 110.265 130.580 ;
        RECT 110.445 130.370 110.705 130.875 ;
        RECT 110.875 130.200 114.385 130.970 ;
        RECT 115.245 130.950 115.765 131.490 ;
        RECT 114.555 130.200 115.765 130.950 ;
        RECT 14.650 130.030 115.850 130.200 ;
        RECT 14.735 129.280 15.945 130.030 ;
        RECT 14.735 128.740 15.255 129.280 ;
        RECT 16.115 129.260 18.705 130.030 ;
        RECT 18.965 129.480 19.135 129.860 ;
        RECT 19.315 129.650 19.645 130.030 ;
        RECT 18.965 129.310 19.630 129.480 ;
        RECT 19.825 129.355 20.085 129.860 ;
        RECT 15.425 128.570 15.945 129.110 ;
        RECT 14.735 127.480 15.945 128.570 ;
        RECT 16.115 128.570 17.325 129.090 ;
        RECT 17.495 128.740 18.705 129.260 ;
        RECT 18.895 128.760 19.225 129.130 ;
        RECT 19.460 129.055 19.630 129.310 ;
        RECT 19.460 128.725 19.745 129.055 ;
        RECT 19.460 128.580 19.630 128.725 ;
        RECT 16.115 127.480 18.705 128.570 ;
        RECT 18.965 128.410 19.630 128.580 ;
        RECT 19.915 128.555 20.085 129.355 ;
        RECT 18.965 127.650 19.135 128.410 ;
        RECT 19.315 127.480 19.645 128.240 ;
        RECT 19.815 127.650 20.085 128.555 ;
        RECT 20.260 129.290 20.515 129.860 ;
        RECT 20.685 129.630 21.015 130.030 ;
        RECT 21.440 129.495 21.970 129.860 ;
        RECT 21.440 129.460 21.615 129.495 ;
        RECT 20.685 129.290 21.615 129.460 ;
        RECT 22.160 129.350 22.435 129.860 ;
        RECT 20.260 128.620 20.430 129.290 ;
        RECT 20.685 129.120 20.855 129.290 ;
        RECT 20.600 128.790 20.855 129.120 ;
        RECT 21.080 128.790 21.275 129.120 ;
        RECT 20.260 127.650 20.595 128.620 ;
        RECT 20.765 127.480 20.935 128.620 ;
        RECT 21.105 127.820 21.275 128.790 ;
        RECT 21.445 128.160 21.615 129.290 ;
        RECT 21.785 128.500 21.955 129.300 ;
        RECT 22.155 129.180 22.435 129.350 ;
        RECT 22.160 128.700 22.435 129.180 ;
        RECT 22.605 128.500 22.795 129.860 ;
        RECT 22.975 129.495 23.485 130.030 ;
        RECT 23.705 129.220 23.950 129.825 ;
        RECT 25.315 129.305 25.605 130.030 ;
        RECT 26.785 129.550 27.085 130.030 ;
        RECT 27.255 129.380 27.515 129.835 ;
        RECT 27.685 129.550 27.945 130.030 ;
        RECT 28.125 129.380 28.385 129.835 ;
        RECT 28.555 129.550 28.805 130.030 ;
        RECT 28.985 129.380 29.245 129.835 ;
        RECT 29.415 129.550 29.665 130.030 ;
        RECT 29.845 129.380 30.105 129.835 ;
        RECT 30.275 129.550 30.520 130.030 ;
        RECT 30.690 129.380 30.965 129.835 ;
        RECT 31.135 129.550 31.380 130.030 ;
        RECT 31.550 129.380 31.810 129.835 ;
        RECT 31.980 129.550 32.240 130.030 ;
        RECT 32.410 129.380 32.670 129.835 ;
        RECT 32.840 129.550 33.100 130.030 ;
        RECT 33.270 129.380 33.530 129.835 ;
        RECT 33.700 129.470 33.960 130.030 ;
        RECT 26.785 129.350 33.530 129.380 ;
        RECT 22.995 129.050 24.225 129.220 ;
        RECT 26.755 129.210 33.530 129.350 ;
        RECT 26.755 129.180 27.950 129.210 ;
        RECT 21.785 128.330 22.795 128.500 ;
        RECT 22.965 128.485 23.715 128.675 ;
        RECT 21.445 127.990 22.570 128.160 ;
        RECT 22.965 127.820 23.135 128.485 ;
        RECT 23.885 128.240 24.225 129.050 ;
        RECT 21.105 127.650 23.135 127.820 ;
        RECT 23.305 127.480 23.475 128.240 ;
        RECT 23.710 127.830 24.225 128.240 ;
        RECT 25.315 127.480 25.605 128.645 ;
        RECT 26.785 128.620 27.950 129.180 ;
        RECT 34.130 129.040 34.380 129.850 ;
        RECT 34.560 129.505 34.820 130.030 ;
        RECT 34.990 129.040 35.240 129.850 ;
        RECT 35.420 129.520 35.725 130.030 ;
        RECT 35.895 129.355 36.155 129.860 ;
        RECT 36.335 129.650 36.665 130.030 ;
        RECT 36.845 129.480 37.015 129.860 ;
        RECT 28.120 128.790 35.240 129.040 ;
        RECT 35.410 128.790 35.725 129.350 ;
        RECT 26.785 128.395 33.530 128.620 ;
        RECT 26.785 127.480 27.055 128.225 ;
        RECT 27.225 127.655 27.515 128.395 ;
        RECT 28.125 128.380 33.530 128.395 ;
        RECT 27.685 127.485 27.940 128.210 ;
        RECT 28.125 127.655 28.385 128.380 ;
        RECT 28.555 127.485 28.800 128.210 ;
        RECT 28.985 127.655 29.245 128.380 ;
        RECT 29.415 127.485 29.660 128.210 ;
        RECT 29.845 127.655 30.105 128.380 ;
        RECT 30.275 127.485 30.520 128.210 ;
        RECT 30.690 127.655 30.950 128.380 ;
        RECT 31.120 127.485 31.380 128.210 ;
        RECT 31.550 127.655 31.810 128.380 ;
        RECT 31.980 127.485 32.240 128.210 ;
        RECT 32.410 127.655 32.670 128.380 ;
        RECT 32.840 127.485 33.100 128.210 ;
        RECT 33.270 127.655 33.530 128.380 ;
        RECT 33.700 127.485 33.960 128.280 ;
        RECT 34.130 127.655 34.380 128.790 ;
        RECT 27.685 127.480 33.960 127.485 ;
        RECT 34.560 127.480 34.820 128.290 ;
        RECT 34.995 127.650 35.240 128.790 ;
        RECT 35.895 128.555 36.065 129.355 ;
        RECT 36.350 129.310 37.015 129.480 ;
        RECT 36.350 129.055 36.520 129.310 ;
        RECT 37.550 129.220 37.795 129.825 ;
        RECT 38.015 129.495 38.525 130.030 ;
        RECT 36.235 128.725 36.520 129.055 ;
        RECT 36.755 128.760 37.085 129.130 ;
        RECT 37.275 129.050 38.505 129.220 ;
        RECT 36.350 128.580 36.520 128.725 ;
        RECT 35.420 127.480 35.715 128.290 ;
        RECT 35.895 127.650 36.165 128.555 ;
        RECT 36.350 128.410 37.015 128.580 ;
        RECT 36.335 127.480 36.665 128.240 ;
        RECT 36.845 127.650 37.015 128.410 ;
        RECT 37.275 128.240 37.615 129.050 ;
        RECT 37.785 128.485 38.535 128.675 ;
        RECT 37.275 127.830 37.790 128.240 ;
        RECT 38.025 127.480 38.195 128.240 ;
        RECT 38.365 127.820 38.535 128.485 ;
        RECT 38.705 128.500 38.895 129.860 ;
        RECT 39.065 129.010 39.340 129.860 ;
        RECT 39.530 129.495 40.060 129.860 ;
        RECT 40.485 129.630 40.815 130.030 ;
        RECT 39.885 129.460 40.060 129.495 ;
        RECT 39.065 128.840 39.345 129.010 ;
        RECT 39.065 128.700 39.340 128.840 ;
        RECT 39.545 128.500 39.715 129.300 ;
        RECT 38.705 128.330 39.715 128.500 ;
        RECT 39.885 129.290 40.815 129.460 ;
        RECT 40.985 129.290 41.240 129.860 ;
        RECT 41.415 129.520 41.720 130.030 ;
        RECT 39.885 128.160 40.055 129.290 ;
        RECT 40.645 129.120 40.815 129.290 ;
        RECT 38.930 127.990 40.055 128.160 ;
        RECT 40.225 128.790 40.420 129.120 ;
        RECT 40.645 128.790 40.900 129.120 ;
        RECT 40.225 127.820 40.395 128.790 ;
        RECT 41.070 128.620 41.240 129.290 ;
        RECT 41.415 128.790 41.730 129.350 ;
        RECT 41.900 129.040 42.150 129.850 ;
        RECT 42.320 129.505 42.580 130.030 ;
        RECT 42.760 129.040 43.010 129.850 ;
        RECT 43.180 129.470 43.440 130.030 ;
        RECT 43.610 129.380 43.870 129.835 ;
        RECT 44.040 129.550 44.300 130.030 ;
        RECT 44.470 129.380 44.730 129.835 ;
        RECT 44.900 129.550 45.160 130.030 ;
        RECT 45.330 129.380 45.590 129.835 ;
        RECT 45.760 129.550 46.005 130.030 ;
        RECT 46.175 129.380 46.450 129.835 ;
        RECT 46.620 129.550 46.865 130.030 ;
        RECT 47.035 129.380 47.295 129.835 ;
        RECT 47.475 129.550 47.725 130.030 ;
        RECT 47.895 129.380 48.155 129.835 ;
        RECT 48.335 129.550 48.585 130.030 ;
        RECT 48.755 129.380 49.015 129.835 ;
        RECT 49.195 129.550 49.455 130.030 ;
        RECT 49.625 129.380 49.885 129.835 ;
        RECT 50.055 129.550 50.355 130.030 ;
        RECT 43.610 129.210 50.355 129.380 ;
        RECT 51.075 129.305 51.365 130.030 ;
        RECT 51.535 129.260 53.205 130.030 ;
        RECT 53.750 129.690 54.005 129.850 ;
        RECT 53.665 129.520 54.005 129.690 ;
        RECT 54.185 129.570 54.470 130.030 ;
        RECT 41.900 128.790 49.020 129.040 ;
        RECT 38.365 127.650 40.395 127.820 ;
        RECT 40.565 127.480 40.735 128.620 ;
        RECT 40.905 127.650 41.240 128.620 ;
        RECT 41.425 127.480 41.720 128.290 ;
        RECT 41.900 127.650 42.145 128.790 ;
        RECT 42.320 127.480 42.580 128.290 ;
        RECT 42.760 127.655 43.010 128.790 ;
        RECT 49.190 128.620 50.355 129.210 ;
        RECT 43.610 128.395 50.355 128.620 ;
        RECT 43.610 128.380 49.015 128.395 ;
        RECT 43.180 127.485 43.440 128.280 ;
        RECT 43.610 127.655 43.870 128.380 ;
        RECT 44.040 127.485 44.300 128.210 ;
        RECT 44.470 127.655 44.730 128.380 ;
        RECT 44.900 127.485 45.160 128.210 ;
        RECT 45.330 127.655 45.590 128.380 ;
        RECT 45.760 127.485 46.020 128.210 ;
        RECT 46.190 127.655 46.450 128.380 ;
        RECT 46.620 127.485 46.865 128.210 ;
        RECT 47.035 127.655 47.295 128.380 ;
        RECT 47.480 127.485 47.725 128.210 ;
        RECT 47.895 127.655 48.155 128.380 ;
        RECT 48.340 127.485 48.585 128.210 ;
        RECT 48.755 127.655 49.015 128.380 ;
        RECT 49.200 127.485 49.455 128.210 ;
        RECT 49.625 127.655 49.915 128.395 ;
        RECT 43.180 127.480 49.455 127.485 ;
        RECT 50.085 127.480 50.355 128.225 ;
        RECT 51.075 127.480 51.365 128.645 ;
        RECT 51.535 128.570 52.285 129.090 ;
        RECT 52.455 128.740 53.205 129.260 ;
        RECT 53.750 129.320 54.005 129.520 ;
        RECT 51.535 127.480 53.205 128.570 ;
        RECT 53.750 128.460 53.930 129.320 ;
        RECT 54.650 129.120 54.900 129.770 ;
        RECT 54.100 128.790 54.900 129.120 ;
        RECT 53.750 127.790 54.005 128.460 ;
        RECT 54.185 127.480 54.470 128.280 ;
        RECT 54.650 128.200 54.900 128.790 ;
        RECT 55.100 129.435 55.420 129.765 ;
        RECT 55.600 129.550 56.260 130.030 ;
        RECT 56.460 129.640 57.310 129.810 ;
        RECT 55.100 128.540 55.290 129.435 ;
        RECT 55.610 129.110 56.270 129.380 ;
        RECT 55.940 129.050 56.270 129.110 ;
        RECT 55.460 128.880 55.790 128.940 ;
        RECT 56.460 128.880 56.630 129.640 ;
        RECT 57.870 129.570 58.190 130.030 ;
        RECT 58.390 129.390 58.640 129.820 ;
        RECT 58.930 129.590 59.340 130.030 ;
        RECT 59.510 129.650 60.525 129.850 ;
        RECT 56.800 129.220 58.050 129.390 ;
        RECT 56.800 129.100 57.130 129.220 ;
        RECT 55.460 128.710 57.360 128.880 ;
        RECT 55.100 128.370 57.020 128.540 ;
        RECT 55.100 128.350 55.420 128.370 ;
        RECT 54.650 127.690 54.980 128.200 ;
        RECT 55.250 127.740 55.420 128.350 ;
        RECT 57.190 128.200 57.360 128.710 ;
        RECT 57.530 128.640 57.710 129.050 ;
        RECT 57.880 128.460 58.050 129.220 ;
        RECT 55.590 127.480 55.920 128.170 ;
        RECT 56.150 128.030 57.360 128.200 ;
        RECT 57.530 128.150 58.050 128.460 ;
        RECT 58.220 129.050 58.640 129.390 ;
        RECT 58.930 129.050 59.340 129.380 ;
        RECT 58.220 128.280 58.410 129.050 ;
        RECT 59.510 128.920 59.680 129.650 ;
        RECT 60.825 129.480 60.995 129.810 ;
        RECT 61.165 129.650 61.495 130.030 ;
        RECT 59.850 129.100 60.200 129.470 ;
        RECT 59.510 128.880 59.930 128.920 ;
        RECT 58.580 128.710 59.930 128.880 ;
        RECT 58.580 128.550 58.830 128.710 ;
        RECT 59.340 128.280 59.590 128.540 ;
        RECT 58.220 128.030 59.590 128.280 ;
        RECT 56.150 127.740 56.390 128.030 ;
        RECT 57.190 127.950 57.360 128.030 ;
        RECT 56.590 127.480 57.010 127.860 ;
        RECT 57.190 127.700 57.820 127.950 ;
        RECT 58.290 127.480 58.620 127.860 ;
        RECT 58.790 127.740 58.960 128.030 ;
        RECT 59.760 127.865 59.930 128.710 ;
        RECT 60.380 128.540 60.600 129.410 ;
        RECT 60.825 129.290 61.520 129.480 ;
        RECT 60.100 128.160 60.600 128.540 ;
        RECT 60.770 128.490 61.180 129.110 ;
        RECT 61.350 128.320 61.520 129.290 ;
        RECT 60.825 128.150 61.520 128.320 ;
        RECT 59.140 127.480 59.520 127.860 ;
        RECT 59.760 127.695 60.590 127.865 ;
        RECT 60.825 127.650 60.995 128.150 ;
        RECT 61.165 127.480 61.495 127.980 ;
        RECT 61.710 127.650 61.935 129.770 ;
        RECT 62.105 129.650 62.435 130.030 ;
        RECT 62.605 129.480 62.775 129.770 ;
        RECT 63.095 129.550 63.375 130.030 ;
        RECT 62.110 129.310 62.775 129.480 ;
        RECT 63.545 129.380 63.805 129.770 ;
        RECT 63.980 129.550 64.235 130.030 ;
        RECT 64.405 129.380 64.700 129.770 ;
        RECT 64.880 129.550 65.155 130.030 ;
        RECT 65.325 129.530 65.625 129.860 ;
        RECT 62.110 128.320 62.340 129.310 ;
        RECT 63.050 129.210 64.700 129.380 ;
        RECT 62.510 128.490 62.860 129.140 ;
        RECT 63.050 128.700 63.455 129.210 ;
        RECT 63.625 128.870 64.765 129.040 ;
        RECT 63.050 128.530 63.805 128.700 ;
        RECT 62.110 128.150 62.775 128.320 ;
        RECT 62.105 127.480 62.435 127.980 ;
        RECT 62.605 127.650 62.775 128.150 ;
        RECT 63.090 127.480 63.375 128.350 ;
        RECT 63.545 128.280 63.805 128.530 ;
        RECT 64.595 128.620 64.765 128.870 ;
        RECT 64.935 128.790 65.285 129.360 ;
        RECT 65.455 128.620 65.625 129.530 ;
        RECT 64.595 128.450 65.625 128.620 ;
        RECT 63.545 128.110 64.665 128.280 ;
        RECT 63.545 127.650 63.805 128.110 ;
        RECT 63.980 127.480 64.235 127.940 ;
        RECT 64.405 127.650 64.665 128.110 ;
        RECT 64.835 127.480 65.145 128.280 ;
        RECT 65.315 127.650 65.625 128.450 ;
        RECT 65.795 129.530 66.095 129.860 ;
        RECT 66.265 129.550 66.540 130.030 ;
        RECT 65.795 128.620 65.965 129.530 ;
        RECT 66.720 129.380 67.015 129.770 ;
        RECT 67.185 129.550 67.440 130.030 ;
        RECT 67.615 129.380 67.875 129.770 ;
        RECT 68.045 129.550 68.325 130.030 ;
        RECT 66.135 128.790 66.485 129.360 ;
        RECT 66.720 129.210 68.370 129.380 ;
        RECT 68.555 129.260 70.225 130.030 ;
        RECT 66.655 128.870 67.795 129.040 ;
        RECT 66.655 128.620 66.825 128.870 ;
        RECT 67.965 128.700 68.370 129.210 ;
        RECT 65.795 128.450 66.825 128.620 ;
        RECT 67.615 128.530 68.370 128.700 ;
        RECT 68.555 128.570 69.305 129.090 ;
        RECT 69.475 128.740 70.225 129.260 ;
        RECT 70.395 129.570 70.955 129.860 ;
        RECT 71.125 129.570 71.375 130.030 ;
        RECT 65.795 127.650 66.105 128.450 ;
        RECT 67.615 128.280 67.875 128.530 ;
        RECT 66.275 127.480 66.585 128.280 ;
        RECT 66.755 128.110 67.875 128.280 ;
        RECT 66.755 127.650 67.015 128.110 ;
        RECT 67.185 127.480 67.440 127.940 ;
        RECT 67.615 127.650 67.875 128.110 ;
        RECT 68.045 127.480 68.330 128.350 ;
        RECT 68.555 127.480 70.225 128.570 ;
        RECT 70.395 128.200 70.645 129.570 ;
        RECT 71.995 129.400 72.325 129.760 ;
        RECT 70.935 129.210 72.325 129.400 ;
        RECT 72.970 129.220 73.215 129.825 ;
        RECT 73.435 129.495 73.945 130.030 ;
        RECT 70.935 129.120 71.105 129.210 ;
        RECT 70.815 128.790 71.105 129.120 ;
        RECT 72.695 129.050 73.925 129.220 ;
        RECT 71.275 128.790 71.615 129.040 ;
        RECT 71.835 128.790 72.510 129.040 ;
        RECT 70.935 128.540 71.105 128.790 ;
        RECT 70.935 128.370 71.875 128.540 ;
        RECT 72.245 128.430 72.510 128.790 ;
        RECT 70.395 127.650 70.855 128.200 ;
        RECT 71.045 127.480 71.375 128.200 ;
        RECT 71.575 127.820 71.875 128.370 ;
        RECT 72.695 128.240 73.035 129.050 ;
        RECT 73.205 128.485 73.955 128.675 ;
        RECT 72.045 127.480 72.325 128.150 ;
        RECT 72.695 127.830 73.210 128.240 ;
        RECT 73.445 127.480 73.615 128.240 ;
        RECT 73.785 127.820 73.955 128.485 ;
        RECT 74.125 128.500 74.315 129.860 ;
        RECT 74.485 129.690 74.760 129.860 ;
        RECT 74.485 129.520 74.765 129.690 ;
        RECT 74.485 128.700 74.760 129.520 ;
        RECT 74.950 129.495 75.480 129.860 ;
        RECT 75.905 129.630 76.235 130.030 ;
        RECT 75.305 129.460 75.480 129.495 ;
        RECT 74.965 128.500 75.135 129.300 ;
        RECT 74.125 128.330 75.135 128.500 ;
        RECT 75.305 129.290 76.235 129.460 ;
        RECT 76.405 129.290 76.660 129.860 ;
        RECT 76.835 129.305 77.125 130.030 ;
        RECT 77.295 129.570 77.855 129.860 ;
        RECT 78.025 129.570 78.275 130.030 ;
        RECT 75.305 128.160 75.475 129.290 ;
        RECT 76.065 129.120 76.235 129.290 ;
        RECT 74.350 127.990 75.475 128.160 ;
        RECT 75.645 128.790 75.840 129.120 ;
        RECT 76.065 128.790 76.320 129.120 ;
        RECT 75.645 127.820 75.815 128.790 ;
        RECT 76.490 128.620 76.660 129.290 ;
        RECT 73.785 127.650 75.815 127.820 ;
        RECT 75.985 127.480 76.155 128.620 ;
        RECT 76.325 127.650 76.660 128.620 ;
        RECT 76.835 127.480 77.125 128.645 ;
        RECT 77.295 128.200 77.545 129.570 ;
        RECT 78.895 129.400 79.225 129.760 ;
        RECT 77.835 129.210 79.225 129.400 ;
        RECT 79.595 129.260 83.105 130.030 ;
        RECT 83.365 129.480 83.535 129.770 ;
        RECT 83.705 129.650 84.035 130.030 ;
        RECT 83.365 129.310 84.030 129.480 ;
        RECT 77.835 129.120 78.005 129.210 ;
        RECT 77.715 128.790 78.005 129.120 ;
        RECT 78.175 128.790 78.515 129.040 ;
        RECT 78.735 128.790 79.410 129.040 ;
        RECT 77.835 128.540 78.005 128.790 ;
        RECT 77.835 128.370 78.775 128.540 ;
        RECT 79.145 128.430 79.410 128.790 ;
        RECT 79.595 128.570 81.285 129.090 ;
        RECT 81.455 128.740 83.105 129.260 ;
        RECT 77.295 127.650 77.755 128.200 ;
        RECT 77.945 127.480 78.275 128.200 ;
        RECT 78.475 127.820 78.775 128.370 ;
        RECT 78.945 127.480 79.225 128.150 ;
        RECT 79.595 127.480 83.105 128.570 ;
        RECT 83.280 128.490 83.630 129.140 ;
        RECT 83.800 128.320 84.030 129.310 ;
        RECT 83.365 128.150 84.030 128.320 ;
        RECT 83.365 127.650 83.535 128.150 ;
        RECT 83.705 127.480 84.035 127.980 ;
        RECT 84.205 127.650 84.430 129.770 ;
        RECT 84.645 129.650 84.975 130.030 ;
        RECT 85.145 129.480 85.315 129.810 ;
        RECT 85.615 129.650 86.630 129.850 ;
        RECT 84.620 129.290 85.315 129.480 ;
        RECT 84.620 128.320 84.790 129.290 ;
        RECT 84.960 128.490 85.370 129.110 ;
        RECT 85.540 128.540 85.760 129.410 ;
        RECT 85.940 129.100 86.290 129.470 ;
        RECT 86.460 128.920 86.630 129.650 ;
        RECT 86.800 129.590 87.210 130.030 ;
        RECT 87.500 129.390 87.750 129.820 ;
        RECT 87.950 129.570 88.270 130.030 ;
        RECT 88.830 129.640 89.680 129.810 ;
        RECT 86.800 129.050 87.210 129.380 ;
        RECT 87.500 129.050 87.920 129.390 ;
        RECT 86.210 128.880 86.630 128.920 ;
        RECT 86.210 128.710 87.560 128.880 ;
        RECT 84.620 128.150 85.315 128.320 ;
        RECT 85.540 128.160 86.040 128.540 ;
        RECT 84.645 127.480 84.975 127.980 ;
        RECT 85.145 127.650 85.315 128.150 ;
        RECT 86.210 127.865 86.380 128.710 ;
        RECT 87.310 128.550 87.560 128.710 ;
        RECT 86.550 128.280 86.800 128.540 ;
        RECT 87.730 128.280 87.920 129.050 ;
        RECT 86.550 128.030 87.920 128.280 ;
        RECT 88.090 129.220 89.340 129.390 ;
        RECT 88.090 128.460 88.260 129.220 ;
        RECT 89.010 129.100 89.340 129.220 ;
        RECT 88.430 128.640 88.610 129.050 ;
        RECT 89.510 128.880 89.680 129.640 ;
        RECT 89.880 129.550 90.540 130.030 ;
        RECT 90.720 129.435 91.040 129.765 ;
        RECT 89.870 129.110 90.530 129.380 ;
        RECT 89.870 129.050 90.200 129.110 ;
        RECT 90.350 128.880 90.680 128.940 ;
        RECT 88.780 128.710 90.680 128.880 ;
        RECT 88.090 128.150 88.610 128.460 ;
        RECT 88.780 128.200 88.950 128.710 ;
        RECT 90.850 128.540 91.040 129.435 ;
        RECT 89.120 128.370 91.040 128.540 ;
        RECT 90.720 128.350 91.040 128.370 ;
        RECT 91.240 129.120 91.490 129.770 ;
        RECT 91.670 129.570 91.955 130.030 ;
        RECT 92.135 129.350 92.390 129.850 ;
        RECT 92.135 129.320 92.475 129.350 ;
        RECT 92.210 129.180 92.475 129.320 ;
        RECT 92.935 129.260 94.605 130.030 ;
        RECT 91.240 128.790 92.040 129.120 ;
        RECT 88.780 128.030 89.990 128.200 ;
        RECT 85.550 127.695 86.380 127.865 ;
        RECT 86.620 127.480 87.000 127.860 ;
        RECT 87.180 127.740 87.350 128.030 ;
        RECT 88.780 127.950 88.950 128.030 ;
        RECT 87.520 127.480 87.850 127.860 ;
        RECT 88.320 127.700 88.950 127.950 ;
        RECT 89.130 127.480 89.550 127.860 ;
        RECT 89.750 127.740 89.990 128.030 ;
        RECT 90.220 127.480 90.550 128.170 ;
        RECT 90.720 127.740 90.890 128.350 ;
        RECT 91.240 128.200 91.490 128.790 ;
        RECT 92.210 128.460 92.390 129.180 ;
        RECT 91.160 127.690 91.490 128.200 ;
        RECT 91.670 127.480 91.955 128.280 ;
        RECT 92.135 127.790 92.390 128.460 ;
        RECT 92.935 128.570 93.685 129.090 ;
        RECT 93.855 128.740 94.605 129.260 ;
        RECT 94.775 129.570 95.335 129.860 ;
        RECT 95.505 129.570 95.755 130.030 ;
        RECT 92.935 127.480 94.605 128.570 ;
        RECT 94.775 128.200 95.025 129.570 ;
        RECT 96.375 129.400 96.705 129.760 ;
        RECT 95.315 129.210 96.705 129.400 ;
        RECT 97.075 129.280 98.285 130.030 ;
        RECT 95.315 129.120 95.485 129.210 ;
        RECT 95.195 128.790 95.485 129.120 ;
        RECT 95.655 128.790 95.995 129.040 ;
        RECT 96.215 128.790 96.890 129.040 ;
        RECT 95.315 128.540 95.485 128.790 ;
        RECT 95.315 128.370 96.255 128.540 ;
        RECT 96.625 128.430 96.890 128.790 ;
        RECT 97.075 128.570 97.595 129.110 ;
        RECT 97.765 128.740 98.285 129.280 ;
        RECT 98.730 129.220 98.975 129.825 ;
        RECT 99.195 129.495 99.705 130.030 ;
        RECT 98.455 129.050 99.685 129.220 ;
        RECT 94.775 127.650 95.235 128.200 ;
        RECT 95.425 127.480 95.755 128.200 ;
        RECT 95.955 127.820 96.255 128.370 ;
        RECT 96.425 127.480 96.705 128.150 ;
        RECT 97.075 127.480 98.285 128.570 ;
        RECT 98.455 128.240 98.795 129.050 ;
        RECT 98.965 128.485 99.715 128.675 ;
        RECT 98.455 127.830 98.970 128.240 ;
        RECT 99.205 127.480 99.375 128.240 ;
        RECT 99.545 127.820 99.715 128.485 ;
        RECT 99.885 128.500 100.075 129.860 ;
        RECT 100.245 129.010 100.520 129.860 ;
        RECT 100.710 129.495 101.240 129.860 ;
        RECT 101.665 129.630 101.995 130.030 ;
        RECT 101.065 129.460 101.240 129.495 ;
        RECT 100.245 128.840 100.525 129.010 ;
        RECT 100.245 128.700 100.520 128.840 ;
        RECT 100.725 128.500 100.895 129.300 ;
        RECT 99.885 128.330 100.895 128.500 ;
        RECT 101.065 129.290 101.995 129.460 ;
        RECT 102.165 129.290 102.420 129.860 ;
        RECT 102.595 129.305 102.885 130.030 ;
        RECT 101.065 128.160 101.235 129.290 ;
        RECT 101.825 129.120 101.995 129.290 ;
        RECT 100.110 127.990 101.235 128.160 ;
        RECT 101.405 128.790 101.600 129.120 ;
        RECT 101.825 128.790 102.080 129.120 ;
        RECT 101.405 127.820 101.575 128.790 ;
        RECT 102.250 128.620 102.420 129.290 ;
        RECT 103.575 129.210 103.785 130.030 ;
        RECT 103.955 129.230 104.285 129.860 ;
        RECT 99.545 127.650 101.575 127.820 ;
        RECT 101.745 127.480 101.915 128.620 ;
        RECT 102.085 127.650 102.420 128.620 ;
        RECT 102.595 127.480 102.885 128.645 ;
        RECT 103.955 128.630 104.205 129.230 ;
        RECT 104.455 129.210 104.685 130.030 ;
        RECT 105.270 129.320 105.525 129.850 ;
        RECT 105.705 129.570 105.990 130.030 ;
        RECT 104.375 128.790 104.705 129.040 ;
        RECT 103.575 127.480 103.785 128.620 ;
        RECT 103.955 127.650 104.285 128.630 ;
        RECT 104.455 127.480 104.685 128.620 ;
        RECT 105.270 128.460 105.450 129.320 ;
        RECT 106.170 129.120 106.420 129.770 ;
        RECT 105.620 128.790 106.420 129.120 ;
        RECT 105.270 128.330 105.525 128.460 ;
        RECT 105.185 128.160 105.525 128.330 ;
        RECT 105.270 127.790 105.525 128.160 ;
        RECT 105.705 127.480 105.990 128.280 ;
        RECT 106.170 128.200 106.420 128.790 ;
        RECT 106.620 129.435 106.940 129.765 ;
        RECT 107.120 129.550 107.780 130.030 ;
        RECT 107.980 129.640 108.830 129.810 ;
        RECT 106.620 128.540 106.810 129.435 ;
        RECT 107.130 129.110 107.790 129.380 ;
        RECT 107.460 129.050 107.790 129.110 ;
        RECT 106.980 128.880 107.310 128.940 ;
        RECT 107.980 128.880 108.150 129.640 ;
        RECT 109.390 129.570 109.710 130.030 ;
        RECT 109.910 129.390 110.160 129.820 ;
        RECT 110.450 129.590 110.860 130.030 ;
        RECT 111.030 129.650 112.045 129.850 ;
        RECT 108.320 129.220 109.570 129.390 ;
        RECT 108.320 129.100 108.650 129.220 ;
        RECT 106.980 128.710 108.880 128.880 ;
        RECT 106.620 128.370 108.540 128.540 ;
        RECT 106.620 128.350 106.940 128.370 ;
        RECT 106.170 127.690 106.500 128.200 ;
        RECT 106.770 127.740 106.940 128.350 ;
        RECT 108.710 128.200 108.880 128.710 ;
        RECT 109.050 128.640 109.230 129.050 ;
        RECT 109.400 128.460 109.570 129.220 ;
        RECT 107.110 127.480 107.440 128.170 ;
        RECT 107.670 128.030 108.880 128.200 ;
        RECT 109.050 128.150 109.570 128.460 ;
        RECT 109.740 129.050 110.160 129.390 ;
        RECT 110.450 129.050 110.860 129.380 ;
        RECT 109.740 128.280 109.930 129.050 ;
        RECT 111.030 128.920 111.200 129.650 ;
        RECT 112.345 129.480 112.515 129.810 ;
        RECT 112.685 129.650 113.015 130.030 ;
        RECT 111.370 129.100 111.720 129.470 ;
        RECT 111.030 128.880 111.450 128.920 ;
        RECT 110.100 128.710 111.450 128.880 ;
        RECT 110.100 128.550 110.350 128.710 ;
        RECT 110.860 128.280 111.110 128.540 ;
        RECT 109.740 128.030 111.110 128.280 ;
        RECT 107.670 127.740 107.910 128.030 ;
        RECT 108.710 127.950 108.880 128.030 ;
        RECT 108.110 127.480 108.530 127.860 ;
        RECT 108.710 127.700 109.340 127.950 ;
        RECT 109.810 127.480 110.140 127.860 ;
        RECT 110.310 127.740 110.480 128.030 ;
        RECT 111.280 127.865 111.450 128.710 ;
        RECT 111.900 128.540 112.120 129.410 ;
        RECT 112.345 129.290 113.040 129.480 ;
        RECT 111.620 128.160 112.120 128.540 ;
        RECT 112.290 128.490 112.700 129.110 ;
        RECT 112.870 128.320 113.040 129.290 ;
        RECT 112.345 128.150 113.040 128.320 ;
        RECT 110.660 127.480 111.040 127.860 ;
        RECT 111.280 127.695 112.110 127.865 ;
        RECT 112.345 127.650 112.515 128.150 ;
        RECT 112.685 127.480 113.015 127.980 ;
        RECT 113.230 127.650 113.455 129.770 ;
        RECT 113.625 129.650 113.955 130.030 ;
        RECT 114.125 129.480 114.295 129.770 ;
        RECT 113.630 129.310 114.295 129.480 ;
        RECT 113.630 128.320 113.860 129.310 ;
        RECT 114.555 129.280 115.765 130.030 ;
        RECT 114.030 128.490 114.380 129.140 ;
        RECT 114.555 128.570 115.075 129.110 ;
        RECT 115.245 128.740 115.765 129.280 ;
        RECT 113.630 128.150 114.295 128.320 ;
        RECT 113.625 127.480 113.955 127.980 ;
        RECT 114.125 127.650 114.295 128.150 ;
        RECT 114.555 127.480 115.765 128.570 ;
        RECT 14.650 127.310 115.850 127.480 ;
        RECT 14.735 126.220 15.945 127.310 ;
        RECT 14.735 125.510 15.255 126.050 ;
        RECT 15.425 125.680 15.945 126.220 ;
        RECT 16.950 126.330 17.205 127.000 ;
        RECT 17.385 126.510 17.670 127.310 ;
        RECT 17.850 126.590 18.180 127.100 ;
        RECT 14.735 124.760 15.945 125.510 ;
        RECT 16.950 125.470 17.130 126.330 ;
        RECT 17.850 126.000 18.100 126.590 ;
        RECT 18.450 126.440 18.620 127.050 ;
        RECT 18.790 126.620 19.120 127.310 ;
        RECT 19.350 126.760 19.590 127.050 ;
        RECT 19.790 126.930 20.210 127.310 ;
        RECT 20.390 126.840 21.020 127.090 ;
        RECT 21.490 126.930 21.820 127.310 ;
        RECT 20.390 126.760 20.560 126.840 ;
        RECT 21.990 126.760 22.160 127.050 ;
        RECT 22.340 126.930 22.720 127.310 ;
        RECT 22.960 126.925 23.790 127.095 ;
        RECT 19.350 126.590 20.560 126.760 ;
        RECT 17.300 125.670 18.100 126.000 ;
        RECT 16.950 125.270 17.205 125.470 ;
        RECT 16.865 125.100 17.205 125.270 ;
        RECT 16.950 124.940 17.205 125.100 ;
        RECT 17.385 124.760 17.670 125.220 ;
        RECT 17.850 125.020 18.100 125.670 ;
        RECT 18.300 126.420 18.620 126.440 ;
        RECT 18.300 126.250 20.220 126.420 ;
        RECT 18.300 125.355 18.490 126.250 ;
        RECT 20.390 126.080 20.560 126.590 ;
        RECT 20.730 126.330 21.250 126.640 ;
        RECT 18.660 125.910 20.560 126.080 ;
        RECT 18.660 125.850 18.990 125.910 ;
        RECT 19.140 125.680 19.470 125.740 ;
        RECT 18.810 125.410 19.470 125.680 ;
        RECT 18.300 125.025 18.620 125.355 ;
        RECT 18.800 124.760 19.460 125.240 ;
        RECT 19.660 125.150 19.830 125.910 ;
        RECT 20.730 125.740 20.910 126.150 ;
        RECT 20.000 125.570 20.330 125.690 ;
        RECT 21.080 125.570 21.250 126.330 ;
        RECT 20.000 125.400 21.250 125.570 ;
        RECT 21.420 126.510 22.790 126.760 ;
        RECT 21.420 125.740 21.610 126.510 ;
        RECT 22.540 126.250 22.790 126.510 ;
        RECT 21.780 126.080 22.030 126.240 ;
        RECT 22.960 126.080 23.130 126.925 ;
        RECT 24.025 126.640 24.195 127.140 ;
        RECT 24.365 126.810 24.695 127.310 ;
        RECT 23.300 126.250 23.800 126.630 ;
        RECT 24.025 126.470 24.720 126.640 ;
        RECT 21.780 125.910 23.130 126.080 ;
        RECT 22.710 125.870 23.130 125.910 ;
        RECT 21.420 125.400 21.840 125.740 ;
        RECT 22.130 125.410 22.540 125.740 ;
        RECT 19.660 124.980 20.510 125.150 ;
        RECT 21.070 124.760 21.390 125.220 ;
        RECT 21.590 124.970 21.840 125.400 ;
        RECT 22.130 124.760 22.540 125.200 ;
        RECT 22.710 125.140 22.880 125.870 ;
        RECT 23.050 125.320 23.400 125.690 ;
        RECT 23.580 125.380 23.800 126.250 ;
        RECT 23.970 125.680 24.380 126.300 ;
        RECT 24.550 125.500 24.720 126.470 ;
        RECT 24.025 125.310 24.720 125.500 ;
        RECT 22.710 124.940 23.725 125.140 ;
        RECT 24.025 124.980 24.195 125.310 ;
        RECT 24.365 124.760 24.695 125.140 ;
        RECT 24.910 125.020 25.135 127.140 ;
        RECT 25.305 126.810 25.635 127.310 ;
        RECT 25.805 126.640 25.975 127.140 ;
        RECT 25.310 126.470 25.975 126.640 ;
        RECT 25.310 125.480 25.540 126.470 ;
        RECT 25.710 125.650 26.060 126.300 ;
        RECT 27.155 126.235 27.425 127.140 ;
        RECT 27.595 126.550 27.925 127.310 ;
        RECT 28.105 126.380 28.275 127.140 ;
        RECT 28.625 126.640 28.795 127.140 ;
        RECT 28.965 126.810 29.295 127.310 ;
        RECT 28.625 126.470 29.290 126.640 ;
        RECT 25.310 125.310 25.975 125.480 ;
        RECT 25.305 124.760 25.635 125.140 ;
        RECT 25.805 125.020 25.975 125.310 ;
        RECT 27.155 125.435 27.325 126.235 ;
        RECT 27.610 126.210 28.275 126.380 ;
        RECT 27.610 126.065 27.780 126.210 ;
        RECT 27.495 125.735 27.780 126.065 ;
        RECT 27.610 125.480 27.780 125.735 ;
        RECT 28.015 125.660 28.345 126.030 ;
        RECT 28.540 125.650 28.890 126.300 ;
        RECT 29.060 125.480 29.290 126.470 ;
        RECT 27.155 124.930 27.415 125.435 ;
        RECT 27.610 125.310 28.275 125.480 ;
        RECT 27.595 124.760 27.925 125.140 ;
        RECT 28.105 124.930 28.275 125.310 ;
        RECT 28.625 125.310 29.290 125.480 ;
        RECT 28.625 125.020 28.795 125.310 ;
        RECT 28.965 124.760 29.295 125.140 ;
        RECT 29.465 125.020 29.690 127.140 ;
        RECT 29.905 126.810 30.235 127.310 ;
        RECT 30.405 126.640 30.575 127.140 ;
        RECT 30.810 126.925 31.640 127.095 ;
        RECT 31.880 126.930 32.260 127.310 ;
        RECT 29.880 126.470 30.575 126.640 ;
        RECT 29.880 125.500 30.050 126.470 ;
        RECT 30.220 125.680 30.630 126.300 ;
        RECT 30.800 126.250 31.300 126.630 ;
        RECT 29.880 125.310 30.575 125.500 ;
        RECT 30.800 125.380 31.020 126.250 ;
        RECT 31.470 126.080 31.640 126.925 ;
        RECT 32.440 126.760 32.610 127.050 ;
        RECT 32.780 126.930 33.110 127.310 ;
        RECT 33.580 126.840 34.210 127.090 ;
        RECT 34.390 126.930 34.810 127.310 ;
        RECT 34.040 126.760 34.210 126.840 ;
        RECT 35.010 126.760 35.250 127.050 ;
        RECT 31.810 126.510 33.180 126.760 ;
        RECT 31.810 126.250 32.060 126.510 ;
        RECT 32.570 126.080 32.820 126.240 ;
        RECT 31.470 125.910 32.820 126.080 ;
        RECT 31.470 125.870 31.890 125.910 ;
        RECT 31.200 125.320 31.550 125.690 ;
        RECT 29.905 124.760 30.235 125.140 ;
        RECT 30.405 124.980 30.575 125.310 ;
        RECT 31.720 125.140 31.890 125.870 ;
        RECT 32.990 125.740 33.180 126.510 ;
        RECT 32.060 125.410 32.470 125.740 ;
        RECT 32.760 125.400 33.180 125.740 ;
        RECT 33.350 126.330 33.870 126.640 ;
        RECT 34.040 126.590 35.250 126.760 ;
        RECT 35.480 126.620 35.810 127.310 ;
        RECT 33.350 125.570 33.520 126.330 ;
        RECT 33.690 125.740 33.870 126.150 ;
        RECT 34.040 126.080 34.210 126.590 ;
        RECT 35.980 126.440 36.150 127.050 ;
        RECT 36.420 126.590 36.750 127.100 ;
        RECT 35.980 126.420 36.300 126.440 ;
        RECT 34.380 126.250 36.300 126.420 ;
        RECT 34.040 125.910 35.940 126.080 ;
        RECT 34.270 125.570 34.600 125.690 ;
        RECT 33.350 125.400 34.600 125.570 ;
        RECT 30.875 124.940 31.890 125.140 ;
        RECT 32.060 124.760 32.470 125.200 ;
        RECT 32.760 124.970 33.010 125.400 ;
        RECT 33.210 124.760 33.530 125.220 ;
        RECT 34.770 125.150 34.940 125.910 ;
        RECT 35.610 125.850 35.940 125.910 ;
        RECT 35.130 125.680 35.460 125.740 ;
        RECT 35.130 125.410 35.790 125.680 ;
        RECT 36.110 125.355 36.300 126.250 ;
        RECT 34.090 124.980 34.940 125.150 ;
        RECT 35.140 124.760 35.800 125.240 ;
        RECT 35.980 125.025 36.300 125.355 ;
        RECT 36.500 126.000 36.750 126.590 ;
        RECT 36.930 126.510 37.215 127.310 ;
        RECT 37.395 126.970 37.650 127.000 ;
        RECT 37.395 126.800 37.735 126.970 ;
        RECT 37.395 126.330 37.650 126.800 ;
        RECT 36.500 125.670 37.300 126.000 ;
        RECT 36.500 125.020 36.750 125.670 ;
        RECT 37.470 125.470 37.650 126.330 ;
        RECT 38.195 126.145 38.485 127.310 ;
        RECT 39.685 126.510 39.855 127.310 ;
        RECT 40.025 126.290 40.355 127.140 ;
        RECT 40.525 126.510 40.695 127.310 ;
        RECT 40.865 126.290 41.195 127.140 ;
        RECT 41.365 126.510 41.535 127.310 ;
        RECT 41.705 126.290 42.035 127.140 ;
        RECT 42.205 126.510 42.375 127.310 ;
        RECT 42.545 126.290 42.875 127.140 ;
        RECT 43.045 126.510 43.215 127.310 ;
        RECT 43.385 126.290 43.715 127.140 ;
        RECT 43.885 126.510 44.055 127.310 ;
        RECT 44.225 126.290 44.555 127.140 ;
        RECT 44.725 126.510 44.895 127.310 ;
        RECT 45.065 126.290 45.395 127.140 ;
        RECT 45.565 126.510 45.735 127.310 ;
        RECT 45.905 126.290 46.235 127.140 ;
        RECT 46.405 126.510 46.575 127.310 ;
        RECT 46.745 126.290 47.075 127.140 ;
        RECT 47.245 126.510 47.415 127.310 ;
        RECT 47.585 126.290 47.915 127.140 ;
        RECT 48.085 126.510 48.255 127.310 ;
        RECT 48.425 126.290 48.755 127.140 ;
        RECT 48.925 126.460 49.095 127.310 ;
        RECT 49.265 126.290 49.595 127.140 ;
        RECT 49.765 126.460 49.935 127.310 ;
        RECT 50.105 126.290 50.435 127.140 ;
        RECT 39.575 126.120 46.235 126.290 ;
        RECT 46.405 126.120 48.755 126.290 ;
        RECT 48.925 126.120 50.435 126.290 ;
        RECT 50.615 126.590 51.075 127.140 ;
        RECT 51.265 126.590 51.595 127.310 ;
        RECT 39.575 125.580 39.850 126.120 ;
        RECT 46.405 125.950 46.580 126.120 ;
        RECT 48.925 125.950 49.095 126.120 ;
        RECT 40.020 125.750 46.580 125.950 ;
        RECT 46.785 125.750 49.095 125.950 ;
        RECT 49.265 125.750 50.440 125.950 ;
        RECT 46.405 125.580 46.580 125.750 ;
        RECT 48.925 125.580 49.095 125.750 ;
        RECT 36.930 124.760 37.215 125.220 ;
        RECT 37.395 124.940 37.650 125.470 ;
        RECT 38.195 124.760 38.485 125.485 ;
        RECT 39.575 125.410 46.235 125.580 ;
        RECT 46.405 125.410 48.755 125.580 ;
        RECT 48.925 125.410 50.435 125.580 ;
        RECT 39.685 124.760 39.855 125.240 ;
        RECT 40.025 124.935 40.355 125.410 ;
        RECT 40.525 124.760 40.695 125.240 ;
        RECT 40.865 124.935 41.195 125.410 ;
        RECT 41.365 124.760 41.535 125.240 ;
        RECT 41.705 124.935 42.035 125.410 ;
        RECT 42.205 124.760 42.375 125.240 ;
        RECT 42.545 124.935 42.875 125.410 ;
        RECT 43.045 124.760 43.215 125.240 ;
        RECT 43.385 124.935 43.715 125.410 ;
        RECT 43.885 124.760 44.055 125.240 ;
        RECT 44.225 124.935 44.555 125.410 ;
        RECT 44.305 124.930 44.475 124.935 ;
        RECT 44.725 124.760 44.895 125.240 ;
        RECT 45.065 124.935 45.395 125.410 ;
        RECT 45.145 124.930 45.315 124.935 ;
        RECT 45.565 124.760 45.735 125.240 ;
        RECT 45.905 124.935 46.235 125.410 ;
        RECT 45.985 124.930 46.235 124.935 ;
        RECT 46.405 124.760 46.575 125.240 ;
        RECT 46.745 124.935 47.075 125.410 ;
        RECT 47.245 124.760 47.415 125.240 ;
        RECT 47.585 124.935 47.915 125.410 ;
        RECT 48.085 124.760 48.255 125.240 ;
        RECT 48.425 124.935 48.755 125.410 ;
        RECT 48.925 124.760 49.095 125.240 ;
        RECT 49.265 124.935 49.595 125.410 ;
        RECT 49.765 124.760 49.935 125.240 ;
        RECT 50.105 124.935 50.435 125.410 ;
        RECT 50.615 125.220 50.865 126.590 ;
        RECT 51.795 126.420 52.095 126.970 ;
        RECT 52.265 126.640 52.545 127.310 ;
        RECT 51.155 126.250 52.095 126.420 ;
        RECT 51.155 126.000 51.325 126.250 ;
        RECT 52.465 126.000 52.730 126.360 ;
        RECT 51.035 125.670 51.325 126.000 ;
        RECT 51.495 125.750 51.835 126.000 ;
        RECT 52.055 125.750 52.730 126.000 ;
        RECT 53.375 126.220 56.885 127.310 ;
        RECT 53.375 125.700 55.065 126.220 ;
        RECT 57.115 126.170 57.325 127.310 ;
        RECT 57.495 126.160 57.825 127.140 ;
        RECT 57.995 126.170 58.225 127.310 ;
        RECT 58.525 126.380 58.695 127.140 ;
        RECT 58.875 126.550 59.205 127.310 ;
        RECT 58.525 126.210 59.190 126.380 ;
        RECT 59.375 126.235 59.645 127.140 ;
        RECT 51.155 125.580 51.325 125.670 ;
        RECT 51.155 125.390 52.545 125.580 ;
        RECT 55.235 125.530 56.885 126.050 ;
        RECT 50.615 124.930 51.175 125.220 ;
        RECT 51.345 124.760 51.595 125.220 ;
        RECT 52.215 125.030 52.545 125.390 ;
        RECT 53.375 124.760 56.885 125.530 ;
        RECT 57.115 124.760 57.325 125.580 ;
        RECT 57.495 125.560 57.745 126.160 ;
        RECT 59.020 126.065 59.190 126.210 ;
        RECT 57.915 125.750 58.245 126.000 ;
        RECT 58.455 125.660 58.785 126.030 ;
        RECT 59.020 125.735 59.305 126.065 ;
        RECT 57.495 124.930 57.825 125.560 ;
        RECT 57.995 124.760 58.225 125.580 ;
        RECT 59.020 125.480 59.190 125.735 ;
        RECT 58.525 125.310 59.190 125.480 ;
        RECT 59.475 125.435 59.645 126.235 ;
        RECT 60.275 126.220 63.785 127.310 ;
        RECT 60.275 125.700 61.965 126.220 ;
        RECT 63.955 126.145 64.245 127.310 ;
        RECT 64.415 126.220 67.005 127.310 ;
        RECT 62.135 125.530 63.785 126.050 ;
        RECT 64.415 125.700 65.625 126.220 ;
        RECT 67.180 126.170 67.515 127.140 ;
        RECT 67.685 126.170 67.855 127.310 ;
        RECT 68.025 126.970 70.055 127.140 ;
        RECT 65.795 125.530 67.005 126.050 ;
        RECT 58.525 124.930 58.695 125.310 ;
        RECT 58.875 124.760 59.205 125.140 ;
        RECT 59.385 124.930 59.645 125.435 ;
        RECT 60.275 124.760 63.785 125.530 ;
        RECT 63.955 124.760 64.245 125.485 ;
        RECT 64.415 124.760 67.005 125.530 ;
        RECT 67.180 125.500 67.350 126.170 ;
        RECT 68.025 126.000 68.195 126.970 ;
        RECT 67.520 125.670 67.775 126.000 ;
        RECT 68.000 125.670 68.195 126.000 ;
        RECT 68.365 126.630 69.490 126.800 ;
        RECT 67.605 125.500 67.775 125.670 ;
        RECT 68.365 125.500 68.535 126.630 ;
        RECT 67.180 124.930 67.435 125.500 ;
        RECT 67.605 125.330 68.535 125.500 ;
        RECT 68.705 126.290 69.715 126.460 ;
        RECT 68.705 125.490 68.875 126.290 ;
        RECT 69.080 125.950 69.355 126.090 ;
        RECT 69.075 125.780 69.355 125.950 ;
        RECT 68.360 125.295 68.535 125.330 ;
        RECT 67.605 124.760 67.935 125.160 ;
        RECT 68.360 124.930 68.890 125.295 ;
        RECT 69.080 124.930 69.355 125.780 ;
        RECT 69.525 124.930 69.715 126.290 ;
        RECT 69.885 126.305 70.055 126.970 ;
        RECT 70.225 126.550 70.395 127.310 ;
        RECT 70.630 126.550 71.145 126.960 ;
        RECT 69.885 126.115 70.635 126.305 ;
        RECT 70.805 125.740 71.145 126.550 ;
        RECT 69.915 125.570 71.145 125.740 ;
        RECT 71.315 126.590 71.775 127.140 ;
        RECT 71.965 126.590 72.295 127.310 ;
        RECT 69.895 124.760 70.405 125.295 ;
        RECT 70.625 124.965 70.870 125.570 ;
        RECT 71.315 125.220 71.565 126.590 ;
        RECT 72.495 126.420 72.795 126.970 ;
        RECT 72.965 126.640 73.245 127.310 ;
        RECT 73.990 126.970 74.245 127.000 ;
        RECT 73.905 126.800 74.245 126.970 ;
        RECT 71.855 126.250 72.795 126.420 ;
        RECT 71.855 126.000 72.025 126.250 ;
        RECT 73.165 126.000 73.430 126.360 ;
        RECT 71.735 125.670 72.025 126.000 ;
        RECT 72.195 125.750 72.535 126.000 ;
        RECT 72.755 125.750 73.430 126.000 ;
        RECT 73.990 126.330 74.245 126.800 ;
        RECT 74.425 126.510 74.710 127.310 ;
        RECT 74.890 126.590 75.220 127.100 ;
        RECT 71.855 125.580 72.025 125.670 ;
        RECT 71.855 125.390 73.245 125.580 ;
        RECT 71.315 124.930 71.875 125.220 ;
        RECT 72.045 124.760 72.295 125.220 ;
        RECT 72.915 125.030 73.245 125.390 ;
        RECT 73.990 125.470 74.170 126.330 ;
        RECT 74.890 126.000 75.140 126.590 ;
        RECT 75.490 126.440 75.660 127.050 ;
        RECT 75.830 126.620 76.160 127.310 ;
        RECT 76.390 126.760 76.630 127.050 ;
        RECT 76.830 126.930 77.250 127.310 ;
        RECT 77.430 126.840 78.060 127.090 ;
        RECT 78.530 126.930 78.860 127.310 ;
        RECT 77.430 126.760 77.600 126.840 ;
        RECT 79.030 126.760 79.200 127.050 ;
        RECT 79.380 126.930 79.760 127.310 ;
        RECT 80.000 126.925 80.830 127.095 ;
        RECT 76.390 126.590 77.600 126.760 ;
        RECT 74.340 125.670 75.140 126.000 ;
        RECT 73.990 124.940 74.245 125.470 ;
        RECT 74.425 124.760 74.710 125.220 ;
        RECT 74.890 125.020 75.140 125.670 ;
        RECT 75.340 126.420 75.660 126.440 ;
        RECT 75.340 126.250 77.260 126.420 ;
        RECT 75.340 125.355 75.530 126.250 ;
        RECT 77.430 126.080 77.600 126.590 ;
        RECT 77.770 126.330 78.290 126.640 ;
        RECT 75.700 125.910 77.600 126.080 ;
        RECT 75.700 125.850 76.030 125.910 ;
        RECT 76.180 125.680 76.510 125.740 ;
        RECT 75.850 125.410 76.510 125.680 ;
        RECT 75.340 125.025 75.660 125.355 ;
        RECT 75.840 124.760 76.500 125.240 ;
        RECT 76.700 125.150 76.870 125.910 ;
        RECT 77.770 125.740 77.950 126.150 ;
        RECT 77.040 125.570 77.370 125.690 ;
        RECT 78.120 125.570 78.290 126.330 ;
        RECT 77.040 125.400 78.290 125.570 ;
        RECT 78.460 126.510 79.830 126.760 ;
        RECT 78.460 125.740 78.650 126.510 ;
        RECT 79.580 126.250 79.830 126.510 ;
        RECT 78.820 126.080 79.070 126.240 ;
        RECT 80.000 126.080 80.170 126.925 ;
        RECT 81.065 126.640 81.235 127.140 ;
        RECT 81.405 126.810 81.735 127.310 ;
        RECT 80.340 126.250 80.840 126.630 ;
        RECT 81.065 126.470 81.760 126.640 ;
        RECT 78.820 125.910 80.170 126.080 ;
        RECT 79.750 125.870 80.170 125.910 ;
        RECT 78.460 125.400 78.880 125.740 ;
        RECT 79.170 125.410 79.580 125.740 ;
        RECT 76.700 124.980 77.550 125.150 ;
        RECT 78.110 124.760 78.430 125.220 ;
        RECT 78.630 124.970 78.880 125.400 ;
        RECT 79.170 124.760 79.580 125.200 ;
        RECT 79.750 125.140 79.920 125.870 ;
        RECT 80.090 125.320 80.440 125.690 ;
        RECT 80.620 125.380 80.840 126.250 ;
        RECT 81.010 125.680 81.420 126.300 ;
        RECT 81.590 125.500 81.760 126.470 ;
        RECT 81.065 125.310 81.760 125.500 ;
        RECT 79.750 124.940 80.765 125.140 ;
        RECT 81.065 124.980 81.235 125.310 ;
        RECT 81.405 124.760 81.735 125.140 ;
        RECT 81.950 125.020 82.175 127.140 ;
        RECT 82.345 126.810 82.675 127.310 ;
        RECT 82.845 126.640 83.015 127.140 ;
        RECT 82.350 126.470 83.015 126.640 ;
        RECT 82.350 125.480 82.580 126.470 ;
        RECT 82.750 125.650 83.100 126.300 ;
        RECT 83.275 126.235 83.545 127.140 ;
        RECT 83.715 126.550 84.045 127.310 ;
        RECT 84.225 126.380 84.395 127.140 ;
        RECT 82.350 125.310 83.015 125.480 ;
        RECT 82.345 124.760 82.675 125.140 ;
        RECT 82.845 125.020 83.015 125.310 ;
        RECT 83.275 125.435 83.445 126.235 ;
        RECT 83.730 126.210 84.395 126.380 ;
        RECT 85.115 126.220 86.785 127.310 ;
        RECT 83.730 126.065 83.900 126.210 ;
        RECT 83.615 125.735 83.900 126.065 ;
        RECT 83.730 125.480 83.900 125.735 ;
        RECT 84.135 125.660 84.465 126.030 ;
        RECT 85.115 125.700 85.865 126.220 ;
        RECT 86.995 126.170 87.225 127.310 ;
        RECT 87.395 126.160 87.725 127.140 ;
        RECT 87.895 126.170 88.105 127.310 ;
        RECT 88.335 126.220 89.545 127.310 ;
        RECT 86.035 125.530 86.785 126.050 ;
        RECT 86.975 125.750 87.305 126.000 ;
        RECT 83.275 124.930 83.535 125.435 ;
        RECT 83.730 125.310 84.395 125.480 ;
        RECT 83.715 124.760 84.045 125.140 ;
        RECT 84.225 124.930 84.395 125.310 ;
        RECT 85.115 124.760 86.785 125.530 ;
        RECT 86.995 124.760 87.225 125.580 ;
        RECT 87.475 125.560 87.725 126.160 ;
        RECT 88.335 125.680 88.855 126.220 ;
        RECT 89.715 126.145 90.005 127.310 ;
        RECT 90.180 126.170 90.515 127.140 ;
        RECT 90.685 126.170 90.855 127.310 ;
        RECT 91.025 126.970 93.055 127.140 ;
        RECT 87.395 124.930 87.725 125.560 ;
        RECT 87.895 124.760 88.105 125.580 ;
        RECT 89.025 125.510 89.545 126.050 ;
        RECT 88.335 124.760 89.545 125.510 ;
        RECT 90.180 125.500 90.350 126.170 ;
        RECT 91.025 126.000 91.195 126.970 ;
        RECT 90.520 125.670 90.775 126.000 ;
        RECT 91.000 125.670 91.195 126.000 ;
        RECT 91.365 126.630 92.490 126.800 ;
        RECT 90.605 125.500 90.775 125.670 ;
        RECT 91.365 125.500 91.535 126.630 ;
        RECT 89.715 124.760 90.005 125.485 ;
        RECT 90.180 124.930 90.435 125.500 ;
        RECT 90.605 125.330 91.535 125.500 ;
        RECT 91.705 126.290 92.715 126.460 ;
        RECT 91.705 125.490 91.875 126.290 ;
        RECT 92.080 125.950 92.355 126.090 ;
        RECT 92.075 125.780 92.355 125.950 ;
        RECT 91.360 125.295 91.535 125.330 ;
        RECT 90.605 124.760 90.935 125.160 ;
        RECT 91.360 124.930 91.890 125.295 ;
        RECT 92.080 124.930 92.355 125.780 ;
        RECT 92.525 124.930 92.715 126.290 ;
        RECT 92.885 126.305 93.055 126.970 ;
        RECT 93.225 126.550 93.395 127.310 ;
        RECT 93.630 126.550 94.145 126.960 ;
        RECT 92.885 126.115 93.635 126.305 ;
        RECT 93.805 125.740 94.145 126.550 ;
        RECT 92.915 125.570 94.145 125.740 ;
        RECT 94.315 126.220 95.525 127.310 ;
        RECT 95.695 126.550 96.210 126.960 ;
        RECT 96.445 126.550 96.615 127.310 ;
        RECT 96.785 126.970 98.815 127.140 ;
        RECT 94.315 125.680 94.835 126.220 ;
        RECT 92.895 124.760 93.405 125.295 ;
        RECT 93.625 124.965 93.870 125.570 ;
        RECT 95.005 125.510 95.525 126.050 ;
        RECT 95.695 125.740 96.035 126.550 ;
        RECT 96.785 126.305 96.955 126.970 ;
        RECT 97.350 126.630 98.475 126.800 ;
        RECT 96.205 126.115 96.955 126.305 ;
        RECT 97.125 126.290 98.135 126.460 ;
        RECT 95.695 125.570 96.925 125.740 ;
        RECT 94.315 124.760 95.525 125.510 ;
        RECT 95.970 124.965 96.215 125.570 ;
        RECT 96.435 124.760 96.945 125.295 ;
        RECT 97.125 124.930 97.315 126.290 ;
        RECT 97.485 125.270 97.760 126.090 ;
        RECT 97.965 125.490 98.135 126.290 ;
        RECT 98.305 125.500 98.475 126.630 ;
        RECT 98.645 126.000 98.815 126.970 ;
        RECT 98.985 126.170 99.155 127.310 ;
        RECT 99.325 126.170 99.660 127.140 ;
        RECT 100.210 126.970 100.465 127.000 ;
        RECT 100.125 126.800 100.465 126.970 ;
        RECT 98.645 125.670 98.840 126.000 ;
        RECT 99.065 125.670 99.320 126.000 ;
        RECT 99.065 125.500 99.235 125.670 ;
        RECT 99.490 125.500 99.660 126.170 ;
        RECT 98.305 125.330 99.235 125.500 ;
        RECT 98.305 125.295 98.480 125.330 ;
        RECT 97.485 125.100 97.765 125.270 ;
        RECT 97.485 124.930 97.760 125.100 ;
        RECT 97.950 124.930 98.480 125.295 ;
        RECT 98.905 124.760 99.235 125.160 ;
        RECT 99.405 124.930 99.660 125.500 ;
        RECT 100.210 126.330 100.465 126.800 ;
        RECT 100.645 126.510 100.930 127.310 ;
        RECT 101.110 126.590 101.440 127.100 ;
        RECT 100.210 125.470 100.390 126.330 ;
        RECT 101.110 126.000 101.360 126.590 ;
        RECT 101.710 126.440 101.880 127.050 ;
        RECT 102.050 126.620 102.380 127.310 ;
        RECT 102.610 126.760 102.850 127.050 ;
        RECT 103.050 126.930 103.470 127.310 ;
        RECT 103.650 126.840 104.280 127.090 ;
        RECT 104.750 126.930 105.080 127.310 ;
        RECT 103.650 126.760 103.820 126.840 ;
        RECT 105.250 126.760 105.420 127.050 ;
        RECT 105.600 126.930 105.980 127.310 ;
        RECT 106.220 126.925 107.050 127.095 ;
        RECT 102.610 126.590 103.820 126.760 ;
        RECT 100.560 125.670 101.360 126.000 ;
        RECT 100.210 124.940 100.465 125.470 ;
        RECT 100.645 124.760 100.930 125.220 ;
        RECT 101.110 125.020 101.360 125.670 ;
        RECT 101.560 126.420 101.880 126.440 ;
        RECT 101.560 126.250 103.480 126.420 ;
        RECT 101.560 125.355 101.750 126.250 ;
        RECT 103.650 126.080 103.820 126.590 ;
        RECT 103.990 126.330 104.510 126.640 ;
        RECT 101.920 125.910 103.820 126.080 ;
        RECT 101.920 125.850 102.250 125.910 ;
        RECT 102.400 125.680 102.730 125.740 ;
        RECT 102.070 125.410 102.730 125.680 ;
        RECT 101.560 125.025 101.880 125.355 ;
        RECT 102.060 124.760 102.720 125.240 ;
        RECT 102.920 125.150 103.090 125.910 ;
        RECT 103.990 125.740 104.170 126.150 ;
        RECT 103.260 125.570 103.590 125.690 ;
        RECT 104.340 125.570 104.510 126.330 ;
        RECT 103.260 125.400 104.510 125.570 ;
        RECT 104.680 126.510 106.050 126.760 ;
        RECT 104.680 125.740 104.870 126.510 ;
        RECT 105.800 126.250 106.050 126.510 ;
        RECT 105.040 126.080 105.290 126.240 ;
        RECT 106.220 126.080 106.390 126.925 ;
        RECT 107.285 126.640 107.455 127.140 ;
        RECT 107.625 126.810 107.955 127.310 ;
        RECT 106.560 126.250 107.060 126.630 ;
        RECT 107.285 126.470 107.980 126.640 ;
        RECT 105.040 125.910 106.390 126.080 ;
        RECT 105.970 125.870 106.390 125.910 ;
        RECT 104.680 125.400 105.100 125.740 ;
        RECT 105.390 125.410 105.800 125.740 ;
        RECT 102.920 124.980 103.770 125.150 ;
        RECT 104.330 124.760 104.650 125.220 ;
        RECT 104.850 124.970 105.100 125.400 ;
        RECT 105.390 124.760 105.800 125.200 ;
        RECT 105.970 125.140 106.140 125.870 ;
        RECT 106.310 125.320 106.660 125.690 ;
        RECT 106.840 125.380 107.060 126.250 ;
        RECT 107.230 125.680 107.640 126.300 ;
        RECT 107.810 125.500 107.980 126.470 ;
        RECT 107.285 125.310 107.980 125.500 ;
        RECT 105.970 124.940 106.985 125.140 ;
        RECT 107.285 124.980 107.455 125.310 ;
        RECT 107.625 124.760 107.955 125.140 ;
        RECT 108.170 125.020 108.395 127.140 ;
        RECT 108.565 126.810 108.895 127.310 ;
        RECT 109.065 126.640 109.235 127.140 ;
        RECT 108.570 126.470 109.235 126.640 ;
        RECT 108.570 125.480 108.800 126.470 ;
        RECT 109.585 126.380 109.755 127.140 ;
        RECT 109.935 126.550 110.265 127.310 ;
        RECT 108.970 125.650 109.320 126.300 ;
        RECT 109.585 126.210 110.250 126.380 ;
        RECT 110.435 126.235 110.705 127.140 ;
        RECT 110.080 126.065 110.250 126.210 ;
        RECT 109.515 125.660 109.845 126.030 ;
        RECT 110.080 125.735 110.365 126.065 ;
        RECT 110.080 125.480 110.250 125.735 ;
        RECT 108.570 125.310 109.235 125.480 ;
        RECT 108.565 124.760 108.895 125.140 ;
        RECT 109.065 125.020 109.235 125.310 ;
        RECT 109.585 125.310 110.250 125.480 ;
        RECT 110.535 125.435 110.705 126.235 ;
        RECT 110.875 126.220 114.385 127.310 ;
        RECT 114.555 126.220 115.765 127.310 ;
        RECT 110.875 125.700 112.565 126.220 ;
        RECT 112.735 125.530 114.385 126.050 ;
        RECT 114.555 125.680 115.075 126.220 ;
        RECT 109.585 124.930 109.755 125.310 ;
        RECT 109.935 124.760 110.265 125.140 ;
        RECT 110.445 124.930 110.705 125.435 ;
        RECT 110.875 124.760 114.385 125.530 ;
        RECT 115.245 125.510 115.765 126.050 ;
        RECT 114.555 124.760 115.765 125.510 ;
        RECT 14.650 124.590 115.850 124.760 ;
        RECT 14.735 123.840 15.945 124.590 ;
        RECT 14.735 123.300 15.255 123.840 ;
        RECT 16.635 123.770 16.845 124.590 ;
        RECT 17.015 123.790 17.345 124.420 ;
        RECT 15.425 123.130 15.945 123.670 ;
        RECT 17.015 123.190 17.265 123.790 ;
        RECT 17.515 123.770 17.745 124.590 ;
        RECT 17.995 123.770 18.225 124.590 ;
        RECT 18.395 123.790 18.725 124.420 ;
        RECT 17.435 123.350 17.765 123.600 ;
        RECT 17.975 123.350 18.305 123.600 ;
        RECT 18.475 123.190 18.725 123.790 ;
        RECT 18.895 123.770 19.105 124.590 ;
        RECT 19.425 124.040 19.595 124.420 ;
        RECT 19.775 124.210 20.105 124.590 ;
        RECT 19.425 123.870 20.090 124.040 ;
        RECT 20.285 123.915 20.545 124.420 ;
        RECT 19.355 123.320 19.685 123.690 ;
        RECT 19.920 123.615 20.090 123.870 ;
        RECT 14.735 122.040 15.945 123.130 ;
        RECT 16.635 122.040 16.845 123.180 ;
        RECT 17.015 122.210 17.345 123.190 ;
        RECT 17.515 122.040 17.745 123.180 ;
        RECT 17.995 122.040 18.225 123.180 ;
        RECT 18.395 122.210 18.725 123.190 ;
        RECT 19.920 123.285 20.205 123.615 ;
        RECT 18.895 122.040 19.105 123.180 ;
        RECT 19.920 123.140 20.090 123.285 ;
        RECT 19.425 122.970 20.090 123.140 ;
        RECT 20.375 123.115 20.545 123.915 ;
        RECT 19.425 122.210 19.595 122.970 ;
        RECT 19.775 122.040 20.105 122.800 ;
        RECT 20.275 122.210 20.545 123.115 ;
        RECT 20.720 123.850 20.975 124.420 ;
        RECT 21.145 124.190 21.475 124.590 ;
        RECT 21.900 124.055 22.430 124.420 ;
        RECT 21.900 124.020 22.075 124.055 ;
        RECT 21.145 123.850 22.075 124.020 ;
        RECT 20.720 123.180 20.890 123.850 ;
        RECT 21.145 123.680 21.315 123.850 ;
        RECT 21.060 123.350 21.315 123.680 ;
        RECT 21.540 123.350 21.735 123.680 ;
        RECT 20.720 122.210 21.055 123.180 ;
        RECT 21.225 122.040 21.395 123.180 ;
        RECT 21.565 122.380 21.735 123.350 ;
        RECT 21.905 122.720 22.075 123.850 ;
        RECT 22.245 123.060 22.415 123.860 ;
        RECT 22.620 123.570 22.895 124.420 ;
        RECT 22.615 123.400 22.895 123.570 ;
        RECT 22.620 123.260 22.895 123.400 ;
        RECT 23.065 123.060 23.255 124.420 ;
        RECT 23.435 124.055 23.945 124.590 ;
        RECT 24.165 123.780 24.410 124.385 ;
        RECT 25.315 123.865 25.605 124.590 ;
        RECT 26.700 123.850 26.955 124.420 ;
        RECT 27.125 124.190 27.455 124.590 ;
        RECT 27.880 124.055 28.410 124.420 ;
        RECT 27.880 124.020 28.055 124.055 ;
        RECT 27.125 123.850 28.055 124.020 ;
        RECT 23.455 123.610 24.685 123.780 ;
        RECT 22.245 122.890 23.255 123.060 ;
        RECT 23.425 123.045 24.175 123.235 ;
        RECT 21.905 122.550 23.030 122.720 ;
        RECT 23.425 122.380 23.595 123.045 ;
        RECT 24.345 122.800 24.685 123.610 ;
        RECT 21.565 122.210 23.595 122.380 ;
        RECT 23.765 122.040 23.935 122.800 ;
        RECT 24.170 122.390 24.685 122.800 ;
        RECT 25.315 122.040 25.605 123.205 ;
        RECT 26.700 123.180 26.870 123.850 ;
        RECT 27.125 123.680 27.295 123.850 ;
        RECT 27.040 123.350 27.295 123.680 ;
        RECT 27.520 123.350 27.715 123.680 ;
        RECT 26.700 122.210 27.035 123.180 ;
        RECT 27.205 122.040 27.375 123.180 ;
        RECT 27.545 122.380 27.715 123.350 ;
        RECT 27.885 122.720 28.055 123.850 ;
        RECT 28.225 123.060 28.395 123.860 ;
        RECT 28.600 123.570 28.875 124.420 ;
        RECT 28.595 123.400 28.875 123.570 ;
        RECT 28.600 123.260 28.875 123.400 ;
        RECT 29.045 123.060 29.235 124.420 ;
        RECT 29.415 124.055 29.925 124.590 ;
        RECT 30.145 123.780 30.390 124.385 ;
        RECT 31.755 123.915 32.015 124.420 ;
        RECT 32.195 124.210 32.525 124.590 ;
        RECT 32.705 124.040 32.875 124.420 ;
        RECT 33.140 124.120 33.470 124.590 ;
        RECT 29.435 123.610 30.665 123.780 ;
        RECT 28.225 122.890 29.235 123.060 ;
        RECT 29.405 123.045 30.155 123.235 ;
        RECT 27.885 122.550 29.010 122.720 ;
        RECT 29.405 122.380 29.575 123.045 ;
        RECT 30.325 122.800 30.665 123.610 ;
        RECT 27.545 122.210 29.575 122.380 ;
        RECT 29.745 122.040 29.915 122.800 ;
        RECT 30.150 122.390 30.665 122.800 ;
        RECT 31.755 123.115 31.925 123.915 ;
        RECT 32.210 123.870 32.875 124.040 ;
        RECT 33.640 123.950 33.865 124.395 ;
        RECT 34.035 124.065 34.330 124.590 ;
        RECT 35.350 124.250 35.605 124.410 ;
        RECT 35.265 124.080 35.605 124.250 ;
        RECT 35.785 124.130 36.070 124.590 ;
        RECT 32.210 123.615 32.380 123.870 ;
        RECT 33.135 123.780 33.865 123.950 ;
        RECT 35.350 123.880 35.605 124.080 ;
        RECT 32.095 123.285 32.380 123.615 ;
        RECT 32.615 123.320 32.945 123.690 ;
        RECT 32.210 123.140 32.380 123.285 ;
        RECT 33.135 123.215 33.415 123.780 ;
        RECT 33.585 123.385 34.805 123.610 ;
        RECT 31.755 122.210 32.025 123.115 ;
        RECT 32.210 122.970 32.875 123.140 ;
        RECT 33.135 123.045 34.735 123.215 ;
        RECT 32.195 122.040 32.525 122.800 ;
        RECT 32.705 122.210 32.875 122.970 ;
        RECT 33.195 122.040 33.450 122.875 ;
        RECT 33.620 122.240 33.880 123.045 ;
        RECT 34.050 122.040 34.310 122.875 ;
        RECT 34.480 122.240 34.735 123.045 ;
        RECT 35.350 123.020 35.530 123.880 ;
        RECT 36.250 123.680 36.500 124.330 ;
        RECT 35.700 123.350 36.500 123.680 ;
        RECT 35.350 122.350 35.605 123.020 ;
        RECT 35.785 122.040 36.070 122.840 ;
        RECT 36.250 122.760 36.500 123.350 ;
        RECT 36.700 123.995 37.020 124.325 ;
        RECT 37.200 124.110 37.860 124.590 ;
        RECT 38.060 124.200 38.910 124.370 ;
        RECT 36.700 123.100 36.890 123.995 ;
        RECT 37.210 123.670 37.870 123.940 ;
        RECT 37.540 123.610 37.870 123.670 ;
        RECT 37.060 123.440 37.390 123.500 ;
        RECT 38.060 123.440 38.230 124.200 ;
        RECT 39.470 124.130 39.790 124.590 ;
        RECT 39.990 123.950 40.240 124.380 ;
        RECT 40.530 124.150 40.940 124.590 ;
        RECT 41.110 124.210 42.125 124.410 ;
        RECT 38.400 123.780 39.650 123.950 ;
        RECT 38.400 123.660 38.730 123.780 ;
        RECT 37.060 123.270 38.960 123.440 ;
        RECT 36.700 122.930 38.620 123.100 ;
        RECT 36.700 122.910 37.020 122.930 ;
        RECT 36.250 122.250 36.580 122.760 ;
        RECT 36.850 122.300 37.020 122.910 ;
        RECT 38.790 122.760 38.960 123.270 ;
        RECT 39.130 123.200 39.310 123.610 ;
        RECT 39.480 123.020 39.650 123.780 ;
        RECT 37.190 122.040 37.520 122.730 ;
        RECT 37.750 122.590 38.960 122.760 ;
        RECT 39.130 122.710 39.650 123.020 ;
        RECT 39.820 123.610 40.240 123.950 ;
        RECT 40.530 123.610 40.940 123.940 ;
        RECT 39.820 122.840 40.010 123.610 ;
        RECT 41.110 123.480 41.280 124.210 ;
        RECT 42.425 124.040 42.595 124.370 ;
        RECT 42.765 124.210 43.095 124.590 ;
        RECT 41.450 123.660 41.800 124.030 ;
        RECT 41.110 123.440 41.530 123.480 ;
        RECT 40.180 123.270 41.530 123.440 ;
        RECT 40.180 123.110 40.430 123.270 ;
        RECT 40.940 122.840 41.190 123.100 ;
        RECT 39.820 122.590 41.190 122.840 ;
        RECT 37.750 122.300 37.990 122.590 ;
        RECT 38.790 122.510 38.960 122.590 ;
        RECT 38.190 122.040 38.610 122.420 ;
        RECT 38.790 122.260 39.420 122.510 ;
        RECT 39.890 122.040 40.220 122.420 ;
        RECT 40.390 122.300 40.560 122.590 ;
        RECT 41.360 122.425 41.530 123.270 ;
        RECT 41.980 123.100 42.200 123.970 ;
        RECT 42.425 123.850 43.120 124.040 ;
        RECT 41.700 122.720 42.200 123.100 ;
        RECT 42.370 123.050 42.780 123.670 ;
        RECT 42.950 122.880 43.120 123.850 ;
        RECT 42.425 122.710 43.120 122.880 ;
        RECT 40.740 122.040 41.120 122.420 ;
        RECT 41.360 122.255 42.190 122.425 ;
        RECT 42.425 122.210 42.595 122.710 ;
        RECT 42.765 122.040 43.095 122.540 ;
        RECT 43.310 122.210 43.535 124.330 ;
        RECT 43.705 124.210 44.035 124.590 ;
        RECT 44.205 124.040 44.375 124.330 ;
        RECT 43.710 123.870 44.375 124.040 ;
        RECT 44.635 124.130 45.195 124.420 ;
        RECT 45.365 124.130 45.615 124.590 ;
        RECT 43.710 122.880 43.940 123.870 ;
        RECT 44.110 123.050 44.460 123.700 ;
        RECT 43.710 122.710 44.375 122.880 ;
        RECT 43.705 122.040 44.035 122.540 ;
        RECT 44.205 122.210 44.375 122.710 ;
        RECT 44.635 122.760 44.885 124.130 ;
        RECT 46.235 123.960 46.565 124.320 ;
        RECT 45.175 123.770 46.565 123.960 ;
        RECT 47.210 123.780 47.455 124.385 ;
        RECT 47.675 124.055 48.185 124.590 ;
        RECT 45.175 123.680 45.345 123.770 ;
        RECT 45.055 123.350 45.345 123.680 ;
        RECT 46.935 123.610 48.165 123.780 ;
        RECT 45.515 123.350 45.855 123.600 ;
        RECT 46.075 123.350 46.750 123.600 ;
        RECT 45.175 123.100 45.345 123.350 ;
        RECT 45.175 122.930 46.115 123.100 ;
        RECT 46.485 122.990 46.750 123.350 ;
        RECT 44.635 122.210 45.095 122.760 ;
        RECT 45.285 122.040 45.615 122.760 ;
        RECT 45.815 122.380 46.115 122.930 ;
        RECT 46.935 122.800 47.275 123.610 ;
        RECT 47.445 123.045 48.195 123.235 ;
        RECT 46.285 122.040 46.565 122.710 ;
        RECT 46.935 122.390 47.450 122.800 ;
        RECT 47.685 122.040 47.855 122.800 ;
        RECT 48.025 122.380 48.195 123.045 ;
        RECT 48.365 123.060 48.555 124.420 ;
        RECT 48.725 123.570 49.000 124.420 ;
        RECT 49.190 124.055 49.720 124.420 ;
        RECT 50.145 124.190 50.475 124.590 ;
        RECT 49.545 124.020 49.720 124.055 ;
        RECT 48.725 123.400 49.005 123.570 ;
        RECT 48.725 123.260 49.000 123.400 ;
        RECT 49.205 123.060 49.375 123.860 ;
        RECT 48.365 122.890 49.375 123.060 ;
        RECT 49.545 123.850 50.475 124.020 ;
        RECT 50.645 123.850 50.900 124.420 ;
        RECT 51.075 123.865 51.365 124.590 ;
        RECT 49.545 122.720 49.715 123.850 ;
        RECT 50.305 123.680 50.475 123.850 ;
        RECT 48.590 122.550 49.715 122.720 ;
        RECT 49.885 123.350 50.080 123.680 ;
        RECT 50.305 123.350 50.560 123.680 ;
        RECT 49.885 122.380 50.055 123.350 ;
        RECT 50.730 123.180 50.900 123.850 ;
        RECT 51.995 123.820 53.665 124.590 ;
        RECT 48.025 122.210 50.055 122.380 ;
        RECT 50.225 122.040 50.395 123.180 ;
        RECT 50.565 122.210 50.900 123.180 ;
        RECT 51.075 122.040 51.365 123.205 ;
        RECT 51.995 123.130 52.745 123.650 ;
        RECT 52.915 123.300 53.665 123.820 ;
        RECT 53.875 123.770 54.105 124.590 ;
        RECT 54.275 123.790 54.605 124.420 ;
        RECT 53.855 123.350 54.185 123.600 ;
        RECT 54.355 123.190 54.605 123.790 ;
        RECT 54.775 123.770 54.985 124.590 ;
        RECT 55.365 123.790 55.695 124.590 ;
        RECT 55.865 123.940 56.035 124.420 ;
        RECT 56.205 124.110 56.535 124.590 ;
        RECT 56.705 123.940 56.875 124.420 ;
        RECT 57.125 124.110 57.365 124.590 ;
        RECT 57.545 123.940 57.715 124.420 ;
        RECT 55.865 123.770 56.875 123.940 ;
        RECT 57.080 123.770 57.715 123.940 ;
        RECT 57.975 123.820 61.485 124.590 ;
        RECT 61.745 124.040 61.915 124.330 ;
        RECT 62.085 124.210 62.415 124.590 ;
        RECT 61.745 123.870 62.410 124.040 ;
        RECT 55.865 123.570 56.360 123.770 ;
        RECT 57.080 123.600 57.250 123.770 ;
        RECT 55.865 123.400 56.365 123.570 ;
        RECT 56.750 123.430 57.250 123.600 ;
        RECT 55.865 123.230 56.360 123.400 ;
        RECT 51.995 122.040 53.665 123.130 ;
        RECT 53.875 122.040 54.105 123.180 ;
        RECT 54.275 122.210 54.605 123.190 ;
        RECT 54.775 122.040 54.985 123.180 ;
        RECT 55.365 122.040 55.695 123.190 ;
        RECT 55.865 123.060 56.875 123.230 ;
        RECT 55.865 122.210 56.035 123.060 ;
        RECT 56.205 122.040 56.535 122.840 ;
        RECT 56.705 122.210 56.875 123.060 ;
        RECT 57.080 123.190 57.250 123.430 ;
        RECT 57.420 123.360 57.800 123.600 ;
        RECT 57.080 123.020 57.795 123.190 ;
        RECT 57.055 122.040 57.295 122.840 ;
        RECT 57.465 122.210 57.795 123.020 ;
        RECT 57.975 123.130 59.665 123.650 ;
        RECT 59.835 123.300 61.485 123.820 ;
        RECT 57.975 122.040 61.485 123.130 ;
        RECT 61.660 123.050 62.010 123.700 ;
        RECT 62.180 122.880 62.410 123.870 ;
        RECT 61.745 122.710 62.410 122.880 ;
        RECT 61.745 122.210 61.915 122.710 ;
        RECT 62.085 122.040 62.415 122.540 ;
        RECT 62.585 122.210 62.810 124.330 ;
        RECT 63.025 124.210 63.355 124.590 ;
        RECT 63.525 124.040 63.695 124.370 ;
        RECT 63.995 124.210 65.010 124.410 ;
        RECT 63.000 123.850 63.695 124.040 ;
        RECT 63.000 122.880 63.170 123.850 ;
        RECT 63.340 123.050 63.750 123.670 ;
        RECT 63.920 123.100 64.140 123.970 ;
        RECT 64.320 123.660 64.670 124.030 ;
        RECT 64.840 123.480 65.010 124.210 ;
        RECT 65.180 124.150 65.590 124.590 ;
        RECT 65.880 123.950 66.130 124.380 ;
        RECT 66.330 124.130 66.650 124.590 ;
        RECT 67.210 124.200 68.060 124.370 ;
        RECT 65.180 123.610 65.590 123.940 ;
        RECT 65.880 123.610 66.300 123.950 ;
        RECT 64.590 123.440 65.010 123.480 ;
        RECT 64.590 123.270 65.940 123.440 ;
        RECT 63.000 122.710 63.695 122.880 ;
        RECT 63.920 122.720 64.420 123.100 ;
        RECT 63.025 122.040 63.355 122.540 ;
        RECT 63.525 122.210 63.695 122.710 ;
        RECT 64.590 122.425 64.760 123.270 ;
        RECT 65.690 123.110 65.940 123.270 ;
        RECT 64.930 122.840 65.180 123.100 ;
        RECT 66.110 122.840 66.300 123.610 ;
        RECT 64.930 122.590 66.300 122.840 ;
        RECT 66.470 123.780 67.720 123.950 ;
        RECT 66.470 123.020 66.640 123.780 ;
        RECT 67.390 123.660 67.720 123.780 ;
        RECT 66.810 123.200 66.990 123.610 ;
        RECT 67.890 123.440 68.060 124.200 ;
        RECT 68.260 124.110 68.920 124.590 ;
        RECT 69.100 123.995 69.420 124.325 ;
        RECT 68.250 123.670 68.910 123.940 ;
        RECT 68.250 123.610 68.580 123.670 ;
        RECT 68.730 123.440 69.060 123.500 ;
        RECT 67.160 123.270 69.060 123.440 ;
        RECT 66.470 122.710 66.990 123.020 ;
        RECT 67.160 122.760 67.330 123.270 ;
        RECT 69.230 123.100 69.420 123.995 ;
        RECT 67.500 122.930 69.420 123.100 ;
        RECT 69.100 122.910 69.420 122.930 ;
        RECT 69.620 123.680 69.870 124.330 ;
        RECT 70.050 124.130 70.335 124.590 ;
        RECT 70.515 123.910 70.770 124.410 ;
        RECT 70.515 123.880 70.855 123.910 ;
        RECT 70.590 123.740 70.855 123.880 ;
        RECT 71.590 123.780 71.835 124.385 ;
        RECT 72.055 124.055 72.565 124.590 ;
        RECT 69.620 123.350 70.420 123.680 ;
        RECT 67.160 122.590 68.370 122.760 ;
        RECT 63.930 122.255 64.760 122.425 ;
        RECT 65.000 122.040 65.380 122.420 ;
        RECT 65.560 122.300 65.730 122.590 ;
        RECT 67.160 122.510 67.330 122.590 ;
        RECT 65.900 122.040 66.230 122.420 ;
        RECT 66.700 122.260 67.330 122.510 ;
        RECT 67.510 122.040 67.930 122.420 ;
        RECT 68.130 122.300 68.370 122.590 ;
        RECT 68.600 122.040 68.930 122.730 ;
        RECT 69.100 122.300 69.270 122.910 ;
        RECT 69.620 122.760 69.870 123.350 ;
        RECT 70.590 123.020 70.770 123.740 ;
        RECT 69.540 122.250 69.870 122.760 ;
        RECT 70.050 122.040 70.335 122.840 ;
        RECT 70.515 122.350 70.770 123.020 ;
        RECT 71.315 123.610 72.545 123.780 ;
        RECT 71.315 122.800 71.655 123.610 ;
        RECT 71.825 123.045 72.575 123.235 ;
        RECT 71.315 122.390 71.830 122.800 ;
        RECT 72.065 122.040 72.235 122.800 ;
        RECT 72.405 122.380 72.575 123.045 ;
        RECT 72.745 123.060 72.935 124.420 ;
        RECT 73.105 123.570 73.380 124.420 ;
        RECT 73.570 124.055 74.100 124.420 ;
        RECT 74.525 124.190 74.855 124.590 ;
        RECT 73.925 124.020 74.100 124.055 ;
        RECT 73.105 123.400 73.385 123.570 ;
        RECT 73.105 123.260 73.380 123.400 ;
        RECT 73.585 123.060 73.755 123.860 ;
        RECT 72.745 122.890 73.755 123.060 ;
        RECT 73.925 123.850 74.855 124.020 ;
        RECT 75.025 123.850 75.280 124.420 ;
        RECT 73.925 122.720 74.095 123.850 ;
        RECT 74.685 123.680 74.855 123.850 ;
        RECT 72.970 122.550 74.095 122.720 ;
        RECT 74.265 123.350 74.460 123.680 ;
        RECT 74.685 123.350 74.940 123.680 ;
        RECT 74.265 122.380 74.435 123.350 ;
        RECT 75.110 123.180 75.280 123.850 ;
        RECT 75.455 123.840 76.665 124.590 ;
        RECT 76.835 123.865 77.125 124.590 ;
        RECT 72.405 122.210 74.435 122.380 ;
        RECT 74.605 122.040 74.775 123.180 ;
        RECT 74.945 122.210 75.280 123.180 ;
        RECT 75.455 123.130 75.975 123.670 ;
        RECT 76.145 123.300 76.665 123.840 ;
        RECT 77.355 123.770 77.565 124.590 ;
        RECT 77.735 123.790 78.065 124.420 ;
        RECT 75.455 122.040 76.665 123.130 ;
        RECT 76.835 122.040 77.125 123.205 ;
        RECT 77.735 123.190 77.985 123.790 ;
        RECT 78.235 123.770 78.465 124.590 ;
        RECT 79.870 123.780 80.115 124.385 ;
        RECT 80.335 124.055 80.845 124.590 ;
        RECT 79.595 123.610 80.825 123.780 ;
        RECT 78.155 123.350 78.485 123.600 ;
        RECT 77.355 122.040 77.565 123.180 ;
        RECT 77.735 122.210 78.065 123.190 ;
        RECT 78.235 122.040 78.465 123.180 ;
        RECT 79.595 122.800 79.935 123.610 ;
        RECT 80.105 123.045 80.855 123.235 ;
        RECT 79.595 122.390 80.110 122.800 ;
        RECT 80.345 122.040 80.515 122.800 ;
        RECT 80.685 122.380 80.855 123.045 ;
        RECT 81.025 123.060 81.215 124.420 ;
        RECT 81.385 123.570 81.660 124.420 ;
        RECT 81.850 124.055 82.380 124.420 ;
        RECT 82.805 124.190 83.135 124.590 ;
        RECT 82.205 124.020 82.380 124.055 ;
        RECT 81.385 123.400 81.665 123.570 ;
        RECT 81.385 123.260 81.660 123.400 ;
        RECT 81.865 123.060 82.035 123.860 ;
        RECT 81.025 122.890 82.035 123.060 ;
        RECT 82.205 123.850 83.135 124.020 ;
        RECT 83.305 123.850 83.560 124.420 ;
        RECT 84.110 124.250 84.365 124.410 ;
        RECT 84.025 124.080 84.365 124.250 ;
        RECT 84.545 124.130 84.830 124.590 ;
        RECT 82.205 122.720 82.375 123.850 ;
        RECT 82.965 123.680 83.135 123.850 ;
        RECT 81.250 122.550 82.375 122.720 ;
        RECT 82.545 123.350 82.740 123.680 ;
        RECT 82.965 123.350 83.220 123.680 ;
        RECT 82.545 122.380 82.715 123.350 ;
        RECT 83.390 123.180 83.560 123.850 ;
        RECT 80.685 122.210 82.715 122.380 ;
        RECT 82.885 122.040 83.055 123.180 ;
        RECT 83.225 122.210 83.560 123.180 ;
        RECT 84.110 123.880 84.365 124.080 ;
        RECT 84.110 123.020 84.290 123.880 ;
        RECT 85.010 123.680 85.260 124.330 ;
        RECT 84.460 123.350 85.260 123.680 ;
        RECT 84.110 122.350 84.365 123.020 ;
        RECT 84.545 122.040 84.830 122.840 ;
        RECT 85.010 122.760 85.260 123.350 ;
        RECT 85.460 123.995 85.780 124.325 ;
        RECT 85.960 124.110 86.620 124.590 ;
        RECT 86.820 124.200 87.670 124.370 ;
        RECT 85.460 123.100 85.650 123.995 ;
        RECT 85.970 123.670 86.630 123.940 ;
        RECT 86.300 123.610 86.630 123.670 ;
        RECT 85.820 123.440 86.150 123.500 ;
        RECT 86.820 123.440 86.990 124.200 ;
        RECT 88.230 124.130 88.550 124.590 ;
        RECT 88.750 123.950 89.000 124.380 ;
        RECT 89.290 124.150 89.700 124.590 ;
        RECT 89.870 124.210 90.885 124.410 ;
        RECT 87.160 123.780 88.410 123.950 ;
        RECT 87.160 123.660 87.490 123.780 ;
        RECT 85.820 123.270 87.720 123.440 ;
        RECT 85.460 122.930 87.380 123.100 ;
        RECT 85.460 122.910 85.780 122.930 ;
        RECT 85.010 122.250 85.340 122.760 ;
        RECT 85.610 122.300 85.780 122.910 ;
        RECT 87.550 122.760 87.720 123.270 ;
        RECT 87.890 123.200 88.070 123.610 ;
        RECT 88.240 123.020 88.410 123.780 ;
        RECT 85.950 122.040 86.280 122.730 ;
        RECT 86.510 122.590 87.720 122.760 ;
        RECT 87.890 122.710 88.410 123.020 ;
        RECT 88.580 123.610 89.000 123.950 ;
        RECT 89.290 123.610 89.700 123.940 ;
        RECT 88.580 122.840 88.770 123.610 ;
        RECT 89.870 123.480 90.040 124.210 ;
        RECT 91.185 124.040 91.355 124.370 ;
        RECT 91.525 124.210 91.855 124.590 ;
        RECT 90.210 123.660 90.560 124.030 ;
        RECT 89.870 123.440 90.290 123.480 ;
        RECT 88.940 123.270 90.290 123.440 ;
        RECT 88.940 123.110 89.190 123.270 ;
        RECT 89.700 122.840 89.950 123.100 ;
        RECT 88.580 122.590 89.950 122.840 ;
        RECT 86.510 122.300 86.750 122.590 ;
        RECT 87.550 122.510 87.720 122.590 ;
        RECT 86.950 122.040 87.370 122.420 ;
        RECT 87.550 122.260 88.180 122.510 ;
        RECT 88.650 122.040 88.980 122.420 ;
        RECT 89.150 122.300 89.320 122.590 ;
        RECT 90.120 122.425 90.290 123.270 ;
        RECT 90.740 123.100 90.960 123.970 ;
        RECT 91.185 123.850 91.880 124.040 ;
        RECT 90.460 122.720 90.960 123.100 ;
        RECT 91.130 123.050 91.540 123.670 ;
        RECT 91.710 122.880 91.880 123.850 ;
        RECT 91.185 122.710 91.880 122.880 ;
        RECT 89.500 122.040 89.880 122.420 ;
        RECT 90.120 122.255 90.950 122.425 ;
        RECT 91.185 122.210 91.355 122.710 ;
        RECT 91.525 122.040 91.855 122.540 ;
        RECT 92.070 122.210 92.295 124.330 ;
        RECT 92.465 124.210 92.795 124.590 ;
        RECT 92.965 124.040 93.135 124.330 ;
        RECT 92.470 123.870 93.135 124.040 ;
        RECT 92.470 122.880 92.700 123.870 ;
        RECT 93.395 123.840 94.605 124.590 ;
        RECT 92.870 123.050 93.220 123.700 ;
        RECT 93.395 123.130 93.915 123.670 ;
        RECT 94.085 123.300 94.605 123.840 ;
        RECT 94.815 123.770 95.045 124.590 ;
        RECT 95.215 123.790 95.545 124.420 ;
        RECT 94.795 123.350 95.125 123.600 ;
        RECT 95.295 123.190 95.545 123.790 ;
        RECT 95.715 123.770 95.925 124.590 ;
        RECT 96.430 123.780 96.675 124.385 ;
        RECT 96.895 124.055 97.405 124.590 ;
        RECT 92.470 122.710 93.135 122.880 ;
        RECT 92.465 122.040 92.795 122.540 ;
        RECT 92.965 122.210 93.135 122.710 ;
        RECT 93.395 122.040 94.605 123.130 ;
        RECT 94.815 122.040 95.045 123.180 ;
        RECT 95.215 122.210 95.545 123.190 ;
        RECT 96.155 123.610 97.385 123.780 ;
        RECT 95.715 122.040 95.925 123.180 ;
        RECT 96.155 122.800 96.495 123.610 ;
        RECT 96.665 123.045 97.415 123.235 ;
        RECT 96.155 122.390 96.670 122.800 ;
        RECT 96.905 122.040 97.075 122.800 ;
        RECT 97.245 122.380 97.415 123.045 ;
        RECT 97.585 123.060 97.775 124.420 ;
        RECT 97.945 123.570 98.220 124.420 ;
        RECT 98.410 124.055 98.940 124.420 ;
        RECT 99.365 124.190 99.695 124.590 ;
        RECT 98.765 124.020 98.940 124.055 ;
        RECT 97.945 123.400 98.225 123.570 ;
        RECT 97.945 123.260 98.220 123.400 ;
        RECT 98.425 123.060 98.595 123.860 ;
        RECT 97.585 122.890 98.595 123.060 ;
        RECT 98.765 123.850 99.695 124.020 ;
        RECT 99.865 123.850 100.120 124.420 ;
        RECT 101.305 124.040 101.475 124.420 ;
        RECT 101.655 124.210 101.985 124.590 ;
        RECT 101.305 123.870 101.970 124.040 ;
        RECT 102.165 123.915 102.425 124.420 ;
        RECT 98.765 122.720 98.935 123.850 ;
        RECT 99.525 123.680 99.695 123.850 ;
        RECT 97.810 122.550 98.935 122.720 ;
        RECT 99.105 123.350 99.300 123.680 ;
        RECT 99.525 123.350 99.780 123.680 ;
        RECT 99.105 122.380 99.275 123.350 ;
        RECT 99.950 123.180 100.120 123.850 ;
        RECT 101.235 123.320 101.565 123.690 ;
        RECT 101.800 123.615 101.970 123.870 ;
        RECT 97.245 122.210 99.275 122.380 ;
        RECT 99.445 122.040 99.615 123.180 ;
        RECT 99.785 122.210 100.120 123.180 ;
        RECT 101.800 123.285 102.085 123.615 ;
        RECT 101.800 123.140 101.970 123.285 ;
        RECT 101.305 122.970 101.970 123.140 ;
        RECT 102.255 123.115 102.425 123.915 ;
        RECT 102.595 123.865 102.885 124.590 ;
        RECT 103.430 123.910 103.685 124.410 ;
        RECT 103.865 124.130 104.150 124.590 ;
        RECT 103.345 123.880 103.685 123.910 ;
        RECT 103.345 123.740 103.610 123.880 ;
        RECT 101.305 122.210 101.475 122.970 ;
        RECT 101.655 122.040 101.985 122.800 ;
        RECT 102.155 122.210 102.425 123.115 ;
        RECT 102.595 122.040 102.885 123.205 ;
        RECT 103.430 123.020 103.610 123.740 ;
        RECT 104.330 123.680 104.580 124.330 ;
        RECT 103.780 123.350 104.580 123.680 ;
        RECT 103.430 122.350 103.685 123.020 ;
        RECT 103.865 122.040 104.150 122.840 ;
        RECT 104.330 122.760 104.580 123.350 ;
        RECT 104.780 123.995 105.100 124.325 ;
        RECT 105.280 124.110 105.940 124.590 ;
        RECT 106.140 124.200 106.990 124.370 ;
        RECT 104.780 123.100 104.970 123.995 ;
        RECT 105.290 123.670 105.950 123.940 ;
        RECT 105.620 123.610 105.950 123.670 ;
        RECT 105.140 123.440 105.470 123.500 ;
        RECT 106.140 123.440 106.310 124.200 ;
        RECT 107.550 124.130 107.870 124.590 ;
        RECT 108.070 123.950 108.320 124.380 ;
        RECT 108.610 124.150 109.020 124.590 ;
        RECT 109.190 124.210 110.205 124.410 ;
        RECT 106.480 123.780 107.730 123.950 ;
        RECT 106.480 123.660 106.810 123.780 ;
        RECT 105.140 123.270 107.040 123.440 ;
        RECT 104.780 122.930 106.700 123.100 ;
        RECT 104.780 122.910 105.100 122.930 ;
        RECT 104.330 122.250 104.660 122.760 ;
        RECT 104.930 122.300 105.100 122.910 ;
        RECT 106.870 122.760 107.040 123.270 ;
        RECT 107.210 123.200 107.390 123.610 ;
        RECT 107.560 123.020 107.730 123.780 ;
        RECT 105.270 122.040 105.600 122.730 ;
        RECT 105.830 122.590 107.040 122.760 ;
        RECT 107.210 122.710 107.730 123.020 ;
        RECT 107.900 123.610 108.320 123.950 ;
        RECT 108.610 123.610 109.020 123.940 ;
        RECT 107.900 122.840 108.090 123.610 ;
        RECT 109.190 123.480 109.360 124.210 ;
        RECT 110.505 124.040 110.675 124.370 ;
        RECT 110.845 124.210 111.175 124.590 ;
        RECT 109.530 123.660 109.880 124.030 ;
        RECT 109.190 123.440 109.610 123.480 ;
        RECT 108.260 123.270 109.610 123.440 ;
        RECT 108.260 123.110 108.510 123.270 ;
        RECT 109.020 122.840 109.270 123.100 ;
        RECT 107.900 122.590 109.270 122.840 ;
        RECT 105.830 122.300 106.070 122.590 ;
        RECT 106.870 122.510 107.040 122.590 ;
        RECT 106.270 122.040 106.690 122.420 ;
        RECT 106.870 122.260 107.500 122.510 ;
        RECT 107.970 122.040 108.300 122.420 ;
        RECT 108.470 122.300 108.640 122.590 ;
        RECT 109.440 122.425 109.610 123.270 ;
        RECT 110.060 123.100 110.280 123.970 ;
        RECT 110.505 123.850 111.200 124.040 ;
        RECT 109.780 122.720 110.280 123.100 ;
        RECT 110.450 123.050 110.860 123.670 ;
        RECT 111.030 122.880 111.200 123.850 ;
        RECT 110.505 122.710 111.200 122.880 ;
        RECT 108.820 122.040 109.200 122.420 ;
        RECT 109.440 122.255 110.270 122.425 ;
        RECT 110.505 122.210 110.675 122.710 ;
        RECT 110.845 122.040 111.175 122.540 ;
        RECT 111.390 122.210 111.615 124.330 ;
        RECT 111.785 124.210 112.115 124.590 ;
        RECT 112.285 124.040 112.455 124.330 ;
        RECT 111.790 123.870 112.455 124.040 ;
        RECT 111.790 122.880 112.020 123.870 ;
        RECT 112.715 123.820 114.385 124.590 ;
        RECT 114.555 123.840 115.765 124.590 ;
        RECT 112.190 123.050 112.540 123.700 ;
        RECT 112.715 123.130 113.465 123.650 ;
        RECT 113.635 123.300 114.385 123.820 ;
        RECT 114.555 123.130 115.075 123.670 ;
        RECT 115.245 123.300 115.765 123.840 ;
        RECT 111.790 122.710 112.455 122.880 ;
        RECT 111.785 122.040 112.115 122.540 ;
        RECT 112.285 122.210 112.455 122.710 ;
        RECT 112.715 122.040 114.385 123.130 ;
        RECT 114.555 122.040 115.765 123.130 ;
        RECT 14.650 121.870 115.850 122.040 ;
        RECT 14.735 120.780 15.945 121.870 ;
        RECT 14.735 120.070 15.255 120.610 ;
        RECT 15.425 120.240 15.945 120.780 ;
        RECT 16.115 120.780 17.785 121.870 ;
        RECT 17.960 121.435 23.305 121.870 ;
        RECT 16.115 120.260 16.865 120.780 ;
        RECT 17.035 120.090 17.785 120.610 ;
        RECT 19.550 120.185 19.900 121.435 ;
        RECT 23.565 121.200 23.735 121.700 ;
        RECT 23.905 121.370 24.235 121.870 ;
        RECT 23.565 121.030 24.230 121.200 ;
        RECT 14.735 119.320 15.945 120.070 ;
        RECT 16.115 119.320 17.785 120.090 ;
        RECT 21.380 119.865 21.720 120.695 ;
        RECT 23.480 120.210 23.830 120.860 ;
        RECT 24.000 120.040 24.230 121.030 ;
        RECT 23.565 119.870 24.230 120.040 ;
        RECT 17.960 119.320 23.305 119.865 ;
        RECT 23.565 119.580 23.735 119.870 ;
        RECT 23.905 119.320 24.235 119.700 ;
        RECT 24.405 119.580 24.630 121.700 ;
        RECT 24.845 121.370 25.175 121.870 ;
        RECT 25.345 121.200 25.515 121.700 ;
        RECT 25.750 121.485 26.580 121.655 ;
        RECT 26.820 121.490 27.200 121.870 ;
        RECT 24.820 121.030 25.515 121.200 ;
        RECT 24.820 120.060 24.990 121.030 ;
        RECT 25.160 120.240 25.570 120.860 ;
        RECT 25.740 120.810 26.240 121.190 ;
        RECT 24.820 119.870 25.515 120.060 ;
        RECT 25.740 119.940 25.960 120.810 ;
        RECT 26.410 120.640 26.580 121.485 ;
        RECT 27.380 121.320 27.550 121.610 ;
        RECT 27.720 121.490 28.050 121.870 ;
        RECT 28.520 121.400 29.150 121.650 ;
        RECT 29.330 121.490 29.750 121.870 ;
        RECT 28.980 121.320 29.150 121.400 ;
        RECT 29.950 121.320 30.190 121.610 ;
        RECT 26.750 121.070 28.120 121.320 ;
        RECT 26.750 120.810 27.000 121.070 ;
        RECT 27.510 120.640 27.760 120.800 ;
        RECT 26.410 120.470 27.760 120.640 ;
        RECT 26.410 120.430 26.830 120.470 ;
        RECT 26.140 119.880 26.490 120.250 ;
        RECT 24.845 119.320 25.175 119.700 ;
        RECT 25.345 119.540 25.515 119.870 ;
        RECT 26.660 119.700 26.830 120.430 ;
        RECT 27.930 120.300 28.120 121.070 ;
        RECT 27.000 119.970 27.410 120.300 ;
        RECT 27.700 119.960 28.120 120.300 ;
        RECT 28.290 120.890 28.810 121.200 ;
        RECT 28.980 121.150 30.190 121.320 ;
        RECT 30.420 121.180 30.750 121.870 ;
        RECT 28.290 120.130 28.460 120.890 ;
        RECT 28.630 120.300 28.810 120.710 ;
        RECT 28.980 120.640 29.150 121.150 ;
        RECT 30.920 121.000 31.090 121.610 ;
        RECT 31.360 121.150 31.690 121.660 ;
        RECT 30.920 120.980 31.240 121.000 ;
        RECT 29.320 120.810 31.240 120.980 ;
        RECT 28.980 120.470 30.880 120.640 ;
        RECT 29.210 120.130 29.540 120.250 ;
        RECT 28.290 119.960 29.540 120.130 ;
        RECT 25.815 119.500 26.830 119.700 ;
        RECT 27.000 119.320 27.410 119.760 ;
        RECT 27.700 119.530 27.950 119.960 ;
        RECT 28.150 119.320 28.470 119.780 ;
        RECT 29.710 119.710 29.880 120.470 ;
        RECT 30.550 120.410 30.880 120.470 ;
        RECT 30.070 120.240 30.400 120.300 ;
        RECT 30.070 119.970 30.730 120.240 ;
        RECT 31.050 119.915 31.240 120.810 ;
        RECT 29.030 119.540 29.880 119.710 ;
        RECT 30.080 119.320 30.740 119.800 ;
        RECT 30.920 119.585 31.240 119.915 ;
        RECT 31.440 120.560 31.690 121.150 ;
        RECT 31.870 121.070 32.155 121.870 ;
        RECT 32.335 120.890 32.590 121.560 ;
        RECT 31.440 120.230 32.240 120.560 ;
        RECT 32.410 120.510 32.590 120.890 ;
        RECT 34.060 120.730 34.395 121.700 ;
        RECT 34.565 120.730 34.735 121.870 ;
        RECT 34.905 121.530 36.935 121.700 ;
        RECT 32.410 120.340 32.675 120.510 ;
        RECT 31.440 119.580 31.690 120.230 ;
        RECT 32.410 120.030 32.590 120.340 ;
        RECT 31.870 119.320 32.155 119.780 ;
        RECT 32.335 119.500 32.590 120.030 ;
        RECT 34.060 120.060 34.230 120.730 ;
        RECT 34.905 120.560 35.075 121.530 ;
        RECT 34.400 120.230 34.655 120.560 ;
        RECT 34.880 120.230 35.075 120.560 ;
        RECT 35.245 121.190 36.370 121.360 ;
        RECT 34.485 120.060 34.655 120.230 ;
        RECT 35.245 120.060 35.415 121.190 ;
        RECT 34.060 119.490 34.315 120.060 ;
        RECT 34.485 119.890 35.415 120.060 ;
        RECT 35.585 120.850 36.595 121.020 ;
        RECT 35.585 120.050 35.755 120.850 ;
        RECT 35.960 120.170 36.235 120.650 ;
        RECT 35.955 120.000 36.235 120.170 ;
        RECT 35.240 119.855 35.415 119.890 ;
        RECT 34.485 119.320 34.815 119.720 ;
        RECT 35.240 119.490 35.770 119.855 ;
        RECT 35.960 119.490 36.235 120.000 ;
        RECT 36.405 119.490 36.595 120.850 ;
        RECT 36.765 120.865 36.935 121.530 ;
        RECT 37.105 121.110 37.275 121.870 ;
        RECT 37.510 121.110 38.025 121.520 ;
        RECT 36.765 120.675 37.515 120.865 ;
        RECT 37.685 120.300 38.025 121.110 ;
        RECT 38.195 120.705 38.485 121.870 ;
        RECT 38.855 121.200 39.135 121.870 ;
        RECT 39.305 120.980 39.605 121.530 ;
        RECT 39.805 121.150 40.135 121.870 ;
        RECT 40.325 121.150 40.785 121.700 ;
        RECT 38.670 120.560 38.935 120.920 ;
        RECT 39.305 120.810 40.245 120.980 ;
        RECT 40.075 120.560 40.245 120.810 ;
        RECT 38.670 120.310 39.345 120.560 ;
        RECT 39.565 120.310 39.905 120.560 ;
        RECT 36.795 120.130 38.025 120.300 ;
        RECT 40.075 120.230 40.365 120.560 ;
        RECT 40.075 120.140 40.245 120.230 ;
        RECT 36.775 119.320 37.285 119.855 ;
        RECT 37.505 119.525 37.750 120.130 ;
        RECT 38.195 119.320 38.485 120.045 ;
        RECT 38.855 119.950 40.245 120.140 ;
        RECT 38.855 119.590 39.185 119.950 ;
        RECT 40.535 119.780 40.785 121.150 ;
        RECT 41.330 120.890 41.585 121.560 ;
        RECT 41.765 121.070 42.050 121.870 ;
        RECT 42.230 121.150 42.560 121.660 ;
        RECT 41.330 120.510 41.510 120.890 ;
        RECT 42.230 120.560 42.480 121.150 ;
        RECT 42.830 121.000 43.000 121.610 ;
        RECT 43.170 121.180 43.500 121.870 ;
        RECT 43.730 121.320 43.970 121.610 ;
        RECT 44.170 121.490 44.590 121.870 ;
        RECT 44.770 121.400 45.400 121.650 ;
        RECT 45.870 121.490 46.200 121.870 ;
        RECT 44.770 121.320 44.940 121.400 ;
        RECT 46.370 121.320 46.540 121.610 ;
        RECT 46.720 121.490 47.100 121.870 ;
        RECT 47.340 121.485 48.170 121.655 ;
        RECT 43.730 121.150 44.940 121.320 ;
        RECT 41.245 120.340 41.510 120.510 ;
        RECT 39.805 119.320 40.055 119.780 ;
        RECT 40.225 119.490 40.785 119.780 ;
        RECT 41.330 120.030 41.510 120.340 ;
        RECT 41.680 120.230 42.480 120.560 ;
        RECT 41.330 119.500 41.585 120.030 ;
        RECT 41.765 119.320 42.050 119.780 ;
        RECT 42.230 119.580 42.480 120.230 ;
        RECT 42.680 120.980 43.000 121.000 ;
        RECT 42.680 120.810 44.600 120.980 ;
        RECT 42.680 119.915 42.870 120.810 ;
        RECT 44.770 120.640 44.940 121.150 ;
        RECT 45.110 120.890 45.630 121.200 ;
        RECT 43.040 120.470 44.940 120.640 ;
        RECT 43.040 120.410 43.370 120.470 ;
        RECT 43.520 120.240 43.850 120.300 ;
        RECT 43.190 119.970 43.850 120.240 ;
        RECT 42.680 119.585 43.000 119.915 ;
        RECT 43.180 119.320 43.840 119.800 ;
        RECT 44.040 119.710 44.210 120.470 ;
        RECT 45.110 120.300 45.290 120.710 ;
        RECT 44.380 120.130 44.710 120.250 ;
        RECT 45.460 120.130 45.630 120.890 ;
        RECT 44.380 119.960 45.630 120.130 ;
        RECT 45.800 121.070 47.170 121.320 ;
        RECT 45.800 120.300 45.990 121.070 ;
        RECT 46.920 120.810 47.170 121.070 ;
        RECT 46.160 120.640 46.410 120.800 ;
        RECT 47.340 120.640 47.510 121.485 ;
        RECT 48.405 121.200 48.575 121.700 ;
        RECT 48.745 121.370 49.075 121.870 ;
        RECT 47.680 120.810 48.180 121.190 ;
        RECT 48.405 121.030 49.100 121.200 ;
        RECT 46.160 120.470 47.510 120.640 ;
        RECT 47.090 120.430 47.510 120.470 ;
        RECT 45.800 119.960 46.220 120.300 ;
        RECT 46.510 119.970 46.920 120.300 ;
        RECT 44.040 119.540 44.890 119.710 ;
        RECT 45.450 119.320 45.770 119.780 ;
        RECT 45.970 119.530 46.220 119.960 ;
        RECT 46.510 119.320 46.920 119.760 ;
        RECT 47.090 119.700 47.260 120.430 ;
        RECT 47.430 119.880 47.780 120.250 ;
        RECT 47.960 119.940 48.180 120.810 ;
        RECT 48.350 120.240 48.760 120.860 ;
        RECT 48.930 120.060 49.100 121.030 ;
        RECT 48.405 119.870 49.100 120.060 ;
        RECT 47.090 119.500 48.105 119.700 ;
        RECT 48.405 119.540 48.575 119.870 ;
        RECT 48.745 119.320 49.075 119.700 ;
        RECT 49.290 119.580 49.515 121.700 ;
        RECT 49.685 121.370 50.015 121.870 ;
        RECT 50.185 121.200 50.355 121.700 ;
        RECT 50.990 121.530 51.245 121.560 ;
        RECT 50.905 121.360 51.245 121.530 ;
        RECT 49.690 121.030 50.355 121.200 ;
        RECT 49.690 120.040 49.920 121.030 ;
        RECT 50.990 120.890 51.245 121.360 ;
        RECT 51.425 121.070 51.710 121.870 ;
        RECT 51.890 121.150 52.220 121.660 ;
        RECT 50.090 120.210 50.440 120.860 ;
        RECT 49.690 119.870 50.355 120.040 ;
        RECT 49.685 119.320 50.015 119.700 ;
        RECT 50.185 119.580 50.355 119.870 ;
        RECT 50.990 120.030 51.170 120.890 ;
        RECT 51.890 120.560 52.140 121.150 ;
        RECT 52.490 121.000 52.660 121.610 ;
        RECT 52.830 121.180 53.160 121.870 ;
        RECT 53.390 121.320 53.630 121.610 ;
        RECT 53.830 121.490 54.250 121.870 ;
        RECT 54.430 121.400 55.060 121.650 ;
        RECT 55.530 121.490 55.860 121.870 ;
        RECT 54.430 121.320 54.600 121.400 ;
        RECT 56.030 121.320 56.200 121.610 ;
        RECT 56.380 121.490 56.760 121.870 ;
        RECT 57.000 121.485 57.830 121.655 ;
        RECT 53.390 121.150 54.600 121.320 ;
        RECT 51.340 120.230 52.140 120.560 ;
        RECT 50.990 119.500 51.245 120.030 ;
        RECT 51.425 119.320 51.710 119.780 ;
        RECT 51.890 119.580 52.140 120.230 ;
        RECT 52.340 120.980 52.660 121.000 ;
        RECT 52.340 120.810 54.260 120.980 ;
        RECT 52.340 119.915 52.530 120.810 ;
        RECT 54.430 120.640 54.600 121.150 ;
        RECT 54.770 120.890 55.290 121.200 ;
        RECT 52.700 120.470 54.600 120.640 ;
        RECT 52.700 120.410 53.030 120.470 ;
        RECT 53.180 120.240 53.510 120.300 ;
        RECT 52.850 119.970 53.510 120.240 ;
        RECT 52.340 119.585 52.660 119.915 ;
        RECT 52.840 119.320 53.500 119.800 ;
        RECT 53.700 119.710 53.870 120.470 ;
        RECT 54.770 120.300 54.950 120.710 ;
        RECT 54.040 120.130 54.370 120.250 ;
        RECT 55.120 120.130 55.290 120.890 ;
        RECT 54.040 119.960 55.290 120.130 ;
        RECT 55.460 121.070 56.830 121.320 ;
        RECT 55.460 120.300 55.650 121.070 ;
        RECT 56.580 120.810 56.830 121.070 ;
        RECT 55.820 120.640 56.070 120.800 ;
        RECT 57.000 120.640 57.170 121.485 ;
        RECT 58.065 121.200 58.235 121.700 ;
        RECT 58.405 121.370 58.735 121.870 ;
        RECT 57.340 120.810 57.840 121.190 ;
        RECT 58.065 121.030 58.760 121.200 ;
        RECT 55.820 120.470 57.170 120.640 ;
        RECT 56.750 120.430 57.170 120.470 ;
        RECT 55.460 119.960 55.880 120.300 ;
        RECT 56.170 119.970 56.580 120.300 ;
        RECT 53.700 119.540 54.550 119.710 ;
        RECT 55.110 119.320 55.430 119.780 ;
        RECT 55.630 119.530 55.880 119.960 ;
        RECT 56.170 119.320 56.580 119.760 ;
        RECT 56.750 119.700 56.920 120.430 ;
        RECT 57.090 119.880 57.440 120.250 ;
        RECT 57.620 119.940 57.840 120.810 ;
        RECT 58.010 120.240 58.420 120.860 ;
        RECT 58.590 120.060 58.760 121.030 ;
        RECT 58.065 119.870 58.760 120.060 ;
        RECT 56.750 119.500 57.765 119.700 ;
        RECT 58.065 119.540 58.235 119.870 ;
        RECT 58.405 119.320 58.735 119.700 ;
        RECT 58.950 119.580 59.175 121.700 ;
        RECT 59.345 121.370 59.675 121.870 ;
        RECT 59.845 121.200 60.015 121.700 ;
        RECT 59.350 121.030 60.015 121.200 ;
        RECT 59.350 120.040 59.580 121.030 ;
        RECT 59.750 120.210 60.100 120.860 ;
        RECT 60.275 120.780 63.785 121.870 ;
        RECT 60.275 120.260 61.965 120.780 ;
        RECT 63.955 120.705 64.245 121.870 ;
        RECT 64.455 120.730 64.685 121.870 ;
        RECT 64.855 120.720 65.185 121.700 ;
        RECT 65.355 120.730 65.565 121.870 ;
        RECT 66.170 121.530 66.425 121.560 ;
        RECT 66.085 121.360 66.425 121.530 ;
        RECT 66.170 120.890 66.425 121.360 ;
        RECT 66.605 121.070 66.890 121.870 ;
        RECT 67.070 121.150 67.400 121.660 ;
        RECT 62.135 120.090 63.785 120.610 ;
        RECT 64.435 120.310 64.765 120.560 ;
        RECT 59.350 119.870 60.015 120.040 ;
        RECT 59.345 119.320 59.675 119.700 ;
        RECT 59.845 119.580 60.015 119.870 ;
        RECT 60.275 119.320 63.785 120.090 ;
        RECT 63.955 119.320 64.245 120.045 ;
        RECT 64.455 119.320 64.685 120.140 ;
        RECT 64.935 120.120 65.185 120.720 ;
        RECT 64.855 119.490 65.185 120.120 ;
        RECT 65.355 119.320 65.565 120.140 ;
        RECT 66.170 120.030 66.350 120.890 ;
        RECT 67.070 120.560 67.320 121.150 ;
        RECT 67.670 121.000 67.840 121.610 ;
        RECT 68.010 121.180 68.340 121.870 ;
        RECT 68.570 121.320 68.810 121.610 ;
        RECT 69.010 121.490 69.430 121.870 ;
        RECT 69.610 121.400 70.240 121.650 ;
        RECT 70.710 121.490 71.040 121.870 ;
        RECT 69.610 121.320 69.780 121.400 ;
        RECT 71.210 121.320 71.380 121.610 ;
        RECT 71.560 121.490 71.940 121.870 ;
        RECT 72.180 121.485 73.010 121.655 ;
        RECT 68.570 121.150 69.780 121.320 ;
        RECT 66.520 120.230 67.320 120.560 ;
        RECT 66.170 119.500 66.425 120.030 ;
        RECT 66.605 119.320 66.890 119.780 ;
        RECT 67.070 119.580 67.320 120.230 ;
        RECT 67.520 120.980 67.840 121.000 ;
        RECT 67.520 120.810 69.440 120.980 ;
        RECT 67.520 119.915 67.710 120.810 ;
        RECT 69.610 120.640 69.780 121.150 ;
        RECT 69.950 120.890 70.470 121.200 ;
        RECT 67.880 120.470 69.780 120.640 ;
        RECT 67.880 120.410 68.210 120.470 ;
        RECT 68.360 120.240 68.690 120.300 ;
        RECT 68.030 119.970 68.690 120.240 ;
        RECT 67.520 119.585 67.840 119.915 ;
        RECT 68.020 119.320 68.680 119.800 ;
        RECT 68.880 119.710 69.050 120.470 ;
        RECT 69.950 120.300 70.130 120.710 ;
        RECT 69.220 120.130 69.550 120.250 ;
        RECT 70.300 120.130 70.470 120.890 ;
        RECT 69.220 119.960 70.470 120.130 ;
        RECT 70.640 121.070 72.010 121.320 ;
        RECT 70.640 120.300 70.830 121.070 ;
        RECT 71.760 120.810 72.010 121.070 ;
        RECT 71.000 120.640 71.250 120.800 ;
        RECT 72.180 120.640 72.350 121.485 ;
        RECT 73.245 121.200 73.415 121.700 ;
        RECT 73.585 121.370 73.915 121.870 ;
        RECT 72.520 120.810 73.020 121.190 ;
        RECT 73.245 121.030 73.940 121.200 ;
        RECT 71.000 120.470 72.350 120.640 ;
        RECT 71.930 120.430 72.350 120.470 ;
        RECT 70.640 119.960 71.060 120.300 ;
        RECT 71.350 119.970 71.760 120.300 ;
        RECT 68.880 119.540 69.730 119.710 ;
        RECT 70.290 119.320 70.610 119.780 ;
        RECT 70.810 119.530 71.060 119.960 ;
        RECT 71.350 119.320 71.760 119.760 ;
        RECT 71.930 119.700 72.100 120.430 ;
        RECT 72.270 119.880 72.620 120.250 ;
        RECT 72.800 119.940 73.020 120.810 ;
        RECT 73.190 120.240 73.600 120.860 ;
        RECT 73.770 120.060 73.940 121.030 ;
        RECT 73.245 119.870 73.940 120.060 ;
        RECT 71.930 119.500 72.945 119.700 ;
        RECT 73.245 119.540 73.415 119.870 ;
        RECT 73.585 119.320 73.915 119.700 ;
        RECT 74.130 119.580 74.355 121.700 ;
        RECT 74.525 121.370 74.855 121.870 ;
        RECT 75.025 121.200 75.195 121.700 ;
        RECT 74.530 121.030 75.195 121.200 ;
        RECT 74.530 120.040 74.760 121.030 ;
        RECT 74.930 120.210 75.280 120.860 ;
        RECT 75.455 120.795 75.725 121.700 ;
        RECT 75.895 121.110 76.225 121.870 ;
        RECT 76.405 120.940 76.575 121.700 ;
        RECT 77.210 121.530 77.465 121.560 ;
        RECT 77.125 121.360 77.465 121.530 ;
        RECT 74.530 119.870 75.195 120.040 ;
        RECT 74.525 119.320 74.855 119.700 ;
        RECT 75.025 119.580 75.195 119.870 ;
        RECT 75.455 119.995 75.625 120.795 ;
        RECT 75.910 120.770 76.575 120.940 ;
        RECT 77.210 120.890 77.465 121.360 ;
        RECT 77.645 121.070 77.930 121.870 ;
        RECT 78.110 121.150 78.440 121.660 ;
        RECT 75.910 120.625 76.080 120.770 ;
        RECT 75.795 120.295 76.080 120.625 ;
        RECT 75.910 120.040 76.080 120.295 ;
        RECT 76.315 120.220 76.645 120.590 ;
        RECT 75.455 119.490 75.715 119.995 ;
        RECT 75.910 119.870 76.575 120.040 ;
        RECT 75.895 119.320 76.225 119.700 ;
        RECT 76.405 119.490 76.575 119.870 ;
        RECT 77.210 120.030 77.390 120.890 ;
        RECT 78.110 120.560 78.360 121.150 ;
        RECT 78.710 121.000 78.880 121.610 ;
        RECT 79.050 121.180 79.380 121.870 ;
        RECT 79.610 121.320 79.850 121.610 ;
        RECT 80.050 121.490 80.470 121.870 ;
        RECT 80.650 121.400 81.280 121.650 ;
        RECT 81.750 121.490 82.080 121.870 ;
        RECT 80.650 121.320 80.820 121.400 ;
        RECT 82.250 121.320 82.420 121.610 ;
        RECT 82.600 121.490 82.980 121.870 ;
        RECT 83.220 121.485 84.050 121.655 ;
        RECT 79.610 121.150 80.820 121.320 ;
        RECT 77.560 120.230 78.360 120.560 ;
        RECT 77.210 119.500 77.465 120.030 ;
        RECT 77.645 119.320 77.930 119.780 ;
        RECT 78.110 119.580 78.360 120.230 ;
        RECT 78.560 120.980 78.880 121.000 ;
        RECT 78.560 120.810 80.480 120.980 ;
        RECT 78.560 119.915 78.750 120.810 ;
        RECT 80.650 120.640 80.820 121.150 ;
        RECT 80.990 120.890 81.510 121.200 ;
        RECT 78.920 120.470 80.820 120.640 ;
        RECT 78.920 120.410 79.250 120.470 ;
        RECT 79.400 120.240 79.730 120.300 ;
        RECT 79.070 119.970 79.730 120.240 ;
        RECT 78.560 119.585 78.880 119.915 ;
        RECT 79.060 119.320 79.720 119.800 ;
        RECT 79.920 119.710 80.090 120.470 ;
        RECT 80.990 120.300 81.170 120.710 ;
        RECT 80.260 120.130 80.590 120.250 ;
        RECT 81.340 120.130 81.510 120.890 ;
        RECT 80.260 119.960 81.510 120.130 ;
        RECT 81.680 121.070 83.050 121.320 ;
        RECT 81.680 120.300 81.870 121.070 ;
        RECT 82.800 120.810 83.050 121.070 ;
        RECT 82.040 120.640 82.290 120.800 ;
        RECT 83.220 120.640 83.390 121.485 ;
        RECT 84.285 121.200 84.455 121.700 ;
        RECT 84.625 121.370 84.955 121.870 ;
        RECT 83.560 120.810 84.060 121.190 ;
        RECT 84.285 121.030 84.980 121.200 ;
        RECT 82.040 120.470 83.390 120.640 ;
        RECT 82.970 120.430 83.390 120.470 ;
        RECT 81.680 119.960 82.100 120.300 ;
        RECT 82.390 119.970 82.800 120.300 ;
        RECT 79.920 119.540 80.770 119.710 ;
        RECT 81.330 119.320 81.650 119.780 ;
        RECT 81.850 119.530 82.100 119.960 ;
        RECT 82.390 119.320 82.800 119.760 ;
        RECT 82.970 119.700 83.140 120.430 ;
        RECT 83.310 119.880 83.660 120.250 ;
        RECT 83.840 119.940 84.060 120.810 ;
        RECT 84.230 120.240 84.640 120.860 ;
        RECT 84.810 120.060 84.980 121.030 ;
        RECT 84.285 119.870 84.980 120.060 ;
        RECT 82.970 119.500 83.985 119.700 ;
        RECT 84.285 119.540 84.455 119.870 ;
        RECT 84.625 119.320 84.955 119.700 ;
        RECT 85.170 119.580 85.395 121.700 ;
        RECT 85.565 121.370 85.895 121.870 ;
        RECT 86.065 121.200 86.235 121.700 ;
        RECT 85.570 121.030 86.235 121.200 ;
        RECT 85.570 120.040 85.800 121.030 ;
        RECT 85.970 120.210 86.320 120.860 ;
        RECT 86.495 120.795 86.765 121.700 ;
        RECT 86.935 121.110 87.265 121.870 ;
        RECT 87.445 120.940 87.615 121.700 ;
        RECT 85.570 119.870 86.235 120.040 ;
        RECT 85.565 119.320 85.895 119.700 ;
        RECT 86.065 119.580 86.235 119.870 ;
        RECT 86.495 119.995 86.665 120.795 ;
        RECT 86.950 120.770 87.615 120.940 ;
        RECT 87.875 120.780 89.545 121.870 ;
        RECT 86.950 120.625 87.120 120.770 ;
        RECT 86.835 120.295 87.120 120.625 ;
        RECT 86.950 120.040 87.120 120.295 ;
        RECT 87.355 120.220 87.685 120.590 ;
        RECT 87.875 120.260 88.625 120.780 ;
        RECT 89.715 120.705 90.005 121.870 ;
        RECT 90.725 120.940 90.895 121.700 ;
        RECT 91.075 121.110 91.405 121.870 ;
        RECT 90.725 120.770 91.390 120.940 ;
        RECT 91.575 120.795 91.845 121.700 ;
        RECT 92.390 121.530 92.645 121.560 ;
        RECT 92.305 121.360 92.645 121.530 ;
        RECT 91.220 120.625 91.390 120.770 ;
        RECT 88.795 120.090 89.545 120.610 ;
        RECT 90.655 120.220 90.985 120.590 ;
        RECT 91.220 120.295 91.505 120.625 ;
        RECT 86.495 119.490 86.755 119.995 ;
        RECT 86.950 119.870 87.615 120.040 ;
        RECT 86.935 119.320 87.265 119.700 ;
        RECT 87.445 119.490 87.615 119.870 ;
        RECT 87.875 119.320 89.545 120.090 ;
        RECT 89.715 119.320 90.005 120.045 ;
        RECT 91.220 120.040 91.390 120.295 ;
        RECT 90.725 119.870 91.390 120.040 ;
        RECT 91.675 119.995 91.845 120.795 ;
        RECT 90.725 119.490 90.895 119.870 ;
        RECT 91.075 119.320 91.405 119.700 ;
        RECT 91.585 119.490 91.845 119.995 ;
        RECT 92.390 120.890 92.645 121.360 ;
        RECT 92.825 121.070 93.110 121.870 ;
        RECT 93.290 121.150 93.620 121.660 ;
        RECT 92.390 120.030 92.570 120.890 ;
        RECT 93.290 120.560 93.540 121.150 ;
        RECT 93.890 121.000 94.060 121.610 ;
        RECT 94.230 121.180 94.560 121.870 ;
        RECT 94.790 121.320 95.030 121.610 ;
        RECT 95.230 121.490 95.650 121.870 ;
        RECT 95.830 121.400 96.460 121.650 ;
        RECT 96.930 121.490 97.260 121.870 ;
        RECT 95.830 121.320 96.000 121.400 ;
        RECT 97.430 121.320 97.600 121.610 ;
        RECT 97.780 121.490 98.160 121.870 ;
        RECT 98.400 121.485 99.230 121.655 ;
        RECT 94.790 121.150 96.000 121.320 ;
        RECT 92.740 120.230 93.540 120.560 ;
        RECT 92.390 119.500 92.645 120.030 ;
        RECT 92.825 119.320 93.110 119.780 ;
        RECT 93.290 119.580 93.540 120.230 ;
        RECT 93.740 120.980 94.060 121.000 ;
        RECT 93.740 120.810 95.660 120.980 ;
        RECT 93.740 119.915 93.930 120.810 ;
        RECT 95.830 120.640 96.000 121.150 ;
        RECT 96.170 120.890 96.690 121.200 ;
        RECT 94.100 120.470 96.000 120.640 ;
        RECT 94.100 120.410 94.430 120.470 ;
        RECT 94.580 120.240 94.910 120.300 ;
        RECT 94.250 119.970 94.910 120.240 ;
        RECT 93.740 119.585 94.060 119.915 ;
        RECT 94.240 119.320 94.900 119.800 ;
        RECT 95.100 119.710 95.270 120.470 ;
        RECT 96.170 120.300 96.350 120.710 ;
        RECT 95.440 120.130 95.770 120.250 ;
        RECT 96.520 120.130 96.690 120.890 ;
        RECT 95.440 119.960 96.690 120.130 ;
        RECT 96.860 121.070 98.230 121.320 ;
        RECT 96.860 120.300 97.050 121.070 ;
        RECT 97.980 120.810 98.230 121.070 ;
        RECT 97.220 120.640 97.470 120.800 ;
        RECT 98.400 120.640 98.570 121.485 ;
        RECT 99.465 121.200 99.635 121.700 ;
        RECT 99.805 121.370 100.135 121.870 ;
        RECT 98.740 120.810 99.240 121.190 ;
        RECT 99.465 121.030 100.160 121.200 ;
        RECT 97.220 120.470 98.570 120.640 ;
        RECT 98.150 120.430 98.570 120.470 ;
        RECT 96.860 119.960 97.280 120.300 ;
        RECT 97.570 119.970 97.980 120.300 ;
        RECT 95.100 119.540 95.950 119.710 ;
        RECT 96.510 119.320 96.830 119.780 ;
        RECT 97.030 119.530 97.280 119.960 ;
        RECT 97.570 119.320 97.980 119.760 ;
        RECT 98.150 119.700 98.320 120.430 ;
        RECT 98.490 119.880 98.840 120.250 ;
        RECT 99.020 119.940 99.240 120.810 ;
        RECT 99.410 120.240 99.820 120.860 ;
        RECT 99.990 120.060 100.160 121.030 ;
        RECT 99.465 119.870 100.160 120.060 ;
        RECT 98.150 119.500 99.165 119.700 ;
        RECT 99.465 119.540 99.635 119.870 ;
        RECT 99.805 119.320 100.135 119.700 ;
        RECT 100.350 119.580 100.575 121.700 ;
        RECT 100.745 121.370 101.075 121.870 ;
        RECT 101.245 121.200 101.415 121.700 ;
        RECT 100.750 121.030 101.415 121.200 ;
        RECT 100.750 120.040 100.980 121.030 ;
        RECT 101.150 120.210 101.500 120.860 ;
        RECT 102.135 120.780 105.645 121.870 ;
        RECT 102.135 120.260 103.825 120.780 ;
        RECT 105.855 120.730 106.085 121.870 ;
        RECT 106.255 120.720 106.585 121.700 ;
        RECT 106.755 120.730 106.965 121.870 ;
        RECT 107.195 120.780 108.865 121.870 ;
        RECT 109.040 121.435 114.385 121.870 ;
        RECT 103.995 120.090 105.645 120.610 ;
        RECT 105.835 120.310 106.165 120.560 ;
        RECT 100.750 119.870 101.415 120.040 ;
        RECT 100.745 119.320 101.075 119.700 ;
        RECT 101.245 119.580 101.415 119.870 ;
        RECT 102.135 119.320 105.645 120.090 ;
        RECT 105.855 119.320 106.085 120.140 ;
        RECT 106.335 120.120 106.585 120.720 ;
        RECT 107.195 120.260 107.945 120.780 ;
        RECT 106.255 119.490 106.585 120.120 ;
        RECT 106.755 119.320 106.965 120.140 ;
        RECT 108.115 120.090 108.865 120.610 ;
        RECT 110.630 120.185 110.980 121.435 ;
        RECT 114.555 120.780 115.765 121.870 ;
        RECT 107.195 119.320 108.865 120.090 ;
        RECT 112.460 119.865 112.800 120.695 ;
        RECT 114.555 120.240 115.075 120.780 ;
        RECT 115.245 120.070 115.765 120.610 ;
        RECT 109.040 119.320 114.385 119.865 ;
        RECT 114.555 119.320 115.765 120.070 ;
        RECT 14.650 119.150 115.850 119.320 ;
        RECT 14.735 118.400 15.945 119.150 ;
        RECT 14.735 117.860 15.255 118.400 ;
        RECT 16.115 118.380 19.625 119.150 ;
        RECT 19.800 118.605 25.145 119.150 ;
        RECT 15.425 117.690 15.945 118.230 ;
        RECT 14.735 116.600 15.945 117.690 ;
        RECT 16.115 117.690 17.805 118.210 ;
        RECT 17.975 117.860 19.625 118.380 ;
        RECT 16.115 116.600 19.625 117.690 ;
        RECT 21.390 117.035 21.740 118.285 ;
        RECT 23.220 117.775 23.560 118.605 ;
        RECT 25.315 118.425 25.605 119.150 ;
        RECT 26.700 118.605 32.045 119.150 ;
        RECT 19.800 116.600 25.145 117.035 ;
        RECT 25.315 116.600 25.605 117.765 ;
        RECT 28.290 117.035 28.640 118.285 ;
        RECT 30.120 117.775 30.460 118.605 ;
        RECT 32.275 118.330 32.485 119.150 ;
        RECT 32.655 118.350 32.985 118.980 ;
        RECT 32.655 117.750 32.905 118.350 ;
        RECT 33.155 118.330 33.385 119.150 ;
        RECT 34.515 118.380 38.025 119.150 ;
        RECT 33.075 117.910 33.405 118.160 ;
        RECT 26.700 116.600 32.045 117.035 ;
        RECT 32.275 116.600 32.485 117.740 ;
        RECT 32.655 116.770 32.985 117.750 ;
        RECT 33.155 116.600 33.385 117.740 ;
        RECT 34.515 117.690 36.205 118.210 ;
        RECT 36.375 117.860 38.025 118.380 ;
        RECT 38.235 118.330 38.465 119.150 ;
        RECT 38.635 118.350 38.965 118.980 ;
        RECT 38.215 117.910 38.545 118.160 ;
        RECT 38.715 117.750 38.965 118.350 ;
        RECT 39.135 118.330 39.345 119.150 ;
        RECT 39.665 118.600 39.835 118.980 ;
        RECT 40.015 118.770 40.345 119.150 ;
        RECT 39.665 118.430 40.330 118.600 ;
        RECT 40.525 118.475 40.785 118.980 ;
        RECT 39.595 117.880 39.925 118.250 ;
        RECT 40.160 118.175 40.330 118.430 ;
        RECT 34.515 116.600 38.025 117.690 ;
        RECT 38.235 116.600 38.465 117.740 ;
        RECT 38.635 116.770 38.965 117.750 ;
        RECT 40.160 117.845 40.445 118.175 ;
        RECT 39.135 116.600 39.345 117.740 ;
        RECT 40.160 117.700 40.330 117.845 ;
        RECT 39.665 117.530 40.330 117.700 ;
        RECT 40.615 117.675 40.785 118.475 ;
        RECT 41.415 118.380 44.005 119.150 ;
        RECT 39.665 116.770 39.835 117.530 ;
        RECT 40.015 116.600 40.345 117.360 ;
        RECT 40.515 116.770 40.785 117.675 ;
        RECT 41.415 117.690 42.625 118.210 ;
        RECT 42.795 117.860 44.005 118.380 ;
        RECT 44.215 118.330 44.445 119.150 ;
        RECT 44.615 118.350 44.945 118.980 ;
        RECT 44.195 117.910 44.525 118.160 ;
        RECT 44.695 117.750 44.945 118.350 ;
        RECT 45.115 118.330 45.325 119.150 ;
        RECT 45.645 118.600 45.815 118.980 ;
        RECT 45.995 118.770 46.325 119.150 ;
        RECT 45.645 118.430 46.310 118.600 ;
        RECT 46.505 118.475 46.765 118.980 ;
        RECT 45.575 117.880 45.905 118.250 ;
        RECT 46.140 118.175 46.310 118.430 ;
        RECT 41.415 116.600 44.005 117.690 ;
        RECT 44.215 116.600 44.445 117.740 ;
        RECT 44.615 116.770 44.945 117.750 ;
        RECT 46.140 117.845 46.425 118.175 ;
        RECT 45.115 116.600 45.325 117.740 ;
        RECT 46.140 117.700 46.310 117.845 ;
        RECT 45.645 117.530 46.310 117.700 ;
        RECT 46.595 117.675 46.765 118.475 ;
        RECT 45.645 116.770 45.815 117.530 ;
        RECT 45.995 116.600 46.325 117.360 ;
        RECT 46.495 116.770 46.765 117.675 ;
        RECT 46.940 118.410 47.195 118.980 ;
        RECT 47.365 118.750 47.695 119.150 ;
        RECT 48.120 118.615 48.650 118.980 ;
        RECT 48.120 118.580 48.295 118.615 ;
        RECT 47.365 118.410 48.295 118.580 ;
        RECT 48.840 118.470 49.115 118.980 ;
        RECT 46.940 117.740 47.110 118.410 ;
        RECT 47.365 118.240 47.535 118.410 ;
        RECT 47.280 117.910 47.535 118.240 ;
        RECT 47.760 117.910 47.955 118.240 ;
        RECT 46.940 116.770 47.275 117.740 ;
        RECT 47.445 116.600 47.615 117.740 ;
        RECT 47.785 116.940 47.955 117.910 ;
        RECT 48.125 117.280 48.295 118.410 ;
        RECT 48.465 117.620 48.635 118.420 ;
        RECT 48.835 118.300 49.115 118.470 ;
        RECT 48.840 117.820 49.115 118.300 ;
        RECT 49.285 117.620 49.475 118.980 ;
        RECT 49.655 118.615 50.165 119.150 ;
        RECT 50.385 118.340 50.630 118.945 ;
        RECT 51.075 118.425 51.365 119.150 ;
        RECT 51.995 118.380 55.505 119.150 ;
        RECT 55.765 118.600 55.935 118.980 ;
        RECT 56.115 118.770 56.445 119.150 ;
        RECT 55.765 118.430 56.430 118.600 ;
        RECT 56.625 118.475 56.885 118.980 ;
        RECT 49.675 118.170 50.905 118.340 ;
        RECT 48.465 117.450 49.475 117.620 ;
        RECT 49.645 117.605 50.395 117.795 ;
        RECT 48.125 117.110 49.250 117.280 ;
        RECT 49.645 116.940 49.815 117.605 ;
        RECT 50.565 117.360 50.905 118.170 ;
        RECT 47.785 116.770 49.815 116.940 ;
        RECT 49.985 116.600 50.155 117.360 ;
        RECT 50.390 116.950 50.905 117.360 ;
        RECT 51.075 116.600 51.365 117.765 ;
        RECT 51.995 117.690 53.685 118.210 ;
        RECT 53.855 117.860 55.505 118.380 ;
        RECT 55.695 117.880 56.025 118.250 ;
        RECT 56.260 118.175 56.430 118.430 ;
        RECT 56.260 117.845 56.545 118.175 ;
        RECT 56.260 117.700 56.430 117.845 ;
        RECT 51.995 116.600 55.505 117.690 ;
        RECT 55.765 117.530 56.430 117.700 ;
        RECT 56.715 117.675 56.885 118.475 ;
        RECT 57.055 118.400 58.265 119.150 ;
        RECT 55.765 116.770 55.935 117.530 ;
        RECT 56.115 116.600 56.445 117.360 ;
        RECT 56.615 116.770 56.885 117.675 ;
        RECT 57.055 117.690 57.575 118.230 ;
        RECT 57.745 117.860 58.265 118.400 ;
        RECT 58.435 118.380 61.945 119.150 ;
        RECT 62.120 118.605 67.465 119.150 ;
        RECT 58.435 117.690 60.125 118.210 ;
        RECT 60.295 117.860 61.945 118.380 ;
        RECT 57.055 116.600 58.265 117.690 ;
        RECT 58.435 116.600 61.945 117.690 ;
        RECT 63.710 117.035 64.060 118.285 ;
        RECT 65.540 117.775 65.880 118.605 ;
        RECT 67.635 118.475 67.895 118.980 ;
        RECT 68.075 118.770 68.405 119.150 ;
        RECT 68.585 118.600 68.755 118.980 ;
        RECT 67.635 117.675 67.805 118.475 ;
        RECT 68.090 118.430 68.755 118.600 ;
        RECT 68.090 118.175 68.260 118.430 ;
        RECT 69.055 118.330 69.285 119.150 ;
        RECT 69.455 118.350 69.785 118.980 ;
        RECT 67.975 117.845 68.260 118.175 ;
        RECT 68.495 117.880 68.825 118.250 ;
        RECT 69.035 117.910 69.365 118.160 ;
        RECT 68.090 117.700 68.260 117.845 ;
        RECT 69.535 117.750 69.785 118.350 ;
        RECT 69.955 118.330 70.165 119.150 ;
        RECT 71.320 118.605 76.665 119.150 ;
        RECT 62.120 116.600 67.465 117.035 ;
        RECT 67.635 116.770 67.905 117.675 ;
        RECT 68.090 117.530 68.755 117.700 ;
        RECT 68.075 116.600 68.405 117.360 ;
        RECT 68.585 116.770 68.755 117.530 ;
        RECT 69.055 116.600 69.285 117.740 ;
        RECT 69.455 116.770 69.785 117.750 ;
        RECT 69.955 116.600 70.165 117.740 ;
        RECT 72.910 117.035 73.260 118.285 ;
        RECT 74.740 117.775 75.080 118.605 ;
        RECT 76.835 118.425 77.125 119.150 ;
        RECT 77.755 118.380 80.345 119.150 ;
        RECT 71.320 116.600 76.665 117.035 ;
        RECT 76.835 116.600 77.125 117.765 ;
        RECT 77.755 117.690 78.965 118.210 ;
        RECT 79.135 117.860 80.345 118.380 ;
        RECT 80.575 118.330 80.785 119.150 ;
        RECT 80.955 118.350 81.285 118.980 ;
        RECT 80.955 117.750 81.205 118.350 ;
        RECT 81.455 118.330 81.685 119.150 ;
        RECT 81.895 118.380 83.565 119.150 ;
        RECT 81.375 117.910 81.705 118.160 ;
        RECT 77.755 116.600 80.345 117.690 ;
        RECT 80.575 116.600 80.785 117.740 ;
        RECT 80.955 116.770 81.285 117.750 ;
        RECT 81.455 116.600 81.685 117.740 ;
        RECT 81.895 117.690 82.645 118.210 ;
        RECT 82.815 117.860 83.565 118.380 ;
        RECT 83.775 118.330 84.005 119.150 ;
        RECT 84.175 118.350 84.505 118.980 ;
        RECT 83.755 117.910 84.085 118.160 ;
        RECT 84.255 117.750 84.505 118.350 ;
        RECT 84.675 118.330 84.885 119.150 ;
        RECT 85.115 118.380 87.705 119.150 ;
        RECT 87.880 118.605 93.225 119.150 ;
        RECT 93.400 118.605 98.745 119.150 ;
        RECT 81.895 116.600 83.565 117.690 ;
        RECT 83.775 116.600 84.005 117.740 ;
        RECT 84.175 116.770 84.505 117.750 ;
        RECT 84.675 116.600 84.885 117.740 ;
        RECT 85.115 117.690 86.325 118.210 ;
        RECT 86.495 117.860 87.705 118.380 ;
        RECT 85.115 116.600 87.705 117.690 ;
        RECT 89.470 117.035 89.820 118.285 ;
        RECT 91.300 117.775 91.640 118.605 ;
        RECT 94.990 117.035 95.340 118.285 ;
        RECT 96.820 117.775 97.160 118.605 ;
        RECT 98.915 118.475 99.175 118.980 ;
        RECT 99.355 118.770 99.685 119.150 ;
        RECT 99.865 118.600 100.035 118.980 ;
        RECT 98.915 117.675 99.085 118.475 ;
        RECT 99.370 118.430 100.035 118.600 ;
        RECT 99.370 118.175 99.540 118.430 ;
        RECT 100.755 118.380 102.425 119.150 ;
        RECT 102.595 118.425 102.885 119.150 ;
        RECT 103.055 118.400 104.265 119.150 ;
        RECT 99.255 117.845 99.540 118.175 ;
        RECT 99.775 117.880 100.105 118.250 ;
        RECT 99.370 117.700 99.540 117.845 ;
        RECT 87.880 116.600 93.225 117.035 ;
        RECT 93.400 116.600 98.745 117.035 ;
        RECT 98.915 116.770 99.185 117.675 ;
        RECT 99.370 117.530 100.035 117.700 ;
        RECT 99.355 116.600 99.685 117.360 ;
        RECT 99.865 116.770 100.035 117.530 ;
        RECT 100.755 117.690 101.505 118.210 ;
        RECT 101.675 117.860 102.425 118.380 ;
        RECT 100.755 116.600 102.425 117.690 ;
        RECT 102.595 116.600 102.885 117.765 ;
        RECT 103.055 117.690 103.575 118.230 ;
        RECT 103.745 117.860 104.265 118.400 ;
        RECT 104.435 118.380 107.945 119.150 ;
        RECT 104.435 117.690 106.125 118.210 ;
        RECT 106.295 117.860 107.945 118.380 ;
        RECT 108.155 118.330 108.385 119.150 ;
        RECT 108.555 118.350 108.885 118.980 ;
        RECT 108.135 117.910 108.465 118.160 ;
        RECT 108.635 117.750 108.885 118.350 ;
        RECT 109.055 118.330 109.265 119.150 ;
        RECT 109.495 118.475 109.755 118.980 ;
        RECT 109.935 118.770 110.265 119.150 ;
        RECT 110.445 118.600 110.615 118.980 ;
        RECT 103.055 116.600 104.265 117.690 ;
        RECT 104.435 116.600 107.945 117.690 ;
        RECT 108.155 116.600 108.385 117.740 ;
        RECT 108.555 116.770 108.885 117.750 ;
        RECT 109.055 116.600 109.265 117.740 ;
        RECT 109.495 117.675 109.665 118.475 ;
        RECT 109.950 118.430 110.615 118.600 ;
        RECT 110.875 118.475 111.135 118.980 ;
        RECT 111.315 118.770 111.645 119.150 ;
        RECT 111.825 118.600 111.995 118.980 ;
        RECT 109.950 118.175 110.120 118.430 ;
        RECT 109.835 117.845 110.120 118.175 ;
        RECT 110.355 117.880 110.685 118.250 ;
        RECT 109.950 117.700 110.120 117.845 ;
        RECT 109.495 116.770 109.765 117.675 ;
        RECT 109.950 117.530 110.615 117.700 ;
        RECT 109.935 116.600 110.265 117.360 ;
        RECT 110.445 116.770 110.615 117.530 ;
        RECT 110.875 117.675 111.045 118.475 ;
        RECT 111.330 118.430 111.995 118.600 ;
        RECT 113.175 118.475 113.435 118.980 ;
        RECT 113.615 118.770 113.945 119.150 ;
        RECT 114.125 118.600 114.295 118.980 ;
        RECT 111.330 118.175 111.500 118.430 ;
        RECT 111.215 117.845 111.500 118.175 ;
        RECT 111.735 117.880 112.065 118.250 ;
        RECT 111.330 117.700 111.500 117.845 ;
        RECT 110.875 116.770 111.145 117.675 ;
        RECT 111.330 117.530 111.995 117.700 ;
        RECT 111.315 116.600 111.645 117.360 ;
        RECT 111.825 116.770 111.995 117.530 ;
        RECT 113.175 117.675 113.355 118.475 ;
        RECT 113.630 118.430 114.295 118.600 ;
        RECT 113.630 118.175 113.800 118.430 ;
        RECT 114.555 118.400 115.765 119.150 ;
        RECT 113.525 117.845 113.800 118.175 ;
        RECT 114.025 117.880 114.365 118.250 ;
        RECT 113.630 117.700 113.800 117.845 ;
        RECT 113.175 116.770 113.445 117.675 ;
        RECT 113.630 117.530 114.305 117.700 ;
        RECT 113.615 116.600 113.945 117.360 ;
        RECT 114.125 116.770 114.305 117.530 ;
        RECT 114.555 117.690 115.075 118.230 ;
        RECT 115.245 117.860 115.765 118.400 ;
        RECT 114.555 116.600 115.765 117.690 ;
        RECT 14.650 116.430 115.850 116.600 ;
        RECT 14.735 115.340 15.945 116.430 ;
        RECT 17.345 115.590 17.515 116.430 ;
        RECT 17.725 115.420 17.975 116.260 ;
        RECT 18.185 115.590 18.355 116.430 ;
        RECT 18.525 115.420 18.815 116.260 ;
        RECT 14.735 114.630 15.255 115.170 ;
        RECT 15.425 114.800 15.945 115.340 ;
        RECT 17.090 115.250 18.815 115.420 ;
        RECT 19.025 115.370 19.195 116.430 ;
        RECT 19.490 116.050 19.820 116.430 ;
        RECT 20.000 115.880 20.170 116.170 ;
        RECT 20.340 115.970 20.590 116.430 ;
        RECT 19.370 115.710 20.170 115.880 ;
        RECT 20.760 115.920 21.630 116.260 ;
        RECT 17.090 114.700 17.500 115.250 ;
        RECT 19.370 115.090 19.540 115.710 ;
        RECT 20.760 115.540 20.930 115.920 ;
        RECT 21.865 115.800 22.035 116.260 ;
        RECT 22.205 115.970 22.575 116.430 ;
        RECT 22.870 115.830 23.040 116.170 ;
        RECT 23.210 116.000 23.540 116.430 ;
        RECT 23.775 115.830 23.945 116.170 ;
        RECT 19.710 115.370 20.930 115.540 ;
        RECT 21.100 115.460 21.560 115.750 ;
        RECT 21.865 115.630 22.425 115.800 ;
        RECT 22.870 115.660 23.945 115.830 ;
        RECT 24.115 115.930 24.795 116.260 ;
        RECT 25.010 115.930 25.260 116.260 ;
        RECT 25.430 115.970 25.680 116.430 ;
        RECT 22.255 115.490 22.425 115.630 ;
        RECT 21.100 115.450 22.065 115.460 ;
        RECT 20.760 115.280 20.930 115.370 ;
        RECT 21.390 115.290 22.065 115.450 ;
        RECT 19.370 115.080 19.715 115.090 ;
        RECT 17.685 114.870 19.715 115.080 ;
        RECT 14.735 113.880 15.945 114.630 ;
        RECT 17.090 114.530 18.855 114.700 ;
        RECT 17.345 113.880 17.515 114.350 ;
        RECT 17.685 114.050 18.015 114.530 ;
        RECT 18.185 113.880 18.355 114.350 ;
        RECT 18.525 114.050 18.855 114.530 ;
        RECT 19.025 113.880 19.195 114.690 ;
        RECT 19.390 114.615 19.715 114.870 ;
        RECT 19.395 114.260 19.715 114.615 ;
        RECT 19.885 114.830 20.425 115.200 ;
        RECT 20.760 115.110 21.165 115.280 ;
        RECT 19.885 114.430 20.125 114.830 ;
        RECT 20.605 114.660 20.825 114.940 ;
        RECT 20.295 114.490 20.825 114.660 ;
        RECT 20.295 114.260 20.465 114.490 ;
        RECT 20.995 114.330 21.165 115.110 ;
        RECT 21.335 114.500 21.685 115.120 ;
        RECT 21.855 114.500 22.065 115.290 ;
        RECT 22.255 115.320 23.755 115.490 ;
        RECT 22.255 114.630 22.425 115.320 ;
        RECT 24.115 115.150 24.285 115.930 ;
        RECT 25.090 115.800 25.260 115.930 ;
        RECT 22.595 114.980 24.285 115.150 ;
        RECT 24.455 115.370 24.920 115.760 ;
        RECT 25.090 115.630 25.485 115.800 ;
        RECT 22.595 114.800 22.765 114.980 ;
        RECT 19.395 114.090 20.465 114.260 ;
        RECT 20.635 113.880 20.825 114.320 ;
        RECT 20.995 114.050 21.945 114.330 ;
        RECT 22.255 114.240 22.515 114.630 ;
        RECT 22.935 114.560 23.725 114.810 ;
        RECT 22.165 114.070 22.515 114.240 ;
        RECT 22.725 113.880 23.055 114.340 ;
        RECT 23.930 114.270 24.100 114.980 ;
        RECT 24.455 114.780 24.625 115.370 ;
        RECT 24.270 114.560 24.625 114.780 ;
        RECT 24.795 114.560 25.145 115.180 ;
        RECT 25.315 114.270 25.485 115.630 ;
        RECT 25.850 115.460 26.175 116.245 ;
        RECT 25.655 114.410 26.115 115.460 ;
        RECT 23.930 114.100 24.785 114.270 ;
        RECT 24.990 114.100 25.485 114.270 ;
        RECT 25.655 113.880 25.985 114.240 ;
        RECT 26.345 114.140 26.515 116.260 ;
        RECT 26.685 115.930 27.015 116.430 ;
        RECT 27.185 115.760 27.440 116.260 ;
        RECT 26.690 115.590 27.440 115.760 ;
        RECT 26.690 114.600 26.920 115.590 ;
        RECT 27.090 114.770 27.440 115.420 ;
        RECT 28.115 115.290 28.345 116.430 ;
        RECT 28.515 115.280 28.845 116.260 ;
        RECT 29.015 115.290 29.225 116.430 ;
        RECT 29.455 115.355 29.725 116.260 ;
        RECT 29.895 115.670 30.225 116.430 ;
        RECT 30.405 115.500 30.575 116.260 ;
        RECT 28.095 114.870 28.425 115.120 ;
        RECT 26.690 114.430 27.440 114.600 ;
        RECT 26.685 113.880 27.015 114.260 ;
        RECT 27.185 114.140 27.440 114.430 ;
        RECT 28.115 113.880 28.345 114.700 ;
        RECT 28.595 114.680 28.845 115.280 ;
        RECT 28.515 114.050 28.845 114.680 ;
        RECT 29.015 113.880 29.225 114.700 ;
        RECT 29.455 114.555 29.625 115.355 ;
        RECT 29.910 115.330 30.575 115.500 ;
        RECT 31.295 115.355 31.565 116.260 ;
        RECT 31.735 115.670 32.065 116.430 ;
        RECT 32.245 115.500 32.415 116.260 ;
        RECT 29.910 115.185 30.080 115.330 ;
        RECT 29.795 114.855 30.080 115.185 ;
        RECT 29.910 114.600 30.080 114.855 ;
        RECT 30.315 114.780 30.645 115.150 ;
        RECT 29.455 114.050 29.715 114.555 ;
        RECT 29.910 114.430 30.575 114.600 ;
        RECT 29.895 113.880 30.225 114.260 ;
        RECT 30.405 114.050 30.575 114.430 ;
        RECT 31.295 114.555 31.465 115.355 ;
        RECT 31.750 115.330 32.415 115.500 ;
        RECT 33.225 115.500 33.395 116.260 ;
        RECT 33.575 115.670 33.905 116.430 ;
        RECT 33.225 115.330 33.890 115.500 ;
        RECT 34.075 115.355 34.345 116.260 ;
        RECT 31.750 115.185 31.920 115.330 ;
        RECT 31.635 114.855 31.920 115.185 ;
        RECT 33.720 115.185 33.890 115.330 ;
        RECT 31.750 114.600 31.920 114.855 ;
        RECT 32.155 114.780 32.485 115.150 ;
        RECT 33.155 114.780 33.485 115.150 ;
        RECT 33.720 114.855 34.005 115.185 ;
        RECT 33.720 114.600 33.890 114.855 ;
        RECT 31.295 114.050 31.555 114.555 ;
        RECT 31.750 114.430 32.415 114.600 ;
        RECT 31.735 113.880 32.065 114.260 ;
        RECT 32.245 114.050 32.415 114.430 ;
        RECT 33.225 114.430 33.890 114.600 ;
        RECT 34.175 114.555 34.345 115.355 ;
        RECT 34.515 115.340 38.025 116.430 ;
        RECT 34.515 114.820 36.205 115.340 ;
        RECT 38.195 115.265 38.485 116.430 ;
        RECT 39.115 115.340 41.705 116.430 ;
        RECT 41.880 115.995 47.225 116.430 ;
        RECT 36.375 114.650 38.025 115.170 ;
        RECT 39.115 114.820 40.325 115.340 ;
        RECT 40.495 114.650 41.705 115.170 ;
        RECT 43.470 114.745 43.820 115.995 ;
        RECT 47.485 115.500 47.655 116.260 ;
        RECT 47.835 115.670 48.165 116.430 ;
        RECT 47.485 115.330 48.150 115.500 ;
        RECT 48.335 115.355 48.605 116.260 ;
        RECT 33.225 114.050 33.395 114.430 ;
        RECT 33.575 113.880 33.905 114.260 ;
        RECT 34.085 114.050 34.345 114.555 ;
        RECT 34.515 113.880 38.025 114.650 ;
        RECT 38.195 113.880 38.485 114.605 ;
        RECT 39.115 113.880 41.705 114.650 ;
        RECT 45.300 114.425 45.640 115.255 ;
        RECT 47.980 115.185 48.150 115.330 ;
        RECT 47.415 114.780 47.745 115.150 ;
        RECT 47.980 114.855 48.265 115.185 ;
        RECT 47.980 114.600 48.150 114.855 ;
        RECT 47.485 114.430 48.150 114.600 ;
        RECT 48.435 114.555 48.605 115.355 ;
        RECT 49.235 115.340 51.825 116.430 ;
        RECT 52.000 115.995 57.345 116.430 ;
        RECT 49.235 114.820 50.445 115.340 ;
        RECT 50.615 114.650 51.825 115.170 ;
        RECT 53.590 114.745 53.940 115.995 ;
        RECT 57.525 115.450 57.855 116.260 ;
        RECT 58.025 115.630 58.265 116.430 ;
        RECT 57.525 115.280 58.240 115.450 ;
        RECT 41.880 113.880 47.225 114.425 ;
        RECT 47.485 114.050 47.655 114.430 ;
        RECT 47.835 113.880 48.165 114.260 ;
        RECT 48.345 114.050 48.605 114.555 ;
        RECT 49.235 113.880 51.825 114.650 ;
        RECT 55.420 114.425 55.760 115.255 ;
        RECT 57.520 114.870 57.900 115.110 ;
        RECT 58.070 115.040 58.240 115.280 ;
        RECT 58.445 115.410 58.615 116.260 ;
        RECT 58.785 115.630 59.115 116.430 ;
        RECT 59.285 115.410 59.455 116.260 ;
        RECT 58.445 115.240 59.455 115.410 ;
        RECT 59.625 115.280 59.955 116.430 ;
        RECT 60.275 115.340 63.785 116.430 ;
        RECT 58.070 114.870 58.570 115.040 ;
        RECT 58.070 114.700 58.240 114.870 ;
        RECT 58.960 114.700 59.455 115.240 ;
        RECT 60.275 114.820 61.965 115.340 ;
        RECT 63.955 115.265 64.245 116.430 ;
        RECT 64.875 115.340 68.385 116.430 ;
        RECT 57.605 114.530 58.240 114.700 ;
        RECT 58.445 114.530 59.455 114.700 ;
        RECT 52.000 113.880 57.345 114.425 ;
        RECT 57.605 114.050 57.775 114.530 ;
        RECT 57.955 113.880 58.195 114.360 ;
        RECT 58.445 114.050 58.615 114.530 ;
        RECT 58.785 113.880 59.115 114.360 ;
        RECT 59.285 114.050 59.455 114.530 ;
        RECT 59.625 113.880 59.955 114.680 ;
        RECT 62.135 114.650 63.785 115.170 ;
        RECT 64.875 114.820 66.565 115.340 ;
        RECT 68.615 115.290 68.825 116.430 ;
        RECT 68.995 115.280 69.325 116.260 ;
        RECT 69.495 115.290 69.725 116.430 ;
        RECT 70.025 115.500 70.195 116.260 ;
        RECT 70.375 115.670 70.705 116.430 ;
        RECT 70.025 115.330 70.690 115.500 ;
        RECT 70.875 115.355 71.145 116.260 ;
        RECT 66.735 114.650 68.385 115.170 ;
        RECT 60.275 113.880 63.785 114.650 ;
        RECT 63.955 113.880 64.245 114.605 ;
        RECT 64.875 113.880 68.385 114.650 ;
        RECT 68.615 113.880 68.825 114.700 ;
        RECT 68.995 114.680 69.245 115.280 ;
        RECT 70.520 115.185 70.690 115.330 ;
        RECT 69.415 114.870 69.745 115.120 ;
        RECT 69.955 114.780 70.285 115.150 ;
        RECT 70.520 114.855 70.805 115.185 ;
        RECT 68.995 114.050 69.325 114.680 ;
        RECT 69.495 113.880 69.725 114.700 ;
        RECT 70.520 114.600 70.690 114.855 ;
        RECT 70.025 114.430 70.690 114.600 ;
        RECT 70.975 114.555 71.145 115.355 ;
        RECT 71.375 115.290 71.585 116.430 ;
        RECT 71.755 115.280 72.085 116.260 ;
        RECT 72.255 115.290 72.485 116.430 ;
        RECT 73.625 115.450 73.955 116.260 ;
        RECT 74.125 115.630 74.365 116.430 ;
        RECT 73.625 115.280 74.340 115.450 ;
        RECT 70.025 114.050 70.195 114.430 ;
        RECT 70.375 113.880 70.705 114.260 ;
        RECT 70.885 114.050 71.145 114.555 ;
        RECT 71.375 113.880 71.585 114.700 ;
        RECT 71.755 114.680 72.005 115.280 ;
        RECT 72.175 114.870 72.505 115.120 ;
        RECT 73.620 114.870 74.000 115.110 ;
        RECT 74.170 115.040 74.340 115.280 ;
        RECT 74.545 115.410 74.715 116.260 ;
        RECT 74.885 115.630 75.215 116.430 ;
        RECT 75.385 115.410 75.555 116.260 ;
        RECT 74.545 115.240 75.555 115.410 ;
        RECT 75.725 115.280 76.055 116.430 ;
        RECT 77.295 115.340 80.805 116.430 ;
        RECT 80.980 115.995 86.325 116.430 ;
        RECT 74.170 114.870 74.670 115.040 ;
        RECT 74.170 114.700 74.340 114.870 ;
        RECT 75.060 114.730 75.555 115.240 ;
        RECT 77.295 114.820 78.985 115.340 ;
        RECT 75.055 114.700 75.555 114.730 ;
        RECT 71.755 114.050 72.085 114.680 ;
        RECT 72.255 113.880 72.485 114.700 ;
        RECT 73.705 114.530 74.340 114.700 ;
        RECT 74.545 114.530 75.555 114.700 ;
        RECT 73.705 114.050 73.875 114.530 ;
        RECT 74.055 113.880 74.295 114.360 ;
        RECT 74.545 114.050 74.715 114.530 ;
        RECT 74.885 113.880 75.215 114.360 ;
        RECT 75.385 114.050 75.555 114.530 ;
        RECT 75.725 113.880 76.055 114.680 ;
        RECT 79.155 114.650 80.805 115.170 ;
        RECT 82.570 114.745 82.920 115.995 ;
        RECT 86.585 115.500 86.755 116.260 ;
        RECT 86.935 115.670 87.265 116.430 ;
        RECT 86.585 115.330 87.250 115.500 ;
        RECT 87.435 115.355 87.705 116.260 ;
        RECT 77.295 113.880 80.805 114.650 ;
        RECT 84.400 114.425 84.740 115.255 ;
        RECT 87.080 115.185 87.250 115.330 ;
        RECT 86.515 114.780 86.845 115.150 ;
        RECT 87.080 114.855 87.365 115.185 ;
        RECT 87.080 114.600 87.250 114.855 ;
        RECT 86.585 114.430 87.250 114.600 ;
        RECT 87.535 114.555 87.705 115.355 ;
        RECT 87.875 115.340 89.545 116.430 ;
        RECT 87.875 114.820 88.625 115.340 ;
        RECT 89.715 115.265 90.005 116.430 ;
        RECT 90.175 115.340 91.845 116.430 ;
        RECT 92.105 115.500 92.275 116.260 ;
        RECT 92.455 115.670 92.785 116.430 ;
        RECT 88.795 114.650 89.545 115.170 ;
        RECT 90.175 114.820 90.925 115.340 ;
        RECT 92.105 115.330 92.770 115.500 ;
        RECT 92.955 115.355 93.225 116.260 ;
        RECT 92.600 115.185 92.770 115.330 ;
        RECT 91.095 114.650 91.845 115.170 ;
        RECT 92.035 114.780 92.365 115.150 ;
        RECT 92.600 114.855 92.885 115.185 ;
        RECT 80.980 113.880 86.325 114.425 ;
        RECT 86.585 114.050 86.755 114.430 ;
        RECT 86.935 113.880 87.265 114.260 ;
        RECT 87.445 114.050 87.705 114.555 ;
        RECT 87.875 113.880 89.545 114.650 ;
        RECT 89.715 113.880 90.005 114.605 ;
        RECT 90.175 113.880 91.845 114.650 ;
        RECT 92.600 114.600 92.770 114.855 ;
        RECT 92.105 114.430 92.770 114.600 ;
        RECT 93.055 114.555 93.225 115.355 ;
        RECT 93.395 115.340 96.905 116.430 ;
        RECT 97.165 115.500 97.335 116.260 ;
        RECT 97.515 115.670 97.845 116.430 ;
        RECT 93.395 114.820 95.085 115.340 ;
        RECT 97.165 115.330 97.830 115.500 ;
        RECT 98.015 115.355 98.285 116.260 ;
        RECT 97.660 115.185 97.830 115.330 ;
        RECT 95.255 114.650 96.905 115.170 ;
        RECT 97.095 114.780 97.425 115.150 ;
        RECT 97.660 114.855 97.945 115.185 ;
        RECT 92.105 114.050 92.275 114.430 ;
        RECT 92.455 113.880 92.785 114.260 ;
        RECT 92.965 114.050 93.225 114.555 ;
        RECT 93.395 113.880 96.905 114.650 ;
        RECT 97.660 114.600 97.830 114.855 ;
        RECT 97.165 114.430 97.830 114.600 ;
        RECT 98.115 114.555 98.285 115.355 ;
        RECT 99.005 115.500 99.175 116.260 ;
        RECT 99.355 115.670 99.685 116.430 ;
        RECT 99.005 115.330 99.670 115.500 ;
        RECT 99.855 115.355 100.125 116.260 ;
        RECT 99.500 115.185 99.670 115.330 ;
        RECT 98.935 114.780 99.265 115.150 ;
        RECT 99.500 114.855 99.785 115.185 ;
        RECT 99.500 114.600 99.670 114.855 ;
        RECT 97.165 114.050 97.335 114.430 ;
        RECT 97.515 113.880 97.845 114.260 ;
        RECT 98.025 114.050 98.285 114.555 ;
        RECT 99.005 114.430 99.670 114.600 ;
        RECT 99.955 114.555 100.125 115.355 ;
        RECT 100.385 115.500 100.555 116.260 ;
        RECT 100.735 115.670 101.065 116.430 ;
        RECT 100.385 115.330 101.050 115.500 ;
        RECT 101.235 115.355 101.505 116.260 ;
        RECT 100.880 115.185 101.050 115.330 ;
        RECT 100.315 114.780 100.645 115.150 ;
        RECT 100.880 114.855 101.165 115.185 ;
        RECT 100.880 114.600 101.050 114.855 ;
        RECT 99.005 114.050 99.175 114.430 ;
        RECT 99.355 113.880 99.685 114.260 ;
        RECT 99.865 114.050 100.125 114.555 ;
        RECT 100.385 114.430 101.050 114.600 ;
        RECT 101.335 114.555 101.505 115.355 ;
        RECT 102.135 115.340 103.805 116.430 ;
        RECT 103.980 115.760 104.235 116.260 ;
        RECT 104.405 115.930 104.735 116.430 ;
        RECT 103.980 115.590 104.730 115.760 ;
        RECT 102.135 114.820 102.885 115.340 ;
        RECT 103.055 114.650 103.805 115.170 ;
        RECT 103.980 114.770 104.330 115.420 ;
        RECT 100.385 114.050 100.555 114.430 ;
        RECT 100.735 113.880 101.065 114.260 ;
        RECT 101.245 114.050 101.505 114.555 ;
        RECT 102.135 113.880 103.805 114.650 ;
        RECT 104.500 114.600 104.730 115.590 ;
        RECT 103.980 114.430 104.730 114.600 ;
        RECT 103.980 114.140 104.235 114.430 ;
        RECT 104.405 113.880 104.735 114.260 ;
        RECT 104.905 114.140 105.075 116.260 ;
        RECT 105.245 115.460 105.570 116.245 ;
        RECT 105.740 115.970 105.990 116.430 ;
        RECT 106.160 115.930 106.410 116.260 ;
        RECT 106.625 115.930 107.305 116.260 ;
        RECT 106.160 115.800 106.330 115.930 ;
        RECT 105.935 115.630 106.330 115.800 ;
        RECT 105.305 114.410 105.765 115.460 ;
        RECT 105.935 114.270 106.105 115.630 ;
        RECT 106.500 115.370 106.965 115.760 ;
        RECT 106.275 114.560 106.625 115.180 ;
        RECT 106.795 114.780 106.965 115.370 ;
        RECT 107.135 115.150 107.305 115.930 ;
        RECT 107.475 115.830 107.645 116.170 ;
        RECT 107.880 116.000 108.210 116.430 ;
        RECT 108.380 115.830 108.550 116.170 ;
        RECT 108.845 115.970 109.215 116.430 ;
        RECT 107.475 115.660 108.550 115.830 ;
        RECT 109.385 115.800 109.555 116.260 ;
        RECT 109.790 115.920 110.660 116.260 ;
        RECT 110.830 115.970 111.080 116.430 ;
        RECT 108.995 115.630 109.555 115.800 ;
        RECT 108.995 115.490 109.165 115.630 ;
        RECT 107.665 115.320 109.165 115.490 ;
        RECT 109.860 115.460 110.320 115.750 ;
        RECT 107.135 114.980 108.825 115.150 ;
        RECT 106.795 114.560 107.150 114.780 ;
        RECT 107.320 114.270 107.490 114.980 ;
        RECT 107.695 114.560 108.485 114.810 ;
        RECT 108.655 114.800 108.825 114.980 ;
        RECT 108.995 114.630 109.165 115.320 ;
        RECT 105.435 113.880 105.765 114.240 ;
        RECT 105.935 114.100 106.430 114.270 ;
        RECT 106.635 114.100 107.490 114.270 ;
        RECT 108.365 113.880 108.695 114.340 ;
        RECT 108.905 114.240 109.165 114.630 ;
        RECT 109.355 115.450 110.320 115.460 ;
        RECT 110.490 115.540 110.660 115.920 ;
        RECT 111.250 115.880 111.420 116.170 ;
        RECT 111.600 116.050 111.930 116.430 ;
        RECT 111.250 115.710 112.050 115.880 ;
        RECT 109.355 115.290 110.030 115.450 ;
        RECT 110.490 115.370 111.710 115.540 ;
        RECT 109.355 114.500 109.565 115.290 ;
        RECT 110.490 115.280 110.660 115.370 ;
        RECT 109.735 114.500 110.085 115.120 ;
        RECT 110.255 115.110 110.660 115.280 ;
        RECT 110.255 114.330 110.425 115.110 ;
        RECT 110.595 114.660 110.815 114.940 ;
        RECT 110.995 114.830 111.535 115.200 ;
        RECT 111.880 115.090 112.050 115.710 ;
        RECT 112.225 115.370 112.395 116.430 ;
        RECT 112.605 115.420 112.895 116.260 ;
        RECT 113.065 115.590 113.235 116.430 ;
        RECT 113.445 115.420 113.695 116.260 ;
        RECT 113.905 115.590 114.075 116.430 ;
        RECT 112.605 115.250 114.330 115.420 ;
        RECT 110.595 114.490 111.125 114.660 ;
        RECT 108.905 114.070 109.255 114.240 ;
        RECT 109.475 114.050 110.425 114.330 ;
        RECT 110.595 113.880 110.785 114.320 ;
        RECT 110.955 114.260 111.125 114.490 ;
        RECT 111.295 114.430 111.535 114.830 ;
        RECT 111.705 115.080 112.050 115.090 ;
        RECT 111.705 114.870 113.735 115.080 ;
        RECT 111.705 114.615 112.030 114.870 ;
        RECT 113.920 114.700 114.330 115.250 ;
        RECT 114.555 115.340 115.765 116.430 ;
        RECT 114.555 114.800 115.075 115.340 ;
        RECT 111.705 114.260 112.025 114.615 ;
        RECT 110.955 114.090 112.025 114.260 ;
        RECT 112.225 113.880 112.395 114.690 ;
        RECT 112.565 114.530 114.330 114.700 ;
        RECT 115.245 114.630 115.765 115.170 ;
        RECT 112.565 114.050 112.895 114.530 ;
        RECT 113.065 113.880 113.235 114.350 ;
        RECT 113.405 114.050 113.735 114.530 ;
        RECT 113.905 113.880 114.075 114.350 ;
        RECT 114.555 113.880 115.765 114.630 ;
        RECT 14.650 113.710 115.850 113.880 ;
        RECT 14.735 112.960 15.945 113.710 ;
        RECT 14.735 112.420 15.255 112.960 ;
        RECT 16.115 112.940 19.625 113.710 ;
        RECT 15.425 112.250 15.945 112.790 ;
        RECT 14.735 111.160 15.945 112.250 ;
        RECT 16.115 112.250 17.805 112.770 ;
        RECT 17.975 112.420 19.625 112.940 ;
        RECT 19.855 112.890 20.065 113.710 ;
        RECT 20.235 112.910 20.565 113.540 ;
        RECT 20.235 112.310 20.485 112.910 ;
        RECT 20.735 112.890 20.965 113.710 ;
        RECT 21.235 112.890 21.445 113.710 ;
        RECT 21.615 112.910 21.945 113.540 ;
        RECT 20.655 112.470 20.985 112.720 ;
        RECT 21.615 112.310 21.865 112.910 ;
        RECT 22.115 112.890 22.345 113.710 ;
        RECT 22.615 112.890 22.825 113.710 ;
        RECT 22.995 112.910 23.325 113.540 ;
        RECT 22.035 112.470 22.365 112.720 ;
        RECT 22.995 112.310 23.245 112.910 ;
        RECT 23.495 112.890 23.725 113.710 ;
        RECT 24.025 113.160 24.195 113.540 ;
        RECT 24.375 113.330 24.705 113.710 ;
        RECT 24.025 112.990 24.690 113.160 ;
        RECT 24.885 113.035 25.145 113.540 ;
        RECT 23.415 112.470 23.745 112.720 ;
        RECT 23.955 112.440 24.285 112.810 ;
        RECT 24.520 112.735 24.690 112.990 ;
        RECT 24.520 112.405 24.805 112.735 ;
        RECT 16.115 111.160 19.625 112.250 ;
        RECT 19.855 111.160 20.065 112.300 ;
        RECT 20.235 111.330 20.565 112.310 ;
        RECT 20.735 111.160 20.965 112.300 ;
        RECT 21.235 111.160 21.445 112.300 ;
        RECT 21.615 111.330 21.945 112.310 ;
        RECT 22.115 111.160 22.345 112.300 ;
        RECT 22.615 111.160 22.825 112.300 ;
        RECT 22.995 111.330 23.325 112.310 ;
        RECT 23.495 111.160 23.725 112.300 ;
        RECT 24.520 112.260 24.690 112.405 ;
        RECT 24.025 112.090 24.690 112.260 ;
        RECT 24.975 112.235 25.145 113.035 ;
        RECT 25.315 112.985 25.605 113.710 ;
        RECT 26.545 113.240 26.715 113.710 ;
        RECT 26.885 113.060 27.215 113.540 ;
        RECT 27.385 113.240 27.555 113.710 ;
        RECT 27.725 113.060 28.055 113.540 ;
        RECT 26.290 112.890 28.055 113.060 ;
        RECT 28.225 112.900 28.395 113.710 ;
        RECT 28.595 113.330 29.665 113.500 ;
        RECT 28.595 112.975 28.915 113.330 ;
        RECT 26.290 112.340 26.700 112.890 ;
        RECT 28.590 112.720 28.915 112.975 ;
        RECT 26.885 112.510 28.915 112.720 ;
        RECT 28.570 112.500 28.915 112.510 ;
        RECT 29.085 112.760 29.325 113.160 ;
        RECT 29.495 113.100 29.665 113.330 ;
        RECT 29.835 113.270 30.025 113.710 ;
        RECT 30.195 113.260 31.145 113.540 ;
        RECT 31.365 113.350 31.715 113.520 ;
        RECT 29.495 112.930 30.025 113.100 ;
        RECT 24.025 111.330 24.195 112.090 ;
        RECT 24.375 111.160 24.705 111.920 ;
        RECT 24.875 111.330 25.145 112.235 ;
        RECT 25.315 111.160 25.605 112.325 ;
        RECT 26.290 112.170 28.015 112.340 ;
        RECT 26.545 111.160 26.715 112.000 ;
        RECT 26.925 111.330 27.175 112.170 ;
        RECT 27.385 111.160 27.555 112.000 ;
        RECT 27.725 111.330 28.015 112.170 ;
        RECT 28.225 111.160 28.395 112.220 ;
        RECT 28.570 111.880 28.740 112.500 ;
        RECT 29.085 112.390 29.625 112.760 ;
        RECT 29.805 112.650 30.025 112.930 ;
        RECT 30.195 112.480 30.365 113.260 ;
        RECT 29.960 112.310 30.365 112.480 ;
        RECT 30.535 112.470 30.885 113.090 ;
        RECT 29.960 112.220 30.130 112.310 ;
        RECT 31.055 112.300 31.265 113.090 ;
        RECT 28.910 112.050 30.130 112.220 ;
        RECT 30.590 112.140 31.265 112.300 ;
        RECT 28.570 111.710 29.370 111.880 ;
        RECT 28.690 111.160 29.020 111.540 ;
        RECT 29.200 111.420 29.370 111.710 ;
        RECT 29.960 111.670 30.130 112.050 ;
        RECT 30.300 112.130 31.265 112.140 ;
        RECT 31.455 112.960 31.715 113.350 ;
        RECT 31.925 113.250 32.255 113.710 ;
        RECT 33.130 113.320 33.985 113.490 ;
        RECT 34.190 113.320 34.685 113.490 ;
        RECT 34.855 113.350 35.185 113.710 ;
        RECT 31.455 112.270 31.625 112.960 ;
        RECT 31.795 112.610 31.965 112.790 ;
        RECT 32.135 112.780 32.925 113.030 ;
        RECT 33.130 112.610 33.300 113.320 ;
        RECT 33.470 112.810 33.825 113.030 ;
        RECT 31.795 112.440 33.485 112.610 ;
        RECT 30.300 111.840 30.760 112.130 ;
        RECT 31.455 112.100 32.955 112.270 ;
        RECT 31.455 111.960 31.625 112.100 ;
        RECT 31.065 111.790 31.625 111.960 ;
        RECT 29.540 111.160 29.790 111.620 ;
        RECT 29.960 111.330 30.830 111.670 ;
        RECT 31.065 111.330 31.235 111.790 ;
        RECT 32.070 111.760 33.145 111.930 ;
        RECT 31.405 111.160 31.775 111.620 ;
        RECT 32.070 111.420 32.240 111.760 ;
        RECT 32.410 111.160 32.740 111.590 ;
        RECT 32.975 111.420 33.145 111.760 ;
        RECT 33.315 111.660 33.485 112.440 ;
        RECT 33.655 112.220 33.825 112.810 ;
        RECT 33.995 112.410 34.345 113.030 ;
        RECT 33.655 111.830 34.120 112.220 ;
        RECT 34.515 111.960 34.685 113.320 ;
        RECT 34.855 112.130 35.315 113.180 ;
        RECT 34.290 111.790 34.685 111.960 ;
        RECT 34.290 111.660 34.460 111.790 ;
        RECT 33.315 111.330 33.995 111.660 ;
        RECT 34.210 111.330 34.460 111.660 ;
        RECT 34.630 111.160 34.880 111.620 ;
        RECT 35.050 111.345 35.375 112.130 ;
        RECT 35.545 111.330 35.715 113.450 ;
        RECT 35.885 113.330 36.215 113.710 ;
        RECT 36.385 113.160 36.640 113.450 ;
        RECT 35.890 112.990 36.640 113.160 ;
        RECT 37.735 113.035 37.995 113.540 ;
        RECT 38.175 113.330 38.505 113.710 ;
        RECT 38.685 113.160 38.855 113.540 ;
        RECT 35.890 112.000 36.120 112.990 ;
        RECT 36.290 112.170 36.640 112.820 ;
        RECT 37.735 112.235 37.905 113.035 ;
        RECT 38.190 112.990 38.855 113.160 ;
        RECT 39.205 113.160 39.375 113.540 ;
        RECT 39.555 113.330 39.885 113.710 ;
        RECT 39.205 112.990 39.870 113.160 ;
        RECT 40.065 113.035 40.325 113.540 ;
        RECT 40.805 113.240 40.975 113.710 ;
        RECT 41.145 113.060 41.475 113.540 ;
        RECT 41.645 113.240 41.815 113.710 ;
        RECT 41.985 113.060 42.315 113.540 ;
        RECT 38.190 112.735 38.360 112.990 ;
        RECT 38.075 112.405 38.360 112.735 ;
        RECT 38.595 112.440 38.925 112.810 ;
        RECT 39.135 112.440 39.465 112.810 ;
        RECT 39.700 112.735 39.870 112.990 ;
        RECT 38.190 112.260 38.360 112.405 ;
        RECT 39.700 112.405 39.985 112.735 ;
        RECT 39.700 112.260 39.870 112.405 ;
        RECT 35.890 111.830 36.640 112.000 ;
        RECT 35.885 111.160 36.215 111.660 ;
        RECT 36.385 111.330 36.640 111.830 ;
        RECT 37.735 111.330 38.005 112.235 ;
        RECT 38.190 112.090 38.855 112.260 ;
        RECT 38.175 111.160 38.505 111.920 ;
        RECT 38.685 111.330 38.855 112.090 ;
        RECT 39.205 112.090 39.870 112.260 ;
        RECT 40.155 112.235 40.325 113.035 ;
        RECT 39.205 111.330 39.375 112.090 ;
        RECT 39.555 111.160 39.885 111.920 ;
        RECT 40.055 111.330 40.325 112.235 ;
        RECT 40.550 112.890 42.315 113.060 ;
        RECT 42.485 112.900 42.655 113.710 ;
        RECT 42.855 113.330 43.925 113.500 ;
        RECT 42.855 112.975 43.175 113.330 ;
        RECT 40.550 112.340 40.960 112.890 ;
        RECT 42.850 112.720 43.175 112.975 ;
        RECT 41.145 112.510 43.175 112.720 ;
        RECT 42.830 112.500 43.175 112.510 ;
        RECT 43.345 112.760 43.585 113.160 ;
        RECT 43.755 113.100 43.925 113.330 ;
        RECT 44.095 113.270 44.285 113.710 ;
        RECT 44.455 113.260 45.405 113.540 ;
        RECT 45.625 113.350 45.975 113.520 ;
        RECT 43.755 112.930 44.285 113.100 ;
        RECT 40.550 112.170 42.275 112.340 ;
        RECT 40.805 111.160 40.975 112.000 ;
        RECT 41.185 111.330 41.435 112.170 ;
        RECT 41.645 111.160 41.815 112.000 ;
        RECT 41.985 111.330 42.275 112.170 ;
        RECT 42.485 111.160 42.655 112.220 ;
        RECT 42.830 111.880 43.000 112.500 ;
        RECT 43.345 112.390 43.885 112.760 ;
        RECT 44.065 112.650 44.285 112.930 ;
        RECT 44.455 112.480 44.625 113.260 ;
        RECT 44.220 112.310 44.625 112.480 ;
        RECT 44.795 112.470 45.145 113.090 ;
        RECT 44.220 112.220 44.390 112.310 ;
        RECT 45.315 112.300 45.525 113.090 ;
        RECT 43.170 112.050 44.390 112.220 ;
        RECT 44.850 112.140 45.525 112.300 ;
        RECT 42.830 111.710 43.630 111.880 ;
        RECT 42.950 111.160 43.280 111.540 ;
        RECT 43.460 111.420 43.630 111.710 ;
        RECT 44.220 111.670 44.390 112.050 ;
        RECT 44.560 112.130 45.525 112.140 ;
        RECT 45.715 112.960 45.975 113.350 ;
        RECT 46.185 113.250 46.515 113.710 ;
        RECT 47.390 113.320 48.245 113.490 ;
        RECT 48.450 113.320 48.945 113.490 ;
        RECT 49.115 113.350 49.445 113.710 ;
        RECT 45.715 112.270 45.885 112.960 ;
        RECT 46.055 112.610 46.225 112.790 ;
        RECT 46.395 112.780 47.185 113.030 ;
        RECT 47.390 112.610 47.560 113.320 ;
        RECT 47.730 112.810 48.085 113.030 ;
        RECT 46.055 112.440 47.745 112.610 ;
        RECT 44.560 111.840 45.020 112.130 ;
        RECT 45.715 112.100 47.215 112.270 ;
        RECT 45.715 111.960 45.885 112.100 ;
        RECT 45.325 111.790 45.885 111.960 ;
        RECT 43.800 111.160 44.050 111.620 ;
        RECT 44.220 111.330 45.090 111.670 ;
        RECT 45.325 111.330 45.495 111.790 ;
        RECT 46.330 111.760 47.405 111.930 ;
        RECT 45.665 111.160 46.035 111.620 ;
        RECT 46.330 111.420 46.500 111.760 ;
        RECT 46.670 111.160 47.000 111.590 ;
        RECT 47.235 111.420 47.405 111.760 ;
        RECT 47.575 111.660 47.745 112.440 ;
        RECT 47.915 112.220 48.085 112.810 ;
        RECT 48.255 112.410 48.605 113.030 ;
        RECT 47.915 111.830 48.380 112.220 ;
        RECT 48.775 111.960 48.945 113.320 ;
        RECT 49.115 112.130 49.575 113.180 ;
        RECT 48.550 111.790 48.945 111.960 ;
        RECT 48.550 111.660 48.720 111.790 ;
        RECT 47.575 111.330 48.255 111.660 ;
        RECT 48.470 111.330 48.720 111.660 ;
        RECT 48.890 111.160 49.140 111.620 ;
        RECT 49.310 111.345 49.635 112.130 ;
        RECT 49.805 111.330 49.975 113.450 ;
        RECT 50.145 113.330 50.475 113.710 ;
        RECT 50.645 113.160 50.900 113.450 ;
        RECT 50.150 112.990 50.900 113.160 ;
        RECT 50.150 112.000 50.380 112.990 ;
        RECT 51.075 112.985 51.365 113.710 ;
        RECT 52.545 113.160 52.715 113.540 ;
        RECT 52.895 113.330 53.225 113.710 ;
        RECT 52.545 112.990 53.210 113.160 ;
        RECT 53.405 113.035 53.665 113.540 ;
        RECT 54.145 113.240 54.315 113.710 ;
        RECT 54.485 113.060 54.815 113.540 ;
        RECT 54.985 113.240 55.155 113.710 ;
        RECT 55.325 113.060 55.655 113.540 ;
        RECT 50.550 112.170 50.900 112.820 ;
        RECT 52.475 112.440 52.805 112.810 ;
        RECT 53.040 112.735 53.210 112.990 ;
        RECT 53.040 112.405 53.325 112.735 ;
        RECT 50.150 111.830 50.900 112.000 ;
        RECT 50.145 111.160 50.475 111.660 ;
        RECT 50.645 111.330 50.900 111.830 ;
        RECT 51.075 111.160 51.365 112.325 ;
        RECT 53.040 112.260 53.210 112.405 ;
        RECT 52.545 112.090 53.210 112.260 ;
        RECT 53.495 112.235 53.665 113.035 ;
        RECT 52.545 111.330 52.715 112.090 ;
        RECT 52.895 111.160 53.225 111.920 ;
        RECT 53.395 111.330 53.665 112.235 ;
        RECT 53.890 112.890 55.655 113.060 ;
        RECT 55.825 112.900 55.995 113.710 ;
        RECT 56.195 113.330 57.265 113.500 ;
        RECT 56.195 112.975 56.515 113.330 ;
        RECT 53.890 112.340 54.300 112.890 ;
        RECT 56.190 112.720 56.515 112.975 ;
        RECT 54.485 112.510 56.515 112.720 ;
        RECT 56.170 112.500 56.515 112.510 ;
        RECT 56.685 112.760 56.925 113.160 ;
        RECT 57.095 113.100 57.265 113.330 ;
        RECT 57.435 113.270 57.625 113.710 ;
        RECT 57.795 113.260 58.745 113.540 ;
        RECT 58.965 113.350 59.315 113.520 ;
        RECT 57.095 112.930 57.625 113.100 ;
        RECT 53.890 112.170 55.615 112.340 ;
        RECT 54.145 111.160 54.315 112.000 ;
        RECT 54.525 111.330 54.775 112.170 ;
        RECT 54.985 111.160 55.155 112.000 ;
        RECT 55.325 111.330 55.615 112.170 ;
        RECT 55.825 111.160 55.995 112.220 ;
        RECT 56.170 111.880 56.340 112.500 ;
        RECT 56.685 112.390 57.225 112.760 ;
        RECT 57.405 112.650 57.625 112.930 ;
        RECT 57.795 112.480 57.965 113.260 ;
        RECT 57.560 112.310 57.965 112.480 ;
        RECT 58.135 112.470 58.485 113.090 ;
        RECT 57.560 112.220 57.730 112.310 ;
        RECT 58.655 112.300 58.865 113.090 ;
        RECT 56.510 112.050 57.730 112.220 ;
        RECT 58.190 112.140 58.865 112.300 ;
        RECT 56.170 111.710 56.970 111.880 ;
        RECT 56.290 111.160 56.620 111.540 ;
        RECT 56.800 111.420 56.970 111.710 ;
        RECT 57.560 111.670 57.730 112.050 ;
        RECT 57.900 112.130 58.865 112.140 ;
        RECT 59.055 112.960 59.315 113.350 ;
        RECT 59.525 113.250 59.855 113.710 ;
        RECT 60.730 113.320 61.585 113.490 ;
        RECT 61.790 113.320 62.285 113.490 ;
        RECT 62.455 113.350 62.785 113.710 ;
        RECT 59.055 112.270 59.225 112.960 ;
        RECT 59.395 112.610 59.565 112.790 ;
        RECT 59.735 112.780 60.525 113.030 ;
        RECT 60.730 112.610 60.900 113.320 ;
        RECT 61.070 112.810 61.425 113.030 ;
        RECT 59.395 112.440 61.085 112.610 ;
        RECT 57.900 111.840 58.360 112.130 ;
        RECT 59.055 112.100 60.555 112.270 ;
        RECT 59.055 111.960 59.225 112.100 ;
        RECT 58.665 111.790 59.225 111.960 ;
        RECT 57.140 111.160 57.390 111.620 ;
        RECT 57.560 111.330 58.430 111.670 ;
        RECT 58.665 111.330 58.835 111.790 ;
        RECT 59.670 111.760 60.745 111.930 ;
        RECT 59.005 111.160 59.375 111.620 ;
        RECT 59.670 111.420 59.840 111.760 ;
        RECT 60.010 111.160 60.340 111.590 ;
        RECT 60.575 111.420 60.745 111.760 ;
        RECT 60.915 111.660 61.085 112.440 ;
        RECT 61.255 112.220 61.425 112.810 ;
        RECT 61.595 112.410 61.945 113.030 ;
        RECT 61.255 111.830 61.720 112.220 ;
        RECT 62.115 111.960 62.285 113.320 ;
        RECT 62.455 112.130 62.915 113.180 ;
        RECT 61.890 111.790 62.285 111.960 ;
        RECT 61.890 111.660 62.060 111.790 ;
        RECT 60.915 111.330 61.595 111.660 ;
        RECT 61.810 111.330 62.060 111.660 ;
        RECT 62.230 111.160 62.480 111.620 ;
        RECT 62.650 111.345 62.975 112.130 ;
        RECT 63.145 111.330 63.315 113.450 ;
        RECT 63.485 113.330 63.815 113.710 ;
        RECT 63.985 113.160 64.240 113.450 ;
        RECT 63.490 112.990 64.240 113.160 ;
        RECT 64.505 113.160 64.675 113.540 ;
        RECT 64.855 113.330 65.185 113.710 ;
        RECT 64.505 112.990 65.170 113.160 ;
        RECT 65.365 113.035 65.625 113.540 ;
        RECT 66.105 113.240 66.275 113.710 ;
        RECT 66.445 113.060 66.775 113.540 ;
        RECT 66.945 113.240 67.115 113.710 ;
        RECT 67.285 113.060 67.615 113.540 ;
        RECT 63.490 112.000 63.720 112.990 ;
        RECT 63.890 112.170 64.240 112.820 ;
        RECT 64.435 112.440 64.765 112.810 ;
        RECT 65.000 112.735 65.170 112.990 ;
        RECT 65.000 112.405 65.285 112.735 ;
        RECT 65.000 112.260 65.170 112.405 ;
        RECT 64.505 112.090 65.170 112.260 ;
        RECT 65.455 112.235 65.625 113.035 ;
        RECT 63.490 111.830 64.240 112.000 ;
        RECT 63.485 111.160 63.815 111.660 ;
        RECT 63.985 111.330 64.240 111.830 ;
        RECT 64.505 111.330 64.675 112.090 ;
        RECT 64.855 111.160 65.185 111.920 ;
        RECT 65.355 111.330 65.625 112.235 ;
        RECT 65.850 112.890 67.615 113.060 ;
        RECT 67.785 112.900 67.955 113.710 ;
        RECT 68.155 113.330 69.225 113.500 ;
        RECT 68.155 112.975 68.475 113.330 ;
        RECT 65.850 112.340 66.260 112.890 ;
        RECT 68.150 112.720 68.475 112.975 ;
        RECT 66.445 112.510 68.475 112.720 ;
        RECT 68.130 112.500 68.475 112.510 ;
        RECT 68.645 112.760 68.885 113.160 ;
        RECT 69.055 113.100 69.225 113.330 ;
        RECT 69.395 113.270 69.585 113.710 ;
        RECT 69.755 113.260 70.705 113.540 ;
        RECT 70.925 113.350 71.275 113.520 ;
        RECT 69.055 112.930 69.585 113.100 ;
        RECT 65.850 112.170 67.575 112.340 ;
        RECT 66.105 111.160 66.275 112.000 ;
        RECT 66.485 111.330 66.735 112.170 ;
        RECT 66.945 111.160 67.115 112.000 ;
        RECT 67.285 111.330 67.575 112.170 ;
        RECT 67.785 111.160 67.955 112.220 ;
        RECT 68.130 111.880 68.300 112.500 ;
        RECT 68.645 112.390 69.185 112.760 ;
        RECT 69.365 112.650 69.585 112.930 ;
        RECT 69.755 112.480 69.925 113.260 ;
        RECT 69.520 112.310 69.925 112.480 ;
        RECT 70.095 112.470 70.445 113.090 ;
        RECT 69.520 112.220 69.690 112.310 ;
        RECT 70.615 112.300 70.825 113.090 ;
        RECT 68.470 112.050 69.690 112.220 ;
        RECT 70.150 112.140 70.825 112.300 ;
        RECT 68.130 111.710 68.930 111.880 ;
        RECT 68.250 111.160 68.580 111.540 ;
        RECT 68.760 111.420 68.930 111.710 ;
        RECT 69.520 111.670 69.690 112.050 ;
        RECT 69.860 112.130 70.825 112.140 ;
        RECT 71.015 112.960 71.275 113.350 ;
        RECT 71.485 113.250 71.815 113.710 ;
        RECT 72.690 113.320 73.545 113.490 ;
        RECT 73.750 113.320 74.245 113.490 ;
        RECT 74.415 113.350 74.745 113.710 ;
        RECT 71.015 112.270 71.185 112.960 ;
        RECT 71.355 112.610 71.525 112.790 ;
        RECT 71.695 112.780 72.485 113.030 ;
        RECT 72.690 112.610 72.860 113.320 ;
        RECT 73.030 112.810 73.385 113.030 ;
        RECT 71.355 112.440 73.045 112.610 ;
        RECT 69.860 111.840 70.320 112.130 ;
        RECT 71.015 112.100 72.515 112.270 ;
        RECT 71.015 111.960 71.185 112.100 ;
        RECT 70.625 111.790 71.185 111.960 ;
        RECT 69.100 111.160 69.350 111.620 ;
        RECT 69.520 111.330 70.390 111.670 ;
        RECT 70.625 111.330 70.795 111.790 ;
        RECT 71.630 111.760 72.705 111.930 ;
        RECT 70.965 111.160 71.335 111.620 ;
        RECT 71.630 111.420 71.800 111.760 ;
        RECT 71.970 111.160 72.300 111.590 ;
        RECT 72.535 111.420 72.705 111.760 ;
        RECT 72.875 111.660 73.045 112.440 ;
        RECT 73.215 112.220 73.385 112.810 ;
        RECT 73.555 112.410 73.905 113.030 ;
        RECT 73.215 111.830 73.680 112.220 ;
        RECT 74.075 111.960 74.245 113.320 ;
        RECT 74.415 112.130 74.875 113.180 ;
        RECT 73.850 111.790 74.245 111.960 ;
        RECT 73.850 111.660 74.020 111.790 ;
        RECT 72.875 111.330 73.555 111.660 ;
        RECT 73.770 111.330 74.020 111.660 ;
        RECT 74.190 111.160 74.440 111.620 ;
        RECT 74.610 111.345 74.935 112.130 ;
        RECT 75.105 111.330 75.275 113.450 ;
        RECT 75.445 113.330 75.775 113.710 ;
        RECT 75.945 113.160 76.200 113.450 ;
        RECT 75.450 112.990 76.200 113.160 ;
        RECT 75.450 112.000 75.680 112.990 ;
        RECT 76.835 112.985 77.125 113.710 ;
        RECT 77.295 113.035 77.555 113.540 ;
        RECT 77.735 113.330 78.065 113.710 ;
        RECT 78.245 113.160 78.415 113.540 ;
        RECT 75.850 112.170 76.200 112.820 ;
        RECT 75.450 111.830 76.200 112.000 ;
        RECT 75.445 111.160 75.775 111.660 ;
        RECT 75.945 111.330 76.200 111.830 ;
        RECT 76.835 111.160 77.125 112.325 ;
        RECT 77.295 112.235 77.465 113.035 ;
        RECT 77.750 112.990 78.415 113.160 ;
        RECT 79.685 113.160 79.855 113.540 ;
        RECT 80.035 113.330 80.365 113.710 ;
        RECT 79.685 112.990 80.350 113.160 ;
        RECT 80.545 113.035 80.805 113.540 ;
        RECT 81.285 113.240 81.455 113.710 ;
        RECT 81.625 113.060 81.955 113.540 ;
        RECT 82.125 113.240 82.295 113.710 ;
        RECT 82.465 113.060 82.795 113.540 ;
        RECT 77.750 112.735 77.920 112.990 ;
        RECT 77.635 112.405 77.920 112.735 ;
        RECT 78.155 112.440 78.485 112.810 ;
        RECT 79.615 112.440 79.945 112.810 ;
        RECT 80.180 112.735 80.350 112.990 ;
        RECT 77.750 112.260 77.920 112.405 ;
        RECT 80.180 112.405 80.465 112.735 ;
        RECT 80.180 112.260 80.350 112.405 ;
        RECT 77.295 111.330 77.565 112.235 ;
        RECT 77.750 112.090 78.415 112.260 ;
        RECT 77.735 111.160 78.065 111.920 ;
        RECT 78.245 111.330 78.415 112.090 ;
        RECT 79.685 112.090 80.350 112.260 ;
        RECT 80.635 112.235 80.805 113.035 ;
        RECT 79.685 111.330 79.855 112.090 ;
        RECT 80.035 111.160 80.365 111.920 ;
        RECT 80.535 111.330 80.805 112.235 ;
        RECT 81.030 112.890 82.795 113.060 ;
        RECT 82.965 112.900 83.135 113.710 ;
        RECT 83.335 113.330 84.405 113.500 ;
        RECT 83.335 112.975 83.655 113.330 ;
        RECT 81.030 112.340 81.440 112.890 ;
        RECT 83.330 112.720 83.655 112.975 ;
        RECT 81.625 112.510 83.655 112.720 ;
        RECT 83.310 112.500 83.655 112.510 ;
        RECT 83.825 112.760 84.065 113.160 ;
        RECT 84.235 113.100 84.405 113.330 ;
        RECT 84.575 113.270 84.765 113.710 ;
        RECT 84.935 113.260 85.885 113.540 ;
        RECT 86.105 113.350 86.455 113.520 ;
        RECT 84.235 112.930 84.765 113.100 ;
        RECT 81.030 112.170 82.755 112.340 ;
        RECT 81.285 111.160 81.455 112.000 ;
        RECT 81.665 111.330 81.915 112.170 ;
        RECT 82.125 111.160 82.295 112.000 ;
        RECT 82.465 111.330 82.755 112.170 ;
        RECT 82.965 111.160 83.135 112.220 ;
        RECT 83.310 111.880 83.480 112.500 ;
        RECT 83.825 112.390 84.365 112.760 ;
        RECT 84.545 112.650 84.765 112.930 ;
        RECT 84.935 112.480 85.105 113.260 ;
        RECT 84.700 112.310 85.105 112.480 ;
        RECT 85.275 112.470 85.625 113.090 ;
        RECT 84.700 112.220 84.870 112.310 ;
        RECT 85.795 112.300 86.005 113.090 ;
        RECT 83.650 112.050 84.870 112.220 ;
        RECT 85.330 112.140 86.005 112.300 ;
        RECT 83.310 111.710 84.110 111.880 ;
        RECT 83.430 111.160 83.760 111.540 ;
        RECT 83.940 111.420 84.110 111.710 ;
        RECT 84.700 111.670 84.870 112.050 ;
        RECT 85.040 112.130 86.005 112.140 ;
        RECT 86.195 112.960 86.455 113.350 ;
        RECT 86.665 113.250 86.995 113.710 ;
        RECT 87.870 113.320 88.725 113.490 ;
        RECT 88.930 113.320 89.425 113.490 ;
        RECT 89.595 113.350 89.925 113.710 ;
        RECT 86.195 112.270 86.365 112.960 ;
        RECT 86.535 112.610 86.705 112.790 ;
        RECT 86.875 112.780 87.665 113.030 ;
        RECT 87.870 112.610 88.040 113.320 ;
        RECT 88.210 112.810 88.565 113.030 ;
        RECT 86.535 112.440 88.225 112.610 ;
        RECT 85.040 111.840 85.500 112.130 ;
        RECT 86.195 112.100 87.695 112.270 ;
        RECT 86.195 111.960 86.365 112.100 ;
        RECT 85.805 111.790 86.365 111.960 ;
        RECT 84.280 111.160 84.530 111.620 ;
        RECT 84.700 111.330 85.570 111.670 ;
        RECT 85.805 111.330 85.975 111.790 ;
        RECT 86.810 111.760 87.885 111.930 ;
        RECT 86.145 111.160 86.515 111.620 ;
        RECT 86.810 111.420 86.980 111.760 ;
        RECT 87.150 111.160 87.480 111.590 ;
        RECT 87.715 111.420 87.885 111.760 ;
        RECT 88.055 111.660 88.225 112.440 ;
        RECT 88.395 112.220 88.565 112.810 ;
        RECT 88.735 112.410 89.085 113.030 ;
        RECT 88.395 111.830 88.860 112.220 ;
        RECT 89.255 111.960 89.425 113.320 ;
        RECT 89.595 112.130 90.055 113.180 ;
        RECT 89.030 111.790 89.425 111.960 ;
        RECT 89.030 111.660 89.200 111.790 ;
        RECT 88.055 111.330 88.735 111.660 ;
        RECT 88.950 111.330 89.200 111.660 ;
        RECT 89.370 111.160 89.620 111.620 ;
        RECT 89.790 111.345 90.115 112.130 ;
        RECT 90.285 111.330 90.455 113.450 ;
        RECT 90.625 113.330 90.955 113.710 ;
        RECT 91.125 113.160 91.380 113.450 ;
        RECT 91.865 113.240 92.035 113.710 ;
        RECT 90.630 112.990 91.380 113.160 ;
        RECT 92.205 113.060 92.535 113.540 ;
        RECT 92.705 113.240 92.875 113.710 ;
        RECT 93.045 113.060 93.375 113.540 ;
        RECT 90.630 112.000 90.860 112.990 ;
        RECT 91.610 112.890 93.375 113.060 ;
        RECT 93.545 112.900 93.715 113.710 ;
        RECT 93.915 113.330 94.985 113.500 ;
        RECT 93.915 112.975 94.235 113.330 ;
        RECT 91.030 112.170 91.380 112.820 ;
        RECT 91.610 112.340 92.020 112.890 ;
        RECT 93.910 112.720 94.235 112.975 ;
        RECT 92.205 112.510 94.235 112.720 ;
        RECT 93.890 112.500 94.235 112.510 ;
        RECT 94.405 112.760 94.645 113.160 ;
        RECT 94.815 113.100 94.985 113.330 ;
        RECT 95.155 113.270 95.345 113.710 ;
        RECT 95.515 113.260 96.465 113.540 ;
        RECT 96.685 113.350 97.035 113.520 ;
        RECT 94.815 112.930 95.345 113.100 ;
        RECT 91.610 112.170 93.335 112.340 ;
        RECT 90.630 111.830 91.380 112.000 ;
        RECT 90.625 111.160 90.955 111.660 ;
        RECT 91.125 111.330 91.380 111.830 ;
        RECT 91.865 111.160 92.035 112.000 ;
        RECT 92.245 111.330 92.495 112.170 ;
        RECT 92.705 111.160 92.875 112.000 ;
        RECT 93.045 111.330 93.335 112.170 ;
        RECT 93.545 111.160 93.715 112.220 ;
        RECT 93.890 111.880 94.060 112.500 ;
        RECT 94.405 112.390 94.945 112.760 ;
        RECT 95.125 112.650 95.345 112.930 ;
        RECT 95.515 112.480 95.685 113.260 ;
        RECT 95.280 112.310 95.685 112.480 ;
        RECT 95.855 112.470 96.205 113.090 ;
        RECT 95.280 112.220 95.450 112.310 ;
        RECT 96.375 112.300 96.585 113.090 ;
        RECT 94.230 112.050 95.450 112.220 ;
        RECT 95.910 112.140 96.585 112.300 ;
        RECT 93.890 111.710 94.690 111.880 ;
        RECT 94.010 111.160 94.340 111.540 ;
        RECT 94.520 111.420 94.690 111.710 ;
        RECT 95.280 111.670 95.450 112.050 ;
        RECT 95.620 112.130 96.585 112.140 ;
        RECT 96.775 112.960 97.035 113.350 ;
        RECT 97.245 113.250 97.575 113.710 ;
        RECT 98.450 113.320 99.305 113.490 ;
        RECT 99.510 113.320 100.005 113.490 ;
        RECT 100.175 113.350 100.505 113.710 ;
        RECT 96.775 112.270 96.945 112.960 ;
        RECT 97.115 112.610 97.285 112.790 ;
        RECT 97.455 112.780 98.245 113.030 ;
        RECT 98.450 112.610 98.620 113.320 ;
        RECT 98.790 112.810 99.145 113.030 ;
        RECT 97.115 112.440 98.805 112.610 ;
        RECT 95.620 111.840 96.080 112.130 ;
        RECT 96.775 112.100 98.275 112.270 ;
        RECT 96.775 111.960 96.945 112.100 ;
        RECT 96.385 111.790 96.945 111.960 ;
        RECT 94.860 111.160 95.110 111.620 ;
        RECT 95.280 111.330 96.150 111.670 ;
        RECT 96.385 111.330 96.555 111.790 ;
        RECT 97.390 111.760 98.465 111.930 ;
        RECT 96.725 111.160 97.095 111.620 ;
        RECT 97.390 111.420 97.560 111.760 ;
        RECT 97.730 111.160 98.060 111.590 ;
        RECT 98.295 111.420 98.465 111.760 ;
        RECT 98.635 111.660 98.805 112.440 ;
        RECT 98.975 112.220 99.145 112.810 ;
        RECT 99.315 112.410 99.665 113.030 ;
        RECT 98.975 111.830 99.440 112.220 ;
        RECT 99.835 111.960 100.005 113.320 ;
        RECT 100.175 112.130 100.635 113.180 ;
        RECT 99.610 111.790 100.005 111.960 ;
        RECT 99.610 111.660 99.780 111.790 ;
        RECT 98.635 111.330 99.315 111.660 ;
        RECT 99.530 111.330 99.780 111.660 ;
        RECT 99.950 111.160 100.200 111.620 ;
        RECT 100.370 111.345 100.695 112.130 ;
        RECT 100.865 111.330 101.035 113.450 ;
        RECT 101.205 113.330 101.535 113.710 ;
        RECT 101.705 113.160 101.960 113.450 ;
        RECT 101.210 112.990 101.960 113.160 ;
        RECT 101.210 112.000 101.440 112.990 ;
        RECT 102.595 112.985 102.885 113.710 ;
        RECT 103.060 113.160 103.315 113.450 ;
        RECT 103.485 113.330 103.815 113.710 ;
        RECT 103.060 112.990 103.810 113.160 ;
        RECT 101.610 112.170 101.960 112.820 ;
        RECT 101.210 111.830 101.960 112.000 ;
        RECT 101.205 111.160 101.535 111.660 ;
        RECT 101.705 111.330 101.960 111.830 ;
        RECT 102.595 111.160 102.885 112.325 ;
        RECT 103.060 112.170 103.410 112.820 ;
        RECT 103.580 112.000 103.810 112.990 ;
        RECT 103.060 111.830 103.810 112.000 ;
        RECT 103.060 111.330 103.315 111.830 ;
        RECT 103.485 111.160 103.815 111.660 ;
        RECT 103.985 111.330 104.155 113.450 ;
        RECT 104.515 113.350 104.845 113.710 ;
        RECT 105.015 113.320 105.510 113.490 ;
        RECT 105.715 113.320 106.570 113.490 ;
        RECT 104.385 112.130 104.845 113.180 ;
        RECT 104.325 111.345 104.650 112.130 ;
        RECT 105.015 111.960 105.185 113.320 ;
        RECT 105.355 112.410 105.705 113.030 ;
        RECT 105.875 112.810 106.230 113.030 ;
        RECT 105.875 112.220 106.045 112.810 ;
        RECT 106.400 112.610 106.570 113.320 ;
        RECT 107.445 113.250 107.775 113.710 ;
        RECT 107.985 113.350 108.335 113.520 ;
        RECT 106.775 112.780 107.565 113.030 ;
        RECT 107.985 112.960 108.245 113.350 ;
        RECT 108.555 113.260 109.505 113.540 ;
        RECT 109.675 113.270 109.865 113.710 ;
        RECT 110.035 113.330 111.105 113.500 ;
        RECT 107.735 112.610 107.905 112.790 ;
        RECT 105.015 111.790 105.410 111.960 ;
        RECT 105.580 111.830 106.045 112.220 ;
        RECT 106.215 112.440 107.905 112.610 ;
        RECT 105.240 111.660 105.410 111.790 ;
        RECT 106.215 111.660 106.385 112.440 ;
        RECT 108.075 112.270 108.245 112.960 ;
        RECT 106.745 112.100 108.245 112.270 ;
        RECT 108.435 112.300 108.645 113.090 ;
        RECT 108.815 112.470 109.165 113.090 ;
        RECT 109.335 112.480 109.505 113.260 ;
        RECT 110.035 113.100 110.205 113.330 ;
        RECT 109.675 112.930 110.205 113.100 ;
        RECT 109.675 112.650 109.895 112.930 ;
        RECT 110.375 112.760 110.615 113.160 ;
        RECT 109.335 112.310 109.740 112.480 ;
        RECT 110.075 112.390 110.615 112.760 ;
        RECT 110.785 112.975 111.105 113.330 ;
        RECT 110.785 112.720 111.110 112.975 ;
        RECT 111.305 112.900 111.475 113.710 ;
        RECT 111.645 113.060 111.975 113.540 ;
        RECT 112.145 113.240 112.315 113.710 ;
        RECT 112.485 113.060 112.815 113.540 ;
        RECT 112.985 113.240 113.155 113.710 ;
        RECT 111.645 112.890 113.410 113.060 ;
        RECT 114.555 112.960 115.765 113.710 ;
        RECT 110.785 112.510 112.815 112.720 ;
        RECT 110.785 112.500 111.130 112.510 ;
        RECT 108.435 112.140 109.110 112.300 ;
        RECT 109.570 112.220 109.740 112.310 ;
        RECT 108.435 112.130 109.400 112.140 ;
        RECT 108.075 111.960 108.245 112.100 ;
        RECT 104.820 111.160 105.070 111.620 ;
        RECT 105.240 111.330 105.490 111.660 ;
        RECT 105.705 111.330 106.385 111.660 ;
        RECT 106.555 111.760 107.630 111.930 ;
        RECT 108.075 111.790 108.635 111.960 ;
        RECT 108.940 111.840 109.400 112.130 ;
        RECT 109.570 112.050 110.790 112.220 ;
        RECT 106.555 111.420 106.725 111.760 ;
        RECT 106.960 111.160 107.290 111.590 ;
        RECT 107.460 111.420 107.630 111.760 ;
        RECT 107.925 111.160 108.295 111.620 ;
        RECT 108.465 111.330 108.635 111.790 ;
        RECT 109.570 111.670 109.740 112.050 ;
        RECT 110.960 111.880 111.130 112.500 ;
        RECT 113.000 112.340 113.410 112.890 ;
        RECT 108.870 111.330 109.740 111.670 ;
        RECT 110.330 111.710 111.130 111.880 ;
        RECT 109.910 111.160 110.160 111.620 ;
        RECT 110.330 111.420 110.500 111.710 ;
        RECT 110.680 111.160 111.010 111.540 ;
        RECT 111.305 111.160 111.475 112.220 ;
        RECT 111.685 112.170 113.410 112.340 ;
        RECT 114.555 112.250 115.075 112.790 ;
        RECT 115.245 112.420 115.765 112.960 ;
        RECT 111.685 111.330 111.975 112.170 ;
        RECT 112.145 111.160 112.315 112.000 ;
        RECT 112.525 111.330 112.775 112.170 ;
        RECT 112.985 111.160 113.155 112.000 ;
        RECT 114.555 111.160 115.765 112.250 ;
        RECT 14.650 110.990 115.850 111.160 ;
        RECT 14.735 109.900 15.945 110.990 ;
        RECT 17.345 110.150 17.515 110.990 ;
        RECT 17.725 109.980 17.975 110.820 ;
        RECT 18.185 110.150 18.355 110.990 ;
        RECT 18.525 109.980 18.815 110.820 ;
        RECT 14.735 109.190 15.255 109.730 ;
        RECT 15.425 109.360 15.945 109.900 ;
        RECT 17.090 109.810 18.815 109.980 ;
        RECT 19.025 109.930 19.195 110.990 ;
        RECT 19.490 110.610 19.820 110.990 ;
        RECT 20.000 110.440 20.170 110.730 ;
        RECT 20.340 110.530 20.590 110.990 ;
        RECT 19.370 110.270 20.170 110.440 ;
        RECT 20.760 110.480 21.630 110.820 ;
        RECT 17.090 109.260 17.500 109.810 ;
        RECT 19.370 109.650 19.540 110.270 ;
        RECT 20.760 110.100 20.930 110.480 ;
        RECT 21.865 110.360 22.035 110.820 ;
        RECT 22.205 110.530 22.575 110.990 ;
        RECT 22.870 110.390 23.040 110.730 ;
        RECT 23.210 110.560 23.540 110.990 ;
        RECT 23.775 110.390 23.945 110.730 ;
        RECT 19.710 109.930 20.930 110.100 ;
        RECT 21.100 110.020 21.560 110.310 ;
        RECT 21.865 110.190 22.425 110.360 ;
        RECT 22.870 110.220 23.945 110.390 ;
        RECT 24.115 110.490 24.795 110.820 ;
        RECT 25.010 110.490 25.260 110.820 ;
        RECT 25.430 110.530 25.680 110.990 ;
        RECT 22.255 110.050 22.425 110.190 ;
        RECT 21.100 110.010 22.065 110.020 ;
        RECT 20.760 109.840 20.930 109.930 ;
        RECT 21.390 109.850 22.065 110.010 ;
        RECT 19.370 109.640 19.715 109.650 ;
        RECT 17.685 109.430 19.715 109.640 ;
        RECT 14.735 108.440 15.945 109.190 ;
        RECT 17.090 109.090 18.855 109.260 ;
        RECT 17.345 108.440 17.515 108.910 ;
        RECT 17.685 108.610 18.015 109.090 ;
        RECT 18.185 108.440 18.355 108.910 ;
        RECT 18.525 108.610 18.855 109.090 ;
        RECT 19.025 108.440 19.195 109.250 ;
        RECT 19.390 109.175 19.715 109.430 ;
        RECT 19.395 108.820 19.715 109.175 ;
        RECT 19.885 109.390 20.425 109.760 ;
        RECT 20.760 109.670 21.165 109.840 ;
        RECT 19.885 108.990 20.125 109.390 ;
        RECT 20.605 109.220 20.825 109.500 ;
        RECT 20.295 109.050 20.825 109.220 ;
        RECT 20.295 108.820 20.465 109.050 ;
        RECT 20.995 108.890 21.165 109.670 ;
        RECT 21.335 109.060 21.685 109.680 ;
        RECT 21.855 109.060 22.065 109.850 ;
        RECT 22.255 109.880 23.755 110.050 ;
        RECT 22.255 109.190 22.425 109.880 ;
        RECT 24.115 109.710 24.285 110.490 ;
        RECT 25.090 110.360 25.260 110.490 ;
        RECT 22.595 109.540 24.285 109.710 ;
        RECT 24.455 109.930 24.920 110.320 ;
        RECT 25.090 110.190 25.485 110.360 ;
        RECT 22.595 109.360 22.765 109.540 ;
        RECT 19.395 108.650 20.465 108.820 ;
        RECT 20.635 108.440 20.825 108.880 ;
        RECT 20.995 108.610 21.945 108.890 ;
        RECT 22.255 108.800 22.515 109.190 ;
        RECT 22.935 109.120 23.725 109.370 ;
        RECT 22.165 108.630 22.515 108.800 ;
        RECT 22.725 108.440 23.055 108.900 ;
        RECT 23.930 108.830 24.100 109.540 ;
        RECT 24.455 109.340 24.625 109.930 ;
        RECT 24.270 109.120 24.625 109.340 ;
        RECT 24.795 109.120 25.145 109.740 ;
        RECT 25.315 108.830 25.485 110.190 ;
        RECT 25.850 110.020 26.175 110.805 ;
        RECT 25.655 108.970 26.115 110.020 ;
        RECT 23.930 108.660 24.785 108.830 ;
        RECT 24.990 108.660 25.485 108.830 ;
        RECT 25.655 108.440 25.985 108.800 ;
        RECT 26.345 108.700 26.515 110.820 ;
        RECT 26.685 110.490 27.015 110.990 ;
        RECT 27.185 110.320 27.440 110.820 ;
        RECT 26.690 110.150 27.440 110.320 ;
        RECT 27.925 110.150 28.095 110.990 ;
        RECT 26.690 109.160 26.920 110.150 ;
        RECT 28.305 109.980 28.555 110.820 ;
        RECT 28.765 110.150 28.935 110.990 ;
        RECT 29.105 109.980 29.395 110.820 ;
        RECT 27.090 109.330 27.440 109.980 ;
        RECT 27.670 109.810 29.395 109.980 ;
        RECT 29.605 109.930 29.775 110.990 ;
        RECT 30.070 110.610 30.400 110.990 ;
        RECT 30.580 110.440 30.750 110.730 ;
        RECT 30.920 110.530 31.170 110.990 ;
        RECT 29.950 110.270 30.750 110.440 ;
        RECT 31.340 110.480 32.210 110.820 ;
        RECT 27.670 109.260 28.080 109.810 ;
        RECT 29.950 109.650 30.120 110.270 ;
        RECT 31.340 110.100 31.510 110.480 ;
        RECT 32.445 110.360 32.615 110.820 ;
        RECT 32.785 110.530 33.155 110.990 ;
        RECT 33.450 110.390 33.620 110.730 ;
        RECT 33.790 110.560 34.120 110.990 ;
        RECT 34.355 110.390 34.525 110.730 ;
        RECT 30.290 109.930 31.510 110.100 ;
        RECT 31.680 110.020 32.140 110.310 ;
        RECT 32.445 110.190 33.005 110.360 ;
        RECT 33.450 110.220 34.525 110.390 ;
        RECT 34.695 110.490 35.375 110.820 ;
        RECT 35.590 110.490 35.840 110.820 ;
        RECT 36.010 110.530 36.260 110.990 ;
        RECT 32.835 110.050 33.005 110.190 ;
        RECT 31.680 110.010 32.645 110.020 ;
        RECT 31.340 109.840 31.510 109.930 ;
        RECT 31.970 109.850 32.645 110.010 ;
        RECT 29.950 109.640 30.295 109.650 ;
        RECT 28.265 109.430 30.295 109.640 ;
        RECT 26.690 108.990 27.440 109.160 ;
        RECT 27.670 109.090 29.435 109.260 ;
        RECT 26.685 108.440 27.015 108.820 ;
        RECT 27.185 108.700 27.440 108.990 ;
        RECT 27.925 108.440 28.095 108.910 ;
        RECT 28.265 108.610 28.595 109.090 ;
        RECT 28.765 108.440 28.935 108.910 ;
        RECT 29.105 108.610 29.435 109.090 ;
        RECT 29.605 108.440 29.775 109.250 ;
        RECT 29.970 109.175 30.295 109.430 ;
        RECT 29.975 108.820 30.295 109.175 ;
        RECT 30.465 109.390 31.005 109.760 ;
        RECT 31.340 109.670 31.745 109.840 ;
        RECT 30.465 108.990 30.705 109.390 ;
        RECT 31.185 109.220 31.405 109.500 ;
        RECT 30.875 109.050 31.405 109.220 ;
        RECT 30.875 108.820 31.045 109.050 ;
        RECT 31.575 108.890 31.745 109.670 ;
        RECT 31.915 109.060 32.265 109.680 ;
        RECT 32.435 109.060 32.645 109.850 ;
        RECT 32.835 109.880 34.335 110.050 ;
        RECT 32.835 109.190 33.005 109.880 ;
        RECT 34.695 109.710 34.865 110.490 ;
        RECT 35.670 110.360 35.840 110.490 ;
        RECT 33.175 109.540 34.865 109.710 ;
        RECT 35.035 109.930 35.500 110.320 ;
        RECT 35.670 110.190 36.065 110.360 ;
        RECT 33.175 109.360 33.345 109.540 ;
        RECT 29.975 108.650 31.045 108.820 ;
        RECT 31.215 108.440 31.405 108.880 ;
        RECT 31.575 108.610 32.525 108.890 ;
        RECT 32.835 108.800 33.095 109.190 ;
        RECT 33.515 109.120 34.305 109.370 ;
        RECT 32.745 108.630 33.095 108.800 ;
        RECT 33.305 108.440 33.635 108.900 ;
        RECT 34.510 108.830 34.680 109.540 ;
        RECT 35.035 109.340 35.205 109.930 ;
        RECT 34.850 109.120 35.205 109.340 ;
        RECT 35.375 109.120 35.725 109.740 ;
        RECT 35.895 108.830 36.065 110.190 ;
        RECT 36.430 110.020 36.755 110.805 ;
        RECT 36.235 108.970 36.695 110.020 ;
        RECT 34.510 108.660 35.365 108.830 ;
        RECT 35.570 108.660 36.065 108.830 ;
        RECT 36.235 108.440 36.565 108.800 ;
        RECT 36.925 108.700 37.095 110.820 ;
        RECT 37.265 110.490 37.595 110.990 ;
        RECT 37.765 110.320 38.020 110.820 ;
        RECT 37.270 110.150 38.020 110.320 ;
        RECT 37.270 109.160 37.500 110.150 ;
        RECT 37.670 109.330 38.020 109.980 ;
        RECT 38.195 109.825 38.485 110.990 ;
        RECT 38.715 109.850 38.925 110.990 ;
        RECT 39.095 109.840 39.425 110.820 ;
        RECT 39.595 109.850 39.825 110.990 ;
        RECT 40.995 109.850 41.225 110.990 ;
        RECT 41.395 109.840 41.725 110.820 ;
        RECT 41.895 109.850 42.105 110.990 ;
        RECT 43.255 109.900 46.765 110.990 ;
        RECT 37.270 108.990 38.020 109.160 ;
        RECT 37.265 108.440 37.595 108.820 ;
        RECT 37.765 108.700 38.020 108.990 ;
        RECT 38.195 108.440 38.485 109.165 ;
        RECT 38.715 108.440 38.925 109.260 ;
        RECT 39.095 109.240 39.345 109.840 ;
        RECT 39.515 109.430 39.845 109.680 ;
        RECT 40.975 109.430 41.305 109.680 ;
        RECT 39.095 108.610 39.425 109.240 ;
        RECT 39.595 108.440 39.825 109.260 ;
        RECT 40.995 108.440 41.225 109.260 ;
        RECT 41.475 109.240 41.725 109.840 ;
        RECT 43.255 109.380 44.945 109.900 ;
        RECT 46.995 109.850 47.205 110.990 ;
        RECT 47.375 109.840 47.705 110.820 ;
        RECT 47.875 109.850 48.105 110.990 ;
        RECT 48.625 110.150 48.795 110.990 ;
        RECT 49.005 109.980 49.255 110.820 ;
        RECT 49.465 110.150 49.635 110.990 ;
        RECT 49.805 109.980 50.095 110.820 ;
        RECT 41.395 108.610 41.725 109.240 ;
        RECT 41.895 108.440 42.105 109.260 ;
        RECT 45.115 109.210 46.765 109.730 ;
        RECT 43.255 108.440 46.765 109.210 ;
        RECT 46.995 108.440 47.205 109.260 ;
        RECT 47.375 109.240 47.625 109.840 ;
        RECT 48.370 109.810 50.095 109.980 ;
        RECT 50.305 109.930 50.475 110.990 ;
        RECT 50.770 110.610 51.100 110.990 ;
        RECT 51.280 110.440 51.450 110.730 ;
        RECT 51.620 110.530 51.870 110.990 ;
        RECT 50.650 110.270 51.450 110.440 ;
        RECT 52.040 110.480 52.910 110.820 ;
        RECT 47.795 109.430 48.125 109.680 ;
        RECT 48.370 109.260 48.780 109.810 ;
        RECT 50.650 109.650 50.820 110.270 ;
        RECT 52.040 110.100 52.210 110.480 ;
        RECT 53.145 110.360 53.315 110.820 ;
        RECT 53.485 110.530 53.855 110.990 ;
        RECT 54.150 110.390 54.320 110.730 ;
        RECT 54.490 110.560 54.820 110.990 ;
        RECT 55.055 110.390 55.225 110.730 ;
        RECT 50.990 109.930 52.210 110.100 ;
        RECT 52.380 110.020 52.840 110.310 ;
        RECT 53.145 110.190 53.705 110.360 ;
        RECT 54.150 110.220 55.225 110.390 ;
        RECT 55.395 110.490 56.075 110.820 ;
        RECT 56.290 110.490 56.540 110.820 ;
        RECT 56.710 110.530 56.960 110.990 ;
        RECT 53.535 110.050 53.705 110.190 ;
        RECT 52.380 110.010 53.345 110.020 ;
        RECT 52.040 109.840 52.210 109.930 ;
        RECT 52.670 109.850 53.345 110.010 ;
        RECT 50.650 109.640 50.995 109.650 ;
        RECT 48.965 109.430 50.995 109.640 ;
        RECT 47.375 108.610 47.705 109.240 ;
        RECT 47.875 108.440 48.105 109.260 ;
        RECT 48.370 109.090 50.135 109.260 ;
        RECT 48.625 108.440 48.795 108.910 ;
        RECT 48.965 108.610 49.295 109.090 ;
        RECT 49.465 108.440 49.635 108.910 ;
        RECT 49.805 108.610 50.135 109.090 ;
        RECT 50.305 108.440 50.475 109.250 ;
        RECT 50.670 109.175 50.995 109.430 ;
        RECT 50.675 108.820 50.995 109.175 ;
        RECT 51.165 109.390 51.705 109.760 ;
        RECT 52.040 109.670 52.445 109.840 ;
        RECT 51.165 108.990 51.405 109.390 ;
        RECT 51.885 109.220 52.105 109.500 ;
        RECT 51.575 109.050 52.105 109.220 ;
        RECT 51.575 108.820 51.745 109.050 ;
        RECT 52.275 108.890 52.445 109.670 ;
        RECT 52.615 109.060 52.965 109.680 ;
        RECT 53.135 109.060 53.345 109.850 ;
        RECT 53.535 109.880 55.035 110.050 ;
        RECT 53.535 109.190 53.705 109.880 ;
        RECT 55.395 109.710 55.565 110.490 ;
        RECT 56.370 110.360 56.540 110.490 ;
        RECT 53.875 109.540 55.565 109.710 ;
        RECT 55.735 109.930 56.200 110.320 ;
        RECT 56.370 110.190 56.765 110.360 ;
        RECT 53.875 109.360 54.045 109.540 ;
        RECT 50.675 108.650 51.745 108.820 ;
        RECT 51.915 108.440 52.105 108.880 ;
        RECT 52.275 108.610 53.225 108.890 ;
        RECT 53.535 108.800 53.795 109.190 ;
        RECT 54.215 109.120 55.005 109.370 ;
        RECT 53.445 108.630 53.795 108.800 ;
        RECT 54.005 108.440 54.335 108.900 ;
        RECT 55.210 108.830 55.380 109.540 ;
        RECT 55.735 109.340 55.905 109.930 ;
        RECT 55.550 109.120 55.905 109.340 ;
        RECT 56.075 109.120 56.425 109.740 ;
        RECT 56.595 108.830 56.765 110.190 ;
        RECT 57.130 110.020 57.455 110.805 ;
        RECT 56.935 108.970 57.395 110.020 ;
        RECT 55.210 108.660 56.065 108.830 ;
        RECT 56.270 108.660 56.765 108.830 ;
        RECT 56.935 108.440 57.265 108.800 ;
        RECT 57.625 108.700 57.795 110.820 ;
        RECT 57.965 110.490 58.295 110.990 ;
        RECT 58.465 110.320 58.720 110.820 ;
        RECT 57.970 110.150 58.720 110.320 ;
        RECT 57.970 109.160 58.200 110.150 ;
        RECT 59.905 110.060 60.075 110.820 ;
        RECT 60.255 110.230 60.585 110.990 ;
        RECT 58.370 109.330 58.720 109.980 ;
        RECT 59.905 109.890 60.570 110.060 ;
        RECT 60.755 109.915 61.025 110.820 ;
        RECT 60.400 109.745 60.570 109.890 ;
        RECT 59.835 109.340 60.165 109.710 ;
        RECT 60.400 109.415 60.685 109.745 ;
        RECT 60.400 109.160 60.570 109.415 ;
        RECT 57.970 108.990 58.720 109.160 ;
        RECT 57.965 108.440 58.295 108.820 ;
        RECT 58.465 108.700 58.720 108.990 ;
        RECT 59.905 108.990 60.570 109.160 ;
        RECT 60.855 109.115 61.025 109.915 ;
        RECT 61.235 109.850 61.465 110.990 ;
        RECT 61.635 109.840 61.965 110.820 ;
        RECT 62.135 109.850 62.345 110.990 ;
        RECT 62.575 109.900 63.785 110.990 ;
        RECT 61.215 109.430 61.545 109.680 ;
        RECT 59.905 108.610 60.075 108.990 ;
        RECT 60.255 108.440 60.585 108.820 ;
        RECT 60.765 108.610 61.025 109.115 ;
        RECT 61.235 108.440 61.465 109.260 ;
        RECT 61.715 109.240 61.965 109.840 ;
        RECT 62.575 109.360 63.095 109.900 ;
        RECT 63.955 109.825 64.245 110.990 ;
        RECT 64.725 110.150 64.895 110.990 ;
        RECT 65.105 109.980 65.355 110.820 ;
        RECT 65.565 110.150 65.735 110.990 ;
        RECT 65.905 109.980 66.195 110.820 ;
        RECT 64.470 109.810 66.195 109.980 ;
        RECT 66.405 109.930 66.575 110.990 ;
        RECT 66.870 110.610 67.200 110.990 ;
        RECT 67.380 110.440 67.550 110.730 ;
        RECT 67.720 110.530 67.970 110.990 ;
        RECT 66.750 110.270 67.550 110.440 ;
        RECT 68.140 110.480 69.010 110.820 ;
        RECT 61.635 108.610 61.965 109.240 ;
        RECT 62.135 108.440 62.345 109.260 ;
        RECT 63.265 109.190 63.785 109.730 ;
        RECT 62.575 108.440 63.785 109.190 ;
        RECT 64.470 109.260 64.880 109.810 ;
        RECT 66.750 109.650 66.920 110.270 ;
        RECT 68.140 110.100 68.310 110.480 ;
        RECT 69.245 110.360 69.415 110.820 ;
        RECT 69.585 110.530 69.955 110.990 ;
        RECT 70.250 110.390 70.420 110.730 ;
        RECT 70.590 110.560 70.920 110.990 ;
        RECT 71.155 110.390 71.325 110.730 ;
        RECT 67.090 109.930 68.310 110.100 ;
        RECT 68.480 110.020 68.940 110.310 ;
        RECT 69.245 110.190 69.805 110.360 ;
        RECT 70.250 110.220 71.325 110.390 ;
        RECT 71.495 110.490 72.175 110.820 ;
        RECT 72.390 110.490 72.640 110.820 ;
        RECT 72.810 110.530 73.060 110.990 ;
        RECT 69.635 110.050 69.805 110.190 ;
        RECT 68.480 110.010 69.445 110.020 ;
        RECT 68.140 109.840 68.310 109.930 ;
        RECT 68.770 109.850 69.445 110.010 ;
        RECT 66.750 109.640 67.095 109.650 ;
        RECT 65.065 109.430 67.095 109.640 ;
        RECT 63.955 108.440 64.245 109.165 ;
        RECT 64.470 109.090 66.235 109.260 ;
        RECT 64.725 108.440 64.895 108.910 ;
        RECT 65.065 108.610 65.395 109.090 ;
        RECT 65.565 108.440 65.735 108.910 ;
        RECT 65.905 108.610 66.235 109.090 ;
        RECT 66.405 108.440 66.575 109.250 ;
        RECT 66.770 109.175 67.095 109.430 ;
        RECT 66.775 108.820 67.095 109.175 ;
        RECT 67.265 109.390 67.805 109.760 ;
        RECT 68.140 109.670 68.545 109.840 ;
        RECT 67.265 108.990 67.505 109.390 ;
        RECT 67.985 109.220 68.205 109.500 ;
        RECT 67.675 109.050 68.205 109.220 ;
        RECT 67.675 108.820 67.845 109.050 ;
        RECT 68.375 108.890 68.545 109.670 ;
        RECT 68.715 109.060 69.065 109.680 ;
        RECT 69.235 109.060 69.445 109.850 ;
        RECT 69.635 109.880 71.135 110.050 ;
        RECT 69.635 109.190 69.805 109.880 ;
        RECT 71.495 109.710 71.665 110.490 ;
        RECT 72.470 110.360 72.640 110.490 ;
        RECT 69.975 109.540 71.665 109.710 ;
        RECT 71.835 109.930 72.300 110.320 ;
        RECT 72.470 110.190 72.865 110.360 ;
        RECT 69.975 109.360 70.145 109.540 ;
        RECT 66.775 108.650 67.845 108.820 ;
        RECT 68.015 108.440 68.205 108.880 ;
        RECT 68.375 108.610 69.325 108.890 ;
        RECT 69.635 108.800 69.895 109.190 ;
        RECT 70.315 109.120 71.105 109.370 ;
        RECT 69.545 108.630 69.895 108.800 ;
        RECT 70.105 108.440 70.435 108.900 ;
        RECT 71.310 108.830 71.480 109.540 ;
        RECT 71.835 109.340 72.005 109.930 ;
        RECT 71.650 109.120 72.005 109.340 ;
        RECT 72.175 109.120 72.525 109.740 ;
        RECT 72.695 108.830 72.865 110.190 ;
        RECT 73.230 110.020 73.555 110.805 ;
        RECT 73.035 108.970 73.495 110.020 ;
        RECT 71.310 108.660 72.165 108.830 ;
        RECT 72.370 108.660 72.865 108.830 ;
        RECT 73.035 108.440 73.365 108.800 ;
        RECT 73.725 108.700 73.895 110.820 ;
        RECT 74.065 110.490 74.395 110.990 ;
        RECT 74.565 110.320 74.820 110.820 ;
        RECT 74.070 110.150 74.820 110.320 ;
        RECT 76.225 110.150 76.395 110.990 ;
        RECT 74.070 109.160 74.300 110.150 ;
        RECT 76.605 109.980 76.855 110.820 ;
        RECT 77.065 110.150 77.235 110.990 ;
        RECT 77.405 109.980 77.695 110.820 ;
        RECT 74.470 109.330 74.820 109.980 ;
        RECT 75.970 109.810 77.695 109.980 ;
        RECT 77.905 109.930 78.075 110.990 ;
        RECT 78.370 110.610 78.700 110.990 ;
        RECT 78.880 110.440 79.050 110.730 ;
        RECT 79.220 110.530 79.470 110.990 ;
        RECT 78.250 110.270 79.050 110.440 ;
        RECT 79.640 110.480 80.510 110.820 ;
        RECT 75.970 109.260 76.380 109.810 ;
        RECT 78.250 109.650 78.420 110.270 ;
        RECT 79.640 110.100 79.810 110.480 ;
        RECT 80.745 110.360 80.915 110.820 ;
        RECT 81.085 110.530 81.455 110.990 ;
        RECT 81.750 110.390 81.920 110.730 ;
        RECT 82.090 110.560 82.420 110.990 ;
        RECT 82.655 110.390 82.825 110.730 ;
        RECT 78.590 109.930 79.810 110.100 ;
        RECT 79.980 110.020 80.440 110.310 ;
        RECT 80.745 110.190 81.305 110.360 ;
        RECT 81.750 110.220 82.825 110.390 ;
        RECT 82.995 110.490 83.675 110.820 ;
        RECT 83.890 110.490 84.140 110.820 ;
        RECT 84.310 110.530 84.560 110.990 ;
        RECT 81.135 110.050 81.305 110.190 ;
        RECT 79.980 110.010 80.945 110.020 ;
        RECT 79.640 109.840 79.810 109.930 ;
        RECT 80.270 109.850 80.945 110.010 ;
        RECT 78.250 109.640 78.595 109.650 ;
        RECT 76.565 109.430 78.595 109.640 ;
        RECT 74.070 108.990 74.820 109.160 ;
        RECT 75.970 109.090 77.735 109.260 ;
        RECT 74.065 108.440 74.395 108.820 ;
        RECT 74.565 108.700 74.820 108.990 ;
        RECT 76.225 108.440 76.395 108.910 ;
        RECT 76.565 108.610 76.895 109.090 ;
        RECT 77.065 108.440 77.235 108.910 ;
        RECT 77.405 108.610 77.735 109.090 ;
        RECT 77.905 108.440 78.075 109.250 ;
        RECT 78.270 109.175 78.595 109.430 ;
        RECT 78.275 108.820 78.595 109.175 ;
        RECT 78.765 109.390 79.305 109.760 ;
        RECT 79.640 109.670 80.045 109.840 ;
        RECT 78.765 108.990 79.005 109.390 ;
        RECT 79.485 109.220 79.705 109.500 ;
        RECT 79.175 109.050 79.705 109.220 ;
        RECT 79.175 108.820 79.345 109.050 ;
        RECT 79.875 108.890 80.045 109.670 ;
        RECT 80.215 109.060 80.565 109.680 ;
        RECT 80.735 109.060 80.945 109.850 ;
        RECT 81.135 109.880 82.635 110.050 ;
        RECT 81.135 109.190 81.305 109.880 ;
        RECT 82.995 109.710 83.165 110.490 ;
        RECT 83.970 110.360 84.140 110.490 ;
        RECT 81.475 109.540 83.165 109.710 ;
        RECT 83.335 109.930 83.800 110.320 ;
        RECT 83.970 110.190 84.365 110.360 ;
        RECT 81.475 109.360 81.645 109.540 ;
        RECT 78.275 108.650 79.345 108.820 ;
        RECT 79.515 108.440 79.705 108.880 ;
        RECT 79.875 108.610 80.825 108.890 ;
        RECT 81.135 108.800 81.395 109.190 ;
        RECT 81.815 109.120 82.605 109.370 ;
        RECT 81.045 108.630 81.395 108.800 ;
        RECT 81.605 108.440 81.935 108.900 ;
        RECT 82.810 108.830 82.980 109.540 ;
        RECT 83.335 109.340 83.505 109.930 ;
        RECT 83.150 109.120 83.505 109.340 ;
        RECT 83.675 109.120 84.025 109.740 ;
        RECT 84.195 108.830 84.365 110.190 ;
        RECT 84.730 110.020 85.055 110.805 ;
        RECT 84.535 108.970 84.995 110.020 ;
        RECT 82.810 108.660 83.665 108.830 ;
        RECT 83.870 108.660 84.365 108.830 ;
        RECT 84.535 108.440 84.865 108.800 ;
        RECT 85.225 108.700 85.395 110.820 ;
        RECT 85.565 110.490 85.895 110.990 ;
        RECT 86.065 110.320 86.320 110.820 ;
        RECT 85.570 110.150 86.320 110.320 ;
        RECT 85.570 109.160 85.800 110.150 ;
        RECT 85.970 109.330 86.320 109.980 ;
        RECT 86.555 109.850 86.765 110.990 ;
        RECT 86.935 109.840 87.265 110.820 ;
        RECT 87.435 109.850 87.665 110.990 ;
        RECT 88.375 109.850 88.605 110.990 ;
        RECT 88.775 109.840 89.105 110.820 ;
        RECT 89.275 109.850 89.485 110.990 ;
        RECT 85.570 108.990 86.320 109.160 ;
        RECT 85.565 108.440 85.895 108.820 ;
        RECT 86.065 108.700 86.320 108.990 ;
        RECT 86.555 108.440 86.765 109.260 ;
        RECT 86.935 109.240 87.185 109.840 ;
        RECT 87.355 109.430 87.685 109.680 ;
        RECT 88.355 109.430 88.685 109.680 ;
        RECT 86.935 108.610 87.265 109.240 ;
        RECT 87.435 108.440 87.665 109.260 ;
        RECT 88.375 108.440 88.605 109.260 ;
        RECT 88.855 109.240 89.105 109.840 ;
        RECT 89.715 109.825 90.005 110.990 ;
        RECT 90.485 110.150 90.655 110.990 ;
        RECT 90.865 109.980 91.115 110.820 ;
        RECT 91.325 110.150 91.495 110.990 ;
        RECT 91.665 109.980 91.955 110.820 ;
        RECT 90.230 109.810 91.955 109.980 ;
        RECT 92.165 109.930 92.335 110.990 ;
        RECT 92.630 110.610 92.960 110.990 ;
        RECT 93.140 110.440 93.310 110.730 ;
        RECT 93.480 110.530 93.730 110.990 ;
        RECT 92.510 110.270 93.310 110.440 ;
        RECT 93.900 110.480 94.770 110.820 ;
        RECT 90.230 109.260 90.640 109.810 ;
        RECT 92.510 109.650 92.680 110.270 ;
        RECT 93.900 110.100 94.070 110.480 ;
        RECT 95.005 110.360 95.175 110.820 ;
        RECT 95.345 110.530 95.715 110.990 ;
        RECT 96.010 110.390 96.180 110.730 ;
        RECT 96.350 110.560 96.680 110.990 ;
        RECT 96.915 110.390 97.085 110.730 ;
        RECT 92.850 109.930 94.070 110.100 ;
        RECT 94.240 110.020 94.700 110.310 ;
        RECT 95.005 110.190 95.565 110.360 ;
        RECT 96.010 110.220 97.085 110.390 ;
        RECT 97.255 110.490 97.935 110.820 ;
        RECT 98.150 110.490 98.400 110.820 ;
        RECT 98.570 110.530 98.820 110.990 ;
        RECT 95.395 110.050 95.565 110.190 ;
        RECT 94.240 110.010 95.205 110.020 ;
        RECT 93.900 109.840 94.070 109.930 ;
        RECT 94.530 109.850 95.205 110.010 ;
        RECT 92.510 109.640 92.855 109.650 ;
        RECT 90.825 109.430 92.855 109.640 ;
        RECT 88.775 108.610 89.105 109.240 ;
        RECT 89.275 108.440 89.485 109.260 ;
        RECT 89.715 108.440 90.005 109.165 ;
        RECT 90.230 109.090 91.995 109.260 ;
        RECT 90.485 108.440 90.655 108.910 ;
        RECT 90.825 108.610 91.155 109.090 ;
        RECT 91.325 108.440 91.495 108.910 ;
        RECT 91.665 108.610 91.995 109.090 ;
        RECT 92.165 108.440 92.335 109.250 ;
        RECT 92.530 109.175 92.855 109.430 ;
        RECT 92.535 108.820 92.855 109.175 ;
        RECT 93.025 109.390 93.565 109.760 ;
        RECT 93.900 109.670 94.305 109.840 ;
        RECT 93.025 108.990 93.265 109.390 ;
        RECT 93.745 109.220 93.965 109.500 ;
        RECT 93.435 109.050 93.965 109.220 ;
        RECT 93.435 108.820 93.605 109.050 ;
        RECT 94.135 108.890 94.305 109.670 ;
        RECT 94.475 109.060 94.825 109.680 ;
        RECT 94.995 109.060 95.205 109.850 ;
        RECT 95.395 109.880 96.895 110.050 ;
        RECT 95.395 109.190 95.565 109.880 ;
        RECT 97.255 109.710 97.425 110.490 ;
        RECT 98.230 110.360 98.400 110.490 ;
        RECT 95.735 109.540 97.425 109.710 ;
        RECT 97.595 109.930 98.060 110.320 ;
        RECT 98.230 110.190 98.625 110.360 ;
        RECT 95.735 109.360 95.905 109.540 ;
        RECT 92.535 108.650 93.605 108.820 ;
        RECT 93.775 108.440 93.965 108.880 ;
        RECT 94.135 108.610 95.085 108.890 ;
        RECT 95.395 108.800 95.655 109.190 ;
        RECT 96.075 109.120 96.865 109.370 ;
        RECT 95.305 108.630 95.655 108.800 ;
        RECT 95.865 108.440 96.195 108.900 ;
        RECT 97.070 108.830 97.240 109.540 ;
        RECT 97.595 109.340 97.765 109.930 ;
        RECT 97.410 109.120 97.765 109.340 ;
        RECT 97.935 109.120 98.285 109.740 ;
        RECT 98.455 108.830 98.625 110.190 ;
        RECT 98.990 110.020 99.315 110.805 ;
        RECT 98.795 108.970 99.255 110.020 ;
        RECT 97.070 108.660 97.925 108.830 ;
        RECT 98.130 108.660 98.625 108.830 ;
        RECT 98.795 108.440 99.125 108.800 ;
        RECT 99.485 108.700 99.655 110.820 ;
        RECT 99.825 110.490 100.155 110.990 ;
        RECT 100.325 110.320 100.580 110.820 ;
        RECT 99.830 110.150 100.580 110.320 ;
        RECT 101.065 110.150 101.235 110.990 ;
        RECT 99.830 109.160 100.060 110.150 ;
        RECT 101.445 109.980 101.695 110.820 ;
        RECT 101.905 110.150 102.075 110.990 ;
        RECT 102.245 109.980 102.535 110.820 ;
        RECT 100.230 109.330 100.580 109.980 ;
        RECT 100.810 109.810 102.535 109.980 ;
        RECT 102.745 109.930 102.915 110.990 ;
        RECT 103.210 110.610 103.540 110.990 ;
        RECT 103.720 110.440 103.890 110.730 ;
        RECT 104.060 110.530 104.310 110.990 ;
        RECT 103.090 110.270 103.890 110.440 ;
        RECT 104.480 110.480 105.350 110.820 ;
        RECT 100.810 109.260 101.220 109.810 ;
        RECT 103.090 109.650 103.260 110.270 ;
        RECT 104.480 110.100 104.650 110.480 ;
        RECT 105.585 110.360 105.755 110.820 ;
        RECT 105.925 110.530 106.295 110.990 ;
        RECT 106.590 110.390 106.760 110.730 ;
        RECT 106.930 110.560 107.260 110.990 ;
        RECT 107.495 110.390 107.665 110.730 ;
        RECT 103.430 109.930 104.650 110.100 ;
        RECT 104.820 110.020 105.280 110.310 ;
        RECT 105.585 110.190 106.145 110.360 ;
        RECT 106.590 110.220 107.665 110.390 ;
        RECT 107.835 110.490 108.515 110.820 ;
        RECT 108.730 110.490 108.980 110.820 ;
        RECT 109.150 110.530 109.400 110.990 ;
        RECT 105.975 110.050 106.145 110.190 ;
        RECT 104.820 110.010 105.785 110.020 ;
        RECT 104.480 109.840 104.650 109.930 ;
        RECT 105.110 109.850 105.785 110.010 ;
        RECT 103.090 109.640 103.435 109.650 ;
        RECT 101.405 109.430 103.435 109.640 ;
        RECT 99.830 108.990 100.580 109.160 ;
        RECT 100.810 109.090 102.575 109.260 ;
        RECT 99.825 108.440 100.155 108.820 ;
        RECT 100.325 108.700 100.580 108.990 ;
        RECT 101.065 108.440 101.235 108.910 ;
        RECT 101.405 108.610 101.735 109.090 ;
        RECT 101.905 108.440 102.075 108.910 ;
        RECT 102.245 108.610 102.575 109.090 ;
        RECT 102.745 108.440 102.915 109.250 ;
        RECT 103.110 109.175 103.435 109.430 ;
        RECT 103.115 108.820 103.435 109.175 ;
        RECT 103.605 109.390 104.145 109.760 ;
        RECT 104.480 109.670 104.885 109.840 ;
        RECT 103.605 108.990 103.845 109.390 ;
        RECT 104.325 109.220 104.545 109.500 ;
        RECT 104.015 109.050 104.545 109.220 ;
        RECT 104.015 108.820 104.185 109.050 ;
        RECT 104.715 108.890 104.885 109.670 ;
        RECT 105.055 109.060 105.405 109.680 ;
        RECT 105.575 109.060 105.785 109.850 ;
        RECT 105.975 109.880 107.475 110.050 ;
        RECT 105.975 109.190 106.145 109.880 ;
        RECT 107.835 109.710 108.005 110.490 ;
        RECT 108.810 110.360 108.980 110.490 ;
        RECT 106.315 109.540 108.005 109.710 ;
        RECT 108.175 109.930 108.640 110.320 ;
        RECT 108.810 110.190 109.205 110.360 ;
        RECT 106.315 109.360 106.485 109.540 ;
        RECT 103.115 108.650 104.185 108.820 ;
        RECT 104.355 108.440 104.545 108.880 ;
        RECT 104.715 108.610 105.665 108.890 ;
        RECT 105.975 108.800 106.235 109.190 ;
        RECT 106.655 109.120 107.445 109.370 ;
        RECT 105.885 108.630 106.235 108.800 ;
        RECT 106.445 108.440 106.775 108.900 ;
        RECT 107.650 108.830 107.820 109.540 ;
        RECT 108.175 109.340 108.345 109.930 ;
        RECT 107.990 109.120 108.345 109.340 ;
        RECT 108.515 109.120 108.865 109.740 ;
        RECT 109.035 108.830 109.205 110.190 ;
        RECT 109.570 110.020 109.895 110.805 ;
        RECT 109.375 108.970 109.835 110.020 ;
        RECT 107.650 108.660 108.505 108.830 ;
        RECT 108.710 108.660 109.205 108.830 ;
        RECT 109.375 108.440 109.705 108.800 ;
        RECT 110.065 108.700 110.235 110.820 ;
        RECT 110.405 110.490 110.735 110.990 ;
        RECT 110.905 110.320 111.160 110.820 ;
        RECT 110.410 110.150 111.160 110.320 ;
        RECT 110.410 109.160 110.640 110.150 ;
        RECT 110.810 109.330 111.160 109.980 ;
        RECT 111.395 109.850 111.605 110.990 ;
        RECT 111.775 109.840 112.105 110.820 ;
        RECT 112.275 109.850 112.505 110.990 ;
        RECT 112.755 109.850 112.985 110.990 ;
        RECT 113.155 109.840 113.485 110.820 ;
        RECT 113.655 109.850 113.865 110.990 ;
        RECT 114.555 109.900 115.765 110.990 ;
        RECT 110.410 108.990 111.160 109.160 ;
        RECT 110.405 108.440 110.735 108.820 ;
        RECT 110.905 108.700 111.160 108.990 ;
        RECT 111.395 108.440 111.605 109.260 ;
        RECT 111.775 109.240 112.025 109.840 ;
        RECT 112.195 109.430 112.525 109.680 ;
        RECT 112.735 109.430 113.065 109.680 ;
        RECT 111.775 108.610 112.105 109.240 ;
        RECT 112.275 108.440 112.505 109.260 ;
        RECT 112.755 108.440 112.985 109.260 ;
        RECT 113.235 109.240 113.485 109.840 ;
        RECT 114.555 109.360 115.075 109.900 ;
        RECT 113.155 108.610 113.485 109.240 ;
        RECT 113.655 108.440 113.865 109.260 ;
        RECT 115.245 109.190 115.765 109.730 ;
        RECT 114.555 108.440 115.765 109.190 ;
        RECT 14.650 108.270 115.850 108.440 ;
        RECT 14.735 107.520 15.945 108.270 ;
        RECT 14.735 106.980 15.255 107.520 ;
        RECT 16.115 107.500 19.625 108.270 ;
        RECT 19.800 107.725 25.145 108.270 ;
        RECT 15.425 106.810 15.945 107.350 ;
        RECT 14.735 105.720 15.945 106.810 ;
        RECT 16.115 106.810 17.805 107.330 ;
        RECT 17.975 106.980 19.625 107.500 ;
        RECT 16.115 105.720 19.625 106.810 ;
        RECT 21.390 106.155 21.740 107.405 ;
        RECT 23.220 106.895 23.560 107.725 ;
        RECT 25.315 107.545 25.605 108.270 ;
        RECT 26.085 107.800 26.255 108.270 ;
        RECT 26.425 107.620 26.755 108.100 ;
        RECT 26.925 107.800 27.095 108.270 ;
        RECT 27.265 107.620 27.595 108.100 ;
        RECT 25.830 107.450 27.595 107.620 ;
        RECT 27.765 107.460 27.935 108.270 ;
        RECT 28.135 107.890 29.205 108.060 ;
        RECT 28.135 107.535 28.455 107.890 ;
        RECT 25.830 106.900 26.240 107.450 ;
        RECT 28.130 107.280 28.455 107.535 ;
        RECT 26.425 107.070 28.455 107.280 ;
        RECT 28.110 107.060 28.455 107.070 ;
        RECT 28.625 107.320 28.865 107.720 ;
        RECT 29.035 107.660 29.205 107.890 ;
        RECT 29.375 107.830 29.565 108.270 ;
        RECT 29.735 107.820 30.685 108.100 ;
        RECT 30.905 107.910 31.255 108.080 ;
        RECT 29.035 107.490 29.565 107.660 ;
        RECT 19.800 105.720 25.145 106.155 ;
        RECT 25.315 105.720 25.605 106.885 ;
        RECT 25.830 106.730 27.555 106.900 ;
        RECT 26.085 105.720 26.255 106.560 ;
        RECT 26.465 105.890 26.715 106.730 ;
        RECT 26.925 105.720 27.095 106.560 ;
        RECT 27.265 105.890 27.555 106.730 ;
        RECT 27.765 105.720 27.935 106.780 ;
        RECT 28.110 106.440 28.280 107.060 ;
        RECT 28.625 106.950 29.165 107.320 ;
        RECT 29.345 107.210 29.565 107.490 ;
        RECT 29.735 107.040 29.905 107.820 ;
        RECT 29.500 106.870 29.905 107.040 ;
        RECT 30.075 107.030 30.425 107.650 ;
        RECT 29.500 106.780 29.670 106.870 ;
        RECT 30.595 106.860 30.805 107.650 ;
        RECT 28.450 106.610 29.670 106.780 ;
        RECT 30.130 106.700 30.805 106.860 ;
        RECT 28.110 106.270 28.910 106.440 ;
        RECT 28.230 105.720 28.560 106.100 ;
        RECT 28.740 105.980 28.910 106.270 ;
        RECT 29.500 106.230 29.670 106.610 ;
        RECT 29.840 106.690 30.805 106.700 ;
        RECT 30.995 107.520 31.255 107.910 ;
        RECT 31.465 107.810 31.795 108.270 ;
        RECT 32.670 107.880 33.525 108.050 ;
        RECT 33.730 107.880 34.225 108.050 ;
        RECT 34.395 107.910 34.725 108.270 ;
        RECT 30.995 106.830 31.165 107.520 ;
        RECT 31.335 107.170 31.505 107.350 ;
        RECT 31.675 107.340 32.465 107.590 ;
        RECT 32.670 107.170 32.840 107.880 ;
        RECT 33.010 107.370 33.365 107.590 ;
        RECT 31.335 107.000 33.025 107.170 ;
        RECT 29.840 106.400 30.300 106.690 ;
        RECT 30.995 106.660 32.495 106.830 ;
        RECT 30.995 106.520 31.165 106.660 ;
        RECT 30.605 106.350 31.165 106.520 ;
        RECT 29.080 105.720 29.330 106.180 ;
        RECT 29.500 105.890 30.370 106.230 ;
        RECT 30.605 105.890 30.775 106.350 ;
        RECT 31.610 106.320 32.685 106.490 ;
        RECT 30.945 105.720 31.315 106.180 ;
        RECT 31.610 105.980 31.780 106.320 ;
        RECT 31.950 105.720 32.280 106.150 ;
        RECT 32.515 105.980 32.685 106.320 ;
        RECT 32.855 106.220 33.025 107.000 ;
        RECT 33.195 106.780 33.365 107.370 ;
        RECT 33.535 106.970 33.885 107.590 ;
        RECT 33.195 106.390 33.660 106.780 ;
        RECT 34.055 106.520 34.225 107.880 ;
        RECT 34.395 106.690 34.855 107.740 ;
        RECT 33.830 106.350 34.225 106.520 ;
        RECT 33.830 106.220 34.000 106.350 ;
        RECT 32.855 105.890 33.535 106.220 ;
        RECT 33.750 105.890 34.000 106.220 ;
        RECT 34.170 105.720 34.420 106.180 ;
        RECT 34.590 105.905 34.915 106.690 ;
        RECT 35.085 105.890 35.255 108.010 ;
        RECT 35.425 107.890 35.755 108.270 ;
        RECT 35.925 107.720 36.180 108.010 ;
        RECT 35.430 107.550 36.180 107.720 ;
        RECT 35.430 106.560 35.660 107.550 ;
        RECT 36.355 107.500 38.025 108.270 ;
        RECT 38.195 107.545 38.485 108.270 ;
        RECT 38.965 107.800 39.135 108.270 ;
        RECT 39.305 107.620 39.635 108.100 ;
        RECT 39.805 107.800 39.975 108.270 ;
        RECT 40.145 107.620 40.475 108.100 ;
        RECT 35.830 106.730 36.180 107.380 ;
        RECT 36.355 106.810 37.105 107.330 ;
        RECT 37.275 106.980 38.025 107.500 ;
        RECT 38.710 107.450 40.475 107.620 ;
        RECT 40.645 107.460 40.815 108.270 ;
        RECT 41.015 107.890 42.085 108.060 ;
        RECT 41.015 107.535 41.335 107.890 ;
        RECT 38.710 106.900 39.120 107.450 ;
        RECT 41.010 107.280 41.335 107.535 ;
        RECT 39.305 107.070 41.335 107.280 ;
        RECT 40.990 107.060 41.335 107.070 ;
        RECT 41.505 107.320 41.745 107.720 ;
        RECT 41.915 107.660 42.085 107.890 ;
        RECT 42.255 107.830 42.445 108.270 ;
        RECT 42.615 107.820 43.565 108.100 ;
        RECT 43.785 107.910 44.135 108.080 ;
        RECT 41.915 107.490 42.445 107.660 ;
        RECT 35.430 106.390 36.180 106.560 ;
        RECT 35.425 105.720 35.755 106.220 ;
        RECT 35.925 105.890 36.180 106.390 ;
        RECT 36.355 105.720 38.025 106.810 ;
        RECT 38.195 105.720 38.485 106.885 ;
        RECT 38.710 106.730 40.435 106.900 ;
        RECT 38.965 105.720 39.135 106.560 ;
        RECT 39.345 105.890 39.595 106.730 ;
        RECT 39.805 105.720 39.975 106.560 ;
        RECT 40.145 105.890 40.435 106.730 ;
        RECT 40.645 105.720 40.815 106.780 ;
        RECT 40.990 106.440 41.160 107.060 ;
        RECT 41.505 106.950 42.045 107.320 ;
        RECT 42.225 107.210 42.445 107.490 ;
        RECT 42.615 107.040 42.785 107.820 ;
        RECT 42.380 106.870 42.785 107.040 ;
        RECT 42.955 107.030 43.305 107.650 ;
        RECT 42.380 106.780 42.550 106.870 ;
        RECT 43.475 106.860 43.685 107.650 ;
        RECT 41.330 106.610 42.550 106.780 ;
        RECT 43.010 106.700 43.685 106.860 ;
        RECT 40.990 106.270 41.790 106.440 ;
        RECT 41.110 105.720 41.440 106.100 ;
        RECT 41.620 105.980 41.790 106.270 ;
        RECT 42.380 106.230 42.550 106.610 ;
        RECT 42.720 106.690 43.685 106.700 ;
        RECT 43.875 107.520 44.135 107.910 ;
        RECT 44.345 107.810 44.675 108.270 ;
        RECT 45.550 107.880 46.405 108.050 ;
        RECT 46.610 107.880 47.105 108.050 ;
        RECT 47.275 107.910 47.605 108.270 ;
        RECT 43.875 106.830 44.045 107.520 ;
        RECT 44.215 107.170 44.385 107.350 ;
        RECT 44.555 107.340 45.345 107.590 ;
        RECT 45.550 107.170 45.720 107.880 ;
        RECT 45.890 107.370 46.245 107.590 ;
        RECT 44.215 107.000 45.905 107.170 ;
        RECT 42.720 106.400 43.180 106.690 ;
        RECT 43.875 106.660 45.375 106.830 ;
        RECT 43.875 106.520 44.045 106.660 ;
        RECT 43.485 106.350 44.045 106.520 ;
        RECT 41.960 105.720 42.210 106.180 ;
        RECT 42.380 105.890 43.250 106.230 ;
        RECT 43.485 105.890 43.655 106.350 ;
        RECT 44.490 106.320 45.565 106.490 ;
        RECT 43.825 105.720 44.195 106.180 ;
        RECT 44.490 105.980 44.660 106.320 ;
        RECT 44.830 105.720 45.160 106.150 ;
        RECT 45.395 105.980 45.565 106.320 ;
        RECT 45.735 106.220 45.905 107.000 ;
        RECT 46.075 106.780 46.245 107.370 ;
        RECT 46.415 106.970 46.765 107.590 ;
        RECT 46.075 106.390 46.540 106.780 ;
        RECT 46.935 106.520 47.105 107.880 ;
        RECT 47.275 106.690 47.735 107.740 ;
        RECT 46.710 106.350 47.105 106.520 ;
        RECT 46.710 106.220 46.880 106.350 ;
        RECT 45.735 105.890 46.415 106.220 ;
        RECT 46.630 105.890 46.880 106.220 ;
        RECT 47.050 105.720 47.300 106.180 ;
        RECT 47.470 105.905 47.795 106.690 ;
        RECT 47.965 105.890 48.135 108.010 ;
        RECT 48.305 107.890 48.635 108.270 ;
        RECT 48.805 107.720 49.060 108.010 ;
        RECT 48.310 107.550 49.060 107.720 ;
        RECT 48.310 106.560 48.540 107.550 ;
        RECT 49.235 107.500 50.905 108.270 ;
        RECT 51.075 107.545 51.365 108.270 ;
        RECT 51.535 107.520 52.745 108.270 ;
        RECT 48.710 106.730 49.060 107.380 ;
        RECT 49.235 106.810 49.985 107.330 ;
        RECT 50.155 106.980 50.905 107.500 ;
        RECT 48.310 106.390 49.060 106.560 ;
        RECT 48.305 105.720 48.635 106.220 ;
        RECT 48.805 105.890 49.060 106.390 ;
        RECT 49.235 105.720 50.905 106.810 ;
        RECT 51.075 105.720 51.365 106.885 ;
        RECT 51.535 106.810 52.055 107.350 ;
        RECT 52.225 106.980 52.745 107.520 ;
        RECT 52.975 107.450 53.185 108.270 ;
        RECT 53.355 107.470 53.685 108.100 ;
        RECT 53.355 106.870 53.605 107.470 ;
        RECT 53.855 107.450 54.085 108.270 ;
        RECT 54.295 107.500 57.805 108.270 ;
        RECT 53.775 107.030 54.105 107.280 ;
        RECT 51.535 105.720 52.745 106.810 ;
        RECT 52.975 105.720 53.185 106.860 ;
        RECT 53.355 105.890 53.685 106.870 ;
        RECT 53.855 105.720 54.085 106.860 ;
        RECT 54.295 106.810 55.985 107.330 ;
        RECT 56.155 106.980 57.805 107.500 ;
        RECT 58.035 107.450 58.245 108.270 ;
        RECT 58.415 107.470 58.745 108.100 ;
        RECT 58.415 106.870 58.665 107.470 ;
        RECT 58.915 107.450 59.145 108.270 ;
        RECT 60.275 107.500 63.785 108.270 ;
        RECT 63.955 107.545 64.245 108.270 ;
        RECT 64.415 107.500 66.085 108.270 ;
        RECT 66.565 107.800 66.735 108.270 ;
        RECT 66.905 107.620 67.235 108.100 ;
        RECT 67.405 107.800 67.575 108.270 ;
        RECT 67.745 107.620 68.075 108.100 ;
        RECT 58.835 107.030 59.165 107.280 ;
        RECT 54.295 105.720 57.805 106.810 ;
        RECT 58.035 105.720 58.245 106.860 ;
        RECT 58.415 105.890 58.745 106.870 ;
        RECT 58.915 105.720 59.145 106.860 ;
        RECT 60.275 106.810 61.965 107.330 ;
        RECT 62.135 106.980 63.785 107.500 ;
        RECT 60.275 105.720 63.785 106.810 ;
        RECT 63.955 105.720 64.245 106.885 ;
        RECT 64.415 106.810 65.165 107.330 ;
        RECT 65.335 106.980 66.085 107.500 ;
        RECT 66.310 107.450 68.075 107.620 ;
        RECT 68.245 107.460 68.415 108.270 ;
        RECT 68.615 107.890 69.685 108.060 ;
        RECT 68.615 107.535 68.935 107.890 ;
        RECT 66.310 106.900 66.720 107.450 ;
        RECT 68.610 107.280 68.935 107.535 ;
        RECT 66.905 107.070 68.935 107.280 ;
        RECT 68.590 107.060 68.935 107.070 ;
        RECT 69.105 107.320 69.345 107.720 ;
        RECT 69.515 107.660 69.685 107.890 ;
        RECT 69.855 107.830 70.045 108.270 ;
        RECT 70.215 107.820 71.165 108.100 ;
        RECT 71.385 107.910 71.735 108.080 ;
        RECT 69.515 107.490 70.045 107.660 ;
        RECT 64.415 105.720 66.085 106.810 ;
        RECT 66.310 106.730 68.035 106.900 ;
        RECT 66.565 105.720 66.735 106.560 ;
        RECT 66.945 105.890 67.195 106.730 ;
        RECT 67.405 105.720 67.575 106.560 ;
        RECT 67.745 105.890 68.035 106.730 ;
        RECT 68.245 105.720 68.415 106.780 ;
        RECT 68.590 106.440 68.760 107.060 ;
        RECT 69.105 106.950 69.645 107.320 ;
        RECT 69.825 107.210 70.045 107.490 ;
        RECT 70.215 107.040 70.385 107.820 ;
        RECT 69.980 106.870 70.385 107.040 ;
        RECT 70.555 107.030 70.905 107.650 ;
        RECT 69.980 106.780 70.150 106.870 ;
        RECT 71.075 106.860 71.285 107.650 ;
        RECT 68.930 106.610 70.150 106.780 ;
        RECT 70.610 106.700 71.285 106.860 ;
        RECT 68.590 106.270 69.390 106.440 ;
        RECT 68.710 105.720 69.040 106.100 ;
        RECT 69.220 105.980 69.390 106.270 ;
        RECT 69.980 106.230 70.150 106.610 ;
        RECT 70.320 106.690 71.285 106.700 ;
        RECT 71.475 107.520 71.735 107.910 ;
        RECT 71.945 107.810 72.275 108.270 ;
        RECT 73.150 107.880 74.005 108.050 ;
        RECT 74.210 107.880 74.705 108.050 ;
        RECT 74.875 107.910 75.205 108.270 ;
        RECT 71.475 106.830 71.645 107.520 ;
        RECT 71.815 107.170 71.985 107.350 ;
        RECT 72.155 107.340 72.945 107.590 ;
        RECT 73.150 107.170 73.320 107.880 ;
        RECT 73.490 107.370 73.845 107.590 ;
        RECT 71.815 107.000 73.505 107.170 ;
        RECT 70.320 106.400 70.780 106.690 ;
        RECT 71.475 106.660 72.975 106.830 ;
        RECT 71.475 106.520 71.645 106.660 ;
        RECT 71.085 106.350 71.645 106.520 ;
        RECT 69.560 105.720 69.810 106.180 ;
        RECT 69.980 105.890 70.850 106.230 ;
        RECT 71.085 105.890 71.255 106.350 ;
        RECT 72.090 106.320 73.165 106.490 ;
        RECT 71.425 105.720 71.795 106.180 ;
        RECT 72.090 105.980 72.260 106.320 ;
        RECT 72.430 105.720 72.760 106.150 ;
        RECT 72.995 105.980 73.165 106.320 ;
        RECT 73.335 106.220 73.505 107.000 ;
        RECT 73.675 106.780 73.845 107.370 ;
        RECT 74.015 106.970 74.365 107.590 ;
        RECT 73.675 106.390 74.140 106.780 ;
        RECT 74.535 106.520 74.705 107.880 ;
        RECT 74.875 106.690 75.335 107.740 ;
        RECT 74.310 106.350 74.705 106.520 ;
        RECT 74.310 106.220 74.480 106.350 ;
        RECT 73.335 105.890 74.015 106.220 ;
        RECT 74.230 105.890 74.480 106.220 ;
        RECT 74.650 105.720 74.900 106.180 ;
        RECT 75.070 105.905 75.395 106.690 ;
        RECT 75.565 105.890 75.735 108.010 ;
        RECT 75.905 107.890 76.235 108.270 ;
        RECT 76.405 107.720 76.660 108.010 ;
        RECT 75.910 107.550 76.660 107.720 ;
        RECT 75.910 106.560 76.140 107.550 ;
        RECT 76.835 107.545 77.125 108.270 ;
        RECT 77.355 107.450 77.565 108.270 ;
        RECT 77.735 107.470 78.065 108.100 ;
        RECT 76.310 106.730 76.660 107.380 ;
        RECT 75.910 106.390 76.660 106.560 ;
        RECT 75.905 105.720 76.235 106.220 ;
        RECT 76.405 105.890 76.660 106.390 ;
        RECT 76.835 105.720 77.125 106.885 ;
        RECT 77.735 106.870 77.985 107.470 ;
        RECT 78.235 107.450 78.465 108.270 ;
        RECT 78.675 107.520 79.885 108.270 ;
        RECT 78.155 107.030 78.485 107.280 ;
        RECT 77.355 105.720 77.565 106.860 ;
        RECT 77.735 105.890 78.065 106.870 ;
        RECT 78.235 105.720 78.465 106.860 ;
        RECT 78.675 106.810 79.195 107.350 ;
        RECT 79.365 106.980 79.885 107.520 ;
        RECT 80.115 107.450 80.325 108.270 ;
        RECT 80.495 107.470 80.825 108.100 ;
        RECT 80.495 106.870 80.745 107.470 ;
        RECT 80.995 107.450 81.225 108.270 ;
        RECT 81.435 107.500 84.025 108.270 ;
        RECT 84.200 107.725 89.545 108.270 ;
        RECT 80.915 107.030 81.245 107.280 ;
        RECT 78.675 105.720 79.885 106.810 ;
        RECT 80.115 105.720 80.325 106.860 ;
        RECT 80.495 105.890 80.825 106.870 ;
        RECT 80.995 105.720 81.225 106.860 ;
        RECT 81.435 106.810 82.645 107.330 ;
        RECT 82.815 106.980 84.025 107.500 ;
        RECT 81.435 105.720 84.025 106.810 ;
        RECT 85.790 106.155 86.140 107.405 ;
        RECT 87.620 106.895 87.960 107.725 ;
        RECT 89.715 107.545 90.005 108.270 ;
        RECT 90.180 107.725 95.525 108.270 ;
        RECT 84.200 105.720 89.545 106.155 ;
        RECT 89.715 105.720 90.005 106.885 ;
        RECT 91.770 106.155 92.120 107.405 ;
        RECT 93.600 106.895 93.940 107.725 ;
        RECT 95.755 107.450 95.965 108.270 ;
        RECT 96.135 107.470 96.465 108.100 ;
        RECT 96.135 106.870 96.385 107.470 ;
        RECT 96.635 107.450 96.865 108.270 ;
        RECT 97.535 107.500 100.125 108.270 ;
        RECT 96.555 107.030 96.885 107.280 ;
        RECT 90.180 105.720 95.525 106.155 ;
        RECT 95.755 105.720 95.965 106.860 ;
        RECT 96.135 105.890 96.465 106.870 ;
        RECT 96.635 105.720 96.865 106.860 ;
        RECT 97.535 106.810 98.745 107.330 ;
        RECT 98.915 106.980 100.125 107.500 ;
        RECT 100.335 107.450 100.565 108.270 ;
        RECT 100.735 107.470 101.065 108.100 ;
        RECT 100.315 107.030 100.645 107.280 ;
        RECT 100.815 106.870 101.065 107.470 ;
        RECT 101.235 107.450 101.445 108.270 ;
        RECT 102.595 107.545 102.885 108.270 ;
        RECT 103.980 107.720 104.235 108.010 ;
        RECT 104.405 107.890 104.735 108.270 ;
        RECT 103.980 107.550 104.730 107.720 ;
        RECT 97.535 105.720 100.125 106.810 ;
        RECT 100.335 105.720 100.565 106.860 ;
        RECT 100.735 105.890 101.065 106.870 ;
        RECT 101.235 105.720 101.445 106.860 ;
        RECT 102.595 105.720 102.885 106.885 ;
        RECT 103.980 106.730 104.330 107.380 ;
        RECT 104.500 106.560 104.730 107.550 ;
        RECT 103.980 106.390 104.730 106.560 ;
        RECT 103.980 105.890 104.235 106.390 ;
        RECT 104.405 105.720 104.735 106.220 ;
        RECT 104.905 105.890 105.075 108.010 ;
        RECT 105.435 107.910 105.765 108.270 ;
        RECT 105.935 107.880 106.430 108.050 ;
        RECT 106.635 107.880 107.490 108.050 ;
        RECT 105.305 106.690 105.765 107.740 ;
        RECT 105.245 105.905 105.570 106.690 ;
        RECT 105.935 106.520 106.105 107.880 ;
        RECT 106.275 106.970 106.625 107.590 ;
        RECT 106.795 107.370 107.150 107.590 ;
        RECT 106.795 106.780 106.965 107.370 ;
        RECT 107.320 107.170 107.490 107.880 ;
        RECT 108.365 107.810 108.695 108.270 ;
        RECT 108.905 107.910 109.255 108.080 ;
        RECT 107.695 107.340 108.485 107.590 ;
        RECT 108.905 107.520 109.165 107.910 ;
        RECT 109.475 107.820 110.425 108.100 ;
        RECT 110.595 107.830 110.785 108.270 ;
        RECT 110.955 107.890 112.025 108.060 ;
        RECT 108.655 107.170 108.825 107.350 ;
        RECT 105.935 106.350 106.330 106.520 ;
        RECT 106.500 106.390 106.965 106.780 ;
        RECT 107.135 107.000 108.825 107.170 ;
        RECT 106.160 106.220 106.330 106.350 ;
        RECT 107.135 106.220 107.305 107.000 ;
        RECT 108.995 106.830 109.165 107.520 ;
        RECT 107.665 106.660 109.165 106.830 ;
        RECT 109.355 106.860 109.565 107.650 ;
        RECT 109.735 107.030 110.085 107.650 ;
        RECT 110.255 107.040 110.425 107.820 ;
        RECT 110.955 107.660 111.125 107.890 ;
        RECT 110.595 107.490 111.125 107.660 ;
        RECT 110.595 107.210 110.815 107.490 ;
        RECT 111.295 107.320 111.535 107.720 ;
        RECT 110.255 106.870 110.660 107.040 ;
        RECT 110.995 106.950 111.535 107.320 ;
        RECT 111.705 107.535 112.025 107.890 ;
        RECT 111.705 107.280 112.030 107.535 ;
        RECT 112.225 107.460 112.395 108.270 ;
        RECT 112.565 107.620 112.895 108.100 ;
        RECT 113.065 107.800 113.235 108.270 ;
        RECT 113.405 107.620 113.735 108.100 ;
        RECT 113.905 107.800 114.075 108.270 ;
        RECT 112.565 107.450 114.330 107.620 ;
        RECT 114.555 107.520 115.765 108.270 ;
        RECT 111.705 107.070 113.735 107.280 ;
        RECT 111.705 107.060 112.050 107.070 ;
        RECT 109.355 106.700 110.030 106.860 ;
        RECT 110.490 106.780 110.660 106.870 ;
        RECT 109.355 106.690 110.320 106.700 ;
        RECT 108.995 106.520 109.165 106.660 ;
        RECT 105.740 105.720 105.990 106.180 ;
        RECT 106.160 105.890 106.410 106.220 ;
        RECT 106.625 105.890 107.305 106.220 ;
        RECT 107.475 106.320 108.550 106.490 ;
        RECT 108.995 106.350 109.555 106.520 ;
        RECT 109.860 106.400 110.320 106.690 ;
        RECT 110.490 106.610 111.710 106.780 ;
        RECT 107.475 105.980 107.645 106.320 ;
        RECT 107.880 105.720 108.210 106.150 ;
        RECT 108.380 105.980 108.550 106.320 ;
        RECT 108.845 105.720 109.215 106.180 ;
        RECT 109.385 105.890 109.555 106.350 ;
        RECT 110.490 106.230 110.660 106.610 ;
        RECT 111.880 106.440 112.050 107.060 ;
        RECT 113.920 106.900 114.330 107.450 ;
        RECT 109.790 105.890 110.660 106.230 ;
        RECT 111.250 106.270 112.050 106.440 ;
        RECT 110.830 105.720 111.080 106.180 ;
        RECT 111.250 105.980 111.420 106.270 ;
        RECT 111.600 105.720 111.930 106.100 ;
        RECT 112.225 105.720 112.395 106.780 ;
        RECT 112.605 106.730 114.330 106.900 ;
        RECT 114.555 106.810 115.075 107.350 ;
        RECT 115.245 106.980 115.765 107.520 ;
        RECT 112.605 105.890 112.895 106.730 ;
        RECT 113.065 105.720 113.235 106.560 ;
        RECT 113.445 105.890 113.695 106.730 ;
        RECT 113.905 105.720 114.075 106.560 ;
        RECT 114.555 105.720 115.765 106.810 ;
        RECT 14.650 105.550 115.850 105.720 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 14.650 206.035 115.850 206.515 ;
        RECT 14.650 203.315 115.850 203.795 ;
        RECT 66.715 203.115 67.005 203.160 ;
        RECT 72.220 203.115 72.540 203.175 ;
        RECT 66.715 202.975 72.540 203.115 ;
        RECT 66.715 202.930 67.005 202.975 ;
        RECT 72.220 202.915 72.540 202.975 ;
        RECT 63.035 202.775 63.325 202.820 ;
        RECT 63.480 202.775 63.800 202.835 ;
        RECT 73.255 202.775 73.545 202.820 ;
        RECT 76.375 202.775 76.665 202.820 ;
        RECT 78.265 202.775 78.555 202.820 ;
        RECT 63.035 202.635 63.800 202.775 ;
        RECT 63.035 202.590 63.325 202.635 ;
        RECT 63.480 202.575 63.800 202.635 ;
        RECT 66.790 202.635 72.910 202.775 ;
        RECT 66.790 202.435 66.930 202.635 ;
        RECT 70.395 202.435 70.685 202.480 ;
        RECT 60.810 202.295 66.930 202.435 ;
        RECT 67.250 202.295 70.685 202.435 ;
        RECT 72.770 202.435 72.910 202.635 ;
        RECT 73.255 202.635 78.555 202.775 ;
        RECT 73.255 202.590 73.545 202.635 ;
        RECT 76.375 202.590 76.665 202.635 ;
        RECT 78.265 202.590 78.555 202.635 ;
        RECT 80.500 202.435 80.820 202.495 ;
        RECT 72.770 202.295 80.820 202.435 ;
        RECT 58.880 202.095 59.200 202.155 ;
        RECT 60.810 202.140 60.950 202.295 ;
        RECT 67.250 202.155 67.390 202.295 ;
        RECT 70.395 202.250 70.685 202.295 ;
        RECT 80.500 202.235 80.820 202.295 ;
        RECT 60.735 202.095 61.025 202.140 ;
        RECT 58.880 201.955 61.025 202.095 ;
        RECT 58.880 201.895 59.200 201.955 ;
        RECT 60.735 201.910 61.025 201.955 ;
        RECT 62.115 201.910 62.405 202.140 ;
        RECT 65.335 201.910 65.625 202.140 ;
        RECT 59.340 201.755 59.660 201.815 ;
        RECT 62.190 201.755 62.330 201.910 ;
        RECT 59.340 201.615 62.330 201.755 ;
        RECT 65.410 201.755 65.550 201.910 ;
        RECT 67.160 201.895 67.480 202.155 ;
        RECT 69.000 201.755 69.320 201.815 ;
        RECT 72.175 201.800 72.465 202.115 ;
        RECT 73.255 202.095 73.545 202.140 ;
        RECT 76.835 202.095 77.125 202.140 ;
        RECT 78.670 202.095 78.960 202.140 ;
        RECT 73.255 201.955 78.960 202.095 ;
        RECT 73.255 201.910 73.545 201.955 ;
        RECT 76.835 201.910 77.125 201.955 ;
        RECT 78.670 201.910 78.960 201.955 ;
        RECT 79.135 201.910 79.425 202.140 ;
        RECT 75.440 201.800 75.760 201.815 ;
        RECT 65.410 201.615 69.320 201.755 ;
        RECT 59.340 201.555 59.660 201.615 ;
        RECT 69.000 201.555 69.320 201.615 ;
        RECT 71.875 201.755 72.465 201.800 ;
        RECT 75.115 201.755 75.765 201.800 ;
        RECT 71.875 201.615 75.765 201.755 ;
        RECT 71.875 201.570 72.165 201.615 ;
        RECT 75.115 201.570 75.765 201.615 ;
        RECT 76.360 201.755 76.680 201.815 ;
        RECT 77.755 201.755 78.045 201.800 ;
        RECT 76.360 201.615 78.045 201.755 ;
        RECT 75.440 201.555 75.760 201.570 ;
        RECT 76.360 201.555 76.680 201.615 ;
        RECT 77.755 201.570 78.045 201.615 ;
        RECT 61.180 201.215 61.500 201.475 ;
        RECT 63.020 201.415 63.340 201.475 ;
        RECT 64.415 201.415 64.705 201.460 ;
        RECT 63.020 201.275 64.705 201.415 ;
        RECT 63.020 201.215 63.340 201.275 ;
        RECT 64.415 201.230 64.705 201.275 ;
        RECT 68.080 201.415 68.400 201.475 ;
        RECT 79.210 201.415 79.350 201.910 ;
        RECT 81.880 201.415 82.200 201.475 ;
        RECT 68.080 201.275 82.200 201.415 ;
        RECT 68.080 201.215 68.400 201.275 ;
        RECT 81.880 201.215 82.200 201.275 ;
        RECT 14.650 200.595 115.850 201.075 ;
        RECT 69.475 200.210 69.765 200.440 ;
        RECT 75.915 200.395 76.205 200.440 ;
        RECT 76.360 200.395 76.680 200.455 ;
        RECT 80.055 200.395 80.345 200.440 ;
        RECT 75.915 200.255 76.680 200.395 ;
        RECT 75.915 200.210 76.205 200.255 ;
        RECT 60.835 200.055 61.125 200.100 ;
        RECT 64.075 200.055 64.725 200.100 ;
        RECT 60.835 199.915 64.725 200.055 ;
        RECT 60.835 199.870 61.425 199.915 ;
        RECT 64.075 199.870 64.725 199.915 ;
        RECT 66.715 200.055 67.005 200.100 ;
        RECT 69.550 200.055 69.690 200.210 ;
        RECT 76.360 200.195 76.680 200.255 ;
        RECT 76.910 200.255 80.345 200.395 ;
        RECT 66.715 199.915 69.690 200.055 ;
        RECT 66.715 199.870 67.005 199.915 ;
        RECT 61.135 199.775 61.425 199.870 ;
        RECT 72.680 199.855 73.000 200.115 ;
        RECT 75.440 200.055 75.760 200.115 ;
        RECT 76.910 200.055 77.050 200.255 ;
        RECT 80.055 200.210 80.345 200.255 ;
        RECT 75.440 199.915 77.050 200.055 ;
        RECT 78.135 200.055 78.425 200.100 ;
        RECT 78.660 200.055 78.980 200.115 ;
        RECT 79.135 200.055 79.425 200.100 ;
        RECT 75.440 199.855 75.760 199.915 ;
        RECT 78.135 199.870 78.430 200.055 ;
        RECT 58.880 199.515 59.200 199.775 ;
        RECT 61.135 199.555 61.500 199.775 ;
        RECT 61.180 199.515 61.500 199.555 ;
        RECT 62.215 199.715 62.505 199.760 ;
        RECT 65.795 199.715 66.085 199.760 ;
        RECT 67.630 199.715 67.920 199.760 ;
        RECT 62.215 199.575 67.920 199.715 ;
        RECT 62.215 199.530 62.505 199.575 ;
        RECT 65.795 199.530 66.085 199.575 ;
        RECT 67.630 199.530 67.920 199.575 ;
        RECT 71.300 199.515 71.620 199.775 ;
        RECT 72.220 199.715 72.540 199.775 ;
        RECT 73.615 199.715 73.905 199.760 ;
        RECT 72.220 199.575 73.905 199.715 ;
        RECT 72.220 199.515 72.540 199.575 ;
        RECT 73.615 199.530 73.905 199.575 ;
        RECT 74.995 199.715 75.285 199.760 ;
        RECT 74.995 199.575 77.510 199.715 ;
        RECT 74.995 199.530 75.285 199.575 ;
        RECT 68.080 199.175 68.400 199.435 ;
        RECT 71.775 199.375 72.065 199.420 ;
        RECT 76.820 199.375 77.140 199.435 ;
        RECT 71.775 199.235 77.140 199.375 ;
        RECT 71.775 199.190 72.065 199.235 ;
        RECT 76.820 199.175 77.140 199.235 ;
        RECT 62.215 199.035 62.505 199.080 ;
        RECT 65.335 199.035 65.625 199.080 ;
        RECT 67.225 199.035 67.515 199.080 ;
        RECT 62.215 198.895 67.515 199.035 ;
        RECT 62.215 198.850 62.505 198.895 ;
        RECT 65.335 198.850 65.625 198.895 ;
        RECT 67.225 198.850 67.515 198.895 ;
        RECT 72.680 199.035 73.000 199.095 ;
        RECT 76.360 199.035 76.680 199.095 ;
        RECT 77.370 199.080 77.510 199.575 ;
        RECT 78.290 199.435 78.430 199.870 ;
        RECT 78.660 199.915 79.425 200.055 ;
        RECT 78.660 199.855 78.980 199.915 ;
        RECT 79.135 199.870 79.425 199.915 ;
        RECT 80.590 199.915 83.490 200.055 ;
        RECT 80.590 199.775 80.730 199.915 ;
        RECT 80.500 199.515 80.820 199.775 ;
        RECT 80.960 199.515 81.280 199.775 ;
        RECT 83.350 199.760 83.490 199.915 ;
        RECT 83.275 199.715 83.565 199.760 ;
        RECT 86.020 199.715 86.340 199.775 ;
        RECT 83.275 199.575 86.340 199.715 ;
        RECT 83.275 199.530 83.565 199.575 ;
        RECT 86.020 199.515 86.340 199.575 ;
        RECT 78.200 199.175 78.520 199.435 ;
        RECT 72.680 198.895 76.680 199.035 ;
        RECT 72.680 198.835 73.000 198.895 ;
        RECT 76.360 198.835 76.680 198.895 ;
        RECT 77.295 198.850 77.585 199.080 ;
        RECT 79.120 199.035 79.440 199.095 ;
        RECT 82.815 199.035 83.105 199.080 ;
        RECT 79.120 198.895 83.105 199.035 ;
        RECT 79.120 198.835 79.440 198.895 ;
        RECT 82.815 198.850 83.105 198.895 ;
        RECT 58.420 198.495 58.740 198.755 ;
        RECT 59.340 198.495 59.660 198.755 ;
        RECT 74.535 198.695 74.825 198.740 ;
        RECT 78.215 198.695 78.505 198.740 ;
        RECT 74.535 198.555 78.505 198.695 ;
        RECT 74.535 198.510 74.825 198.555 ;
        RECT 78.215 198.510 78.505 198.555 ;
        RECT 81.435 198.695 81.725 198.740 ;
        RECT 82.340 198.695 82.660 198.755 ;
        RECT 81.435 198.555 82.660 198.695 ;
        RECT 81.435 198.510 81.725 198.555 ;
        RECT 82.340 198.495 82.660 198.555 ;
        RECT 14.650 197.875 115.850 198.355 ;
        RECT 54.245 197.335 54.535 197.380 ;
        RECT 56.135 197.335 56.425 197.380 ;
        RECT 59.255 197.335 59.545 197.380 ;
        RECT 54.245 197.195 59.545 197.335 ;
        RECT 54.245 197.150 54.535 197.195 ;
        RECT 56.135 197.150 56.425 197.195 ;
        RECT 59.255 197.150 59.545 197.195 ;
        RECT 63.480 197.335 63.800 197.395 ;
        RECT 69.015 197.335 69.305 197.380 ;
        RECT 63.480 197.195 69.305 197.335 ;
        RECT 63.480 197.135 63.800 197.195 ;
        RECT 69.015 197.150 69.305 197.195 ;
        RECT 69.920 197.335 70.240 197.395 ;
        RECT 70.395 197.335 70.685 197.380 ;
        RECT 69.920 197.195 70.685 197.335 ;
        RECT 54.755 196.995 55.045 197.040 ;
        RECT 63.020 196.995 63.340 197.055 ;
        RECT 54.755 196.855 63.340 196.995 ;
        RECT 54.755 196.810 55.045 196.855 ;
        RECT 63.020 196.795 63.340 196.855 ;
        RECT 66.715 196.995 67.005 197.040 ;
        RECT 67.160 196.995 67.480 197.055 ;
        RECT 66.715 196.855 67.480 196.995 ;
        RECT 69.090 196.995 69.230 197.150 ;
        RECT 69.920 197.135 70.240 197.195 ;
        RECT 70.395 197.150 70.685 197.195 ;
        RECT 76.015 197.335 76.305 197.380 ;
        RECT 79.135 197.335 79.425 197.380 ;
        RECT 81.025 197.335 81.315 197.380 ;
        RECT 82.340 197.335 82.660 197.395 ;
        RECT 97.535 197.335 97.825 197.380 ;
        RECT 99.360 197.335 99.680 197.395 ;
        RECT 76.015 197.195 81.315 197.335 ;
        RECT 76.015 197.150 76.305 197.195 ;
        RECT 79.135 197.150 79.425 197.195 ;
        RECT 81.025 197.150 81.315 197.195 ;
        RECT 81.510 197.195 82.660 197.335 ;
        RECT 71.300 196.995 71.620 197.055 ;
        RECT 69.090 196.855 71.620 196.995 ;
        RECT 66.715 196.810 67.005 196.855 ;
        RECT 67.160 196.795 67.480 196.855 ;
        RECT 53.360 196.455 53.680 196.715 ;
        RECT 53.840 196.655 54.130 196.700 ;
        RECT 55.675 196.655 55.965 196.700 ;
        RECT 59.255 196.655 59.545 196.700 ;
        RECT 53.840 196.515 59.545 196.655 ;
        RECT 53.840 196.470 54.130 196.515 ;
        RECT 55.675 196.470 55.965 196.515 ;
        RECT 59.255 196.470 59.545 196.515 ;
        RECT 57.035 196.315 57.685 196.360 ;
        RECT 58.420 196.315 58.740 196.375 ;
        RECT 60.335 196.360 60.625 196.675 ;
        RECT 63.940 196.655 64.260 196.715 ;
        RECT 65.335 196.655 65.625 196.700 ;
        RECT 69.460 196.655 69.780 196.715 ;
        RECT 70.470 196.700 70.610 196.855 ;
        RECT 71.300 196.795 71.620 196.855 ;
        RECT 71.760 196.795 72.080 197.055 ;
        RECT 72.220 196.995 72.540 197.055 ;
        RECT 73.155 196.995 73.445 197.040 ;
        RECT 72.220 196.855 73.445 196.995 ;
        RECT 72.220 196.795 72.540 196.855 ;
        RECT 73.155 196.810 73.445 196.855 ;
        RECT 80.515 196.995 80.805 197.040 ;
        RECT 81.510 196.995 81.650 197.195 ;
        RECT 82.340 197.135 82.660 197.195 ;
        RECT 94.390 197.195 99.680 197.335 ;
        RECT 80.515 196.855 81.650 196.995 ;
        RECT 80.515 196.810 80.805 196.855 ;
        RECT 81.880 196.795 82.200 197.055 ;
        RECT 94.390 197.040 94.530 197.195 ;
        RECT 97.535 197.150 97.825 197.195 ;
        RECT 99.360 197.135 99.680 197.195 ;
        RECT 100.395 197.335 100.685 197.380 ;
        RECT 103.515 197.335 103.805 197.380 ;
        RECT 105.405 197.335 105.695 197.380 ;
        RECT 100.395 197.195 105.695 197.335 ;
        RECT 100.395 197.150 100.685 197.195 ;
        RECT 103.515 197.150 103.805 197.195 ;
        RECT 105.405 197.150 105.695 197.195 ;
        RECT 94.315 196.810 94.605 197.040 ;
        RECT 99.820 196.995 100.140 197.055 ;
        RECT 104.895 196.995 105.185 197.040 ;
        RECT 99.820 196.855 105.185 196.995 ;
        RECT 99.820 196.795 100.140 196.855 ;
        RECT 104.895 196.810 105.185 196.855 ;
        RECT 69.935 196.655 70.225 196.700 ;
        RECT 63.940 196.515 65.625 196.655 ;
        RECT 63.940 196.455 64.260 196.515 ;
        RECT 65.335 196.470 65.625 196.515 ;
        RECT 69.090 196.515 70.225 196.655 ;
        RECT 69.090 196.360 69.230 196.515 ;
        RECT 69.460 196.455 69.780 196.515 ;
        RECT 69.935 196.470 70.225 196.515 ;
        RECT 70.395 196.470 70.685 196.700 ;
        RECT 60.335 196.315 60.925 196.360 ;
        RECT 57.035 196.175 60.925 196.315 ;
        RECT 57.035 196.130 57.685 196.175 ;
        RECT 58.420 196.115 58.740 196.175 ;
        RECT 60.635 196.130 60.925 196.175 ;
        RECT 63.495 196.315 63.785 196.360 ;
        RECT 69.015 196.315 69.305 196.360 ;
        RECT 72.220 196.315 72.540 196.375 ;
        RECT 74.935 196.360 75.225 196.675 ;
        RECT 76.015 196.655 76.305 196.700 ;
        RECT 79.595 196.655 79.885 196.700 ;
        RECT 81.430 196.655 81.720 196.700 ;
        RECT 76.015 196.515 81.720 196.655 ;
        RECT 76.015 196.470 76.305 196.515 ;
        RECT 79.595 196.470 79.885 196.515 ;
        RECT 81.430 196.470 81.720 196.515 ;
        RECT 63.495 196.175 69.305 196.315 ;
        RECT 63.495 196.130 63.785 196.175 ;
        RECT 69.015 196.130 69.305 196.175 ;
        RECT 69.550 196.175 72.540 196.315 ;
        RECT 64.400 195.975 64.720 196.035 ;
        RECT 66.255 195.975 66.545 196.020 ;
        RECT 69.550 195.975 69.690 196.175 ;
        RECT 72.220 196.115 72.540 196.175 ;
        RECT 74.635 196.315 75.225 196.360 ;
        RECT 77.875 196.315 78.525 196.360 ;
        RECT 79.120 196.315 79.440 196.375 ;
        RECT 74.635 196.175 79.440 196.315 ;
        RECT 74.635 196.130 74.925 196.175 ;
        RECT 77.875 196.130 78.525 196.175 ;
        RECT 79.120 196.115 79.440 196.175 ;
        RECT 97.520 196.315 97.840 196.375 ;
        RECT 99.315 196.360 99.605 196.675 ;
        RECT 100.395 196.655 100.685 196.700 ;
        RECT 103.975 196.655 104.265 196.700 ;
        RECT 105.810 196.655 106.100 196.700 ;
        RECT 100.395 196.515 106.100 196.655 ;
        RECT 100.395 196.470 100.685 196.515 ;
        RECT 103.975 196.470 104.265 196.515 ;
        RECT 105.810 196.470 106.100 196.515 ;
        RECT 106.275 196.655 106.565 196.700 ;
        RECT 109.480 196.655 109.800 196.715 ;
        RECT 106.275 196.515 109.800 196.655 ;
        RECT 106.275 196.470 106.565 196.515 ;
        RECT 109.480 196.455 109.800 196.515 ;
        RECT 99.015 196.315 99.605 196.360 ;
        RECT 102.255 196.315 102.905 196.360 ;
        RECT 97.520 196.175 102.905 196.315 ;
        RECT 97.520 196.115 97.840 196.175 ;
        RECT 99.015 196.130 99.305 196.175 ;
        RECT 102.255 196.130 102.905 196.175 ;
        RECT 64.400 195.835 69.690 195.975 ;
        RECT 70.855 195.975 71.145 196.020 ;
        RECT 72.680 195.975 73.000 196.035 ;
        RECT 73.140 195.975 73.460 196.035 ;
        RECT 70.855 195.835 73.460 195.975 ;
        RECT 64.400 195.775 64.720 195.835 ;
        RECT 66.255 195.790 66.545 195.835 ;
        RECT 70.855 195.790 71.145 195.835 ;
        RECT 72.680 195.775 73.000 195.835 ;
        RECT 73.140 195.775 73.460 195.835 ;
        RECT 97.075 195.975 97.365 196.020 ;
        RECT 100.280 195.975 100.600 196.035 ;
        RECT 97.075 195.835 100.600 195.975 ;
        RECT 97.075 195.790 97.365 195.835 ;
        RECT 100.280 195.775 100.600 195.835 ;
        RECT 14.650 195.155 115.850 195.635 ;
        RECT 59.340 194.955 59.660 195.015 ;
        RECT 65.795 194.955 66.085 195.000 ;
        RECT 59.340 194.815 66.085 194.955 ;
        RECT 59.340 194.755 59.660 194.815 ;
        RECT 65.795 194.770 66.085 194.815 ;
        RECT 69.000 194.955 69.320 195.015 ;
        RECT 73.155 194.955 73.445 195.000 ;
        RECT 69.000 194.815 73.445 194.955 ;
        RECT 69.000 194.755 69.320 194.815 ;
        RECT 73.155 194.770 73.445 194.815 ;
        RECT 75.915 194.955 76.205 195.000 ;
        RECT 76.820 194.955 77.140 195.015 ;
        RECT 75.915 194.815 77.140 194.955 ;
        RECT 75.915 194.770 76.205 194.815 ;
        RECT 76.820 194.755 77.140 194.815 ;
        RECT 86.020 194.955 86.340 195.015 ;
        RECT 86.020 194.815 97.290 194.955 ;
        RECT 86.020 194.755 86.340 194.815 ;
        RECT 53.820 194.615 54.140 194.675 ;
        RECT 63.480 194.615 63.800 194.675 ;
        RECT 48.850 194.475 54.140 194.615 ;
        RECT 48.850 194.320 48.990 194.475 ;
        RECT 53.820 194.415 54.140 194.475 ;
        RECT 63.110 194.475 63.800 194.615 ;
        RECT 48.775 194.090 49.065 194.320 ;
        RECT 50.155 194.090 50.445 194.320 ;
        RECT 41.415 193.935 41.705 193.980 ;
        RECT 42.780 193.935 43.100 193.995 ;
        RECT 41.415 193.795 43.100 193.935 ;
        RECT 41.415 193.750 41.705 193.795 ;
        RECT 42.780 193.735 43.100 193.795 ;
        RECT 46.460 193.935 46.780 193.995 ;
        RECT 50.230 193.935 50.370 194.090 ;
        RECT 62.100 194.075 62.420 194.335 ;
        RECT 62.560 194.075 62.880 194.335 ;
        RECT 63.110 194.320 63.250 194.475 ;
        RECT 63.480 194.415 63.800 194.475 ;
        RECT 64.860 194.615 65.180 194.675 ;
        RECT 66.255 194.615 66.545 194.660 ;
        RECT 64.860 194.475 66.545 194.615 ;
        RECT 64.860 194.415 65.180 194.475 ;
        RECT 66.255 194.430 66.545 194.475 ;
        RECT 67.620 194.615 67.940 194.675 ;
        RECT 73.915 194.615 74.205 194.660 ;
        RECT 67.620 194.475 74.205 194.615 ;
        RECT 67.620 194.415 67.940 194.475 ;
        RECT 73.915 194.430 74.205 194.475 ;
        RECT 74.980 194.615 75.300 194.675 ;
        RECT 78.200 194.615 78.520 194.675 ;
        RECT 74.980 194.475 78.520 194.615 ;
        RECT 74.980 194.415 75.300 194.475 ;
        RECT 78.200 194.415 78.520 194.475 ;
        RECT 86.495 194.615 86.785 194.660 ;
        RECT 91.075 194.615 91.725 194.660 ;
        RECT 94.675 194.615 94.965 194.660 ;
        RECT 86.495 194.475 94.965 194.615 ;
        RECT 86.495 194.430 86.785 194.475 ;
        RECT 91.075 194.430 91.725 194.475 ;
        RECT 94.375 194.430 94.965 194.475 ;
        RECT 63.035 194.090 63.325 194.320 ;
        RECT 64.415 194.275 64.705 194.320 ;
        RECT 69.935 194.275 70.225 194.320 ;
        RECT 72.220 194.275 72.540 194.335 ;
        RECT 64.415 194.135 66.470 194.275 ;
        RECT 64.415 194.090 64.705 194.135 ;
        RECT 46.460 193.795 50.370 193.935 ;
        RECT 61.655 193.935 61.945 193.980 ;
        RECT 64.490 193.935 64.630 194.090 ;
        RECT 61.655 193.795 64.630 193.935 ;
        RECT 46.460 193.735 46.780 193.795 ;
        RECT 61.655 193.750 61.945 193.795 ;
        RECT 66.330 193.595 66.470 194.135 ;
        RECT 69.935 194.135 72.540 194.275 ;
        RECT 69.935 194.090 70.225 194.135 ;
        RECT 72.220 194.075 72.540 194.135 ;
        RECT 75.455 194.090 75.745 194.320 ;
        RECT 66.700 193.980 67.020 193.995 ;
        RECT 66.700 193.750 67.130 193.980 ;
        RECT 71.760 193.935 72.080 193.995 ;
        RECT 75.530 193.935 75.670 194.090 ;
        RECT 76.360 194.075 76.680 194.335 ;
        RECT 82.340 194.275 82.660 194.335 ;
        RECT 83.275 194.275 83.565 194.320 ;
        RECT 82.340 194.135 83.565 194.275 ;
        RECT 82.340 194.075 82.660 194.135 ;
        RECT 83.275 194.090 83.565 194.135 ;
        RECT 86.020 194.075 86.340 194.335 ;
        RECT 87.880 194.275 88.170 194.320 ;
        RECT 89.715 194.275 90.005 194.320 ;
        RECT 93.295 194.275 93.585 194.320 ;
        RECT 87.880 194.135 93.585 194.275 ;
        RECT 87.880 194.090 88.170 194.135 ;
        RECT 89.715 194.090 90.005 194.135 ;
        RECT 93.295 194.090 93.585 194.135 ;
        RECT 94.375 194.115 94.665 194.430 ;
        RECT 97.150 194.320 97.290 194.815 ;
        RECT 97.520 194.755 97.840 195.015 ;
        RECT 100.280 194.755 100.600 195.015 ;
        RECT 106.275 194.615 106.565 194.660 ;
        RECT 106.275 194.475 108.330 194.615 ;
        RECT 106.275 194.430 106.565 194.475 ;
        RECT 97.075 194.275 97.365 194.320 ;
        RECT 100.740 194.275 101.060 194.335 ;
        RECT 108.190 194.320 108.330 194.475 ;
        RECT 106.735 194.275 107.025 194.320 ;
        RECT 97.075 194.135 107.025 194.275 ;
        RECT 97.075 194.090 97.365 194.135 ;
        RECT 100.740 194.075 101.060 194.135 ;
        RECT 106.735 194.090 107.025 194.135 ;
        RECT 108.115 194.090 108.405 194.320 ;
        RECT 71.760 193.795 75.670 193.935 ;
        RECT 81.880 193.935 82.200 193.995 ;
        RECT 86.480 193.935 86.800 193.995 ;
        RECT 87.415 193.935 87.705 193.980 ;
        RECT 81.880 193.795 87.705 193.935 ;
        RECT 66.700 193.735 67.020 193.750 ;
        RECT 71.760 193.735 72.080 193.795 ;
        RECT 81.880 193.735 82.200 193.795 ;
        RECT 86.480 193.735 86.800 193.795 ;
        RECT 87.415 193.750 87.705 193.795 ;
        RECT 88.780 193.735 89.100 193.995 ;
        RECT 98.900 193.735 99.220 193.995 ;
        RECT 99.835 193.935 100.125 193.980 ;
        RECT 101.660 193.935 101.980 193.995 ;
        RECT 99.835 193.795 101.980 193.935 ;
        RECT 99.835 193.750 100.125 193.795 ;
        RECT 101.660 193.735 101.980 193.795 ;
        RECT 103.055 193.750 103.345 193.980 ;
        RECT 69.460 193.595 69.780 193.655 ;
        RECT 66.330 193.455 69.780 193.595 ;
        RECT 69.460 193.395 69.780 193.455 ;
        RECT 69.920 193.595 70.240 193.655 ;
        RECT 88.285 193.595 88.575 193.640 ;
        RECT 90.175 193.595 90.465 193.640 ;
        RECT 93.295 193.595 93.585 193.640 ;
        RECT 69.920 193.455 74.290 193.595 ;
        RECT 69.920 193.395 70.240 193.455 ;
        RECT 44.160 193.055 44.480 193.315 ;
        RECT 48.300 193.055 48.620 193.315 ;
        RECT 49.220 193.055 49.540 193.315 ;
        RECT 63.955 193.255 64.245 193.300 ;
        RECT 67.160 193.255 67.480 193.315 ;
        RECT 63.955 193.115 67.480 193.255 ;
        RECT 63.955 193.070 64.245 193.115 ;
        RECT 67.160 193.055 67.480 193.115 ;
        RECT 67.635 193.255 67.925 193.300 ;
        RECT 70.380 193.255 70.700 193.315 ;
        RECT 67.635 193.115 70.700 193.255 ;
        RECT 67.635 193.070 67.925 193.115 ;
        RECT 70.380 193.055 70.700 193.115 ;
        RECT 72.680 193.055 73.000 193.315 ;
        RECT 74.150 193.300 74.290 193.455 ;
        RECT 88.285 193.455 93.585 193.595 ;
        RECT 88.285 193.410 88.575 193.455 ;
        RECT 90.175 193.410 90.465 193.455 ;
        RECT 93.295 193.410 93.585 193.455 ;
        RECT 102.135 193.595 102.425 193.640 ;
        RECT 103.130 193.595 103.270 193.750 ;
        RECT 102.135 193.455 103.270 193.595 ;
        RECT 102.135 193.410 102.425 193.455 ;
        RECT 74.075 193.070 74.365 193.300 ;
        RECT 84.180 193.055 84.500 193.315 ;
        RECT 93.840 193.255 94.160 193.315 ;
        RECT 96.155 193.255 96.445 193.300 ;
        RECT 93.840 193.115 96.445 193.255 ;
        RECT 93.840 193.055 94.160 193.115 ;
        RECT 96.155 193.070 96.445 193.115 ;
        RECT 107.180 193.055 107.500 193.315 ;
        RECT 108.560 193.255 108.880 193.315 ;
        RECT 109.035 193.255 109.325 193.300 ;
        RECT 108.560 193.115 109.325 193.255 ;
        RECT 108.560 193.055 108.880 193.115 ;
        RECT 109.035 193.070 109.325 193.115 ;
        RECT 14.650 192.435 115.850 192.915 ;
        RECT 46.000 192.235 46.320 192.295 ;
        RECT 49.695 192.235 49.985 192.280 ;
        RECT 46.000 192.095 49.985 192.235 ;
        RECT 46.000 192.035 46.320 192.095 ;
        RECT 49.695 192.050 49.985 192.095 ;
        RECT 60.720 192.235 61.040 192.295 ;
        RECT 66.715 192.235 67.005 192.280 ;
        RECT 60.720 192.095 67.005 192.235 ;
        RECT 60.720 192.035 61.040 192.095 ;
        RECT 66.715 192.050 67.005 192.095 ;
        RECT 71.300 192.035 71.620 192.295 ;
        RECT 73.140 192.235 73.460 192.295 ;
        RECT 73.615 192.235 73.905 192.280 ;
        RECT 76.360 192.235 76.680 192.295 ;
        RECT 71.850 192.095 76.680 192.235 ;
        RECT 43.355 191.895 43.645 191.940 ;
        RECT 46.475 191.895 46.765 191.940 ;
        RECT 48.365 191.895 48.655 191.940 ;
        RECT 49.220 191.895 49.540 191.955 ;
        RECT 43.355 191.755 48.655 191.895 ;
        RECT 43.355 191.710 43.645 191.755 ;
        RECT 46.475 191.710 46.765 191.755 ;
        RECT 48.365 191.710 48.655 191.755 ;
        RECT 48.850 191.755 49.540 191.895 ;
        RECT 31.740 191.555 32.060 191.615 ;
        RECT 34.515 191.555 34.805 191.600 ;
        RECT 31.740 191.415 34.805 191.555 ;
        RECT 31.740 191.355 32.060 191.415 ;
        RECT 34.515 191.370 34.805 191.415 ;
        RECT 47.855 191.555 48.145 191.600 ;
        RECT 48.850 191.555 48.990 191.755 ;
        RECT 49.220 191.695 49.540 191.755 ;
        RECT 52.555 191.895 52.845 191.940 ;
        RECT 55.675 191.895 55.965 191.940 ;
        RECT 57.565 191.895 57.855 191.940 ;
        RECT 52.555 191.755 57.855 191.895 ;
        RECT 52.555 191.710 52.845 191.755 ;
        RECT 55.675 191.710 55.965 191.755 ;
        RECT 57.565 191.710 57.855 191.755 ;
        RECT 69.015 191.895 69.305 191.940 ;
        RECT 69.015 191.755 71.070 191.895 ;
        RECT 69.015 191.710 69.305 191.755 ;
        RECT 51.980 191.555 52.300 191.615 ;
        RECT 53.360 191.555 53.680 191.615 ;
        RECT 62.100 191.555 62.420 191.615 ;
        RECT 67.635 191.555 67.925 191.600 ;
        RECT 68.540 191.555 68.860 191.615 ;
        RECT 70.930 191.600 71.070 191.755 ;
        RECT 47.855 191.415 48.990 191.555 ;
        RECT 49.310 191.415 58.650 191.555 ;
        RECT 47.855 191.370 48.145 191.415 ;
        RECT 27.155 191.215 27.445 191.260 ;
        RECT 30.820 191.215 31.140 191.275 ;
        RECT 27.155 191.075 31.140 191.215 ;
        RECT 27.155 191.030 27.445 191.075 ;
        RECT 30.820 191.015 31.140 191.075 ;
        RECT 32.675 191.215 32.965 191.260 ;
        RECT 37.260 191.215 37.580 191.275 ;
        RECT 49.310 191.260 49.450 191.415 ;
        RECT 51.980 191.355 52.300 191.415 ;
        RECT 53.360 191.355 53.680 191.415 ;
        RECT 38.655 191.215 38.945 191.260 ;
        RECT 32.675 191.075 37.580 191.215 ;
        RECT 32.675 191.030 32.965 191.075 ;
        RECT 37.260 191.015 37.580 191.075 ;
        RECT 37.810 191.075 38.945 191.215 ;
        RECT 29.915 190.875 30.205 190.920 ;
        RECT 35.895 190.875 36.185 190.920 ;
        RECT 29.915 190.735 36.185 190.875 ;
        RECT 29.915 190.690 30.205 190.735 ;
        RECT 35.895 190.690 36.185 190.735 ;
        RECT 33.120 190.335 33.440 190.595 ;
        RECT 34.040 190.535 34.360 190.595 ;
        RECT 37.810 190.580 37.950 191.075 ;
        RECT 38.655 191.030 38.945 191.075 ;
        RECT 42.275 190.920 42.565 191.235 ;
        RECT 43.355 191.215 43.645 191.260 ;
        RECT 46.935 191.215 47.225 191.260 ;
        RECT 48.770 191.215 49.060 191.260 ;
        RECT 43.355 191.075 49.060 191.215 ;
        RECT 43.355 191.030 43.645 191.075 ;
        RECT 46.935 191.030 47.225 191.075 ;
        RECT 48.770 191.030 49.060 191.075 ;
        RECT 49.235 191.030 49.525 191.260 ;
        RECT 51.520 191.235 51.840 191.275 ;
        RECT 58.510 191.260 58.650 191.415 ;
        RECT 62.100 191.415 70.150 191.555 ;
        RECT 62.100 191.355 62.420 191.415 ;
        RECT 67.635 191.370 67.925 191.415 ;
        RECT 68.540 191.355 68.860 191.415 ;
        RECT 51.475 191.015 51.840 191.235 ;
        RECT 52.555 191.215 52.845 191.260 ;
        RECT 56.135 191.215 56.425 191.260 ;
        RECT 57.970 191.215 58.260 191.260 ;
        RECT 52.555 191.075 58.260 191.215 ;
        RECT 52.555 191.030 52.845 191.075 ;
        RECT 56.135 191.030 56.425 191.075 ;
        RECT 57.970 191.030 58.260 191.075 ;
        RECT 58.435 191.030 58.725 191.260 ;
        RECT 58.880 191.015 59.200 191.275 ;
        RECT 60.720 191.015 61.040 191.275 ;
        RECT 62.560 191.215 62.880 191.275 ;
        RECT 66.255 191.215 66.545 191.260 ;
        RECT 62.560 191.075 66.545 191.215 ;
        RECT 62.560 191.015 62.880 191.075 ;
        RECT 66.255 191.030 66.545 191.075 ;
        RECT 41.975 190.875 42.565 190.920 ;
        RECT 45.215 190.875 45.865 190.920 ;
        RECT 48.300 190.875 48.620 190.935 ;
        RECT 51.475 190.920 51.765 191.015 ;
        RECT 41.975 190.735 48.620 190.875 ;
        RECT 41.975 190.690 42.265 190.735 ;
        RECT 45.215 190.690 45.865 190.735 ;
        RECT 48.300 190.675 48.620 190.735 ;
        RECT 51.175 190.875 51.765 190.920 ;
        RECT 54.415 190.875 55.065 190.920 ;
        RECT 51.175 190.735 55.065 190.875 ;
        RECT 51.175 190.690 51.465 190.735 ;
        RECT 54.415 190.690 55.065 190.735 ;
        RECT 55.660 190.875 55.980 190.935 ;
        RECT 57.055 190.875 57.345 190.920 ;
        RECT 55.660 190.735 57.345 190.875 ;
        RECT 66.330 190.875 66.470 191.030 ;
        RECT 69.460 191.015 69.780 191.275 ;
        RECT 70.010 191.215 70.150 191.415 ;
        RECT 70.855 191.370 71.145 191.600 ;
        RECT 71.850 191.555 71.990 192.095 ;
        RECT 73.140 192.035 73.460 192.095 ;
        RECT 73.615 192.050 73.905 192.095 ;
        RECT 76.360 192.035 76.680 192.095 ;
        RECT 88.335 192.235 88.625 192.280 ;
        RECT 88.780 192.235 89.100 192.295 ;
        RECT 88.335 192.095 89.100 192.235 ;
        RECT 88.335 192.050 88.625 192.095 ;
        RECT 88.780 192.035 89.100 192.095 ;
        RECT 72.235 191.895 72.525 191.940 ;
        RECT 74.980 191.895 75.300 191.955 ;
        RECT 72.235 191.755 75.300 191.895 ;
        RECT 72.235 191.710 72.525 191.755 ;
        RECT 74.980 191.695 75.300 191.755 ;
        RECT 81.850 191.895 82.140 191.940 ;
        RECT 84.630 191.895 84.920 191.940 ;
        RECT 86.490 191.895 86.780 191.940 ;
        RECT 81.850 191.755 86.780 191.895 ;
        RECT 81.850 191.710 82.140 191.755 ;
        RECT 84.630 191.710 84.920 191.755 ;
        RECT 86.490 191.710 86.780 191.755 ;
        RECT 90.175 191.710 90.465 191.940 ;
        RECT 104.075 191.895 104.365 191.940 ;
        RECT 107.195 191.895 107.485 191.940 ;
        RECT 109.085 191.895 109.375 191.940 ;
        RECT 104.075 191.755 109.375 191.895 ;
        RECT 104.075 191.710 104.365 191.755 ;
        RECT 107.195 191.710 107.485 191.755 ;
        RECT 109.085 191.710 109.375 191.755 ;
        RECT 84.180 191.555 84.500 191.615 ;
        RECT 85.115 191.555 85.405 191.600 ;
        RECT 71.850 191.415 72.450 191.555 ;
        RECT 71.760 191.215 72.080 191.275 ;
        RECT 70.010 191.075 72.080 191.215 ;
        RECT 71.760 191.015 72.080 191.075 ;
        RECT 67.620 190.875 67.940 190.935 ;
        RECT 72.310 190.875 72.450 191.415 ;
        RECT 84.180 191.415 85.405 191.555 ;
        RECT 84.180 191.355 84.500 191.415 ;
        RECT 85.115 191.370 85.405 191.415 ;
        RECT 72.680 191.215 73.000 191.275 ;
        RECT 73.155 191.215 73.445 191.260 ;
        RECT 72.680 191.075 73.445 191.215 ;
        RECT 72.680 191.015 73.000 191.075 ;
        RECT 73.155 191.030 73.445 191.075 ;
        RECT 81.850 191.215 82.140 191.260 ;
        RECT 86.480 191.215 86.800 191.275 ;
        RECT 86.955 191.215 87.245 191.260 ;
        RECT 81.850 191.075 84.385 191.215 ;
        RECT 81.850 191.030 82.140 191.075 ;
        RECT 83.260 190.920 83.580 190.935 ;
        RECT 66.330 190.735 72.450 190.875 ;
        RECT 79.990 190.875 80.280 190.920 ;
        RECT 83.250 190.875 83.580 190.920 ;
        RECT 79.990 190.735 83.580 190.875 ;
        RECT 55.660 190.675 55.980 190.735 ;
        RECT 57.055 190.690 57.345 190.735 ;
        RECT 67.620 190.675 67.940 190.735 ;
        RECT 79.990 190.690 80.280 190.735 ;
        RECT 83.250 190.690 83.580 190.735 ;
        RECT 84.170 190.920 84.385 191.075 ;
        RECT 86.480 191.075 87.245 191.215 ;
        RECT 86.480 191.015 86.800 191.075 ;
        RECT 86.955 191.030 87.245 191.075 ;
        RECT 89.255 191.215 89.545 191.260 ;
        RECT 90.250 191.215 90.390 191.710 ;
        RECT 93.380 191.555 93.700 191.615 ;
        RECT 98.900 191.555 99.220 191.615 ;
        RECT 99.835 191.555 100.125 191.600 ;
        RECT 93.380 191.415 100.125 191.555 ;
        RECT 93.380 191.355 93.700 191.415 ;
        RECT 98.900 191.355 99.220 191.415 ;
        RECT 99.835 191.370 100.125 191.415 ;
        RECT 108.560 191.355 108.880 191.615 ;
        RECT 89.255 191.075 90.390 191.215 ;
        RECT 89.255 191.030 89.545 191.075 ;
        RECT 84.170 190.875 84.460 190.920 ;
        RECT 86.030 190.875 86.320 190.920 ;
        RECT 98.915 190.875 99.205 190.920 ;
        RECT 84.170 190.735 86.320 190.875 ;
        RECT 84.170 190.690 84.460 190.735 ;
        RECT 86.030 190.690 86.320 190.735 ;
        RECT 92.550 190.735 99.205 190.875 ;
        RECT 83.260 190.675 83.580 190.690 ;
        RECT 92.550 190.595 92.690 190.735 ;
        RECT 98.915 190.690 99.205 190.735 ;
        RECT 99.375 190.875 99.665 190.920 ;
        RECT 100.280 190.875 100.600 190.935 ;
        RECT 102.995 190.920 103.285 191.235 ;
        RECT 104.075 191.215 104.365 191.260 ;
        RECT 107.655 191.215 107.945 191.260 ;
        RECT 109.490 191.215 109.780 191.260 ;
        RECT 104.075 191.075 109.780 191.215 ;
        RECT 104.075 191.030 104.365 191.075 ;
        RECT 107.655 191.030 107.945 191.075 ;
        RECT 109.490 191.030 109.780 191.075 ;
        RECT 109.940 191.015 110.260 191.275 ;
        RECT 99.375 190.735 100.600 190.875 ;
        RECT 99.375 190.690 99.665 190.735 ;
        RECT 100.280 190.675 100.600 190.735 ;
        RECT 102.695 190.875 103.285 190.920 ;
        RECT 105.935 190.875 106.585 190.920 ;
        RECT 107.180 190.875 107.500 190.935 ;
        RECT 102.695 190.735 107.500 190.875 ;
        RECT 102.695 190.690 102.985 190.735 ;
        RECT 105.935 190.690 106.585 190.735 ;
        RECT 107.180 190.675 107.500 190.735 ;
        RECT 35.435 190.535 35.725 190.580 ;
        RECT 34.040 190.395 35.725 190.535 ;
        RECT 34.040 190.335 34.360 190.395 ;
        RECT 35.435 190.350 35.725 190.395 ;
        RECT 37.735 190.350 38.025 190.580 ;
        RECT 39.100 190.535 39.420 190.595 ;
        RECT 39.575 190.535 39.865 190.580 ;
        RECT 39.100 190.395 39.865 190.535 ;
        RECT 39.100 190.335 39.420 190.395 ;
        RECT 39.575 190.350 39.865 190.395 ;
        RECT 40.495 190.535 40.785 190.580 ;
        RECT 42.780 190.535 43.100 190.595 ;
        RECT 40.495 190.395 43.100 190.535 ;
        RECT 40.495 190.350 40.785 190.395 ;
        RECT 42.780 190.335 43.100 190.395 ;
        RECT 59.340 190.335 59.660 190.595 ;
        RECT 63.480 190.335 63.800 190.595 ;
        RECT 77.280 190.535 77.600 190.595 ;
        RECT 77.985 190.535 78.275 190.580 ;
        RECT 92.015 190.535 92.305 190.580 ;
        RECT 77.280 190.395 92.305 190.535 ;
        RECT 77.280 190.335 77.600 190.395 ;
        RECT 77.985 190.350 78.275 190.395 ;
        RECT 92.015 190.350 92.305 190.395 ;
        RECT 92.460 190.335 92.780 190.595 ;
        RECT 97.060 190.335 97.380 190.595 ;
        RECT 101.215 190.535 101.505 190.580 ;
        RECT 101.660 190.535 101.980 190.595 ;
        RECT 101.215 190.395 101.980 190.535 ;
        RECT 101.215 190.350 101.505 190.395 ;
        RECT 101.660 190.335 101.980 190.395 ;
        RECT 14.650 189.715 115.850 190.195 ;
        RECT 32.750 189.375 42.550 189.515 ;
        RECT 31.295 189.175 31.585 189.220 ;
        RECT 32.750 189.175 32.890 189.375 ;
        RECT 31.295 189.035 32.890 189.175 ;
        RECT 33.120 189.175 33.440 189.235 ;
        RECT 33.990 189.175 34.280 189.220 ;
        RECT 37.250 189.175 37.540 189.220 ;
        RECT 33.120 189.035 37.540 189.175 ;
        RECT 31.295 188.990 31.585 189.035 ;
        RECT 33.120 188.975 33.440 189.035 ;
        RECT 33.990 188.990 34.280 189.035 ;
        RECT 37.250 188.990 37.540 189.035 ;
        RECT 38.170 189.175 38.460 189.220 ;
        RECT 40.030 189.175 40.320 189.220 ;
        RECT 38.170 189.035 40.320 189.175 ;
        RECT 38.170 188.990 38.460 189.035 ;
        RECT 40.030 188.990 40.320 189.035 ;
        RECT 27.600 188.635 27.920 188.895 ;
        RECT 35.850 188.835 36.140 188.880 ;
        RECT 38.170 188.835 38.385 188.990 ;
        RECT 35.850 188.695 38.385 188.835 ;
        RECT 35.850 188.650 36.140 188.695 ;
        RECT 39.100 188.635 39.420 188.895 ;
        RECT 39.560 188.835 39.880 188.895 ;
        RECT 42.410 188.880 42.550 189.375 ;
        RECT 46.460 189.315 46.780 189.575 ;
        RECT 51.520 189.515 51.840 189.575 ;
        RECT 53.375 189.515 53.665 189.560 ;
        RECT 51.520 189.375 53.665 189.515 ;
        RECT 51.520 189.315 51.840 189.375 ;
        RECT 53.375 189.330 53.665 189.375 ;
        RECT 55.660 189.315 55.980 189.575 ;
        RECT 67.635 189.515 67.925 189.560 ;
        RECT 65.870 189.375 67.925 189.515 ;
        RECT 44.160 189.175 44.480 189.235 ;
        RECT 48.775 189.175 49.065 189.220 ;
        RECT 44.160 189.035 49.065 189.175 ;
        RECT 44.160 188.975 44.480 189.035 ;
        RECT 48.775 188.990 49.065 189.035 ;
        RECT 59.340 189.175 59.660 189.235 ;
        RECT 65.870 189.220 66.010 189.375 ;
        RECT 67.635 189.330 67.925 189.375 ;
        RECT 77.280 189.515 77.600 189.575 ;
        RECT 80.055 189.515 80.345 189.560 ;
        RECT 77.280 189.375 80.345 189.515 ;
        RECT 77.280 189.315 77.600 189.375 ;
        RECT 80.055 189.330 80.345 189.375 ;
        RECT 82.340 189.315 82.660 189.575 ;
        RECT 83.260 189.315 83.580 189.575 ;
        RECT 90.635 189.515 90.925 189.560 ;
        RECT 92.460 189.515 92.780 189.575 ;
        RECT 90.635 189.375 92.780 189.515 ;
        RECT 90.635 189.330 90.925 189.375 ;
        RECT 92.460 189.315 92.780 189.375 ;
        RECT 95.695 189.515 95.985 189.560 ;
        RECT 99.820 189.515 100.140 189.575 ;
        RECT 95.695 189.375 100.140 189.515 ;
        RECT 95.695 189.330 95.985 189.375 ;
        RECT 99.820 189.315 100.140 189.375 ;
        RECT 59.915 189.175 60.205 189.220 ;
        RECT 63.155 189.175 63.805 189.220 ;
        RECT 59.340 189.035 63.805 189.175 ;
        RECT 59.340 188.975 59.660 189.035 ;
        RECT 59.915 188.990 60.505 189.035 ;
        RECT 63.155 188.990 63.805 189.035 ;
        RECT 65.795 188.990 66.085 189.220 ;
        RECT 75.440 189.175 75.760 189.235 ;
        RECT 80.515 189.175 80.805 189.220 ;
        RECT 75.440 189.035 80.805 189.175 ;
        RECT 39.560 188.695 42.090 188.835 ;
        RECT 39.560 188.635 39.880 188.695 ;
        RECT 28.535 188.495 28.825 188.540 ;
        RECT 38.180 188.495 38.500 188.555 ;
        RECT 28.535 188.355 38.500 188.495 ;
        RECT 28.535 188.310 28.825 188.355 ;
        RECT 38.180 188.295 38.500 188.355 ;
        RECT 40.955 188.310 41.245 188.540 ;
        RECT 41.950 188.495 42.090 188.695 ;
        RECT 42.335 188.650 42.625 188.880 ;
        RECT 44.635 188.835 44.925 188.880 ;
        RECT 42.870 188.695 44.925 188.835 ;
        RECT 42.870 188.495 43.010 188.695 ;
        RECT 44.635 188.650 44.925 188.695 ;
        RECT 53.820 188.635 54.140 188.895 ;
        RECT 54.755 188.650 55.045 188.880 ;
        RECT 60.215 188.675 60.505 188.990 ;
        RECT 75.440 188.975 75.760 189.035 ;
        RECT 80.515 188.990 80.805 189.035 ;
        RECT 61.295 188.835 61.585 188.880 ;
        RECT 64.875 188.835 65.165 188.880 ;
        RECT 66.710 188.835 67.000 188.880 ;
        RECT 61.295 188.695 67.000 188.835 ;
        RECT 61.295 188.650 61.585 188.695 ;
        RECT 64.875 188.650 65.165 188.695 ;
        RECT 66.710 188.650 67.000 188.695 ;
        RECT 67.175 188.835 67.465 188.880 ;
        RECT 68.080 188.835 68.400 188.895 ;
        RECT 67.175 188.695 68.400 188.835 ;
        RECT 67.175 188.650 67.465 188.695 ;
        RECT 41.950 188.355 43.010 188.495 ;
        RECT 43.715 188.495 44.005 188.540 ;
        RECT 47.380 188.495 47.700 188.555 ;
        RECT 43.715 188.355 47.700 188.495 ;
        RECT 43.715 188.310 44.005 188.355 ;
        RECT 35.850 188.155 36.140 188.200 ;
        RECT 38.630 188.155 38.920 188.200 ;
        RECT 40.490 188.155 40.780 188.200 ;
        RECT 35.850 188.015 40.780 188.155 ;
        RECT 41.030 188.155 41.170 188.310 ;
        RECT 47.380 188.295 47.700 188.355 ;
        RECT 48.315 188.495 48.605 188.540 ;
        RECT 48.760 188.495 49.080 188.555 ;
        RECT 54.830 188.495 54.970 188.650 ;
        RECT 68.080 188.635 68.400 188.695 ;
        RECT 69.475 188.650 69.765 188.880 ;
        RECT 78.200 188.835 78.520 188.895 ;
        RECT 83.735 188.835 84.025 188.880 ;
        RECT 85.100 188.835 85.420 188.895 ;
        RECT 89.255 188.835 89.545 188.880 ;
        RECT 78.200 188.695 89.545 188.835 ;
        RECT 48.315 188.355 49.080 188.495 ;
        RECT 48.315 188.310 48.605 188.355 ;
        RECT 48.760 188.295 49.080 188.355 ;
        RECT 50.690 188.355 54.970 188.495 ;
        RECT 63.480 188.495 63.800 188.555 ;
        RECT 69.550 188.495 69.690 188.650 ;
        RECT 78.200 188.635 78.520 188.695 ;
        RECT 83.735 188.650 84.025 188.695 ;
        RECT 85.100 188.635 85.420 188.695 ;
        RECT 89.255 188.650 89.545 188.695 ;
        RECT 94.775 188.835 95.065 188.880 ;
        RECT 97.060 188.835 97.380 188.895 ;
        RECT 94.775 188.695 97.380 188.835 ;
        RECT 94.775 188.650 95.065 188.695 ;
        RECT 97.060 188.635 97.380 188.695 ;
        RECT 99.835 188.835 100.125 188.880 ;
        RECT 100.740 188.835 101.060 188.895 ;
        RECT 101.215 188.835 101.505 188.880 ;
        RECT 99.835 188.695 101.505 188.835 ;
        RECT 99.835 188.650 100.125 188.695 ;
        RECT 100.740 188.635 101.060 188.695 ;
        RECT 101.215 188.650 101.505 188.695 ;
        RECT 63.480 188.355 69.690 188.495 ;
        RECT 42.320 188.155 42.640 188.215 ;
        RECT 50.690 188.200 50.830 188.355 ;
        RECT 63.480 188.295 63.800 188.355 ;
        RECT 69.920 188.295 70.240 188.555 ;
        RECT 78.660 188.495 78.980 188.555 ;
        RECT 79.135 188.495 79.425 188.540 ;
        RECT 78.660 188.355 79.425 188.495 ;
        RECT 78.660 188.295 78.980 188.355 ;
        RECT 79.135 188.310 79.425 188.355 ;
        RECT 93.840 188.295 94.160 188.555 ;
        RECT 98.900 188.295 99.220 188.555 ;
        RECT 101.660 188.495 101.980 188.555 ;
        RECT 106.275 188.495 106.565 188.540 ;
        RECT 107.180 188.495 107.500 188.555 ;
        RECT 101.660 188.355 107.500 188.495 ;
        RECT 101.660 188.295 101.980 188.355 ;
        RECT 106.275 188.310 106.565 188.355 ;
        RECT 107.180 188.295 107.500 188.355 ;
        RECT 41.030 188.015 42.640 188.155 ;
        RECT 35.850 187.970 36.140 188.015 ;
        RECT 38.630 187.970 38.920 188.015 ;
        RECT 40.490 187.970 40.780 188.015 ;
        RECT 42.320 187.955 42.640 188.015 ;
        RECT 50.615 187.970 50.905 188.200 ;
        RECT 61.295 188.155 61.585 188.200 ;
        RECT 64.415 188.155 64.705 188.200 ;
        RECT 66.305 188.155 66.595 188.200 ;
        RECT 61.295 188.015 66.595 188.155 ;
        RECT 61.295 187.970 61.585 188.015 ;
        RECT 64.415 187.970 64.705 188.015 ;
        RECT 66.305 187.970 66.595 188.015 ;
        RECT 25.760 187.815 26.080 187.875 ;
        RECT 26.695 187.815 26.985 187.860 ;
        RECT 25.760 187.675 26.985 187.815 ;
        RECT 25.760 187.615 26.080 187.675 ;
        RECT 26.695 187.630 26.985 187.675 ;
        RECT 31.985 187.815 32.275 187.860 ;
        RECT 34.040 187.815 34.360 187.875 ;
        RECT 39.560 187.815 39.880 187.875 ;
        RECT 31.985 187.675 39.880 187.815 ;
        RECT 31.985 187.630 32.275 187.675 ;
        RECT 34.040 187.615 34.360 187.675 ;
        RECT 39.560 187.615 39.880 187.675 ;
        RECT 40.940 187.815 41.260 187.875 ;
        RECT 41.415 187.815 41.705 187.860 ;
        RECT 40.940 187.675 41.705 187.815 ;
        RECT 40.940 187.615 41.260 187.675 ;
        RECT 41.415 187.630 41.705 187.675 ;
        RECT 58.435 187.815 58.725 187.860 ;
        RECT 60.720 187.815 61.040 187.875 ;
        RECT 62.560 187.815 62.880 187.875 ;
        RECT 58.435 187.675 62.880 187.815 ;
        RECT 58.435 187.630 58.725 187.675 ;
        RECT 60.720 187.615 61.040 187.675 ;
        RECT 62.560 187.615 62.880 187.675 ;
        RECT 77.740 187.615 78.060 187.875 ;
        RECT 89.700 187.615 90.020 187.875 ;
        RECT 96.155 187.815 96.445 187.860 ;
        RECT 97.060 187.815 97.380 187.875 ;
        RECT 96.155 187.675 97.380 187.815 ;
        RECT 96.155 187.630 96.445 187.675 ;
        RECT 97.060 187.615 97.380 187.675 ;
        RECT 100.295 187.815 100.585 187.860 ;
        RECT 100.740 187.815 101.060 187.875 ;
        RECT 100.295 187.675 101.060 187.815 ;
        RECT 100.295 187.630 100.585 187.675 ;
        RECT 100.740 187.615 101.060 187.675 ;
        RECT 101.660 187.615 101.980 187.875 ;
        RECT 103.055 187.815 103.345 187.860 ;
        RECT 103.960 187.815 104.280 187.875 ;
        RECT 103.055 187.675 104.280 187.815 ;
        RECT 103.055 187.630 103.345 187.675 ;
        RECT 103.960 187.615 104.280 187.675 ;
        RECT 14.650 186.995 115.850 187.475 ;
        RECT 23.935 186.795 24.225 186.840 ;
        RECT 27.600 186.795 27.920 186.855 ;
        RECT 23.935 186.655 27.920 186.795 ;
        RECT 23.935 186.610 24.225 186.655 ;
        RECT 27.600 186.595 27.920 186.655 ;
        RECT 38.180 186.795 38.500 186.855 ;
        RECT 39.115 186.795 39.405 186.840 ;
        RECT 38.180 186.655 39.405 186.795 ;
        RECT 38.180 186.595 38.500 186.655 ;
        RECT 39.115 186.610 39.405 186.655 ;
        RECT 25.265 186.455 25.555 186.500 ;
        RECT 27.155 186.455 27.445 186.500 ;
        RECT 30.275 186.455 30.565 186.500 ;
        RECT 25.265 186.315 30.565 186.455 ;
        RECT 25.265 186.270 25.555 186.315 ;
        RECT 27.155 186.270 27.445 186.315 ;
        RECT 30.275 186.270 30.565 186.315 ;
        RECT 30.820 186.455 31.140 186.515 ;
        RECT 33.135 186.455 33.425 186.500 ;
        RECT 33.580 186.455 33.900 186.515 ;
        RECT 30.820 186.315 33.900 186.455 ;
        RECT 30.820 186.255 31.140 186.315 ;
        RECT 33.135 186.270 33.425 186.315 ;
        RECT 33.580 186.255 33.900 186.315 ;
        RECT 34.500 186.455 34.820 186.515 ;
        RECT 43.240 186.455 43.560 186.515 ;
        RECT 34.500 186.315 43.560 186.455 ;
        RECT 34.500 186.255 34.820 186.315 ;
        RECT 43.240 186.255 43.560 186.315 ;
        RECT 46.115 186.455 46.405 186.500 ;
        RECT 49.235 186.455 49.525 186.500 ;
        RECT 51.125 186.455 51.415 186.500 ;
        RECT 46.115 186.315 51.415 186.455 ;
        RECT 46.115 186.270 46.405 186.315 ;
        RECT 49.235 186.270 49.525 186.315 ;
        RECT 51.125 186.270 51.415 186.315 ;
        RECT 79.550 186.455 79.840 186.500 ;
        RECT 82.330 186.455 82.620 186.500 ;
        RECT 84.190 186.455 84.480 186.500 ;
        RECT 79.550 186.315 84.480 186.455 ;
        RECT 79.550 186.270 79.840 186.315 ;
        RECT 82.330 186.270 82.620 186.315 ;
        RECT 84.190 186.270 84.480 186.315 ;
        RECT 85.100 186.455 85.420 186.515 ;
        RECT 93.035 186.455 93.325 186.500 ;
        RECT 96.155 186.455 96.445 186.500 ;
        RECT 98.045 186.455 98.335 186.500 ;
        RECT 85.100 186.315 87.170 186.455 ;
        RECT 85.100 186.255 85.420 186.315 ;
        RECT 25.760 185.915 26.080 186.175 ;
        RECT 26.220 186.115 26.540 186.175 ;
        RECT 42.335 186.115 42.625 186.160 ;
        RECT 47.380 186.115 47.700 186.175 ;
        RECT 26.220 185.975 41.170 186.115 ;
        RECT 26.220 185.915 26.540 185.975 ;
        RECT 19.335 185.590 19.625 185.820 ;
        RECT 21.175 185.775 21.465 185.820 ;
        RECT 21.620 185.775 21.940 185.835 ;
        RECT 21.175 185.635 21.940 185.775 ;
        RECT 21.175 185.590 21.465 185.635 ;
        RECT 19.410 185.095 19.550 185.590 ;
        RECT 21.620 185.575 21.940 185.635 ;
        RECT 24.380 185.575 24.700 185.835 ;
        RECT 24.860 185.775 25.150 185.820 ;
        RECT 26.695 185.775 26.985 185.820 ;
        RECT 30.275 185.775 30.565 185.820 ;
        RECT 24.860 185.635 30.565 185.775 ;
        RECT 24.860 185.590 25.150 185.635 ;
        RECT 26.695 185.590 26.985 185.635 ;
        RECT 30.275 185.590 30.565 185.635 ;
        RECT 31.355 185.480 31.645 185.795 ;
        RECT 34.500 185.575 34.820 185.835 ;
        RECT 35.435 185.590 35.725 185.820 ;
        RECT 19.795 185.435 20.085 185.480 ;
        RECT 28.055 185.435 28.705 185.480 ;
        RECT 31.355 185.435 31.945 185.480 ;
        RECT 19.795 185.295 31.945 185.435 ;
        RECT 19.795 185.250 20.085 185.295 ;
        RECT 28.055 185.250 28.705 185.295 ;
        RECT 31.655 185.250 31.945 185.295 ;
        RECT 33.120 185.435 33.440 185.495 ;
        RECT 35.510 185.435 35.650 185.590 ;
        RECT 35.880 185.575 36.200 185.835 ;
        RECT 36.340 185.575 36.660 185.835 ;
        RECT 41.030 185.820 41.170 185.975 ;
        RECT 42.335 185.975 47.700 186.115 ;
        RECT 42.335 185.930 42.625 185.975 ;
        RECT 47.380 185.915 47.700 185.975 ;
        RECT 84.655 186.115 84.945 186.160 ;
        RECT 86.480 186.115 86.800 186.175 ;
        RECT 84.655 185.975 86.800 186.115 ;
        RECT 84.655 185.930 84.945 185.975 ;
        RECT 86.480 185.915 86.800 185.975 ;
        RECT 40.955 185.590 41.245 185.820 ;
        RECT 41.415 185.435 41.705 185.480 ;
        RECT 33.120 185.295 41.705 185.435 ;
        RECT 33.120 185.235 33.440 185.295 ;
        RECT 41.415 185.250 41.705 185.295 ;
        RECT 43.700 185.435 44.020 185.495 ;
        RECT 45.035 185.480 45.325 185.795 ;
        RECT 46.115 185.775 46.405 185.820 ;
        RECT 49.695 185.775 49.985 185.820 ;
        RECT 51.530 185.775 51.820 185.820 ;
        RECT 46.115 185.635 51.820 185.775 ;
        RECT 46.115 185.590 46.405 185.635 ;
        RECT 49.695 185.590 49.985 185.635 ;
        RECT 51.530 185.590 51.820 185.635 ;
        RECT 51.980 185.575 52.300 185.835 ;
        RECT 79.550 185.775 79.840 185.820 ;
        RECT 82.815 185.775 83.105 185.820 ;
        RECT 79.550 185.635 82.085 185.775 ;
        RECT 79.550 185.590 79.840 185.635 ;
        RECT 77.740 185.480 78.060 185.495 ;
        RECT 81.870 185.480 82.085 185.635 ;
        RECT 82.815 185.635 84.410 185.775 ;
        RECT 82.815 185.590 83.105 185.635 ;
        RECT 44.735 185.435 45.325 185.480 ;
        RECT 47.975 185.435 48.625 185.480 ;
        RECT 43.700 185.295 48.625 185.435 ;
        RECT 43.700 185.235 44.020 185.295 ;
        RECT 44.735 185.250 45.025 185.295 ;
        RECT 47.975 185.250 48.625 185.295 ;
        RECT 50.615 185.250 50.905 185.480 ;
        RECT 77.690 185.435 78.060 185.480 ;
        RECT 80.950 185.435 81.240 185.480 ;
        RECT 77.690 185.295 81.240 185.435 ;
        RECT 77.690 185.250 78.060 185.295 ;
        RECT 80.950 185.250 81.240 185.295 ;
        RECT 81.870 185.435 82.160 185.480 ;
        RECT 83.730 185.435 84.020 185.480 ;
        RECT 81.870 185.295 84.020 185.435 ;
        RECT 81.870 185.250 82.160 185.295 ;
        RECT 83.730 185.250 84.020 185.295 ;
        RECT 23.920 185.095 24.240 185.155 ;
        RECT 19.410 184.955 24.240 185.095 ;
        RECT 23.920 184.895 24.240 184.955 ;
        RECT 24.840 185.095 25.160 185.155 ;
        RECT 30.820 185.095 31.140 185.155 ;
        RECT 24.840 184.955 31.140 185.095 ;
        RECT 24.840 184.895 25.160 184.955 ;
        RECT 30.820 184.895 31.140 184.955 ;
        RECT 32.200 185.095 32.520 185.155 ;
        RECT 36.340 185.095 36.660 185.155 ;
        RECT 32.200 184.955 36.660 185.095 ;
        RECT 32.200 184.895 32.520 184.955 ;
        RECT 36.340 184.895 36.660 184.955 ;
        RECT 37.735 185.095 38.025 185.140 ;
        RECT 38.180 185.095 38.500 185.155 ;
        RECT 37.735 184.955 38.500 185.095 ;
        RECT 37.735 184.910 38.025 184.955 ;
        RECT 38.180 184.895 38.500 184.955 ;
        RECT 43.255 185.095 43.545 185.140 ;
        RECT 44.160 185.095 44.480 185.155 ;
        RECT 43.255 184.955 44.480 185.095 ;
        RECT 43.255 184.910 43.545 184.955 ;
        RECT 44.160 184.895 44.480 184.955 ;
        RECT 45.540 185.095 45.860 185.155 ;
        RECT 50.690 185.095 50.830 185.250 ;
        RECT 77.740 185.235 78.060 185.250 ;
        RECT 45.540 184.955 50.830 185.095 ;
        RECT 75.440 185.140 75.760 185.155 ;
        RECT 45.540 184.895 45.860 184.955 ;
        RECT 75.440 184.910 75.975 185.140 ;
        RECT 84.270 185.095 84.410 185.635 ;
        RECT 86.020 185.575 86.340 185.835 ;
        RECT 87.030 185.775 87.170 186.315 ;
        RECT 93.035 186.315 98.335 186.455 ;
        RECT 93.035 186.270 93.325 186.315 ;
        RECT 96.155 186.270 96.445 186.315 ;
        RECT 98.045 186.270 98.335 186.315 ;
        RECT 106.835 186.455 107.125 186.500 ;
        RECT 109.955 186.455 110.245 186.500 ;
        RECT 111.845 186.455 112.135 186.500 ;
        RECT 106.835 186.315 112.135 186.455 ;
        RECT 106.835 186.270 107.125 186.315 ;
        RECT 109.955 186.270 110.245 186.315 ;
        RECT 111.845 186.270 112.135 186.315 ;
        RECT 87.400 186.115 87.720 186.175 ;
        RECT 90.175 186.115 90.465 186.160 ;
        RECT 87.400 185.975 90.465 186.115 ;
        RECT 87.400 185.915 87.720 185.975 ;
        RECT 90.175 185.930 90.465 185.975 ;
        RECT 102.595 186.115 102.885 186.160 ;
        RECT 103.500 186.115 103.820 186.175 ;
        RECT 103.975 186.115 104.265 186.160 ;
        RECT 102.595 185.975 104.265 186.115 ;
        RECT 102.595 185.930 102.885 185.975 ;
        RECT 103.500 185.915 103.820 185.975 ;
        RECT 103.975 185.930 104.265 185.975 ;
        RECT 87.875 185.775 88.165 185.820 ;
        RECT 87.030 185.635 88.165 185.775 ;
        RECT 87.875 185.590 88.165 185.635 ;
        RECT 89.700 185.435 90.020 185.495 ;
        RECT 91.955 185.480 92.245 185.795 ;
        RECT 93.035 185.775 93.325 185.820 ;
        RECT 96.615 185.775 96.905 185.820 ;
        RECT 98.450 185.775 98.740 185.820 ;
        RECT 93.035 185.635 98.740 185.775 ;
        RECT 93.035 185.590 93.325 185.635 ;
        RECT 96.615 185.590 96.905 185.635 ;
        RECT 98.450 185.590 98.740 185.635 ;
        RECT 98.915 185.590 99.205 185.820 ;
        RECT 91.655 185.435 92.245 185.480 ;
        RECT 94.895 185.435 95.545 185.480 ;
        RECT 89.700 185.295 95.545 185.435 ;
        RECT 89.700 185.235 90.020 185.295 ;
        RECT 91.655 185.250 91.945 185.295 ;
        RECT 94.895 185.250 95.545 185.295 ;
        RECT 97.520 185.235 97.840 185.495 ;
        RECT 85.115 185.095 85.405 185.140 ;
        RECT 84.270 184.955 85.405 185.095 ;
        RECT 85.115 184.910 85.405 184.955 ;
        RECT 88.335 185.095 88.625 185.140 ;
        RECT 88.780 185.095 89.100 185.155 ;
        RECT 88.335 184.955 89.100 185.095 ;
        RECT 98.990 185.095 99.130 185.590 ;
        RECT 99.375 185.435 99.665 185.480 ;
        RECT 100.280 185.435 100.600 185.495 ;
        RECT 99.375 185.295 100.600 185.435 ;
        RECT 99.375 185.250 99.665 185.295 ;
        RECT 100.280 185.235 100.600 185.295 ;
        RECT 101.660 185.435 101.980 185.495 ;
        RECT 105.755 185.480 106.045 185.795 ;
        RECT 106.835 185.775 107.125 185.820 ;
        RECT 110.415 185.775 110.705 185.820 ;
        RECT 112.250 185.775 112.540 185.820 ;
        RECT 106.835 185.635 112.540 185.775 ;
        RECT 106.835 185.590 107.125 185.635 ;
        RECT 110.415 185.590 110.705 185.635 ;
        RECT 112.250 185.590 112.540 185.635 ;
        RECT 112.715 185.590 113.005 185.820 ;
        RECT 105.455 185.435 106.045 185.480 ;
        RECT 108.695 185.435 109.345 185.480 ;
        RECT 101.660 185.295 109.345 185.435 ;
        RECT 101.660 185.235 101.980 185.295 ;
        RECT 105.455 185.250 105.745 185.295 ;
        RECT 108.695 185.250 109.345 185.295 ;
        RECT 111.320 185.235 111.640 185.495 ;
        RECT 109.480 185.095 109.800 185.155 ;
        RECT 111.780 185.095 112.100 185.155 ;
        RECT 112.790 185.095 112.930 185.590 ;
        RECT 98.990 184.955 112.930 185.095 ;
        RECT 88.335 184.910 88.625 184.955 ;
        RECT 75.440 184.895 75.760 184.910 ;
        RECT 88.780 184.895 89.100 184.955 ;
        RECT 109.480 184.895 109.800 184.955 ;
        RECT 111.780 184.895 112.100 184.955 ;
        RECT 14.650 184.275 115.850 184.755 ;
        RECT 21.620 184.075 21.940 184.135 ;
        RECT 28.535 184.075 28.825 184.120 ;
        RECT 21.620 183.935 28.825 184.075 ;
        RECT 21.620 183.875 21.940 183.935 ;
        RECT 28.535 183.890 28.825 183.935 ;
        RECT 30.835 184.075 31.125 184.120 ;
        RECT 33.580 184.075 33.900 184.135 ;
        RECT 30.835 183.935 33.900 184.075 ;
        RECT 30.835 183.890 31.125 183.935 ;
        RECT 33.580 183.875 33.900 183.935 ;
        RECT 43.700 183.875 44.020 184.135 ;
        RECT 45.540 183.875 45.860 184.135 ;
        RECT 48.760 184.075 49.080 184.135 ;
        RECT 49.235 184.075 49.525 184.120 ;
        RECT 48.760 183.935 49.525 184.075 ;
        RECT 48.760 183.875 49.080 183.935 ;
        RECT 49.235 183.890 49.525 183.935 ;
        RECT 76.375 184.075 76.665 184.120 ;
        RECT 86.020 184.075 86.340 184.135 ;
        RECT 76.375 183.935 86.340 184.075 ;
        RECT 76.375 183.890 76.665 183.935 ;
        RECT 86.020 183.875 86.340 183.935 ;
        RECT 96.155 184.075 96.445 184.120 ;
        RECT 97.060 184.075 97.380 184.135 ;
        RECT 99.835 184.075 100.125 184.120 ;
        RECT 96.155 183.935 100.125 184.075 ;
        RECT 96.155 183.890 96.445 183.935 ;
        RECT 97.060 183.875 97.380 183.935 ;
        RECT 99.835 183.890 100.125 183.935 ;
        RECT 100.280 183.875 100.600 184.135 ;
        RECT 21.175 183.735 21.465 183.780 ;
        RECT 30.375 183.735 30.665 183.780 ;
        RECT 21.175 183.595 30.665 183.735 ;
        RECT 21.175 183.550 21.465 183.595 ;
        RECT 30.375 183.550 30.665 183.595 ;
        RECT 34.500 183.735 34.820 183.795 ;
        RECT 35.075 183.735 35.365 183.780 ;
        RECT 38.315 183.735 38.965 183.780 ;
        RECT 34.500 183.595 38.965 183.735 ;
        RECT 34.500 183.535 34.820 183.595 ;
        RECT 35.075 183.550 35.665 183.595 ;
        RECT 38.315 183.550 38.965 183.595 ;
        RECT 22.095 183.395 22.385 183.440 ;
        RECT 24.855 183.395 25.145 183.440 ;
        RECT 25.760 183.395 26.080 183.455 ;
        RECT 22.095 183.255 24.150 183.395 ;
        RECT 22.095 183.210 22.385 183.255 ;
        RECT 18.415 183.055 18.705 183.100 ;
        RECT 22.540 183.055 22.860 183.115 ;
        RECT 18.415 182.915 22.860 183.055 ;
        RECT 18.415 182.870 18.705 182.915 ;
        RECT 22.540 182.855 22.860 182.915 ;
        RECT 24.010 182.715 24.150 183.255 ;
        RECT 24.855 183.255 26.080 183.395 ;
        RECT 24.855 183.210 25.145 183.255 ;
        RECT 25.760 183.195 26.080 183.255 ;
        RECT 26.680 183.195 27.000 183.455 ;
        RECT 35.375 183.235 35.665 183.550 ;
        RECT 40.940 183.535 41.260 183.795 ;
        RECT 51.535 183.735 51.825 183.780 ;
        RECT 68.540 183.735 68.860 183.795 ;
        RECT 71.300 183.735 71.620 183.795 ;
        RECT 88.780 183.780 89.100 183.795 ;
        RECT 88.775 183.735 89.425 183.780 ;
        RECT 92.375 183.735 92.665 183.780 ;
        RECT 45.630 183.595 51.825 183.735 ;
        RECT 36.455 183.395 36.745 183.440 ;
        RECT 40.035 183.395 40.325 183.440 ;
        RECT 41.870 183.395 42.160 183.440 ;
        RECT 36.455 183.255 42.160 183.395 ;
        RECT 36.455 183.210 36.745 183.255 ;
        RECT 40.035 183.210 40.325 183.255 ;
        RECT 41.870 183.210 42.160 183.255 ;
        RECT 42.320 183.195 42.640 183.455 ;
        RECT 44.175 183.395 44.465 183.440 ;
        RECT 43.330 183.255 44.465 183.395 ;
        RECT 24.380 183.055 24.700 183.115 ;
        RECT 26.235 183.055 26.525 183.100 ;
        RECT 24.380 182.915 26.525 183.055 ;
        RECT 24.380 182.855 24.700 182.915 ;
        RECT 26.235 182.870 26.525 182.915 ;
        RECT 31.740 182.855 32.060 183.115 ;
        RECT 37.260 183.055 37.580 183.115 ;
        RECT 42.410 183.055 42.550 183.195 ;
        RECT 32.290 182.915 42.550 183.055 ;
        RECT 30.820 182.715 31.140 182.775 ;
        RECT 32.290 182.715 32.430 182.915 ;
        RECT 37.260 182.855 37.580 182.915 ;
        RECT 36.455 182.715 36.745 182.760 ;
        RECT 39.575 182.715 39.865 182.760 ;
        RECT 41.465 182.715 41.755 182.760 ;
        RECT 24.010 182.575 30.590 182.715 ;
        RECT 23.920 182.375 24.240 182.435 ;
        RECT 26.680 182.375 27.000 182.435 ;
        RECT 23.920 182.235 27.000 182.375 ;
        RECT 30.450 182.375 30.590 182.575 ;
        RECT 30.820 182.575 32.430 182.715 ;
        RECT 32.750 182.575 36.110 182.715 ;
        RECT 30.820 182.515 31.140 182.575 ;
        RECT 32.750 182.375 32.890 182.575 ;
        RECT 30.450 182.235 32.890 182.375 ;
        RECT 33.120 182.375 33.440 182.435 ;
        RECT 33.595 182.375 33.885 182.420 ;
        RECT 33.120 182.235 33.885 182.375 ;
        RECT 35.970 182.375 36.110 182.575 ;
        RECT 36.455 182.575 41.755 182.715 ;
        RECT 43.330 182.715 43.470 183.255 ;
        RECT 44.175 183.210 44.465 183.255 ;
        RECT 44.635 183.385 44.925 183.440 ;
        RECT 45.630 183.395 45.770 183.595 ;
        RECT 51.535 183.550 51.825 183.595 ;
        RECT 67.250 183.595 71.620 183.735 ;
        RECT 49.695 183.395 49.985 183.440 ;
        RECT 53.820 183.395 54.140 183.455 ;
        RECT 56.120 183.395 56.440 183.455 ;
        RECT 67.250 183.440 67.390 183.595 ;
        RECT 68.540 183.535 68.860 183.595 ;
        RECT 71.300 183.535 71.620 183.595 ;
        RECT 74.610 183.595 78.890 183.735 ;
        RECT 45.170 183.385 45.770 183.395 ;
        RECT 44.635 183.255 45.770 183.385 ;
        RECT 46.550 183.255 56.440 183.395 ;
        RECT 44.635 183.245 45.310 183.255 ;
        RECT 44.635 183.210 44.925 183.245 ;
        RECT 43.700 183.055 44.020 183.115 ;
        RECT 46.000 183.055 46.320 183.115 ;
        RECT 43.700 182.915 46.320 183.055 ;
        RECT 43.700 182.855 44.020 182.915 ;
        RECT 46.000 182.855 46.320 182.915 ;
        RECT 46.550 182.715 46.690 183.255 ;
        RECT 49.695 183.210 49.985 183.255 ;
        RECT 53.820 183.195 54.140 183.255 ;
        RECT 56.120 183.195 56.440 183.255 ;
        RECT 67.175 183.210 67.465 183.440 ;
        RECT 67.620 183.195 67.940 183.455 ;
        RECT 68.080 183.195 68.400 183.455 ;
        RECT 73.140 183.395 73.460 183.455 ;
        RECT 74.610 183.440 74.750 183.595 ;
        RECT 74.535 183.395 74.825 183.440 ;
        RECT 73.140 183.255 74.825 183.395 ;
        RECT 73.140 183.195 73.460 183.255 ;
        RECT 74.535 183.210 74.825 183.255 ;
        RECT 78.200 183.195 78.520 183.455 ;
        RECT 78.750 183.395 78.890 183.595 ;
        RECT 88.775 183.595 92.665 183.735 ;
        RECT 88.775 183.550 89.425 183.595 ;
        RECT 92.075 183.550 92.665 183.595 ;
        RECT 100.740 183.735 101.060 183.795 ;
        RECT 104.535 183.735 104.825 183.780 ;
        RECT 107.775 183.735 108.425 183.780 ;
        RECT 100.740 183.595 108.425 183.735 ;
        RECT 88.780 183.535 89.100 183.550 ;
        RECT 80.055 183.395 80.345 183.440 ;
        RECT 78.750 183.255 80.345 183.395 ;
        RECT 80.055 183.210 80.345 183.255 ;
        RECT 80.515 183.395 80.805 183.440 ;
        RECT 81.880 183.395 82.200 183.455 ;
        RECT 80.515 183.255 82.200 183.395 ;
        RECT 80.515 183.210 80.805 183.255 ;
        RECT 81.880 183.195 82.200 183.255 ;
        RECT 82.800 183.195 83.120 183.455 ;
        RECT 85.580 183.395 85.870 183.440 ;
        RECT 87.415 183.395 87.705 183.440 ;
        RECT 90.995 183.395 91.285 183.440 ;
        RECT 85.580 183.255 91.285 183.395 ;
        RECT 85.580 183.210 85.870 183.255 ;
        RECT 87.415 183.210 87.705 183.255 ;
        RECT 90.995 183.210 91.285 183.255 ;
        RECT 92.075 183.235 92.365 183.550 ;
        RECT 100.740 183.535 101.060 183.595 ;
        RECT 104.535 183.550 105.125 183.595 ;
        RECT 107.775 183.550 108.425 183.595 ;
        RECT 92.920 183.395 93.240 183.455 ;
        RECT 95.695 183.395 95.985 183.440 ;
        RECT 92.920 183.255 95.985 183.395 ;
        RECT 92.920 183.195 93.240 183.255 ;
        RECT 95.695 183.210 95.985 183.255 ;
        RECT 104.835 183.235 105.125 183.550 ;
        RECT 105.915 183.395 106.205 183.440 ;
        RECT 109.495 183.395 109.785 183.440 ;
        RECT 111.330 183.395 111.620 183.440 ;
        RECT 105.915 183.255 111.620 183.395 ;
        RECT 105.915 183.210 106.205 183.255 ;
        RECT 109.495 183.210 109.785 183.255 ;
        RECT 111.330 183.210 111.620 183.255 ;
        RECT 111.780 183.395 112.100 183.455 ;
        RECT 113.160 183.395 113.480 183.455 ;
        RECT 111.780 183.255 113.480 183.395 ;
        RECT 111.780 183.195 112.100 183.255 ;
        RECT 113.160 183.195 113.480 183.255 ;
        RECT 49.220 183.055 49.540 183.115 ;
        RECT 50.155 183.055 50.445 183.100 ;
        RECT 54.295 183.055 54.585 183.100 ;
        RECT 49.220 182.915 50.445 183.055 ;
        RECT 49.220 182.855 49.540 182.915 ;
        RECT 50.155 182.870 50.445 182.915 ;
        RECT 51.150 182.915 54.585 183.055 ;
        RECT 43.330 182.575 46.690 182.715 ;
        RECT 46.920 182.715 47.240 182.775 ;
        RECT 51.150 182.715 51.290 182.915 ;
        RECT 54.295 182.870 54.585 182.915 ;
        RECT 63.940 183.055 64.260 183.115 ;
        RECT 66.255 183.055 66.545 183.100 ;
        RECT 63.940 182.915 66.545 183.055 ;
        RECT 63.940 182.855 64.260 182.915 ;
        RECT 66.255 182.870 66.545 182.915 ;
        RECT 66.700 183.055 67.020 183.115 ;
        RECT 68.555 183.055 68.845 183.100 ;
        RECT 69.460 183.055 69.780 183.115 ;
        RECT 71.300 183.055 71.620 183.115 ;
        RECT 66.700 182.915 71.620 183.055 ;
        RECT 66.700 182.855 67.020 182.915 ;
        RECT 68.555 182.870 68.845 182.915 ;
        RECT 69.460 182.855 69.780 182.915 ;
        RECT 71.300 182.855 71.620 182.915 ;
        RECT 73.615 182.870 73.905 183.100 ;
        RECT 74.075 183.055 74.365 183.100 ;
        RECT 75.440 183.055 75.760 183.115 ;
        RECT 74.075 182.915 75.760 183.055 ;
        RECT 74.075 182.870 74.365 182.915 ;
        RECT 46.920 182.575 51.290 182.715 ;
        RECT 72.220 182.715 72.540 182.775 ;
        RECT 73.690 182.715 73.830 182.870 ;
        RECT 75.440 182.855 75.760 182.915 ;
        RECT 77.740 182.855 78.060 183.115 ;
        RECT 78.660 183.055 78.980 183.115 ;
        RECT 79.135 183.055 79.425 183.100 ;
        RECT 78.660 182.915 79.425 183.055 ;
        RECT 78.660 182.855 78.980 182.915 ;
        RECT 79.135 182.870 79.425 182.915 ;
        RECT 79.580 183.055 79.900 183.115 ;
        RECT 85.115 183.055 85.405 183.100 ;
        RECT 86.480 183.055 86.800 183.115 ;
        RECT 79.580 182.915 82.570 183.055 ;
        RECT 79.210 182.715 79.350 182.870 ;
        RECT 79.580 182.855 79.900 182.915 ;
        RECT 82.430 182.760 82.570 182.915 ;
        RECT 85.115 182.915 86.800 183.055 ;
        RECT 85.115 182.870 85.405 182.915 ;
        RECT 86.480 182.855 86.800 182.915 ;
        RECT 92.460 183.055 92.780 183.115 ;
        RECT 93.855 183.055 94.145 183.100 ;
        RECT 92.460 182.915 94.145 183.055 ;
        RECT 92.460 182.855 92.780 182.915 ;
        RECT 93.855 182.870 94.145 182.915 ;
        RECT 94.775 183.055 95.065 183.100 ;
        RECT 99.375 183.055 99.665 183.100 ;
        RECT 103.055 183.055 103.345 183.100 ;
        RECT 94.775 182.915 99.665 183.055 ;
        RECT 94.775 182.870 95.065 182.915 ;
        RECT 99.375 182.870 99.665 182.915 ;
        RECT 99.910 182.915 103.345 183.055 ;
        RECT 72.220 182.575 79.350 182.715 ;
        RECT 36.455 182.530 36.745 182.575 ;
        RECT 39.575 182.530 39.865 182.575 ;
        RECT 41.465 182.530 41.755 182.575 ;
        RECT 46.920 182.515 47.240 182.575 ;
        RECT 72.220 182.515 72.540 182.575 ;
        RECT 82.355 182.530 82.645 182.760 ;
        RECT 85.985 182.715 86.275 182.760 ;
        RECT 87.875 182.715 88.165 182.760 ;
        RECT 90.995 182.715 91.285 182.760 ;
        RECT 85.985 182.575 91.285 182.715 ;
        RECT 85.985 182.530 86.275 182.575 ;
        RECT 87.875 182.530 88.165 182.575 ;
        RECT 90.995 182.530 91.285 182.575 ;
        RECT 93.380 182.715 93.700 182.775 ;
        RECT 94.850 182.715 94.990 182.870 ;
        RECT 93.380 182.575 94.990 182.715 ;
        RECT 97.060 182.715 97.380 182.775 ;
        RECT 98.900 182.715 99.220 182.775 ;
        RECT 99.910 182.715 100.050 182.915 ;
        RECT 103.055 182.870 103.345 182.915 ;
        RECT 97.060 182.575 100.050 182.715 ;
        RECT 105.915 182.715 106.205 182.760 ;
        RECT 109.035 182.715 109.325 182.760 ;
        RECT 110.925 182.715 111.215 182.760 ;
        RECT 105.915 182.575 111.215 182.715 ;
        RECT 93.380 182.515 93.700 182.575 ;
        RECT 97.060 182.515 97.380 182.575 ;
        RECT 98.900 182.515 99.220 182.575 ;
        RECT 105.915 182.530 106.205 182.575 ;
        RECT 109.035 182.530 109.325 182.575 ;
        RECT 110.925 182.530 111.215 182.575 ;
        RECT 44.620 182.375 44.940 182.435 ;
        RECT 35.970 182.235 44.940 182.375 ;
        RECT 23.920 182.175 24.240 182.235 ;
        RECT 26.680 182.175 27.000 182.235 ;
        RECT 33.120 182.175 33.440 182.235 ;
        RECT 33.595 182.190 33.885 182.235 ;
        RECT 44.620 182.175 44.940 182.235 ;
        RECT 57.960 182.375 58.280 182.435 ;
        RECT 72.680 182.375 73.000 182.435 ;
        RECT 57.960 182.235 73.000 182.375 ;
        RECT 57.960 182.175 58.280 182.235 ;
        RECT 72.680 182.175 73.000 182.235 ;
        RECT 83.735 182.375 84.025 182.420 ;
        RECT 84.180 182.375 84.500 182.435 ;
        RECT 83.735 182.235 84.500 182.375 ;
        RECT 83.735 182.190 84.025 182.235 ;
        RECT 84.180 182.175 84.500 182.235 ;
        RECT 85.560 182.375 85.880 182.435 ;
        RECT 86.405 182.375 86.695 182.420 ;
        RECT 85.560 182.235 86.695 182.375 ;
        RECT 85.560 182.175 85.880 182.235 ;
        RECT 86.405 182.190 86.695 182.235 ;
        RECT 97.995 182.375 98.285 182.420 ;
        RECT 99.820 182.375 100.140 182.435 ;
        RECT 97.995 182.235 100.140 182.375 ;
        RECT 97.995 182.190 98.285 182.235 ;
        RECT 99.820 182.175 100.140 182.235 ;
        RECT 102.135 182.375 102.425 182.420 ;
        RECT 104.420 182.375 104.740 182.435 ;
        RECT 102.135 182.235 104.740 182.375 ;
        RECT 102.135 182.190 102.425 182.235 ;
        RECT 104.420 182.175 104.740 182.235 ;
        RECT 110.510 182.375 110.800 182.420 ;
        RECT 112.700 182.375 113.020 182.435 ;
        RECT 110.510 182.235 113.020 182.375 ;
        RECT 110.510 182.190 110.800 182.235 ;
        RECT 112.700 182.175 113.020 182.235 ;
        RECT 14.650 181.555 115.850 182.035 ;
        RECT 33.595 181.355 33.885 181.400 ;
        RECT 34.500 181.355 34.820 181.415 ;
        RECT 33.595 181.215 34.820 181.355 ;
        RECT 33.595 181.170 33.885 181.215 ;
        RECT 34.500 181.155 34.820 181.215 ;
        RECT 37.735 181.355 38.025 181.400 ;
        RECT 45.080 181.355 45.400 181.415 ;
        RECT 37.735 181.215 45.400 181.355 ;
        RECT 37.735 181.170 38.025 181.215 ;
        RECT 45.080 181.155 45.400 181.215 ;
        RECT 46.920 181.155 47.240 181.415 ;
        RECT 68.080 181.355 68.400 181.415 ;
        RECT 62.650 181.215 68.400 181.355 ;
        RECT 24.955 181.015 25.245 181.060 ;
        RECT 28.075 181.015 28.365 181.060 ;
        RECT 29.965 181.015 30.255 181.060 ;
        RECT 33.120 181.015 33.440 181.075 ;
        RECT 47.395 181.015 47.685 181.060 ;
        RECT 48.300 181.015 48.620 181.075 ;
        RECT 24.955 180.875 30.255 181.015 ;
        RECT 24.955 180.830 25.245 180.875 ;
        RECT 28.075 180.830 28.365 180.875 ;
        RECT 29.965 180.830 30.255 180.875 ;
        RECT 30.450 180.875 33.440 181.015 ;
        RECT 18.875 180.675 19.165 180.720 ;
        RECT 30.450 180.675 30.590 180.875 ;
        RECT 33.120 180.815 33.440 180.875 ;
        RECT 35.050 180.875 48.620 181.015 ;
        RECT 18.875 180.535 30.590 180.675 ;
        RECT 18.875 180.490 19.165 180.535 ;
        RECT 30.820 180.475 31.140 180.735 ;
        RECT 35.050 180.720 35.190 180.875 ;
        RECT 47.395 180.830 47.685 180.875 ;
        RECT 48.300 180.815 48.620 180.875 ;
        RECT 50.255 181.015 50.545 181.060 ;
        RECT 53.375 181.015 53.665 181.060 ;
        RECT 55.265 181.015 55.555 181.060 ;
        RECT 50.255 180.875 55.555 181.015 ;
        RECT 50.255 180.830 50.545 180.875 ;
        RECT 53.375 180.830 53.665 180.875 ;
        RECT 55.265 180.830 55.555 180.875 ;
        RECT 34.975 180.490 35.265 180.720 ;
        RECT 44.175 180.675 44.465 180.720 ;
        RECT 46.920 180.675 47.240 180.735 ;
        RECT 41.950 180.535 43.930 180.675 ;
        RECT 23.875 180.040 24.165 180.355 ;
        RECT 24.955 180.335 25.245 180.380 ;
        RECT 28.535 180.335 28.825 180.380 ;
        RECT 30.370 180.335 30.660 180.380 ;
        RECT 24.955 180.195 30.660 180.335 ;
        RECT 24.955 180.150 25.245 180.195 ;
        RECT 28.535 180.150 28.825 180.195 ;
        RECT 30.370 180.150 30.660 180.195 ;
        RECT 33.120 180.335 33.440 180.395 ;
        RECT 36.800 180.335 37.120 180.395 ;
        RECT 33.120 180.195 37.120 180.335 ;
        RECT 33.120 180.135 33.440 180.195 ;
        RECT 36.800 180.135 37.120 180.195 ;
        RECT 40.940 180.135 41.260 180.395 ;
        RECT 41.950 180.380 42.090 180.535 ;
        RECT 41.415 180.150 41.705 180.380 ;
        RECT 41.875 180.150 42.165 180.380 ;
        RECT 42.795 180.335 43.085 180.380 ;
        RECT 43.790 180.335 43.930 180.535 ;
        RECT 44.175 180.535 47.240 180.675 ;
        RECT 44.175 180.490 44.465 180.535 ;
        RECT 46.920 180.475 47.240 180.535 ;
        RECT 51.980 180.675 52.300 180.735 ;
        RECT 51.980 180.535 56.350 180.675 ;
        RECT 51.980 180.475 52.300 180.535 ;
        RECT 44.620 180.335 44.940 180.395 ;
        RECT 42.795 180.195 43.470 180.335 ;
        RECT 43.790 180.195 44.940 180.335 ;
        RECT 42.795 180.150 43.085 180.195 ;
        RECT 23.575 179.995 24.165 180.040 ;
        RECT 24.380 179.995 24.700 180.055 ;
        RECT 26.815 179.995 27.465 180.040 ;
        RECT 23.575 179.855 27.465 179.995 ;
        RECT 23.575 179.810 23.865 179.855 ;
        RECT 24.380 179.795 24.700 179.855 ;
        RECT 26.815 179.810 27.465 179.855 ;
        RECT 29.455 179.810 29.745 180.040 ;
        RECT 41.490 179.995 41.630 180.150 ;
        RECT 41.490 179.855 42.550 179.995 ;
        RECT 21.620 179.455 21.940 179.715 ;
        RECT 22.095 179.655 22.385 179.700 ;
        RECT 22.540 179.655 22.860 179.715 ;
        RECT 22.095 179.515 22.860 179.655 ;
        RECT 22.095 179.470 22.385 179.515 ;
        RECT 22.540 179.455 22.860 179.515 ;
        RECT 26.220 179.655 26.540 179.715 ;
        RECT 29.530 179.655 29.670 179.810 ;
        RECT 42.410 179.715 42.550 179.855 ;
        RECT 43.330 179.715 43.470 180.195 ;
        RECT 44.620 180.135 44.940 180.195 ;
        RECT 45.080 180.135 45.400 180.395 ;
        RECT 49.220 180.355 49.540 180.395 ;
        RECT 56.210 180.380 56.350 180.535 ;
        RECT 58.880 180.475 59.200 180.735 ;
        RECT 60.735 180.675 61.025 180.720 ;
        RECT 61.180 180.675 61.500 180.735 ;
        RECT 62.650 180.720 62.790 181.215 ;
        RECT 68.080 181.155 68.400 181.215 ;
        RECT 72.220 181.155 72.540 181.415 ;
        RECT 73.140 181.155 73.460 181.415 ;
        RECT 78.660 181.355 78.980 181.415 ;
        RECT 97.520 181.355 97.840 181.415 ;
        RECT 98.915 181.355 99.205 181.400 ;
        RECT 78.660 181.215 89.930 181.355 ;
        RECT 78.660 181.155 78.980 181.215 ;
        RECT 66.255 181.015 66.545 181.060 ;
        RECT 67.620 181.015 67.940 181.075 ;
        RECT 66.255 180.875 67.940 181.015 ;
        RECT 66.255 180.830 66.545 180.875 ;
        RECT 60.735 180.535 61.500 180.675 ;
        RECT 60.735 180.490 61.025 180.535 ;
        RECT 61.180 180.475 61.500 180.535 ;
        RECT 62.575 180.490 62.865 180.720 ;
        RECT 63.035 180.675 63.325 180.720 ;
        RECT 64.400 180.675 64.720 180.735 ;
        RECT 66.330 180.675 66.470 180.830 ;
        RECT 67.620 180.815 67.940 180.875 ;
        RECT 79.695 181.015 79.985 181.060 ;
        RECT 82.815 181.015 83.105 181.060 ;
        RECT 84.705 181.015 84.995 181.060 ;
        RECT 79.695 180.875 84.995 181.015 ;
        RECT 79.695 180.830 79.985 180.875 ;
        RECT 82.815 180.830 83.105 180.875 ;
        RECT 84.705 180.830 84.995 180.875 ;
        RECT 63.035 180.535 66.470 180.675 ;
        RECT 63.035 180.490 63.325 180.535 ;
        RECT 64.400 180.475 64.720 180.535 ;
        RECT 68.540 180.475 68.860 180.735 ;
        RECT 76.835 180.490 77.125 180.720 ;
        RECT 49.175 180.135 49.540 180.355 ;
        RECT 50.255 180.335 50.545 180.380 ;
        RECT 53.835 180.335 54.125 180.380 ;
        RECT 55.670 180.335 55.960 180.380 ;
        RECT 50.255 180.195 55.960 180.335 ;
        RECT 50.255 180.150 50.545 180.195 ;
        RECT 53.835 180.150 54.125 180.195 ;
        RECT 55.670 180.150 55.960 180.195 ;
        RECT 56.135 180.150 56.425 180.380 ;
        RECT 49.175 180.040 49.465 180.135 ;
        RECT 48.875 179.995 49.465 180.040 ;
        RECT 52.115 179.995 52.765 180.040 ;
        RECT 48.875 179.855 52.765 179.995 ;
        RECT 48.875 179.810 49.165 179.855 ;
        RECT 52.115 179.810 52.765 179.855 ;
        RECT 54.755 179.810 55.045 180.040 ;
        RECT 56.210 179.995 56.350 180.150 ;
        RECT 57.960 180.135 58.280 180.395 ;
        RECT 61.655 180.150 61.945 180.380 ;
        RECT 62.115 180.335 62.405 180.380 ;
        RECT 67.620 180.335 67.940 180.395 ;
        RECT 68.630 180.335 68.770 180.475 ;
        RECT 72.220 180.335 72.540 180.395 ;
        RECT 62.115 180.195 72.540 180.335 ;
        RECT 62.115 180.150 62.405 180.195 ;
        RECT 60.720 179.995 61.040 180.055 ;
        RECT 56.210 179.855 61.040 179.995 ;
        RECT 61.730 179.995 61.870 180.150 ;
        RECT 67.620 180.135 67.940 180.195 ;
        RECT 72.220 180.135 72.540 180.195 ;
        RECT 75.900 180.335 76.220 180.395 ;
        RECT 76.910 180.335 77.050 180.490 ;
        RECT 84.180 180.475 84.500 180.735 ;
        RECT 85.575 180.675 85.865 180.720 ;
        RECT 86.020 180.675 86.340 180.735 ;
        RECT 85.575 180.535 86.340 180.675 ;
        RECT 89.790 180.675 89.930 181.215 ;
        RECT 97.520 181.215 99.205 181.355 ;
        RECT 97.520 181.155 97.840 181.215 ;
        RECT 98.915 181.170 99.205 181.215 ;
        RECT 111.335 181.355 111.625 181.400 ;
        RECT 112.240 181.355 112.560 181.415 ;
        RECT 111.335 181.215 112.560 181.355 ;
        RECT 111.335 181.170 111.625 181.215 ;
        RECT 112.240 181.155 112.560 181.215 ;
        RECT 110.875 181.015 111.165 181.060 ;
        RECT 112.700 181.015 113.020 181.075 ;
        RECT 93.470 180.875 102.810 181.015 ;
        RECT 93.470 180.735 93.610 180.875 ;
        RECT 93.380 180.675 93.700 180.735 ;
        RECT 89.790 180.535 93.700 180.675 ;
        RECT 85.575 180.490 85.865 180.535 ;
        RECT 86.020 180.475 86.340 180.535 ;
        RECT 93.380 180.475 93.700 180.535 ;
        RECT 93.840 180.675 94.160 180.735 ;
        RECT 102.670 180.720 102.810 180.875 ;
        RECT 110.875 180.875 113.020 181.015 ;
        RECT 110.875 180.830 111.165 180.875 ;
        RECT 112.700 180.815 113.020 180.875 ;
        RECT 93.840 180.535 97.750 180.675 ;
        RECT 93.840 180.475 94.160 180.535 ;
        RECT 75.900 180.195 77.050 180.335 ;
        RECT 75.900 180.135 76.220 180.195 ;
        RECT 66.255 179.995 66.545 180.040 ;
        RECT 66.700 179.995 67.020 180.055 ;
        RECT 61.730 179.855 67.020 179.995 ;
        RECT 26.220 179.515 29.670 179.655 ;
        RECT 39.575 179.655 39.865 179.700 ;
        RECT 41.400 179.655 41.720 179.715 ;
        RECT 39.575 179.515 41.720 179.655 ;
        RECT 26.220 179.455 26.540 179.515 ;
        RECT 39.575 179.470 39.865 179.515 ;
        RECT 41.400 179.455 41.720 179.515 ;
        RECT 42.320 179.455 42.640 179.715 ;
        RECT 43.240 179.455 43.560 179.715 ;
        RECT 54.830 179.655 54.970 179.810 ;
        RECT 60.720 179.795 61.040 179.855 ;
        RECT 66.255 179.810 66.545 179.855 ;
        RECT 66.700 179.795 67.020 179.855 ;
        RECT 68.080 179.995 68.400 180.055 ;
        RECT 69.015 179.995 69.305 180.040 ;
        RECT 68.080 179.855 69.305 179.995 ;
        RECT 68.080 179.795 68.400 179.855 ;
        RECT 69.015 179.810 69.305 179.855 ;
        RECT 70.840 179.795 71.160 180.055 ;
        RECT 77.740 179.995 78.060 180.055 ;
        RECT 78.615 180.040 78.905 180.355 ;
        RECT 79.695 180.335 79.985 180.380 ;
        RECT 83.275 180.335 83.565 180.380 ;
        RECT 85.110 180.335 85.400 180.380 ;
        RECT 79.695 180.195 85.400 180.335 ;
        RECT 79.695 180.150 79.985 180.195 ;
        RECT 83.275 180.150 83.565 180.195 ;
        RECT 85.110 180.150 85.400 180.195 ;
        RECT 86.495 180.335 86.785 180.380 ;
        RECT 87.400 180.335 87.720 180.395 ;
        RECT 86.495 180.195 87.720 180.335 ;
        RECT 86.495 180.150 86.785 180.195 ;
        RECT 87.400 180.135 87.720 180.195 ;
        RECT 89.255 180.335 89.545 180.380 ;
        RECT 92.015 180.335 92.305 180.380 ;
        RECT 92.920 180.335 93.240 180.395 ;
        RECT 89.255 180.195 93.240 180.335 ;
        RECT 89.255 180.150 89.545 180.195 ;
        RECT 92.015 180.150 92.305 180.195 ;
        RECT 92.920 180.135 93.240 180.195 ;
        RECT 94.300 180.335 94.620 180.395 ;
        RECT 97.610 180.380 97.750 180.535 ;
        RECT 98.530 180.535 100.510 180.675 ;
        RECT 98.530 180.395 98.670 180.535 ;
        RECT 96.615 180.335 96.905 180.380 ;
        RECT 94.300 180.195 96.905 180.335 ;
        RECT 94.300 180.135 94.620 180.195 ;
        RECT 96.615 180.150 96.905 180.195 ;
        RECT 97.075 180.150 97.365 180.380 ;
        RECT 97.535 180.150 97.825 180.380 ;
        RECT 78.315 179.995 78.905 180.040 ;
        RECT 81.555 179.995 82.205 180.040 ;
        RECT 77.740 179.855 82.205 179.995 ;
        RECT 97.150 179.995 97.290 180.150 ;
        RECT 98.440 180.135 98.760 180.395 ;
        RECT 99.820 180.135 100.140 180.395 ;
        RECT 100.370 180.335 100.510 180.535 ;
        RECT 102.595 180.490 102.885 180.720 ;
        RECT 104.420 180.675 104.740 180.735 ;
        RECT 104.420 180.535 110.170 180.675 ;
        RECT 104.420 180.475 104.740 180.535 ;
        RECT 106.275 180.335 106.565 180.380 ;
        RECT 100.370 180.195 106.565 180.335 ;
        RECT 106.275 180.150 106.565 180.195 ;
        RECT 107.180 180.135 107.500 180.395 ;
        RECT 107.655 180.150 107.945 180.380 ;
        RECT 97.980 179.995 98.300 180.055 ;
        RECT 107.730 179.995 107.870 180.150 ;
        RECT 108.100 180.135 108.420 180.395 ;
        RECT 110.030 180.380 110.170 180.535 ;
        RECT 109.955 180.150 110.245 180.380 ;
        RECT 112.240 180.135 112.560 180.395 ;
        RECT 97.150 179.855 107.870 179.995 ;
        RECT 77.740 179.795 78.060 179.855 ;
        RECT 78.315 179.810 78.605 179.855 ;
        RECT 81.555 179.810 82.205 179.855 ;
        RECT 97.980 179.795 98.300 179.855 ;
        RECT 57.960 179.655 58.280 179.715 ;
        RECT 54.830 179.515 58.280 179.655 ;
        RECT 57.960 179.455 58.280 179.515 ;
        RECT 68.540 179.655 68.860 179.715 ;
        RECT 69.935 179.655 70.225 179.700 ;
        RECT 68.540 179.515 70.225 179.655 ;
        RECT 68.540 179.455 68.860 179.515 ;
        RECT 69.935 179.470 70.225 179.515 ;
        RECT 90.160 179.455 90.480 179.715 ;
        RECT 92.460 179.455 92.780 179.715 ;
        RECT 92.920 179.655 93.240 179.715 ;
        RECT 95.235 179.655 95.525 179.700 ;
        RECT 92.920 179.515 95.525 179.655 ;
        RECT 92.920 179.455 93.240 179.515 ;
        RECT 95.235 179.470 95.525 179.515 ;
        RECT 103.500 179.455 103.820 179.715 ;
        RECT 103.960 179.455 104.280 179.715 ;
        RECT 105.800 179.455 106.120 179.715 ;
        RECT 109.480 179.455 109.800 179.715 ;
        RECT 14.650 178.835 115.850 179.315 ;
        RECT 26.220 178.635 26.540 178.695 ;
        RECT 26.695 178.635 26.985 178.680 ;
        RECT 26.220 178.495 26.985 178.635 ;
        RECT 26.220 178.435 26.540 178.495 ;
        RECT 26.695 178.450 26.985 178.495 ;
        RECT 48.300 178.435 48.620 178.695 ;
        RECT 57.960 178.435 58.280 178.695 ;
        RECT 66.700 178.435 67.020 178.695 ;
        RECT 67.620 178.635 67.940 178.695 ;
        RECT 67.260 178.495 67.940 178.635 ;
        RECT 21.620 178.295 21.940 178.355 ;
        RECT 34.975 178.295 35.265 178.340 ;
        RECT 55.215 178.295 55.505 178.340 ;
        RECT 21.620 178.155 35.265 178.295 ;
        RECT 21.620 178.095 21.940 178.155 ;
        RECT 34.975 178.110 35.265 178.155 ;
        RECT 47.930 178.155 55.505 178.295 ;
        RECT 24.855 177.955 25.145 178.000 ;
        RECT 25.775 177.955 26.065 178.000 ;
        RECT 24.855 177.815 26.065 177.955 ;
        RECT 24.855 177.770 25.145 177.815 ;
        RECT 25.775 177.770 26.065 177.815 ;
        RECT 26.680 177.955 27.000 178.015 ;
        RECT 27.155 177.955 27.445 178.000 ;
        RECT 26.680 177.815 27.445 177.955 ;
        RECT 26.680 177.755 27.000 177.815 ;
        RECT 27.155 177.770 27.445 177.815 ;
        RECT 30.360 177.955 30.680 178.015 ;
        RECT 34.515 177.955 34.805 178.000 ;
        RECT 30.360 177.815 34.805 177.955 ;
        RECT 30.360 177.755 30.680 177.815 ;
        RECT 34.515 177.770 34.805 177.815 ;
        RECT 40.940 177.955 41.260 178.015 ;
        RECT 41.860 177.955 42.180 178.015 ;
        RECT 40.940 177.815 42.180 177.955 ;
        RECT 40.940 177.755 41.260 177.815 ;
        RECT 41.860 177.755 42.180 177.815 ;
        RECT 42.320 177.755 42.640 178.015 ;
        RECT 42.780 177.755 43.100 178.015 ;
        RECT 43.240 177.955 43.560 178.015 ;
        RECT 43.715 177.955 44.005 178.000 ;
        RECT 43.240 177.815 44.005 177.955 ;
        RECT 43.240 177.755 43.560 177.815 ;
        RECT 43.715 177.770 44.005 177.815 ;
        RECT 22.095 177.430 22.385 177.660 ;
        RECT 22.540 177.615 22.860 177.675 ;
        RECT 30.835 177.615 31.125 177.660 ;
        RECT 22.540 177.475 31.125 177.615 ;
        RECT 22.170 177.275 22.310 177.430 ;
        RECT 22.540 177.415 22.860 177.475 ;
        RECT 30.835 177.430 31.125 177.475 ;
        RECT 31.740 177.615 32.060 177.675 ;
        RECT 34.055 177.615 34.345 177.660 ;
        RECT 46.920 177.615 47.240 177.675 ;
        RECT 47.930 177.660 48.070 178.155 ;
        RECT 55.215 178.110 55.505 178.155 ;
        RECT 57.055 178.295 57.345 178.340 ;
        RECT 66.790 178.295 66.930 178.435 ;
        RECT 57.055 178.155 66.930 178.295 ;
        RECT 57.055 178.110 57.345 178.155 ;
        RECT 48.300 177.955 48.620 178.015 ;
        RECT 48.775 177.955 49.065 178.000 ;
        RECT 48.300 177.815 49.065 177.955 ;
        RECT 48.300 177.755 48.620 177.815 ;
        RECT 48.775 177.770 49.065 177.815 ;
        RECT 54.755 177.955 55.045 178.000 ;
        RECT 58.895 177.955 59.185 178.000 ;
        RECT 54.755 177.815 59.185 177.955 ;
        RECT 54.755 177.770 55.045 177.815 ;
        RECT 58.895 177.770 59.185 177.815 ;
        RECT 62.560 177.755 62.880 178.015 ;
        RECT 63.940 177.955 64.260 178.015 ;
        RECT 65.335 177.955 65.625 178.000 ;
        RECT 63.940 177.815 65.625 177.955 ;
        RECT 63.940 177.755 64.260 177.815 ;
        RECT 65.335 177.770 65.625 177.815 ;
        RECT 66.240 177.955 66.560 178.015 ;
        RECT 67.260 178.000 67.400 178.495 ;
        RECT 67.620 178.435 67.940 178.495 ;
        RECT 82.355 178.635 82.645 178.680 ;
        RECT 82.800 178.635 83.120 178.695 ;
        RECT 82.355 178.495 83.120 178.635 ;
        RECT 82.355 178.450 82.645 178.495 ;
        RECT 82.800 178.435 83.120 178.495 ;
        RECT 85.560 178.635 85.880 178.695 ;
        RECT 86.495 178.635 86.785 178.680 ;
        RECT 85.560 178.495 86.785 178.635 ;
        RECT 85.560 178.435 85.880 178.495 ;
        RECT 86.495 178.450 86.785 178.495 ;
        RECT 107.195 178.635 107.485 178.680 ;
        RECT 112.240 178.635 112.560 178.695 ;
        RECT 107.195 178.495 112.560 178.635 ;
        RECT 107.195 178.450 107.485 178.495 ;
        RECT 112.240 178.435 112.560 178.495 ;
        RECT 68.080 178.295 68.400 178.355 ;
        RECT 72.680 178.295 73.000 178.355 ;
        RECT 87.400 178.295 87.720 178.355 ;
        RECT 97.980 178.295 98.300 178.355 ;
        RECT 108.100 178.295 108.420 178.355 ;
        RECT 68.080 178.155 71.990 178.295 ;
        RECT 68.080 178.095 68.400 178.155 ;
        RECT 66.715 177.955 67.005 178.000 ;
        RECT 66.240 177.815 67.005 177.955 ;
        RECT 66.240 177.755 66.560 177.815 ;
        RECT 66.715 177.770 67.005 177.815 ;
        RECT 67.185 177.770 67.475 178.000 ;
        RECT 67.635 177.770 67.925 178.000 ;
        RECT 47.855 177.615 48.145 177.660 ;
        RECT 31.740 177.475 48.145 177.615 ;
        RECT 31.740 177.415 32.060 177.475 ;
        RECT 34.055 177.430 34.345 177.475 ;
        RECT 46.920 177.415 47.240 177.475 ;
        RECT 47.855 177.430 48.145 177.475 ;
        RECT 51.535 177.430 51.825 177.660 ;
        RECT 64.400 177.615 64.720 177.675 ;
        RECT 67.710 177.615 67.850 177.770 ;
        RECT 71.300 177.755 71.620 178.015 ;
        RECT 71.850 178.000 71.990 178.155 ;
        RECT 72.680 178.155 83.030 178.295 ;
        RECT 72.680 178.095 73.000 178.155 ;
        RECT 71.775 177.770 72.065 178.000 ;
        RECT 72.220 177.755 72.540 178.015 ;
        RECT 74.520 177.755 74.840 178.015 ;
        RECT 74.995 177.770 75.285 178.000 ;
        RECT 75.455 177.955 75.745 178.000 ;
        RECT 75.900 177.955 76.220 178.015 ;
        RECT 75.455 177.815 76.220 177.955 ;
        RECT 75.455 177.770 75.745 177.815 ;
        RECT 64.400 177.475 67.850 177.615 ;
        RECT 28.535 177.275 28.825 177.320 ;
        RECT 22.170 177.135 28.825 177.275 ;
        RECT 28.535 177.090 28.825 177.135 ;
        RECT 50.615 177.275 50.905 177.320 ;
        RECT 51.610 177.275 51.750 177.430 ;
        RECT 64.400 177.415 64.720 177.475 ;
        RECT 68.080 177.415 68.400 177.675 ;
        RECT 69.460 177.615 69.780 177.675 ;
        RECT 70.855 177.615 71.145 177.660 ;
        RECT 69.460 177.475 71.145 177.615 ;
        RECT 75.070 177.615 75.210 177.770 ;
        RECT 75.900 177.755 76.220 177.815 ;
        RECT 76.360 177.755 76.680 178.015 ;
        RECT 79.120 177.755 79.440 178.015 ;
        RECT 82.890 178.000 83.030 178.155 ;
        RECT 87.400 178.155 93.150 178.295 ;
        RECT 87.400 178.095 87.720 178.155 ;
        RECT 82.815 177.770 83.105 178.000 ;
        RECT 85.575 177.955 85.865 178.000 ;
        RECT 86.955 177.955 87.245 178.000 ;
        RECT 85.575 177.815 87.245 177.955 ;
        RECT 85.575 177.770 85.865 177.815 ;
        RECT 86.955 177.770 87.245 177.815 ;
        RECT 90.160 177.755 90.480 178.015 ;
        RECT 93.010 178.000 93.150 178.155 ;
        RECT 96.230 178.155 100.510 178.295 ;
        RECT 92.015 177.955 92.305 178.000 ;
        RECT 90.710 177.815 92.305 177.955 ;
        RECT 78.660 177.615 78.980 177.675 ;
        RECT 75.070 177.475 78.980 177.615 ;
        RECT 69.460 177.415 69.780 177.475 ;
        RECT 70.855 177.430 71.145 177.475 ;
        RECT 78.660 177.415 78.980 177.475 ;
        RECT 84.180 177.415 84.500 177.675 ;
        RECT 87.860 177.615 88.180 177.675 ;
        RECT 90.710 177.615 90.850 177.815 ;
        RECT 92.015 177.770 92.305 177.815 ;
        RECT 92.475 177.770 92.765 178.000 ;
        RECT 92.935 177.770 93.225 178.000 ;
        RECT 93.855 177.955 94.145 178.000 ;
        RECT 94.300 177.955 94.620 178.015 ;
        RECT 93.855 177.815 94.620 177.955 ;
        RECT 93.855 177.770 94.145 177.815 ;
        RECT 87.860 177.475 90.850 177.615 ;
        RECT 87.860 177.415 88.180 177.475 ;
        RECT 50.615 177.135 51.750 177.275 ;
        RECT 63.035 177.275 63.325 177.320 ;
        RECT 65.320 177.275 65.640 177.335 ;
        RECT 63.035 177.135 65.640 177.275 ;
        RECT 50.615 177.090 50.905 177.135 ;
        RECT 63.035 177.090 63.325 177.135 ;
        RECT 65.320 177.075 65.640 177.135 ;
        RECT 65.795 177.275 66.085 177.320 ;
        RECT 69.000 177.275 69.320 177.335 ;
        RECT 65.795 177.135 67.055 177.275 ;
        RECT 65.795 177.090 66.085 177.135 ;
        RECT 27.600 176.735 27.920 176.995 ;
        RECT 36.815 176.935 37.105 176.980 ;
        RECT 37.720 176.935 38.040 176.995 ;
        RECT 36.815 176.795 38.040 176.935 ;
        RECT 36.815 176.750 37.105 176.795 ;
        RECT 37.720 176.735 38.040 176.795 ;
        RECT 40.020 176.935 40.340 176.995 ;
        RECT 40.495 176.935 40.785 176.980 ;
        RECT 40.020 176.795 40.785 176.935 ;
        RECT 40.020 176.735 40.340 176.795 ;
        RECT 40.495 176.750 40.785 176.795 ;
        RECT 64.415 176.935 64.705 176.980 ;
        RECT 64.860 176.935 65.180 176.995 ;
        RECT 64.415 176.795 65.180 176.935 ;
        RECT 66.915 176.935 67.055 177.135 ;
        RECT 67.710 177.135 69.320 177.275 ;
        RECT 90.710 177.275 90.850 177.475 ;
        RECT 91.540 177.615 91.860 177.675 ;
        RECT 92.550 177.615 92.690 177.770 ;
        RECT 94.300 177.755 94.620 177.815 ;
        RECT 95.680 177.755 96.000 178.015 ;
        RECT 96.230 178.000 96.370 178.155 ;
        RECT 97.980 178.095 98.300 178.155 ;
        RECT 100.370 178.015 100.510 178.155 ;
        RECT 100.830 178.155 108.420 178.295 ;
        RECT 96.155 177.770 96.445 178.000 ;
        RECT 96.615 177.955 96.905 178.000 ;
        RECT 97.060 177.955 97.380 178.015 ;
        RECT 96.615 177.815 97.380 177.955 ;
        RECT 96.615 177.770 96.905 177.815 ;
        RECT 96.230 177.615 96.370 177.770 ;
        RECT 97.060 177.755 97.380 177.815 ;
        RECT 97.520 177.955 97.840 178.015 ;
        RECT 98.440 177.955 98.760 178.015 ;
        RECT 98.915 177.955 99.205 178.000 ;
        RECT 97.520 177.815 99.205 177.955 ;
        RECT 97.520 177.755 97.840 177.815 ;
        RECT 98.440 177.755 98.760 177.815 ;
        RECT 98.915 177.770 99.205 177.815 ;
        RECT 99.360 177.955 99.680 178.015 ;
        RECT 99.835 177.955 100.125 178.000 ;
        RECT 99.360 177.815 100.125 177.955 ;
        RECT 99.360 177.755 99.680 177.815 ;
        RECT 99.835 177.770 100.125 177.815 ;
        RECT 100.280 177.755 100.600 178.015 ;
        RECT 100.830 178.000 100.970 178.155 ;
        RECT 108.100 178.095 108.420 178.155 ;
        RECT 100.755 177.770 101.045 178.000 ;
        RECT 104.435 177.955 104.725 178.000 ;
        RECT 105.800 177.955 106.120 178.015 ;
        RECT 104.435 177.815 106.120 177.955 ;
        RECT 104.435 177.770 104.725 177.815 ;
        RECT 91.540 177.475 96.370 177.615 ;
        RECT 91.540 177.415 91.860 177.475 ;
        RECT 93.840 177.275 94.160 177.335 ;
        RECT 95.680 177.275 96.000 177.335 ;
        RECT 98.900 177.275 99.220 177.335 ;
        RECT 100.830 177.275 100.970 177.770 ;
        RECT 105.800 177.755 106.120 177.815 ;
        RECT 109.020 177.755 109.340 178.015 ;
        RECT 90.710 177.135 100.970 177.275 ;
        RECT 67.710 176.935 67.850 177.135 ;
        RECT 69.000 177.075 69.320 177.135 ;
        RECT 93.840 177.075 94.160 177.135 ;
        RECT 95.680 177.075 96.000 177.135 ;
        RECT 98.900 177.075 99.220 177.135 ;
        RECT 66.915 176.795 67.850 176.935 ;
        RECT 68.080 176.935 68.400 176.995 ;
        RECT 69.935 176.935 70.225 176.980 ;
        RECT 68.080 176.795 70.225 176.935 ;
        RECT 64.415 176.750 64.705 176.795 ;
        RECT 64.860 176.735 65.180 176.795 ;
        RECT 68.080 176.735 68.400 176.795 ;
        RECT 69.935 176.750 70.225 176.795 ;
        RECT 73.140 176.735 73.460 176.995 ;
        RECT 88.780 176.935 89.100 176.995 ;
        RECT 90.635 176.935 90.925 176.980 ;
        RECT 88.780 176.795 90.925 176.935 ;
        RECT 88.780 176.735 89.100 176.795 ;
        RECT 90.635 176.750 90.925 176.795 ;
        RECT 94.315 176.935 94.605 176.980 ;
        RECT 98.440 176.935 98.760 176.995 ;
        RECT 94.315 176.795 98.760 176.935 ;
        RECT 94.315 176.750 94.605 176.795 ;
        RECT 98.440 176.735 98.760 176.795 ;
        RECT 102.135 176.935 102.425 176.980 ;
        RECT 103.040 176.935 103.360 176.995 ;
        RECT 102.135 176.795 103.360 176.935 ;
        RECT 102.135 176.750 102.425 176.795 ;
        RECT 103.040 176.735 103.360 176.795 ;
        RECT 109.955 176.935 110.245 176.980 ;
        RECT 112.240 176.935 112.560 176.995 ;
        RECT 109.955 176.795 112.560 176.935 ;
        RECT 109.955 176.750 110.245 176.795 ;
        RECT 112.240 176.735 112.560 176.795 ;
        RECT 14.650 176.115 115.850 176.595 ;
        RECT 50.600 175.915 50.920 175.975 ;
        RECT 65.320 175.915 65.640 175.975 ;
        RECT 50.600 175.775 65.640 175.915 ;
        RECT 50.600 175.715 50.920 175.775 ;
        RECT 65.320 175.715 65.640 175.775 ;
        RECT 66.700 175.915 67.020 175.975 ;
        RECT 67.635 175.915 67.925 175.960 ;
        RECT 70.840 175.915 71.160 175.975 ;
        RECT 66.700 175.775 71.160 175.915 ;
        RECT 66.700 175.715 67.020 175.775 ;
        RECT 67.635 175.730 67.925 175.775 ;
        RECT 70.840 175.715 71.160 175.775 ;
        RECT 73.140 175.915 73.460 175.975 ;
        RECT 74.520 175.915 74.840 175.975 ;
        RECT 73.140 175.775 78.430 175.915 ;
        RECT 73.140 175.715 73.460 175.775 ;
        RECT 74.520 175.715 74.840 175.775 ;
        RECT 22.540 175.375 22.860 175.635 ;
        RECT 27.615 175.575 27.905 175.620 ;
        RECT 30.360 175.575 30.680 175.635 ;
        RECT 27.615 175.435 30.680 175.575 ;
        RECT 27.615 175.390 27.905 175.435 ;
        RECT 30.360 175.375 30.680 175.435 ;
        RECT 30.935 175.575 31.225 175.620 ;
        RECT 34.055 175.575 34.345 175.620 ;
        RECT 35.945 175.575 36.235 175.620 ;
        RECT 43.240 175.575 43.560 175.635 ;
        RECT 49.680 175.575 50.000 175.635 ;
        RECT 51.995 175.575 52.285 175.620 ;
        RECT 30.935 175.435 36.235 175.575 ;
        RECT 30.935 175.390 31.225 175.435 ;
        RECT 34.055 175.390 34.345 175.435 ;
        RECT 35.945 175.390 36.235 175.435 ;
        RECT 40.570 175.435 43.560 175.575 ;
        RECT 22.630 175.235 22.770 175.375 ;
        RECT 32.660 175.235 32.980 175.295 ;
        RECT 21.710 175.095 22.770 175.235 ;
        RECT 24.470 175.095 32.980 175.235 ;
        RECT 20.700 174.695 21.020 174.955 ;
        RECT 21.710 174.940 21.850 175.095 ;
        RECT 21.635 174.710 21.925 174.940 ;
        RECT 22.095 174.710 22.385 174.940 ;
        RECT 22.555 174.895 22.845 174.940 ;
        RECT 24.470 174.895 24.610 175.095 ;
        RECT 32.660 175.035 32.980 175.095 ;
        RECT 36.815 175.235 37.105 175.280 ;
        RECT 37.260 175.235 37.580 175.295 ;
        RECT 36.815 175.095 37.580 175.235 ;
        RECT 36.815 175.050 37.105 175.095 ;
        RECT 37.260 175.035 37.580 175.095 ;
        RECT 22.555 174.755 24.610 174.895 ;
        RECT 22.555 174.710 22.845 174.755 ;
        RECT 24.855 174.710 25.145 174.940 ;
        RECT 22.170 174.555 22.310 174.710 ;
        RECT 24.380 174.555 24.700 174.615 ;
        RECT 22.170 174.415 24.700 174.555 ;
        RECT 24.380 174.355 24.700 174.415 ;
        RECT 22.080 174.215 22.400 174.275 ;
        RECT 23.935 174.215 24.225 174.260 ;
        RECT 22.080 174.075 24.225 174.215 ;
        RECT 24.930 174.215 25.070 174.710 ;
        RECT 27.600 174.555 27.920 174.615 ;
        RECT 29.855 174.600 30.145 174.915 ;
        RECT 30.935 174.895 31.225 174.940 ;
        RECT 34.515 174.895 34.805 174.940 ;
        RECT 36.350 174.895 36.640 174.940 ;
        RECT 30.935 174.755 36.640 174.895 ;
        RECT 30.935 174.710 31.225 174.755 ;
        RECT 34.515 174.710 34.805 174.755 ;
        RECT 36.350 174.710 36.640 174.755 ;
        RECT 37.720 174.895 38.040 174.955 ;
        RECT 40.570 174.940 40.710 175.435 ;
        RECT 43.240 175.375 43.560 175.435 ;
        RECT 44.710 175.435 52.285 175.575 ;
        RECT 43.700 175.235 44.020 175.295 ;
        RECT 44.710 175.280 44.850 175.435 ;
        RECT 49.680 175.375 50.000 175.435 ;
        RECT 51.995 175.390 52.285 175.435 ;
        RECT 54.855 175.575 55.145 175.620 ;
        RECT 57.975 175.575 58.265 175.620 ;
        RECT 59.865 175.575 60.155 175.620 ;
        RECT 62.575 175.575 62.865 175.620 ;
        RECT 72.680 175.575 73.000 175.635 ;
        RECT 77.280 175.575 77.600 175.635 ;
        RECT 54.855 175.435 60.155 175.575 ;
        RECT 54.855 175.390 55.145 175.435 ;
        RECT 57.975 175.390 58.265 175.435 ;
        RECT 59.865 175.390 60.155 175.435 ;
        RECT 60.350 175.435 71.070 175.575 ;
        RECT 41.490 175.095 44.020 175.235 ;
        RECT 41.490 174.940 41.630 175.095 ;
        RECT 43.700 175.035 44.020 175.095 ;
        RECT 44.635 175.050 44.925 175.280 ;
        RECT 46.920 175.235 47.240 175.295 ;
        RECT 48.775 175.235 49.065 175.280 ;
        RECT 46.920 175.095 49.065 175.235 ;
        RECT 46.920 175.035 47.240 175.095 ;
        RECT 48.775 175.050 49.065 175.095 ;
        RECT 50.140 175.235 50.460 175.295 ;
        RECT 60.350 175.235 60.490 175.435 ;
        RECT 62.575 175.390 62.865 175.435 ;
        RECT 50.140 175.095 60.490 175.235 ;
        RECT 50.140 175.035 50.460 175.095 ;
        RECT 60.720 175.035 61.040 175.295 ;
        RECT 63.940 175.235 64.260 175.295 ;
        RECT 67.175 175.235 67.465 175.280 ;
        RECT 63.940 175.095 67.465 175.235 ;
        RECT 63.940 175.035 64.260 175.095 ;
        RECT 67.175 175.050 67.465 175.095 ;
        RECT 70.930 174.955 71.070 175.435 ;
        RECT 72.680 175.435 77.600 175.575 ;
        RECT 72.680 175.375 73.000 175.435 ;
        RECT 77.280 175.375 77.600 175.435 ;
        RECT 72.220 175.235 72.540 175.295 ;
        RECT 73.140 175.235 73.460 175.295 ;
        RECT 72.220 175.095 73.460 175.235 ;
        RECT 72.220 175.035 72.540 175.095 ;
        RECT 73.140 175.035 73.460 175.095 ;
        RECT 39.575 174.895 39.865 174.940 ;
        RECT 37.720 174.755 39.865 174.895 ;
        RECT 37.720 174.695 38.040 174.755 ;
        RECT 39.575 174.710 39.865 174.755 ;
        RECT 40.495 174.710 40.785 174.940 ;
        RECT 41.415 174.710 41.705 174.940 ;
        RECT 41.875 174.710 42.165 174.940 ;
        RECT 42.320 174.895 42.640 174.955 ;
        RECT 46.460 174.895 46.780 174.955 ;
        RECT 42.320 174.755 46.780 174.895 ;
        RECT 29.555 174.555 30.145 174.600 ;
        RECT 32.795 174.555 33.445 174.600 ;
        RECT 27.600 174.415 33.445 174.555 ;
        RECT 27.600 174.355 27.920 174.415 ;
        RECT 29.555 174.370 29.845 174.415 ;
        RECT 32.795 174.370 33.445 174.415 ;
        RECT 35.435 174.370 35.725 174.600 ;
        RECT 41.950 174.555 42.090 174.710 ;
        RECT 42.320 174.695 42.640 174.755 ;
        RECT 46.460 174.695 46.780 174.755 ;
        RECT 47.395 174.895 47.685 174.940 ;
        RECT 48.300 174.895 48.620 174.955 ;
        RECT 49.235 174.895 49.525 174.940 ;
        RECT 47.395 174.755 49.525 174.895 ;
        RECT 47.395 174.710 47.685 174.755 ;
        RECT 48.300 174.695 48.620 174.755 ;
        RECT 49.235 174.710 49.525 174.755 ;
        RECT 42.780 174.555 43.100 174.615 ;
        RECT 45.540 174.555 45.860 174.615 ;
        RECT 41.950 174.415 45.860 174.555 ;
        RECT 28.075 174.215 28.365 174.260 ;
        RECT 31.740 174.215 32.060 174.275 ;
        RECT 24.930 174.075 32.060 174.215 ;
        RECT 35.510 174.215 35.650 174.370 ;
        RECT 42.780 174.355 43.100 174.415 ;
        RECT 45.540 174.355 45.860 174.415 ;
        RECT 48.760 174.555 49.080 174.615 ;
        RECT 53.775 174.600 54.065 174.915 ;
        RECT 54.855 174.895 55.145 174.940 ;
        RECT 58.435 174.895 58.725 174.940 ;
        RECT 60.270 174.895 60.560 174.940 ;
        RECT 54.855 174.755 60.560 174.895 ;
        RECT 54.855 174.710 55.145 174.755 ;
        RECT 58.435 174.710 58.725 174.755 ;
        RECT 60.270 174.710 60.560 174.755 ;
        RECT 61.180 174.895 61.500 174.955 ;
        RECT 63.495 174.895 63.785 174.940 ;
        RECT 64.400 174.895 64.720 174.955 ;
        RECT 61.180 174.755 64.720 174.895 ;
        RECT 61.180 174.695 61.500 174.755 ;
        RECT 63.495 174.710 63.785 174.755 ;
        RECT 64.400 174.695 64.720 174.755 ;
        RECT 66.240 174.695 66.560 174.955 ;
        RECT 66.715 174.895 67.005 174.940 ;
        RECT 67.620 174.895 67.940 174.955 ;
        RECT 68.095 174.895 68.385 174.940 ;
        RECT 66.715 174.755 67.390 174.895 ;
        RECT 66.715 174.710 67.005 174.755 ;
        RECT 49.695 174.555 49.985 174.600 ;
        RECT 48.760 174.415 49.985 174.555 ;
        RECT 48.760 174.355 49.080 174.415 ;
        RECT 49.695 174.370 49.985 174.415 ;
        RECT 53.475 174.555 54.065 174.600 ;
        RECT 55.660 174.555 55.980 174.615 ;
        RECT 56.715 174.555 57.365 174.600 ;
        RECT 53.475 174.415 57.365 174.555 ;
        RECT 53.475 174.370 53.765 174.415 ;
        RECT 55.660 174.355 55.980 174.415 ;
        RECT 56.715 174.370 57.365 174.415 ;
        RECT 59.340 174.355 59.660 174.615 ;
        RECT 64.490 174.555 64.630 174.695 ;
        RECT 67.250 174.555 67.390 174.755 ;
        RECT 67.620 174.755 68.385 174.895 ;
        RECT 67.620 174.695 67.940 174.755 ;
        RECT 68.095 174.710 68.385 174.755 ;
        RECT 68.555 174.895 68.845 174.940 ;
        RECT 69.460 174.895 69.780 174.955 ;
        RECT 68.555 174.755 69.780 174.895 ;
        RECT 68.555 174.710 68.845 174.755 ;
        RECT 69.460 174.695 69.780 174.755 ;
        RECT 70.840 174.695 71.160 174.955 ;
        RECT 71.300 174.695 71.620 174.955 ;
        RECT 71.760 174.695 72.080 174.955 ;
        RECT 72.695 174.895 72.985 174.940 ;
        RECT 72.585 174.755 72.985 174.895 ;
        RECT 73.230 174.895 73.370 175.035 ;
        RECT 74.435 174.895 74.725 174.940 ;
        RECT 73.230 174.755 74.725 174.895 ;
        RECT 72.695 174.710 72.985 174.755 ;
        RECT 74.435 174.710 74.725 174.755 ;
        RECT 72.770 174.555 72.910 174.710 ;
        RECT 74.980 174.695 75.300 174.955 ;
        RECT 75.440 174.695 75.760 174.955 ;
        RECT 76.360 174.940 76.680 174.955 ;
        RECT 78.290 174.940 78.430 175.775 ;
        RECT 98.070 175.775 99.130 175.915 ;
        RECT 81.880 175.235 82.200 175.295 ;
        RECT 92.460 175.235 92.780 175.295 ;
        RECT 79.210 175.095 92.780 175.235 ;
        RECT 76.345 174.895 76.680 174.940 ;
        RECT 75.925 174.755 76.680 174.895 ;
        RECT 76.345 174.710 76.680 174.755 ;
        RECT 78.215 174.710 78.505 174.940 ;
        RECT 76.360 174.695 76.680 174.710 ;
        RECT 78.660 174.695 78.980 174.955 ;
        RECT 79.210 174.940 79.350 175.095 ;
        RECT 81.880 175.035 82.200 175.095 ;
        RECT 92.460 175.035 92.780 175.095 ;
        RECT 94.300 175.235 94.620 175.295 ;
        RECT 97.520 175.235 97.840 175.295 ;
        RECT 94.300 175.095 97.840 175.235 ;
        RECT 94.300 175.035 94.620 175.095 ;
        RECT 79.135 174.710 79.425 174.940 ;
        RECT 80.055 174.710 80.345 174.940 ;
        RECT 84.180 174.895 84.500 174.955 ;
        RECT 87.875 174.895 88.165 174.940 ;
        RECT 84.180 174.755 88.165 174.895 ;
        RECT 76.450 174.555 76.590 174.695 ;
        RECT 80.130 174.555 80.270 174.710 ;
        RECT 84.180 174.695 84.500 174.755 ;
        RECT 87.875 174.710 88.165 174.755 ;
        RECT 91.095 174.895 91.385 174.940 ;
        RECT 93.840 174.895 94.160 174.955 ;
        RECT 97.150 174.940 97.290 175.095 ;
        RECT 97.520 175.035 97.840 175.095 ;
        RECT 98.070 174.940 98.210 175.775 ;
        RECT 98.990 175.575 99.130 175.775 ;
        RECT 103.500 175.575 103.820 175.635 ;
        RECT 98.990 175.435 103.820 175.575 ;
        RECT 103.500 175.375 103.820 175.435 ;
        RECT 107.295 175.575 107.585 175.620 ;
        RECT 110.415 175.575 110.705 175.620 ;
        RECT 112.305 175.575 112.595 175.620 ;
        RECT 107.295 175.435 112.595 175.575 ;
        RECT 107.295 175.390 107.585 175.435 ;
        RECT 110.415 175.390 110.705 175.435 ;
        RECT 112.305 175.390 112.595 175.435 ;
        RECT 100.280 175.235 100.600 175.295 ;
        RECT 98.530 175.095 100.600 175.235 ;
        RECT 98.530 174.940 98.670 175.095 ;
        RECT 100.280 175.035 100.600 175.095 ;
        RECT 104.435 175.050 104.725 175.280 ;
        RECT 91.095 174.755 94.160 174.895 ;
        RECT 91.095 174.710 91.385 174.755 ;
        RECT 64.490 174.415 67.390 174.555 ;
        RECT 69.090 174.415 80.270 174.555 ;
        RECT 87.950 174.555 88.090 174.710 ;
        RECT 93.840 174.695 94.160 174.755 ;
        RECT 95.695 174.710 95.985 174.940 ;
        RECT 97.075 174.710 97.365 174.940 ;
        RECT 97.995 174.710 98.285 174.940 ;
        RECT 98.455 174.710 98.745 174.940 ;
        RECT 95.770 174.555 95.910 174.710 ;
        RECT 98.900 174.695 99.220 174.955 ;
        RECT 99.820 174.895 100.140 174.955 ;
        RECT 101.215 174.895 101.505 174.940 ;
        RECT 104.510 174.895 104.650 175.050 ;
        RECT 113.160 175.035 113.480 175.295 ;
        RECT 99.820 174.755 104.650 174.895 ;
        RECT 99.820 174.695 100.140 174.755 ;
        RECT 101.215 174.710 101.505 174.755 ;
        RECT 106.215 174.600 106.505 174.915 ;
        RECT 107.295 174.895 107.585 174.940 ;
        RECT 110.875 174.895 111.165 174.940 ;
        RECT 112.710 174.895 113.000 174.940 ;
        RECT 107.295 174.755 113.000 174.895 ;
        RECT 107.295 174.710 107.585 174.755 ;
        RECT 110.875 174.710 111.165 174.755 ;
        RECT 112.710 174.710 113.000 174.755 ;
        RECT 87.950 174.415 95.910 174.555 ;
        RECT 38.655 174.215 38.945 174.260 ;
        RECT 35.510 174.075 38.945 174.215 ;
        RECT 22.080 174.015 22.400 174.075 ;
        RECT 23.935 174.030 24.225 174.075 ;
        RECT 28.075 174.030 28.365 174.075 ;
        RECT 31.740 174.015 32.060 174.075 ;
        RECT 38.655 174.030 38.945 174.075 ;
        RECT 43.700 174.015 44.020 174.275 ;
        RECT 51.520 174.015 51.840 174.275 ;
        RECT 65.320 174.215 65.640 174.275 ;
        RECT 69.090 174.215 69.230 174.415 ;
        RECT 65.320 174.075 69.230 174.215 ;
        RECT 69.475 174.215 69.765 174.260 ;
        RECT 69.920 174.215 70.240 174.275 ;
        RECT 69.475 174.075 70.240 174.215 ;
        RECT 65.320 174.015 65.640 174.075 ;
        RECT 69.475 174.030 69.765 174.075 ;
        RECT 69.920 174.015 70.240 174.075 ;
        RECT 73.140 174.015 73.460 174.275 ;
        RECT 75.900 174.215 76.220 174.275 ;
        RECT 76.835 174.215 77.125 174.260 ;
        RECT 75.900 174.075 77.125 174.215 ;
        RECT 75.900 174.015 76.220 174.075 ;
        RECT 76.835 174.030 77.125 174.075 ;
        RECT 88.320 174.015 88.640 174.275 ;
        RECT 92.460 174.215 92.780 174.275 ;
        RECT 93.855 174.215 94.145 174.260 ;
        RECT 92.460 174.075 94.145 174.215 ;
        RECT 95.770 174.215 95.910 174.415 ;
        RECT 96.155 174.555 96.445 174.600 ;
        RECT 105.915 174.555 106.505 174.600 ;
        RECT 109.155 174.555 109.805 174.600 ;
        RECT 96.155 174.415 109.805 174.555 ;
        RECT 96.155 174.370 96.445 174.415 ;
        RECT 105.915 174.370 106.205 174.415 ;
        RECT 109.155 174.370 109.805 174.415 ;
        RECT 111.795 174.555 112.085 174.600 ;
        RECT 111.795 174.415 112.930 174.555 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 111.795 174.370 112.085 174.415 ;
        RECT 112.790 174.275 112.930 174.415 ;
        RECT 97.060 174.215 97.380 174.275 ;
        RECT 95.770 174.075 97.380 174.215 ;
        RECT 92.460 174.015 92.780 174.075 ;
        RECT 93.855 174.030 94.145 174.075 ;
        RECT 97.060 174.015 97.380 174.075 ;
        RECT 100.295 174.215 100.585 174.260 ;
        RECT 102.580 174.215 102.900 174.275 ;
        RECT 100.295 174.075 102.900 174.215 ;
        RECT 100.295 174.030 100.585 174.075 ;
        RECT 102.580 174.015 102.900 174.075 ;
        RECT 103.960 174.015 104.280 174.275 ;
        RECT 112.700 174.015 113.020 174.275 ;
        RECT 14.650 173.395 115.850 173.875 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 34.040 173.195 34.360 173.255 ;
        RECT 28.150 173.055 34.360 173.195 ;
        RECT 20.700 172.855 21.020 172.915 ;
        RECT 20.700 172.715 27.370 172.855 ;
        RECT 20.700 172.655 21.020 172.715 ;
        RECT 26.680 172.315 27.000 172.575 ;
        RECT 27.230 172.560 27.370 172.715 ;
        RECT 27.155 172.515 27.445 172.560 ;
        RECT 27.600 172.515 27.920 172.575 ;
        RECT 28.150 172.560 28.290 173.055 ;
        RECT 34.040 172.995 34.360 173.055 ;
        RECT 43.240 173.195 43.560 173.255 ;
        RECT 46.920 173.195 47.240 173.255 ;
        RECT 50.600 173.195 50.920 173.255 ;
        RECT 43.240 173.055 50.920 173.195 ;
        RECT 43.240 172.995 43.560 173.055 ;
        RECT 46.920 172.995 47.240 173.055 ;
        RECT 50.600 172.995 50.920 173.055 ;
        RECT 55.660 172.995 55.980 173.255 ;
        RECT 57.975 173.195 58.265 173.240 ;
        RECT 59.340 173.195 59.660 173.255 ;
        RECT 57.975 173.055 59.660 173.195 ;
        RECT 57.975 173.010 58.265 173.055 ;
        RECT 59.340 172.995 59.660 173.055 ;
        RECT 63.020 173.195 63.340 173.255 ;
        RECT 91.540 173.195 91.860 173.255 ;
        RECT 63.020 173.055 91.860 173.195 ;
        RECT 63.020 172.995 63.340 173.055 ;
        RECT 91.540 172.995 91.860 173.055 ;
        RECT 92.460 173.195 92.780 173.255 ;
        RECT 92.460 173.055 95.450 173.195 ;
        RECT 92.460 172.995 92.780 173.055 ;
        RECT 33.580 172.855 33.900 172.915 ;
        RECT 42.780 172.855 43.100 172.915 ;
        RECT 47.840 172.855 48.160 172.915 ;
        RECT 50.140 172.855 50.460 172.915 ;
        RECT 29.070 172.715 32.890 172.855 ;
        RECT 29.070 172.560 29.210 172.715 ;
        RECT 32.750 172.575 32.890 172.715 ;
        RECT 33.580 172.715 35.650 172.855 ;
        RECT 33.580 172.655 33.900 172.715 ;
        RECT 27.155 172.375 27.920 172.515 ;
        RECT 27.155 172.330 27.445 172.375 ;
        RECT 27.600 172.315 27.920 172.375 ;
        RECT 28.075 172.330 28.365 172.560 ;
        RECT 28.535 172.330 28.825 172.560 ;
        RECT 28.995 172.330 29.285 172.560 ;
        RECT 30.835 172.515 31.125 172.560 ;
        RECT 31.280 172.515 31.600 172.575 ;
        RECT 30.835 172.375 31.600 172.515 ;
        RECT 30.835 172.330 31.125 172.375 ;
        RECT 23.460 171.975 23.780 172.235 ;
        RECT 24.380 172.175 24.700 172.235 ;
        RECT 28.610 172.175 28.750 172.330 ;
        RECT 31.280 172.315 31.600 172.375 ;
        RECT 31.740 172.315 32.060 172.575 ;
        RECT 32.200 172.315 32.520 172.575 ;
        RECT 32.660 172.315 32.980 172.575 ;
        RECT 34.500 172.315 34.820 172.575 ;
        RECT 35.510 172.560 35.650 172.715 ;
        RECT 35.970 172.715 43.100 172.855 ;
        RECT 35.970 172.560 36.110 172.715 ;
        RECT 42.780 172.655 43.100 172.715 ;
        RECT 46.090 172.715 48.160 172.855 ;
        RECT 35.435 172.330 35.725 172.560 ;
        RECT 35.895 172.330 36.185 172.560 ;
        RECT 36.355 172.515 36.645 172.560 ;
        RECT 45.095 172.515 45.385 172.560 ;
        RECT 36.355 172.375 45.385 172.515 ;
        RECT 36.355 172.330 36.645 172.375 ;
        RECT 45.095 172.330 45.385 172.375 ;
        RECT 32.290 172.175 32.430 172.315 ;
        RECT 24.380 172.035 32.430 172.175 ;
        RECT 34.960 172.175 35.280 172.235 ;
        RECT 38.195 172.175 38.485 172.220 ;
        RECT 34.960 172.035 38.485 172.175 ;
        RECT 24.380 171.975 24.700 172.035 ;
        RECT 34.960 171.975 35.280 172.035 ;
        RECT 38.195 171.990 38.485 172.035 ;
        RECT 27.600 171.835 27.920 171.895 ;
        RECT 31.280 171.835 31.600 171.895 ;
        RECT 27.600 171.695 31.600 171.835 ;
        RECT 27.600 171.635 27.920 171.695 ;
        RECT 31.280 171.635 31.600 171.695 ;
        RECT 18.860 171.495 19.180 171.555 ;
        RECT 20.255 171.495 20.545 171.540 ;
        RECT 18.860 171.355 20.545 171.495 ;
        RECT 18.860 171.295 19.180 171.355 ;
        RECT 20.255 171.310 20.545 171.355 ;
        RECT 26.235 171.495 26.525 171.540 ;
        RECT 26.680 171.495 27.000 171.555 ;
        RECT 26.235 171.355 27.000 171.495 ;
        RECT 26.235 171.310 26.525 171.355 ;
        RECT 26.680 171.295 27.000 171.355 ;
        RECT 29.440 171.495 29.760 171.555 ;
        RECT 30.375 171.495 30.665 171.540 ;
        RECT 29.440 171.355 30.665 171.495 ;
        RECT 29.440 171.295 29.760 171.355 ;
        RECT 30.375 171.310 30.665 171.355 ;
        RECT 34.040 171.295 34.360 171.555 ;
        RECT 37.735 171.495 38.025 171.540 ;
        RECT 38.180 171.495 38.500 171.555 ;
        RECT 37.735 171.355 38.500 171.495 ;
        RECT 37.735 171.310 38.025 171.355 ;
        RECT 38.180 171.295 38.500 171.355 ;
        RECT 40.480 171.495 40.800 171.555 ;
        RECT 41.415 171.495 41.705 171.540 ;
        RECT 40.480 171.355 41.705 171.495 ;
        RECT 40.480 171.295 40.800 171.355 ;
        RECT 41.415 171.310 41.705 171.355 ;
        RECT 43.715 171.495 44.005 171.540 ;
        RECT 44.620 171.495 44.940 171.555 ;
        RECT 43.715 171.355 44.940 171.495 ;
        RECT 45.170 171.495 45.310 172.330 ;
        RECT 45.540 172.315 45.860 172.575 ;
        RECT 46.090 172.560 46.230 172.715 ;
        RECT 47.840 172.655 48.160 172.715 ;
        RECT 48.850 172.715 50.460 172.855 ;
        RECT 46.015 172.330 46.305 172.560 ;
        RECT 46.920 172.315 47.240 172.575 ;
        RECT 48.850 172.560 48.990 172.715 ;
        RECT 50.140 172.655 50.460 172.715 ;
        RECT 48.775 172.330 49.065 172.560 ;
        RECT 45.630 171.835 45.770 172.315 ;
        RECT 46.460 172.175 46.780 172.235 ;
        RECT 48.850 172.175 48.990 172.330 ;
        RECT 49.220 172.315 49.540 172.575 ;
        RECT 49.680 172.315 50.000 172.575 ;
        RECT 50.690 172.560 50.830 172.995 ;
        RECT 51.520 172.855 51.840 172.915 ;
        RECT 73.600 172.855 73.920 172.915 ;
        RECT 79.530 172.855 79.820 172.900 ;
        RECT 82.790 172.855 83.080 172.900 ;
        RECT 51.520 172.715 57.270 172.855 ;
        RECT 51.520 172.655 51.840 172.715 ;
        RECT 50.615 172.330 50.905 172.560 ;
        RECT 56.120 172.315 56.440 172.575 ;
        RECT 57.130 172.560 57.270 172.715 ;
        RECT 73.600 172.715 83.080 172.855 ;
        RECT 73.600 172.655 73.920 172.715 ;
        RECT 79.530 172.670 79.820 172.715 ;
        RECT 82.790 172.670 83.080 172.715 ;
        RECT 83.710 172.855 84.000 172.900 ;
        RECT 85.570 172.855 85.860 172.900 ;
        RECT 87.860 172.855 88.180 172.915 ;
        RECT 83.710 172.715 85.860 172.855 ;
        RECT 83.710 172.670 84.000 172.715 ;
        RECT 85.570 172.670 85.860 172.715 ;
        RECT 86.110 172.715 88.180 172.855 ;
        RECT 57.055 172.330 57.345 172.560 ;
        RECT 63.940 172.315 64.260 172.575 ;
        RECT 64.400 172.315 64.720 172.575 ;
        RECT 81.390 172.515 81.680 172.560 ;
        RECT 83.710 172.515 83.925 172.670 ;
        RECT 86.110 172.515 86.250 172.715 ;
        RECT 87.860 172.655 88.180 172.715 ;
        RECT 88.320 172.855 88.640 172.915 ;
        RECT 90.615 172.855 91.265 172.900 ;
        RECT 94.215 172.855 94.505 172.900 ;
        RECT 88.320 172.715 94.505 172.855 ;
        RECT 95.310 172.855 95.450 173.055 ;
        RECT 100.295 172.855 100.585 172.900 ;
        RECT 95.310 172.715 100.585 172.855 ;
        RECT 88.320 172.655 88.640 172.715 ;
        RECT 90.615 172.670 91.265 172.715 ;
        RECT 93.915 172.670 94.505 172.715 ;
        RECT 100.295 172.670 100.585 172.715 ;
        RECT 103.515 172.855 103.805 172.900 ;
        RECT 105.915 172.855 106.205 172.900 ;
        RECT 109.155 172.855 109.805 172.900 ;
        RECT 103.515 172.715 109.805 172.855 ;
        RECT 103.515 172.670 103.805 172.715 ;
        RECT 105.915 172.670 106.505 172.715 ;
        RECT 109.155 172.670 109.805 172.715 ;
        RECT 111.795 172.855 112.085 172.900 ;
        RECT 112.240 172.855 112.560 172.915 ;
        RECT 111.795 172.715 112.560 172.855 ;
        RECT 111.795 172.670 112.085 172.715 ;
        RECT 81.390 172.375 83.925 172.515 ;
        RECT 84.270 172.375 86.250 172.515 ;
        RECT 86.480 172.515 86.800 172.575 ;
        RECT 86.955 172.515 87.245 172.560 ;
        RECT 86.480 172.375 87.245 172.515 ;
        RECT 81.390 172.330 81.680 172.375 ;
        RECT 46.460 172.035 48.990 172.175 ;
        RECT 46.460 171.975 46.780 172.035 ;
        RECT 49.310 171.835 49.450 172.315 ;
        RECT 56.210 172.175 56.350 172.315 ;
        RECT 62.100 172.175 62.420 172.235 ;
        RECT 84.270 172.175 84.410 172.375 ;
        RECT 86.480 172.315 86.800 172.375 ;
        RECT 86.955 172.330 87.245 172.375 ;
        RECT 87.420 172.515 87.710 172.560 ;
        RECT 89.255 172.515 89.545 172.560 ;
        RECT 92.835 172.515 93.125 172.560 ;
        RECT 87.420 172.375 93.125 172.515 ;
        RECT 87.420 172.330 87.710 172.375 ;
        RECT 89.255 172.330 89.545 172.375 ;
        RECT 92.835 172.330 93.125 172.375 ;
        RECT 93.915 172.355 94.205 172.670 ;
        RECT 97.060 172.515 97.380 172.575 ;
        RECT 101.660 172.515 101.980 172.575 ;
        RECT 103.055 172.515 103.345 172.560 ;
        RECT 97.060 172.375 103.345 172.515 ;
        RECT 97.060 172.315 97.380 172.375 ;
        RECT 101.660 172.315 101.980 172.375 ;
        RECT 103.055 172.330 103.345 172.375 ;
        RECT 106.215 172.355 106.505 172.670 ;
        RECT 112.240 172.655 112.560 172.715 ;
        RECT 107.295 172.515 107.585 172.560 ;
        RECT 110.875 172.515 111.165 172.560 ;
        RECT 112.710 172.515 113.000 172.560 ;
        RECT 107.295 172.375 113.000 172.515 ;
        RECT 107.295 172.330 107.585 172.375 ;
        RECT 110.875 172.330 111.165 172.375 ;
        RECT 112.710 172.330 113.000 172.375 ;
        RECT 113.160 172.315 113.480 172.575 ;
        RECT 56.210 172.035 62.420 172.175 ;
        RECT 62.100 171.975 62.420 172.035 ;
        RECT 65.410 172.035 84.410 172.175 ;
        RECT 45.630 171.695 49.450 171.835 ;
        RECT 57.960 171.835 58.280 171.895 ;
        RECT 65.410 171.880 65.550 172.035 ;
        RECT 84.640 171.975 84.960 172.235 ;
        RECT 88.320 171.975 88.640 172.235 ;
        RECT 93.380 172.175 93.700 172.235 ;
        RECT 98.915 172.175 99.205 172.220 ;
        RECT 93.380 172.035 99.205 172.175 ;
        RECT 93.380 171.975 93.700 172.035 ;
        RECT 98.915 171.990 99.205 172.035 ;
        RECT 99.835 172.175 100.125 172.220 ;
        RECT 103.960 172.175 104.280 172.235 ;
        RECT 99.835 172.035 104.280 172.175 ;
        RECT 99.835 171.990 100.125 172.035 ;
        RECT 103.960 171.975 104.280 172.035 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 65.335 171.835 65.625 171.880 ;
        RECT 57.960 171.695 65.625 171.835 ;
        RECT 57.960 171.635 58.280 171.695 ;
        RECT 65.335 171.650 65.625 171.695 ;
        RECT 74.060 171.835 74.380 171.895 ;
        RECT 77.525 171.835 77.815 171.880 ;
        RECT 78.200 171.835 78.520 171.895 ;
        RECT 74.060 171.695 78.520 171.835 ;
        RECT 74.060 171.635 74.380 171.695 ;
        RECT 77.525 171.650 77.815 171.695 ;
        RECT 78.200 171.635 78.520 171.695 ;
        RECT 81.390 171.835 81.680 171.880 ;
        RECT 84.170 171.835 84.460 171.880 ;
        RECT 86.030 171.835 86.320 171.880 ;
        RECT 81.390 171.695 86.320 171.835 ;
        RECT 81.390 171.650 81.680 171.695 ;
        RECT 84.170 171.650 84.460 171.695 ;
        RECT 86.030 171.650 86.320 171.695 ;
        RECT 87.825 171.835 88.115 171.880 ;
        RECT 89.715 171.835 90.005 171.880 ;
        RECT 92.835 171.835 93.125 171.880 ;
        RECT 87.825 171.695 93.125 171.835 ;
        RECT 87.825 171.650 88.115 171.695 ;
        RECT 89.715 171.650 90.005 171.695 ;
        RECT 92.835 171.650 93.125 171.695 ;
        RECT 104.435 171.835 104.725 171.880 ;
        RECT 105.800 171.835 106.120 171.895 ;
        RECT 104.435 171.695 106.120 171.835 ;
        RECT 104.435 171.650 104.725 171.695 ;
        RECT 105.800 171.635 106.120 171.695 ;
        RECT 107.295 171.835 107.585 171.880 ;
        RECT 110.415 171.835 110.705 171.880 ;
        RECT 112.305 171.835 112.595 171.880 ;
        RECT 107.295 171.695 112.595 171.835 ;
        RECT 107.295 171.650 107.585 171.695 ;
        RECT 110.415 171.650 110.705 171.695 ;
        RECT 112.305 171.650 112.595 171.695 ;
        RECT 46.460 171.495 46.780 171.555 ;
        RECT 45.170 171.355 46.780 171.495 ;
        RECT 43.715 171.310 44.005 171.355 ;
        RECT 44.620 171.295 44.940 171.355 ;
        RECT 46.460 171.295 46.780 171.355 ;
        RECT 47.380 171.295 47.700 171.555 ;
        RECT 71.300 171.495 71.620 171.555 ;
        RECT 74.980 171.495 75.300 171.555 ;
        RECT 78.660 171.495 78.980 171.555 ;
        RECT 71.300 171.355 78.980 171.495 ;
        RECT 71.300 171.295 71.620 171.355 ;
        RECT 74.980 171.295 75.300 171.355 ;
        RECT 78.660 171.295 78.980 171.355 ;
        RECT 93.840 171.495 94.160 171.555 ;
        RECT 95.695 171.495 95.985 171.540 ;
        RECT 97.060 171.495 97.380 171.555 ;
        RECT 93.840 171.355 97.380 171.495 ;
        RECT 93.840 171.295 94.160 171.355 ;
        RECT 95.695 171.310 95.985 171.355 ;
        RECT 97.060 171.295 97.380 171.355 ;
        RECT 97.535 171.495 97.825 171.540 ;
        RECT 98.900 171.495 99.220 171.555 ;
        RECT 97.535 171.355 99.220 171.495 ;
        RECT 97.535 171.310 97.825 171.355 ;
        RECT 98.900 171.295 99.220 171.355 ;
        RECT 102.135 171.495 102.425 171.540 ;
        RECT 114.080 171.495 114.400 171.555 ;
        RECT 102.135 171.355 114.400 171.495 ;
        RECT 102.135 171.310 102.425 171.355 ;
        RECT 114.080 171.295 114.400 171.355 ;
        RECT 14.650 170.675 115.850 171.155 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 27.140 170.475 27.460 170.535 ;
        RECT 34.500 170.475 34.820 170.535 ;
        RECT 60.260 170.475 60.580 170.535 ;
        RECT 64.875 170.475 65.165 170.520 ;
        RECT 82.815 170.475 83.105 170.520 ;
        RECT 84.640 170.475 84.960 170.535 ;
        RECT 17.570 170.335 32.430 170.475 ;
        RECT 17.570 169.500 17.710 170.335 ;
        RECT 27.140 170.275 27.460 170.335 ;
        RECT 23.000 170.135 23.320 170.195 ;
        RECT 19.870 169.995 23.320 170.135 ;
        RECT 19.870 169.840 20.010 169.995 ;
        RECT 23.000 169.935 23.320 169.995 ;
        RECT 25.875 170.135 26.165 170.180 ;
        RECT 28.995 170.135 29.285 170.180 ;
        RECT 30.885 170.135 31.175 170.180 ;
        RECT 25.875 169.995 31.175 170.135 ;
        RECT 25.875 169.950 26.165 169.995 ;
        RECT 28.995 169.950 29.285 169.995 ;
        RECT 30.885 169.950 31.175 169.995 ;
        RECT 32.290 170.135 32.430 170.335 ;
        RECT 34.500 170.335 65.165 170.475 ;
        RECT 34.500 170.275 34.820 170.335 ;
        RECT 60.260 170.275 60.580 170.335 ;
        RECT 64.875 170.290 65.165 170.335 ;
        RECT 75.990 170.335 82.570 170.475 ;
        RECT 33.120 170.135 33.440 170.195 ;
        RECT 44.160 170.135 44.480 170.195 ;
        RECT 32.290 169.995 44.480 170.135 ;
        RECT 19.795 169.610 20.085 169.840 ;
        RECT 22.555 169.795 22.845 169.840 ;
        RECT 24.380 169.795 24.700 169.855 ;
        RECT 22.555 169.655 24.700 169.795 ;
        RECT 22.555 169.610 22.845 169.655 ;
        RECT 24.380 169.595 24.700 169.655 ;
        RECT 17.495 169.270 17.785 169.500 ;
        RECT 18.860 169.255 19.180 169.515 ;
        RECT 17.020 168.915 17.340 169.175 ;
        RECT 24.795 169.160 25.085 169.475 ;
        RECT 25.875 169.455 26.165 169.500 ;
        RECT 29.455 169.455 29.745 169.500 ;
        RECT 31.290 169.455 31.580 169.500 ;
        RECT 25.875 169.315 31.580 169.455 ;
        RECT 25.875 169.270 26.165 169.315 ;
        RECT 29.455 169.270 29.745 169.315 ;
        RECT 31.290 169.270 31.580 169.315 ;
        RECT 31.755 169.270 32.045 169.500 ;
        RECT 32.290 169.455 32.430 169.995 ;
        RECT 33.120 169.935 33.440 169.995 ;
        RECT 44.160 169.935 44.480 169.995 ;
        RECT 44.735 170.135 45.025 170.180 ;
        RECT 47.855 170.135 48.145 170.180 ;
        RECT 49.745 170.135 50.035 170.180 ;
        RECT 57.960 170.135 58.280 170.195 ;
        RECT 75.990 170.135 76.130 170.335 ;
        RECT 44.735 169.995 50.035 170.135 ;
        RECT 44.735 169.950 45.025 169.995 ;
        RECT 47.855 169.950 48.145 169.995 ;
        RECT 49.745 169.950 50.035 169.995 ;
        RECT 50.230 169.995 58.280 170.135 ;
        RECT 32.660 169.795 32.980 169.855 ;
        RECT 50.230 169.795 50.370 169.995 ;
        RECT 57.960 169.935 58.280 169.995 ;
        RECT 64.490 169.995 76.130 170.135 ;
        RECT 76.330 170.135 76.620 170.180 ;
        RECT 79.110 170.135 79.400 170.180 ;
        RECT 80.970 170.135 81.260 170.180 ;
        RECT 76.330 169.995 81.260 170.135 ;
        RECT 82.430 170.135 82.570 170.335 ;
        RECT 82.815 170.335 84.960 170.475 ;
        RECT 82.815 170.290 83.105 170.335 ;
        RECT 84.640 170.275 84.960 170.335 ;
        RECT 88.320 170.275 88.640 170.535 ;
        RECT 93.840 170.475 94.160 170.535 ;
        RECT 89.790 170.335 94.160 170.475 ;
        RECT 89.790 170.135 89.930 170.335 ;
        RECT 93.840 170.275 94.160 170.335 ;
        RECT 109.020 170.475 109.340 170.535 ;
        RECT 110.875 170.475 111.165 170.520 ;
        RECT 109.020 170.335 111.165 170.475 ;
        RECT 109.020 170.275 109.340 170.335 ;
        RECT 110.875 170.290 111.165 170.335 ;
        RECT 112.700 170.475 113.020 170.535 ;
        RECT 113.175 170.475 113.465 170.520 ;
        RECT 112.700 170.335 113.465 170.475 ;
        RECT 112.700 170.275 113.020 170.335 ;
        RECT 113.175 170.290 113.465 170.335 ;
        RECT 82.430 169.995 89.930 170.135 ;
        RECT 64.490 169.855 64.630 169.995 ;
        RECT 76.330 169.950 76.620 169.995 ;
        RECT 79.110 169.950 79.400 169.995 ;
        RECT 80.970 169.950 81.260 169.995 ;
        RECT 90.175 169.950 90.465 170.180 ;
        RECT 91.080 170.135 91.400 170.195 ;
        RECT 94.315 170.135 94.605 170.180 ;
        RECT 91.080 169.995 94.605 170.135 ;
        RECT 64.400 169.795 64.720 169.855 ;
        RECT 32.660 169.655 50.370 169.795 ;
        RECT 55.750 169.655 64.720 169.795 ;
        RECT 32.660 169.595 32.980 169.655 ;
        RECT 33.135 169.455 33.425 169.500 ;
        RECT 32.290 169.315 33.425 169.455 ;
        RECT 33.135 169.270 33.425 169.315 ;
        RECT 34.975 169.455 35.265 169.500 ;
        RECT 37.260 169.455 37.580 169.515 ;
        RECT 34.975 169.315 37.580 169.455 ;
        RECT 34.975 169.270 35.265 169.315 ;
        RECT 24.495 169.115 25.085 169.160 ;
        RECT 26.680 169.115 27.000 169.175 ;
        RECT 27.735 169.115 28.385 169.160 ;
        RECT 24.495 168.975 28.385 169.115 ;
        RECT 24.495 168.930 24.785 168.975 ;
        RECT 26.680 168.915 27.000 168.975 ;
        RECT 27.735 168.930 28.385 168.975 ;
        RECT 29.900 169.115 30.220 169.175 ;
        RECT 30.375 169.115 30.665 169.160 ;
        RECT 29.900 168.975 30.665 169.115 ;
        RECT 29.900 168.915 30.220 168.975 ;
        RECT 30.375 168.930 30.665 168.975 ;
        RECT 30.820 169.115 31.140 169.175 ;
        RECT 31.830 169.115 31.970 169.270 ;
        RECT 37.260 169.255 37.580 169.315 ;
        RECT 30.820 168.975 31.970 169.115 ;
        RECT 30.820 168.915 31.140 168.975 ;
        RECT 33.580 168.915 33.900 169.175 ;
        RECT 37.720 168.915 38.040 169.175 ;
        RECT 43.655 169.160 43.945 169.475 ;
        RECT 44.735 169.455 45.025 169.500 ;
        RECT 48.315 169.455 48.605 169.500 ;
        RECT 50.150 169.455 50.440 169.500 ;
        RECT 44.735 169.315 50.440 169.455 ;
        RECT 44.735 169.270 45.025 169.315 ;
        RECT 48.315 169.270 48.605 169.315 ;
        RECT 50.150 169.270 50.440 169.315 ;
        RECT 50.600 169.255 50.920 169.515 ;
        RECT 51.060 169.455 51.380 169.515 ;
        RECT 51.995 169.455 52.285 169.500 ;
        RECT 52.455 169.455 52.745 169.500 ;
        RECT 54.755 169.455 55.045 169.500 ;
        RECT 51.060 169.315 55.045 169.455 ;
        RECT 51.060 169.255 51.380 169.315 ;
        RECT 51.995 169.270 52.285 169.315 ;
        RECT 52.455 169.270 52.745 169.315 ;
        RECT 54.755 169.270 55.045 169.315 ;
        RECT 43.355 169.115 43.945 169.160 ;
        RECT 46.595 169.115 47.245 169.160 ;
        RECT 43.355 168.975 47.610 169.115 ;
        RECT 43.355 168.930 43.645 168.975 ;
        RECT 46.595 168.930 47.245 168.975 ;
        RECT 17.940 168.575 18.260 168.835 ;
        RECT 31.280 168.775 31.600 168.835 ;
        RECT 33.120 168.775 33.440 168.835 ;
        RECT 39.560 168.775 39.880 168.835 ;
        RECT 31.280 168.635 39.880 168.775 ;
        RECT 31.280 168.575 31.600 168.635 ;
        RECT 33.120 168.575 33.440 168.635 ;
        RECT 39.560 168.575 39.880 168.635 ;
        RECT 41.860 168.575 42.180 168.835 ;
        RECT 47.470 168.775 47.610 168.975 ;
        RECT 49.220 168.915 49.540 169.175 ;
        RECT 51.535 169.115 51.825 169.160 ;
        RECT 51.150 168.975 51.825 169.115 ;
        RECT 51.150 168.775 51.290 168.975 ;
        RECT 51.535 168.930 51.825 168.975 ;
        RECT 52.915 169.115 53.205 169.160 ;
        RECT 53.360 169.115 53.680 169.175 ;
        RECT 52.915 168.975 53.680 169.115 ;
        RECT 52.915 168.930 53.205 168.975 ;
        RECT 53.360 168.915 53.680 168.975 ;
        RECT 47.470 168.635 51.290 168.775 ;
        RECT 51.980 168.775 52.300 168.835 ;
        RECT 55.750 168.775 55.890 169.655 ;
        RECT 64.400 169.595 64.720 169.655 ;
        RECT 68.095 169.795 68.385 169.840 ;
        RECT 73.140 169.795 73.460 169.855 ;
        RECT 68.095 169.655 73.460 169.795 ;
        RECT 68.095 169.610 68.385 169.655 ;
        RECT 73.140 169.595 73.460 169.655 ;
        RECT 78.660 169.795 78.980 169.855 ;
        RECT 79.595 169.795 79.885 169.840 ;
        RECT 78.660 169.655 79.885 169.795 ;
        RECT 78.660 169.595 78.980 169.655 ;
        RECT 79.595 169.610 79.885 169.655 ;
        RECT 81.435 169.795 81.725 169.840 ;
        RECT 86.480 169.795 86.800 169.855 ;
        RECT 81.435 169.655 88.090 169.795 ;
        RECT 81.435 169.610 81.725 169.655 ;
        RECT 86.480 169.595 86.800 169.655 ;
        RECT 56.135 169.455 56.425 169.500 ;
        RECT 65.795 169.455 66.085 169.500 ;
        RECT 69.460 169.455 69.780 169.515 ;
        RECT 56.135 169.315 59.340 169.455 ;
        RECT 56.135 169.270 56.425 169.315 ;
        RECT 51.980 168.635 55.890 168.775 ;
        RECT 59.200 168.775 59.340 169.315 ;
        RECT 65.795 169.315 69.780 169.455 ;
        RECT 65.795 169.270 66.085 169.315 ;
        RECT 69.460 169.255 69.780 169.315 ;
        RECT 76.330 169.455 76.620 169.500 ;
        RECT 79.120 169.455 79.440 169.515 ;
        RECT 87.950 169.500 88.090 169.655 ;
        RECT 81.895 169.455 82.185 169.500 ;
        RECT 76.330 169.315 78.865 169.455 ;
        RECT 76.330 169.270 76.620 169.315 ;
        RECT 66.715 169.115 67.005 169.160 ;
        RECT 67.160 169.115 67.480 169.175 ;
        RECT 66.715 168.975 67.480 169.115 ;
        RECT 66.715 168.930 67.005 168.975 ;
        RECT 67.160 168.915 67.480 168.975 ;
        RECT 71.300 169.115 71.620 169.175 ;
        RECT 77.740 169.160 78.060 169.175 ;
        RECT 72.465 169.115 72.755 169.160 ;
        RECT 71.300 168.975 72.755 169.115 ;
        RECT 71.300 168.915 71.620 168.975 ;
        RECT 72.465 168.930 72.755 168.975 ;
        RECT 74.470 169.115 74.760 169.160 ;
        RECT 77.730 169.115 78.060 169.160 ;
        RECT 74.470 168.975 78.060 169.115 ;
        RECT 74.470 168.930 74.760 168.975 ;
        RECT 77.730 168.930 78.060 168.975 ;
        RECT 78.650 169.160 78.865 169.315 ;
        RECT 79.120 169.315 82.185 169.455 ;
        RECT 79.120 169.255 79.440 169.315 ;
        RECT 81.895 169.270 82.185 169.315 ;
        RECT 87.875 169.270 88.165 169.500 ;
        RECT 89.255 169.455 89.545 169.500 ;
        RECT 90.250 169.455 90.390 169.950 ;
        RECT 91.080 169.935 91.400 169.995 ;
        RECT 94.315 169.950 94.605 169.995 ;
        RECT 102.120 169.935 102.440 170.195 ;
        RECT 107.195 170.135 107.485 170.180 ;
        RECT 107.195 169.995 107.870 170.135 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 107.195 169.950 107.485 169.995 ;
        RECT 92.460 169.595 92.780 169.855 ;
        RECT 93.380 169.795 93.700 169.855 ;
        RECT 97.075 169.795 97.365 169.840 ;
        RECT 98.915 169.795 99.205 169.840 ;
        RECT 104.435 169.795 104.725 169.840 ;
        RECT 104.880 169.795 105.200 169.855 ;
        RECT 107.730 169.840 107.870 169.995 ;
        RECT 93.380 169.655 105.200 169.795 ;
        RECT 93.380 169.595 93.700 169.655 ;
        RECT 97.075 169.610 97.365 169.655 ;
        RECT 98.915 169.610 99.205 169.655 ;
        RECT 104.435 169.610 104.725 169.655 ;
        RECT 104.880 169.595 105.200 169.655 ;
        RECT 107.655 169.610 107.945 169.840 ;
        RECT 96.615 169.455 96.905 169.500 ;
        RECT 89.255 169.315 90.390 169.455 ;
        RECT 92.550 169.315 96.905 169.455 ;
        RECT 89.255 169.270 89.545 169.315 ;
        RECT 92.550 169.175 92.690 169.315 ;
        RECT 96.615 169.270 96.905 169.315 ;
        RECT 103.960 169.455 104.280 169.515 ;
        RECT 105.355 169.455 105.645 169.500 ;
        RECT 103.960 169.315 105.645 169.455 ;
        RECT 103.960 169.255 104.280 169.315 ;
        RECT 105.355 169.270 105.645 169.315 ;
        RECT 114.080 169.255 114.400 169.515 ;
        RECT 78.650 169.115 78.940 169.160 ;
        RECT 80.510 169.115 80.800 169.160 ;
        RECT 92.015 169.115 92.305 169.160 ;
        RECT 78.650 168.975 80.800 169.115 ;
        RECT 78.650 168.930 78.940 168.975 ;
        RECT 80.510 168.930 80.800 168.975 ;
        RECT 81.050 168.975 92.305 169.115 ;
        RECT 77.740 168.915 78.060 168.930 ;
        RECT 62.560 168.775 62.880 168.835 ;
        RECT 59.200 168.635 62.880 168.775 ;
        RECT 51.980 168.575 52.300 168.635 ;
        RECT 62.560 168.575 62.880 168.635 ;
        RECT 78.200 168.775 78.520 168.835 ;
        RECT 81.050 168.775 81.190 168.975 ;
        RECT 92.015 168.930 92.305 168.975 ;
        RECT 92.460 168.915 92.780 169.175 ;
        RECT 94.300 169.115 94.620 169.175 ;
        RECT 96.155 169.115 96.445 169.160 ;
        RECT 99.835 169.115 100.125 169.160 ;
        RECT 94.300 168.975 100.125 169.115 ;
        RECT 94.300 168.915 94.620 168.975 ;
        RECT 96.155 168.930 96.445 168.975 ;
        RECT 99.835 168.930 100.125 168.975 ;
        RECT 100.295 169.115 100.585 169.160 ;
        RECT 104.420 169.115 104.740 169.175 ;
        RECT 100.295 168.975 104.740 169.115 ;
        RECT 100.295 168.930 100.585 168.975 ;
        RECT 104.420 168.915 104.740 168.975 ;
        RECT 104.895 169.115 105.185 169.160 ;
        RECT 105.800 169.115 106.120 169.175 ;
        RECT 104.895 168.975 106.120 169.115 ;
        RECT 104.895 168.930 105.185 168.975 ;
        RECT 105.800 168.915 106.120 168.975 ;
        RECT 108.100 169.115 108.420 169.175 ;
        RECT 111.335 169.115 111.625 169.160 ;
        RECT 108.100 168.975 111.625 169.115 ;
        RECT 108.100 168.915 108.420 168.975 ;
        RECT 111.335 168.930 111.625 168.975 ;
        RECT 112.255 169.115 112.545 169.160 ;
        RECT 116.380 169.115 116.700 169.175 ;
        RECT 112.255 168.975 116.700 169.115 ;
        RECT 112.255 168.930 112.545 168.975 ;
        RECT 116.380 168.915 116.700 168.975 ;
        RECT 78.200 168.635 81.190 168.775 ;
        RECT 78.200 168.575 78.520 168.635 ;
        RECT 14.650 167.955 115.850 168.435 ;
        RECT 17.020 167.755 17.340 167.815 ;
        RECT 17.020 167.615 18.630 167.755 ;
        RECT 17.020 167.555 17.340 167.615 ;
        RECT 17.495 167.415 17.785 167.460 ;
        RECT 17.940 167.415 18.260 167.475 ;
        RECT 17.495 167.275 18.260 167.415 ;
        RECT 18.490 167.415 18.630 167.615 ;
        RECT 29.900 167.555 30.220 167.815 ;
        RECT 31.755 167.755 32.045 167.800 ;
        RECT 34.500 167.755 34.820 167.815 ;
        RECT 39.560 167.755 39.880 167.815 ;
        RECT 51.980 167.755 52.300 167.815 ;
        RECT 31.755 167.615 39.330 167.755 ;
        RECT 31.755 167.570 32.045 167.615 ;
        RECT 34.500 167.555 34.820 167.615 ;
        RECT 19.775 167.415 20.425 167.460 ;
        RECT 23.375 167.415 23.665 167.460 ;
        RECT 18.490 167.275 23.665 167.415 ;
        RECT 17.495 167.230 17.785 167.275 ;
        RECT 17.940 167.215 18.260 167.275 ;
        RECT 19.775 167.230 20.425 167.275 ;
        RECT 23.075 167.230 23.665 167.275 ;
        RECT 33.235 167.415 33.525 167.460 ;
        RECT 36.475 167.415 37.125 167.460 ;
        RECT 33.235 167.275 37.125 167.415 ;
        RECT 39.190 167.415 39.330 167.615 ;
        RECT 39.560 167.615 52.300 167.755 ;
        RECT 39.560 167.555 39.880 167.615 ;
        RECT 51.980 167.555 52.300 167.615 ;
        RECT 52.440 167.755 52.760 167.815 ;
        RECT 71.775 167.755 72.065 167.800 ;
        RECT 73.600 167.755 73.920 167.815 ;
        RECT 52.440 167.615 61.410 167.755 ;
        RECT 52.440 167.555 52.760 167.615 ;
        RECT 42.320 167.415 42.640 167.475 ;
        RECT 39.190 167.275 42.640 167.415 ;
        RECT 33.235 167.230 33.825 167.275 ;
        RECT 36.475 167.230 37.125 167.275 ;
        RECT 16.580 167.075 16.870 167.120 ;
        RECT 18.415 167.075 18.705 167.120 ;
        RECT 21.995 167.075 22.285 167.120 ;
        RECT 16.580 166.935 22.285 167.075 ;
        RECT 16.580 166.890 16.870 166.935 ;
        RECT 18.415 166.890 18.705 166.935 ;
        RECT 21.995 166.890 22.285 166.935 ;
        RECT 23.075 166.915 23.365 167.230 ;
        RECT 33.535 167.135 33.825 167.230 ;
        RECT 42.320 167.215 42.640 167.275 ;
        RECT 53.015 167.415 53.305 167.460 ;
        RECT 56.255 167.415 56.905 167.460 ;
        RECT 53.015 167.275 56.905 167.415 ;
        RECT 53.015 167.230 53.605 167.275 ;
        RECT 56.255 167.230 56.905 167.275 ;
        RECT 58.420 167.415 58.740 167.475 ;
        RECT 60.735 167.415 61.025 167.460 ;
        RECT 58.420 167.275 61.025 167.415 ;
        RECT 53.315 167.135 53.605 167.230 ;
        RECT 58.420 167.215 58.740 167.275 ;
        RECT 60.735 167.230 61.025 167.275 ;
        RECT 24.380 167.075 24.700 167.135 ;
        RECT 27.615 167.075 27.905 167.120 ;
        RECT 24.380 166.935 27.905 167.075 ;
        RECT 24.380 166.875 24.700 166.935 ;
        RECT 27.615 166.890 27.905 166.935 ;
        RECT 30.360 167.075 30.680 167.135 ;
        RECT 30.835 167.075 31.125 167.120 ;
        RECT 30.360 166.935 31.125 167.075 ;
        RECT 30.360 166.875 30.680 166.935 ;
        RECT 30.835 166.890 31.125 166.935 ;
        RECT 33.535 166.915 33.900 167.135 ;
        RECT 33.580 166.875 33.900 166.915 ;
        RECT 34.615 167.075 34.905 167.120 ;
        RECT 38.195 167.075 38.485 167.120 ;
        RECT 40.030 167.075 40.320 167.120 ;
        RECT 34.615 166.935 40.320 167.075 ;
        RECT 34.615 166.890 34.905 166.935 ;
        RECT 38.195 166.890 38.485 166.935 ;
        RECT 40.030 166.890 40.320 166.935 ;
        RECT 40.940 166.875 41.260 167.135 ;
        RECT 53.315 166.915 53.680 167.135 ;
        RECT 53.360 166.875 53.680 166.915 ;
        RECT 54.395 167.075 54.685 167.120 ;
        RECT 57.975 167.075 58.265 167.120 ;
        RECT 59.810 167.075 60.100 167.120 ;
        RECT 54.395 166.935 60.100 167.075 ;
        RECT 54.395 166.890 54.685 166.935 ;
        RECT 57.975 166.890 58.265 166.935 ;
        RECT 59.810 166.890 60.100 166.935 ;
        RECT 60.275 166.890 60.565 167.120 ;
        RECT 61.270 167.075 61.410 167.615 ;
        RECT 71.775 167.615 73.920 167.755 ;
        RECT 71.775 167.570 72.065 167.615 ;
        RECT 73.600 167.555 73.920 167.615 ;
        RECT 76.375 167.570 76.665 167.800 ;
        RECT 62.560 167.215 62.880 167.475 ;
        RECT 65.335 167.415 65.625 167.460 ;
        RECT 67.160 167.415 67.480 167.475 ;
        RECT 68.555 167.415 68.845 167.460 ;
        RECT 65.335 167.275 68.845 167.415 ;
        RECT 65.335 167.230 65.625 167.275 ;
        RECT 67.160 167.215 67.480 167.275 ;
        RECT 68.555 167.230 68.845 167.275 ;
        RECT 71.300 167.415 71.620 167.475 ;
        RECT 74.535 167.415 74.825 167.460 ;
        RECT 71.300 167.275 74.825 167.415 ;
        RECT 76.450 167.415 76.590 167.570 ;
        RECT 77.740 167.555 78.060 167.815 ;
        RECT 79.120 167.555 79.440 167.815 ;
        RECT 86.480 167.555 86.800 167.815 ;
        RECT 79.210 167.415 79.350 167.555 ;
        RECT 76.450 167.275 79.350 167.415 ;
        RECT 101.660 167.415 101.980 167.475 ;
        RECT 103.975 167.415 104.265 167.460 ;
        RECT 106.375 167.415 106.665 167.460 ;
        RECT 109.615 167.415 110.265 167.460 ;
        RECT 101.660 167.275 103.730 167.415 ;
        RECT 71.300 167.215 71.620 167.275 ;
        RECT 74.535 167.230 74.825 167.275 ;
        RECT 101.660 167.215 101.980 167.275 ;
        RECT 63.495 167.075 63.785 167.120 ;
        RECT 61.270 166.935 63.785 167.075 ;
        RECT 63.495 166.890 63.785 166.935 ;
        RECT 66.255 166.890 66.545 167.120 ;
        RECT 16.100 166.535 16.420 166.795 ;
        RECT 24.855 166.735 25.145 166.780 ;
        RECT 28.075 166.735 28.365 166.780 ;
        RECT 24.855 166.595 28.365 166.735 ;
        RECT 24.855 166.550 25.145 166.595 ;
        RECT 28.075 166.550 28.365 166.595 ;
        RECT 16.985 166.395 17.275 166.440 ;
        RECT 18.875 166.395 19.165 166.440 ;
        RECT 21.995 166.395 22.285 166.440 ;
        RECT 16.985 166.255 22.285 166.395 ;
        RECT 16.985 166.210 17.275 166.255 ;
        RECT 18.875 166.210 19.165 166.255 ;
        RECT 21.995 166.210 22.285 166.255 ;
        RECT 23.460 166.395 23.780 166.455 ;
        RECT 25.775 166.395 26.065 166.440 ;
        RECT 23.460 166.255 26.065 166.395 ;
        RECT 23.460 166.195 23.780 166.255 ;
        RECT 25.775 166.210 26.065 166.255 ;
        RECT 28.150 166.055 28.290 166.550 ;
        RECT 28.980 166.535 29.300 166.795 ;
        RECT 39.100 166.535 39.420 166.795 ;
        RECT 40.495 166.735 40.785 166.780 ;
        RECT 42.780 166.735 43.100 166.795 ;
        RECT 40.495 166.595 43.100 166.735 ;
        RECT 40.495 166.550 40.785 166.595 ;
        RECT 42.780 166.535 43.100 166.595 ;
        RECT 57.040 166.735 57.360 166.795 ;
        RECT 58.895 166.735 59.185 166.780 ;
        RECT 57.040 166.595 59.185 166.735 ;
        RECT 57.040 166.535 57.360 166.595 ;
        RECT 58.895 166.550 59.185 166.595 ;
        RECT 34.615 166.395 34.905 166.440 ;
        RECT 37.735 166.395 38.025 166.440 ;
        RECT 39.625 166.395 39.915 166.440 ;
        RECT 48.760 166.395 49.080 166.455 ;
        RECT 34.615 166.255 39.915 166.395 ;
        RECT 34.615 166.210 34.905 166.255 ;
        RECT 37.735 166.210 38.025 166.255 ;
        RECT 39.625 166.210 39.915 166.255 ;
        RECT 47.470 166.255 49.080 166.395 ;
        RECT 47.470 166.055 47.610 166.255 ;
        RECT 48.760 166.195 49.080 166.255 ;
        RECT 51.535 166.395 51.825 166.440 ;
        RECT 51.980 166.395 52.300 166.455 ;
        RECT 51.535 166.255 52.300 166.395 ;
        RECT 51.535 166.210 51.825 166.255 ;
        RECT 51.980 166.195 52.300 166.255 ;
        RECT 54.395 166.395 54.685 166.440 ;
        RECT 57.515 166.395 57.805 166.440 ;
        RECT 59.405 166.395 59.695 166.440 ;
        RECT 54.395 166.255 59.695 166.395 ;
        RECT 54.395 166.210 54.685 166.255 ;
        RECT 57.515 166.210 57.805 166.255 ;
        RECT 59.405 166.210 59.695 166.255 ;
        RECT 60.350 166.395 60.490 166.890 ;
        RECT 66.330 166.735 66.470 166.890 ;
        RECT 67.620 166.875 67.940 167.135 ;
        RECT 68.095 167.075 68.385 167.120 ;
        RECT 69.460 167.075 69.780 167.135 ;
        RECT 68.095 166.935 69.780 167.075 ;
        RECT 68.095 166.890 68.385 166.935 ;
        RECT 69.460 166.875 69.780 166.935 ;
        RECT 72.235 167.075 72.525 167.120 ;
        RECT 78.200 167.075 78.520 167.135 ;
        RECT 72.235 166.935 78.520 167.075 ;
        RECT 72.235 166.890 72.525 166.935 ;
        RECT 78.200 166.875 78.520 166.935 ;
        RECT 79.120 166.875 79.440 167.135 ;
        RECT 89.255 166.890 89.545 167.120 ;
        RECT 67.160 166.735 67.480 166.795 ;
        RECT 69.000 166.735 69.320 166.795 ;
        RECT 66.330 166.595 69.320 166.735 ;
        RECT 67.160 166.535 67.480 166.595 ;
        RECT 69.000 166.535 69.320 166.595 ;
        RECT 73.140 166.535 73.460 166.795 ;
        RECT 74.060 166.535 74.380 166.795 ;
        RECT 78.290 166.735 78.430 166.875 ;
        RECT 89.330 166.735 89.470 166.890 ;
        RECT 90.620 166.875 90.940 167.135 ;
        RECT 103.590 167.120 103.730 167.275 ;
        RECT 103.975 167.275 110.265 167.415 ;
        RECT 103.975 167.230 104.265 167.275 ;
        RECT 106.375 167.230 106.965 167.275 ;
        RECT 109.615 167.230 110.265 167.275 ;
        RECT 102.135 166.890 102.425 167.120 ;
        RECT 103.515 166.890 103.805 167.120 ;
        RECT 106.675 166.915 106.965 167.230 ;
        RECT 112.240 167.215 112.560 167.475 ;
        RECT 107.755 167.075 108.045 167.120 ;
        RECT 111.335 167.075 111.625 167.120 ;
        RECT 113.170 167.075 113.460 167.120 ;
        RECT 107.755 166.935 113.460 167.075 ;
        RECT 107.755 166.890 108.045 166.935 ;
        RECT 111.335 166.890 111.625 166.935 ;
        RECT 113.170 166.890 113.460 166.935 ;
        RECT 78.290 166.595 89.470 166.735 ;
        RECT 99.360 166.735 99.680 166.795 ;
        RECT 102.210 166.735 102.350 166.890 ;
        RECT 113.620 166.875 113.940 167.135 ;
        RECT 113.710 166.735 113.850 166.875 ;
        RECT 99.360 166.595 113.850 166.735 ;
        RECT 99.360 166.535 99.680 166.595 ;
        RECT 60.720 166.395 61.040 166.455 ;
        RECT 60.350 166.255 61.040 166.395 ;
        RECT 28.150 165.915 47.610 166.055 ;
        RECT 47.840 166.055 48.160 166.115 ;
        RECT 48.315 166.055 48.605 166.100 ;
        RECT 50.600 166.055 50.920 166.115 ;
        RECT 60.350 166.055 60.490 166.255 ;
        RECT 60.720 166.195 61.040 166.255 ;
        RECT 63.020 166.395 63.340 166.455 ;
        RECT 66.715 166.395 67.005 166.440 ;
        RECT 70.380 166.395 70.700 166.455 ;
        RECT 63.020 166.255 70.700 166.395 ;
        RECT 63.020 166.195 63.340 166.255 ;
        RECT 66.715 166.210 67.005 166.255 ;
        RECT 70.380 166.195 70.700 166.255 ;
        RECT 107.755 166.395 108.045 166.440 ;
        RECT 110.875 166.395 111.165 166.440 ;
        RECT 112.765 166.395 113.055 166.440 ;
        RECT 107.755 166.255 113.055 166.395 ;
        RECT 107.755 166.210 108.045 166.255 ;
        RECT 110.875 166.210 111.165 166.255 ;
        RECT 112.765 166.210 113.055 166.255 ;
        RECT 47.840 165.915 60.490 166.055 ;
        RECT 47.840 165.855 48.160 165.915 ;
        RECT 48.315 165.870 48.605 165.915 ;
        RECT 50.600 165.855 50.920 165.915 ;
        RECT 89.700 165.855 90.020 166.115 ;
        RECT 103.960 166.055 104.280 166.115 ;
        RECT 104.895 166.055 105.185 166.100 ;
        RECT 103.960 165.915 105.185 166.055 ;
        RECT 103.960 165.855 104.280 165.915 ;
        RECT 104.895 165.870 105.185 165.915 ;
        RECT 14.650 165.235 115.850 165.715 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 39.100 164.835 39.420 165.095 ;
        RECT 49.220 165.035 49.540 165.095 ;
        RECT 54.755 165.035 55.045 165.080 ;
        RECT 49.220 164.895 55.045 165.035 ;
        RECT 49.220 164.835 49.540 164.895 ;
        RECT 54.755 164.850 55.045 164.895 ;
        RECT 57.040 164.835 57.360 165.095 ;
        RECT 64.400 165.035 64.720 165.095 ;
        RECT 65.795 165.035 66.085 165.080 ;
        RECT 64.400 164.895 66.085 165.035 ;
        RECT 64.400 164.835 64.720 164.895 ;
        RECT 65.795 164.850 66.085 164.895 ;
        RECT 78.660 164.835 78.980 165.095 ;
        RECT 90.405 165.035 90.695 165.080 ;
        RECT 92.460 165.035 92.780 165.095 ;
        RECT 88.870 164.895 92.780 165.035 ;
        RECT 16.580 164.695 16.870 164.740 ;
        RECT 18.440 164.695 18.730 164.740 ;
        RECT 21.220 164.695 21.510 164.740 ;
        RECT 16.580 164.555 21.510 164.695 ;
        RECT 16.580 164.510 16.870 164.555 ;
        RECT 18.440 164.510 18.730 164.555 ;
        RECT 21.220 164.510 21.510 164.555 ;
        RECT 37.260 164.695 37.580 164.755 ;
        RECT 40.495 164.695 40.785 164.740 ;
        RECT 37.260 164.555 40.785 164.695 ;
        RECT 37.260 164.495 37.580 164.555 ;
        RECT 40.495 164.510 40.785 164.555 ;
        RECT 50.155 164.695 50.445 164.740 ;
        RECT 50.155 164.555 55.890 164.695 ;
        RECT 50.155 164.510 50.445 164.555 ;
        RECT 17.940 164.155 18.260 164.415 ;
        RECT 25.760 164.355 26.080 164.415 ;
        RECT 28.980 164.355 29.300 164.415 ;
        RECT 43.715 164.355 44.005 164.400 ;
        RECT 47.395 164.355 47.685 164.400 ;
        RECT 51.535 164.355 51.825 164.400 ;
        RECT 52.440 164.355 52.760 164.415 ;
        RECT 18.490 164.215 27.830 164.355 ;
        RECT 16.100 164.015 16.420 164.075 ;
        RECT 18.490 164.015 18.630 164.215 ;
        RECT 25.760 164.155 26.080 164.215 ;
        RECT 27.690 164.060 27.830 164.215 ;
        RECT 28.980 164.215 52.760 164.355 ;
        RECT 28.980 164.155 29.300 164.215 ;
        RECT 37.350 164.075 37.490 164.215 ;
        RECT 43.715 164.170 44.005 164.215 ;
        RECT 47.395 164.170 47.685 164.215 ;
        RECT 51.535 164.170 51.825 164.215 ;
        RECT 52.440 164.155 52.760 164.215 ;
        RECT 21.220 164.015 21.510 164.060 ;
        RECT 16.100 163.875 18.630 164.015 ;
        RECT 18.975 163.875 21.510 164.015 ;
        RECT 16.100 163.815 16.420 163.875 ;
        RECT 18.975 163.720 19.190 163.875 ;
        RECT 21.220 163.830 21.510 163.875 ;
        RECT 27.615 164.015 27.905 164.060 ;
        RECT 30.820 164.015 31.140 164.075 ;
        RECT 36.800 164.015 37.120 164.075 ;
        RECT 27.615 163.875 37.120 164.015 ;
        RECT 27.615 163.830 27.905 163.875 ;
        RECT 30.820 163.815 31.140 163.875 ;
        RECT 36.800 163.815 37.120 163.875 ;
        RECT 37.260 163.815 37.580 164.075 ;
        RECT 37.720 164.015 38.040 164.075 ;
        RECT 40.035 164.015 40.325 164.060 ;
        RECT 37.720 163.875 40.325 164.015 ;
        RECT 37.720 163.815 38.040 163.875 ;
        RECT 40.035 163.830 40.325 163.875 ;
        RECT 41.860 164.015 42.180 164.075 ;
        RECT 55.750 164.060 55.890 164.555 ;
        RECT 61.655 164.355 61.945 164.400 ;
        RECT 62.100 164.355 62.420 164.415 ;
        RECT 69.460 164.355 69.780 164.415 ;
        RECT 61.655 164.215 62.420 164.355 ;
        RECT 61.655 164.170 61.945 164.215 ;
        RECT 62.100 164.155 62.420 164.215 ;
        RECT 66.790 164.215 69.780 164.355 ;
        RECT 42.335 164.015 42.625 164.060 ;
        RECT 51.995 164.015 52.285 164.060 ;
        RECT 41.860 163.875 42.625 164.015 ;
        RECT 41.860 163.815 42.180 163.875 ;
        RECT 42.335 163.830 42.625 163.875 ;
        RECT 48.390 163.875 52.285 164.015 ;
        RECT 17.040 163.675 17.330 163.720 ;
        RECT 18.900 163.675 19.190 163.720 ;
        RECT 17.040 163.535 19.190 163.675 ;
        RECT 17.040 163.490 17.330 163.535 ;
        RECT 18.900 163.490 19.190 163.535 ;
        RECT 19.780 163.720 20.100 163.735 ;
        RECT 19.780 163.675 20.110 163.720 ;
        RECT 23.080 163.675 23.370 163.720 ;
        RECT 19.780 163.535 23.370 163.675 ;
        RECT 19.780 163.490 20.110 163.535 ;
        RECT 23.080 163.490 23.370 163.535 ;
        RECT 35.435 163.675 35.725 163.720 ;
        RECT 40.940 163.675 41.260 163.735 ;
        RECT 35.435 163.535 41.260 163.675 ;
        RECT 35.435 163.490 35.725 163.535 ;
        RECT 19.780 163.475 20.100 163.490 ;
        RECT 40.940 163.475 41.260 163.535 ;
        RECT 48.390 163.395 48.530 163.875 ;
        RECT 51.995 163.830 52.285 163.875 ;
        RECT 55.675 163.830 55.965 164.060 ;
        RECT 56.120 163.815 56.440 164.075 ;
        RECT 57.975 164.015 58.265 164.060 ;
        RECT 58.420 164.015 58.740 164.075 ;
        RECT 57.975 163.875 61.870 164.015 ;
        RECT 57.975 163.830 58.265 163.875 ;
        RECT 58.420 163.815 58.740 163.875 ;
        RECT 61.730 163.735 61.870 163.875 ;
        RECT 62.560 163.815 62.880 164.075 ;
        RECT 64.400 164.015 64.720 164.075 ;
        RECT 66.790 164.060 66.930 164.215 ;
        RECT 69.460 164.155 69.780 164.215 ;
        RECT 73.140 164.355 73.460 164.415 ;
        RECT 74.075 164.355 74.365 164.400 ;
        RECT 86.035 164.355 86.325 164.400 ;
        RECT 73.140 164.215 87.170 164.355 ;
        RECT 73.140 164.155 73.460 164.215 ;
        RECT 74.075 164.170 74.365 164.215 ;
        RECT 86.035 164.170 86.325 164.215 ;
        RECT 66.715 164.015 67.005 164.060 ;
        RECT 64.400 163.875 67.005 164.015 ;
        RECT 64.400 163.815 64.720 163.875 ;
        RECT 66.715 163.830 67.005 163.875 ;
        RECT 67.160 163.815 67.480 164.075 ;
        RECT 75.440 164.015 75.760 164.075 ;
        RECT 77.755 164.015 78.045 164.060 ;
        RECT 68.170 163.875 75.760 164.015 ;
        RECT 48.760 163.675 49.080 163.735 ;
        RECT 52.455 163.675 52.745 163.720 ;
        RECT 48.760 163.535 52.745 163.675 ;
        RECT 48.760 163.475 49.080 163.535 ;
        RECT 52.455 163.490 52.745 163.535 ;
        RECT 61.640 163.475 61.960 163.735 ;
        RECT 62.650 163.675 62.790 163.815 ;
        RECT 68.170 163.675 68.310 163.875 ;
        RECT 75.440 163.815 75.760 163.875 ;
        RECT 77.370 163.875 78.045 164.015 ;
        RECT 62.650 163.535 68.310 163.675 ;
        RECT 71.300 163.675 71.620 163.735 ;
        RECT 74.995 163.675 75.285 163.720 ;
        RECT 71.300 163.535 75.285 163.675 ;
        RECT 25.085 163.335 25.375 163.380 ;
        RECT 29.900 163.335 30.220 163.395 ;
        RECT 25.085 163.195 30.220 163.335 ;
        RECT 25.085 163.150 25.375 163.195 ;
        RECT 29.900 163.135 30.220 163.195 ;
        RECT 40.480 163.335 40.800 163.395 ;
        RECT 42.795 163.335 43.085 163.380 ;
        RECT 40.480 163.195 43.085 163.335 ;
        RECT 40.480 163.135 40.800 163.195 ;
        RECT 42.795 163.150 43.085 163.195 ;
        RECT 46.920 163.335 47.240 163.395 ;
        RECT 47.855 163.335 48.145 163.380 ;
        RECT 46.920 163.195 48.145 163.335 ;
        RECT 46.920 163.135 47.240 163.195 ;
        RECT 47.855 163.150 48.145 163.195 ;
        RECT 48.300 163.135 48.620 163.395 ;
        RECT 51.980 163.335 52.300 163.395 ;
        RECT 54.295 163.335 54.585 163.380 ;
        RECT 51.980 163.195 54.585 163.335 ;
        RECT 51.980 163.135 52.300 163.195 ;
        RECT 54.295 163.150 54.585 163.195 ;
        RECT 58.420 163.135 58.740 163.395 ;
        RECT 59.800 163.335 60.120 163.395 ;
        RECT 62.650 163.335 62.790 163.535 ;
        RECT 71.300 163.475 71.620 163.535 ;
        RECT 74.995 163.490 75.285 163.535 ;
        RECT 59.800 163.195 62.790 163.335 ;
        RECT 68.095 163.335 68.385 163.380 ;
        RECT 70.380 163.335 70.700 163.395 ;
        RECT 68.095 163.195 70.700 163.335 ;
        RECT 59.800 163.135 60.120 163.195 ;
        RECT 68.095 163.150 68.385 163.195 ;
        RECT 70.380 163.135 70.700 163.195 ;
        RECT 74.520 163.335 74.840 163.395 ;
        RECT 77.370 163.380 77.510 163.875 ;
        RECT 77.755 163.830 78.045 163.875 ;
        RECT 87.030 163.675 87.170 164.215 ;
        RECT 87.415 164.015 87.705 164.060 ;
        RECT 88.870 164.015 89.010 164.895 ;
        RECT 90.405 164.850 90.695 164.895 ;
        RECT 92.460 164.835 92.780 164.895 ;
        RECT 104.420 165.035 104.740 165.095 ;
        RECT 109.035 165.035 109.325 165.080 ;
        RECT 104.420 164.895 109.325 165.035 ;
        RECT 104.420 164.835 104.740 164.895 ;
        RECT 109.035 164.850 109.325 164.895 ;
        RECT 94.270 164.695 94.560 164.740 ;
        RECT 97.050 164.695 97.340 164.740 ;
        RECT 98.910 164.695 99.200 164.740 ;
        RECT 94.270 164.555 99.200 164.695 ;
        RECT 94.270 164.510 94.560 164.555 ;
        RECT 97.050 164.510 97.340 164.555 ;
        RECT 98.910 164.510 99.200 164.555 ;
        RECT 102.695 164.695 102.985 164.740 ;
        RECT 105.815 164.695 106.105 164.740 ;
        RECT 107.705 164.695 107.995 164.740 ;
        RECT 102.695 164.555 107.995 164.695 ;
        RECT 102.695 164.510 102.985 164.555 ;
        RECT 105.815 164.510 106.105 164.555 ;
        RECT 107.705 164.510 107.995 164.555 ;
        RECT 89.240 164.355 89.560 164.415 ;
        RECT 97.535 164.355 97.825 164.400 ;
        RECT 89.240 164.215 97.825 164.355 ;
        RECT 89.240 164.155 89.560 164.215 ;
        RECT 97.535 164.170 97.825 164.215 ;
        RECT 99.360 164.155 99.680 164.415 ;
        RECT 103.960 164.355 104.280 164.415 ;
        RECT 111.795 164.355 112.085 164.400 ;
        RECT 103.960 164.215 112.085 164.355 ;
        RECT 103.960 164.155 104.280 164.215 ;
        RECT 111.795 164.170 112.085 164.215 ;
        RECT 93.380 164.015 93.700 164.075 ;
        RECT 87.415 163.875 89.010 164.015 ;
        RECT 89.330 163.875 93.700 164.015 ;
        RECT 87.415 163.830 87.705 163.875 ;
        RECT 89.330 163.675 89.470 163.875 ;
        RECT 93.380 163.815 93.700 163.875 ;
        RECT 94.270 164.015 94.560 164.060 ;
        RECT 94.270 163.875 96.805 164.015 ;
        RECT 94.270 163.830 94.560 163.875 ;
        RECT 87.030 163.535 89.470 163.675 ;
        RECT 89.700 163.675 90.020 163.735 ;
        RECT 96.590 163.720 96.805 163.875 ;
        RECT 92.410 163.675 92.700 163.720 ;
        RECT 95.670 163.675 95.960 163.720 ;
        RECT 89.700 163.535 95.960 163.675 ;
        RECT 89.700 163.475 90.020 163.535 ;
        RECT 92.410 163.490 92.700 163.535 ;
        RECT 95.670 163.490 95.960 163.535 ;
        RECT 96.590 163.675 96.880 163.720 ;
        RECT 98.450 163.675 98.740 163.720 ;
        RECT 96.590 163.535 98.740 163.675 ;
        RECT 96.590 163.490 96.880 163.535 ;
        RECT 98.450 163.490 98.740 163.535 ;
        RECT 98.900 163.675 99.220 163.735 ;
        RECT 101.615 163.720 101.905 164.035 ;
        RECT 102.695 164.015 102.985 164.060 ;
        RECT 106.275 164.015 106.565 164.060 ;
        RECT 108.110 164.015 108.400 164.060 ;
        RECT 102.695 163.875 108.400 164.015 ;
        RECT 102.695 163.830 102.985 163.875 ;
        RECT 106.275 163.830 106.565 163.875 ;
        RECT 108.110 163.830 108.400 163.875 ;
        RECT 108.575 164.015 108.865 164.060 ;
        RECT 113.160 164.015 113.480 164.075 ;
        RECT 108.575 163.875 113.480 164.015 ;
        RECT 108.575 163.830 108.865 163.875 ;
        RECT 113.160 163.815 113.480 163.875 ;
        RECT 101.315 163.675 101.905 163.720 ;
        RECT 104.555 163.675 105.205 163.720 ;
        RECT 98.900 163.535 105.205 163.675 ;
        RECT 98.900 163.475 99.220 163.535 ;
        RECT 101.315 163.490 101.605 163.535 ;
        RECT 104.555 163.490 105.205 163.535 ;
        RECT 107.180 163.475 107.500 163.735 ;
        RECT 75.455 163.335 75.745 163.380 ;
        RECT 74.520 163.195 75.745 163.335 ;
        RECT 74.520 163.135 74.840 163.195 ;
        RECT 75.455 163.150 75.745 163.195 ;
        RECT 77.295 163.150 77.585 163.380 ;
        RECT 84.180 163.335 84.500 163.395 ;
        RECT 86.955 163.335 87.245 163.380 ;
        RECT 84.180 163.195 87.245 163.335 ;
        RECT 84.180 163.135 84.500 163.195 ;
        RECT 86.955 163.150 87.245 163.195 ;
        RECT 89.255 163.335 89.545 163.380 ;
        RECT 93.380 163.335 93.700 163.395 ;
        RECT 89.255 163.195 93.700 163.335 ;
        RECT 89.255 163.150 89.545 163.195 ;
        RECT 93.380 163.135 93.700 163.195 ;
        RECT 97.980 163.335 98.300 163.395 ;
        RECT 99.835 163.335 100.125 163.380 ;
        RECT 97.980 163.195 100.125 163.335 ;
        RECT 97.980 163.135 98.300 163.195 ;
        RECT 99.835 163.150 100.125 163.195 ;
        RECT 14.650 162.515 115.850 162.995 ;
        RECT 18.415 162.315 18.705 162.360 ;
        RECT 19.780 162.315 20.100 162.375 ;
        RECT 18.415 162.175 20.100 162.315 ;
        RECT 18.415 162.130 18.705 162.175 ;
        RECT 19.780 162.115 20.100 162.175 ;
        RECT 24.380 162.315 24.700 162.375 ;
        RECT 28.995 162.315 29.285 162.360 ;
        RECT 24.380 162.175 29.285 162.315 ;
        RECT 24.380 162.115 24.700 162.175 ;
        RECT 28.995 162.130 29.285 162.175 ;
        RECT 30.360 162.315 30.680 162.375 ;
        RECT 31.295 162.315 31.585 162.360 ;
        RECT 30.360 162.175 31.585 162.315 ;
        RECT 30.360 162.115 30.680 162.175 ;
        RECT 31.295 162.130 31.585 162.175 ;
        RECT 41.860 162.115 42.180 162.375 ;
        RECT 46.920 162.115 47.240 162.375 ;
        RECT 47.395 162.315 47.685 162.360 ;
        RECT 48.300 162.315 48.620 162.375 ;
        RECT 47.395 162.175 48.620 162.315 ;
        RECT 47.395 162.130 47.685 162.175 ;
        RECT 48.300 162.115 48.620 162.175 ;
        RECT 55.215 162.315 55.505 162.360 ;
        RECT 56.120 162.315 56.440 162.375 ;
        RECT 55.215 162.175 56.440 162.315 ;
        RECT 55.215 162.130 55.505 162.175 ;
        RECT 56.120 162.115 56.440 162.175 ;
        RECT 61.655 162.130 61.945 162.360 ;
        RECT 21.175 161.975 21.465 162.020 ;
        RECT 22.540 161.975 22.860 162.035 ;
        RECT 21.175 161.835 22.860 161.975 ;
        RECT 21.175 161.790 21.465 161.835 ;
        RECT 22.540 161.775 22.860 161.835 ;
        RECT 30.820 161.975 31.140 162.035 ;
        RECT 35.895 161.975 36.185 162.020 ;
        RECT 40.480 161.975 40.800 162.035 ;
        RECT 30.820 161.835 34.730 161.975 ;
        RECT 30.820 161.775 31.140 161.835 ;
        RECT 18.400 161.635 18.720 161.695 ;
        RECT 18.875 161.635 19.165 161.680 ;
        RECT 18.400 161.495 19.165 161.635 ;
        RECT 18.400 161.435 18.720 161.495 ;
        RECT 18.875 161.450 19.165 161.495 ;
        RECT 21.635 161.635 21.925 161.680 ;
        RECT 29.455 161.635 29.745 161.680 ;
        RECT 29.900 161.635 30.220 161.695 ;
        RECT 21.635 161.495 30.220 161.635 ;
        RECT 21.635 161.450 21.925 161.495 ;
        RECT 29.455 161.450 29.745 161.495 ;
        RECT 29.900 161.435 30.220 161.495 ;
        RECT 32.675 161.635 32.965 161.680 ;
        RECT 34.590 161.635 34.730 161.835 ;
        RECT 35.895 161.835 40.800 161.975 ;
        RECT 41.950 161.975 42.090 162.115 ;
        RECT 57.500 161.975 57.820 162.035 ;
        RECT 61.730 161.975 61.870 162.130 ;
        RECT 67.160 162.115 67.480 162.375 ;
        RECT 69.460 162.315 69.780 162.375 ;
        RECT 67.710 162.175 69.780 162.315 ;
        RECT 67.250 161.975 67.390 162.115 ;
        RECT 41.950 161.835 43.930 161.975 ;
        RECT 35.895 161.790 36.185 161.835 ;
        RECT 40.480 161.775 40.800 161.835 ;
        RECT 36.355 161.635 36.645 161.680 ;
        RECT 41.315 161.635 41.605 161.680 ;
        RECT 32.675 161.495 34.270 161.635 ;
        RECT 34.590 161.495 36.645 161.635 ;
        RECT 32.675 161.450 32.965 161.495 ;
        RECT 22.555 161.295 22.845 161.340 ;
        RECT 28.535 161.295 28.825 161.340 ;
        RECT 28.980 161.295 29.300 161.355 ;
        RECT 22.555 161.155 29.300 161.295 ;
        RECT 22.555 161.110 22.845 161.155 ;
        RECT 28.535 161.110 28.825 161.155 ;
        RECT 28.980 161.095 29.300 161.155 ;
        RECT 34.130 161.000 34.270 161.495 ;
        RECT 36.355 161.450 36.645 161.495 ;
        RECT 41.260 161.450 41.605 161.635 ;
        RECT 41.875 161.450 42.165 161.680 ;
        RECT 37.260 161.095 37.580 161.355 ;
        RECT 34.055 160.770 34.345 161.000 ;
        RECT 41.260 160.955 41.400 161.450 ;
        RECT 41.950 160.955 42.090 161.450 ;
        RECT 42.320 161.435 42.640 161.695 ;
        RECT 43.240 161.435 43.560 161.695 ;
        RECT 43.790 161.680 43.930 161.835 ;
        RECT 57.500 161.835 61.870 161.975 ;
        RECT 62.650 161.835 67.390 161.975 ;
        RECT 57.500 161.775 57.820 161.835 ;
        RECT 43.715 161.635 44.005 161.680 ;
        RECT 44.160 161.635 44.480 161.695 ;
        RECT 43.715 161.495 44.480 161.635 ;
        RECT 43.715 161.450 44.005 161.495 ;
        RECT 44.160 161.435 44.480 161.495 ;
        RECT 50.615 161.635 50.905 161.680 ;
        RECT 51.520 161.635 51.840 161.695 ;
        RECT 50.615 161.495 51.840 161.635 ;
        RECT 50.615 161.450 50.905 161.495 ;
        RECT 51.520 161.435 51.840 161.495 ;
        RECT 51.980 161.435 52.300 161.695 ;
        RECT 57.975 161.635 58.265 161.680 ;
        RECT 59.800 161.635 60.120 161.695 ;
        RECT 62.650 161.680 62.790 161.835 ;
        RECT 57.975 161.495 60.120 161.635 ;
        RECT 57.975 161.450 58.265 161.495 ;
        RECT 59.800 161.435 60.120 161.495 ;
        RECT 60.735 161.450 61.025 161.680 ;
        RECT 62.575 161.450 62.865 161.680 ;
        RECT 46.920 161.295 47.240 161.355 ;
        RECT 56.595 161.295 56.885 161.340 ;
        RECT 46.920 161.155 56.885 161.295 ;
        RECT 60.810 161.295 60.950 161.450 ;
        RECT 63.020 161.435 63.340 161.695 ;
        RECT 66.715 161.635 67.005 161.680 ;
        RECT 67.160 161.635 67.480 161.695 ;
        RECT 66.715 161.495 67.480 161.635 ;
        RECT 66.715 161.450 67.005 161.495 ;
        RECT 67.160 161.435 67.480 161.495 ;
        RECT 63.110 161.295 63.250 161.435 ;
        RECT 60.810 161.155 63.250 161.295 ;
        RECT 46.920 161.095 47.240 161.155 ;
        RECT 56.595 161.110 56.885 161.155 ;
        RECT 57.960 160.955 58.280 161.015 ;
        RECT 65.795 160.955 66.085 161.000 ;
        RECT 67.710 160.955 67.850 162.175 ;
        RECT 69.460 162.115 69.780 162.175 ;
        RECT 112.240 162.315 112.560 162.375 ;
        RECT 112.715 162.315 113.005 162.360 ;
        RECT 112.240 162.175 113.005 162.315 ;
        RECT 112.240 162.115 112.560 162.175 ;
        RECT 112.715 162.130 113.005 162.175 ;
        RECT 72.680 161.975 73.000 162.035 ;
        RECT 74.535 161.975 74.825 162.020 ;
        RECT 83.045 161.975 83.335 162.020 ;
        RECT 84.180 161.975 84.500 162.035 ;
        RECT 72.680 161.835 84.500 161.975 ;
        RECT 72.680 161.775 73.000 161.835 ;
        RECT 74.535 161.790 74.825 161.835 ;
        RECT 83.045 161.790 83.335 161.835 ;
        RECT 84.180 161.775 84.500 161.835 ;
        RECT 85.050 161.975 85.340 162.020 ;
        RECT 86.020 161.975 86.340 162.035 ;
        RECT 88.310 161.975 88.600 162.020 ;
        RECT 85.050 161.835 88.600 161.975 ;
        RECT 85.050 161.790 85.340 161.835 ;
        RECT 86.020 161.775 86.340 161.835 ;
        RECT 88.310 161.790 88.600 161.835 ;
        RECT 89.230 161.975 89.520 162.020 ;
        RECT 91.090 161.975 91.380 162.020 ;
        RECT 89.230 161.835 91.380 161.975 ;
        RECT 89.230 161.790 89.520 161.835 ;
        RECT 91.090 161.790 91.380 161.835 ;
        RECT 94.300 161.975 94.620 162.035 ;
        RECT 94.775 161.975 95.065 162.020 ;
        RECT 103.960 161.975 104.280 162.035 ;
        RECT 94.300 161.835 95.065 161.975 ;
        RECT 70.380 161.435 70.700 161.695 ;
        RECT 70.840 161.435 71.160 161.695 ;
        RECT 71.300 161.435 71.620 161.695 ;
        RECT 72.235 161.635 72.525 161.680 ;
        RECT 73.600 161.635 73.920 161.695 ;
        RECT 72.235 161.495 73.920 161.635 ;
        RECT 72.235 161.450 72.525 161.495 ;
        RECT 72.310 160.955 72.450 161.450 ;
        RECT 73.600 161.435 73.920 161.495 ;
        RECT 78.200 161.635 78.520 161.695 ;
        RECT 80.055 161.635 80.345 161.680 ;
        RECT 78.200 161.495 80.345 161.635 ;
        RECT 78.200 161.435 78.520 161.495 ;
        RECT 80.055 161.450 80.345 161.495 ;
        RECT 80.515 161.450 80.805 161.680 ;
        RECT 86.910 161.635 87.200 161.680 ;
        RECT 89.230 161.635 89.445 161.790 ;
        RECT 94.300 161.775 94.620 161.835 ;
        RECT 94.775 161.790 95.065 161.835 ;
        RECT 99.450 161.835 104.280 161.975 ;
        RECT 86.910 161.495 89.445 161.635 ;
        RECT 90.175 161.635 90.465 161.680 ;
        RECT 90.175 161.495 92.690 161.635 ;
        RECT 86.910 161.450 87.200 161.495 ;
        RECT 90.175 161.450 90.465 161.495 ;
        RECT 73.140 161.095 73.460 161.355 ;
        RECT 74.075 161.295 74.365 161.340 ;
        RECT 74.520 161.295 74.840 161.355 ;
        RECT 80.590 161.295 80.730 161.450 ;
        RECT 74.075 161.155 74.840 161.295 ;
        RECT 74.075 161.110 74.365 161.155 ;
        RECT 74.520 161.095 74.840 161.155 ;
        RECT 76.450 161.155 80.730 161.295 ;
        RECT 86.480 161.295 86.800 161.355 ;
        RECT 92.015 161.295 92.305 161.340 ;
        RECT 86.480 161.155 92.305 161.295 ;
        RECT 76.450 161.000 76.590 161.155 ;
        RECT 86.480 161.095 86.800 161.155 ;
        RECT 92.015 161.110 92.305 161.155 ;
        RECT 92.550 161.000 92.690 161.495 ;
        RECT 93.380 161.435 93.700 161.695 ;
        RECT 97.980 161.435 98.300 161.695 ;
        RECT 98.455 161.635 98.745 161.680 ;
        RECT 98.900 161.635 99.220 161.695 ;
        RECT 99.450 161.680 99.590 161.835 ;
        RECT 103.960 161.775 104.280 161.835 ;
        RECT 104.420 161.975 104.740 162.035 ;
        RECT 105.355 161.975 105.645 162.020 ;
        RECT 104.420 161.835 105.645 161.975 ;
        RECT 104.420 161.775 104.740 161.835 ;
        RECT 105.355 161.790 105.645 161.835 ;
        RECT 109.020 161.975 109.340 162.035 ;
        RECT 109.955 161.975 110.245 162.020 ;
        RECT 109.020 161.835 110.245 161.975 ;
        RECT 109.020 161.775 109.340 161.835 ;
        RECT 109.955 161.790 110.245 161.835 ;
        RECT 98.455 161.495 99.220 161.635 ;
        RECT 98.455 161.450 98.745 161.495 ;
        RECT 98.900 161.435 99.220 161.495 ;
        RECT 99.375 161.450 99.665 161.680 ;
        RECT 99.835 161.450 100.125 161.680 ;
        RECT 99.910 161.295 100.050 161.450 ;
        RECT 100.280 161.435 100.600 161.695 ;
        RECT 105.800 161.435 106.120 161.695 ;
        RECT 108.100 161.635 108.420 161.695 ;
        RECT 111.335 161.635 111.625 161.680 ;
        RECT 108.100 161.495 111.625 161.635 ;
        RECT 108.100 161.435 108.420 161.495 ;
        RECT 111.335 161.450 111.625 161.495 ;
        RECT 111.795 161.450 112.085 161.680 ;
        RECT 99.450 161.155 100.050 161.295 ;
        RECT 99.450 161.015 99.590 161.155 ;
        RECT 104.880 161.095 105.200 161.355 ;
        RECT 108.560 161.295 108.880 161.355 ;
        RECT 111.870 161.295 112.010 161.450 ;
        RECT 108.560 161.155 112.010 161.295 ;
        RECT 108.560 161.095 108.880 161.155 ;
        RECT 41.260 160.815 41.630 160.955 ;
        RECT 41.950 160.815 46.690 160.955 ;
        RECT 19.320 160.415 19.640 160.675 ;
        RECT 33.595 160.615 33.885 160.660 ;
        RECT 35.880 160.615 36.200 160.675 ;
        RECT 33.595 160.475 36.200 160.615 ;
        RECT 33.595 160.430 33.885 160.475 ;
        RECT 35.880 160.415 36.200 160.475 ;
        RECT 39.560 160.615 39.880 160.675 ;
        RECT 40.035 160.615 40.325 160.660 ;
        RECT 39.560 160.475 40.325 160.615 ;
        RECT 41.490 160.615 41.630 160.815 ;
        RECT 46.550 160.675 46.690 160.815 ;
        RECT 57.960 160.815 67.850 160.955 ;
        RECT 68.630 160.815 72.450 160.955 ;
        RECT 57.960 160.755 58.280 160.815 ;
        RECT 65.795 160.770 66.085 160.815 ;
        RECT 42.780 160.615 43.100 160.675 ;
        RECT 41.490 160.475 43.100 160.615 ;
        RECT 39.560 160.415 39.880 160.475 ;
        RECT 40.035 160.430 40.325 160.475 ;
        RECT 42.780 160.415 43.100 160.475 ;
        RECT 46.460 160.615 46.780 160.675 ;
        RECT 49.220 160.615 49.540 160.675 ;
        RECT 59.800 160.615 60.120 160.675 ;
        RECT 46.460 160.475 60.120 160.615 ;
        RECT 46.460 160.415 46.780 160.475 ;
        RECT 49.220 160.415 49.540 160.475 ;
        RECT 59.800 160.415 60.120 160.475 ;
        RECT 63.940 160.415 64.260 160.675 ;
        RECT 67.160 160.615 67.480 160.675 ;
        RECT 68.095 160.615 68.385 160.660 ;
        RECT 68.630 160.615 68.770 160.815 ;
        RECT 76.375 160.770 76.665 161.000 ;
        RECT 86.910 160.955 87.200 161.000 ;
        RECT 89.690 160.955 89.980 161.000 ;
        RECT 91.550 160.955 91.840 161.000 ;
        RECT 86.910 160.815 91.840 160.955 ;
        RECT 86.910 160.770 87.200 160.815 ;
        RECT 89.690 160.770 89.980 160.815 ;
        RECT 91.550 160.770 91.840 160.815 ;
        RECT 92.475 160.770 92.765 161.000 ;
        RECT 99.360 160.755 99.680 161.015 ;
        RECT 67.160 160.475 68.770 160.615 ;
        RECT 67.160 160.415 67.480 160.475 ;
        RECT 68.095 160.430 68.385 160.475 ;
        RECT 69.000 160.415 69.320 160.675 ;
        RECT 69.460 160.615 69.780 160.675 ;
        RECT 78.200 160.615 78.520 160.675 ;
        RECT 69.460 160.475 78.520 160.615 ;
        RECT 69.460 160.415 69.780 160.475 ;
        RECT 78.200 160.415 78.520 160.475 ;
        RECT 78.660 160.615 78.980 160.675 ;
        RECT 79.595 160.615 79.885 160.660 ;
        RECT 78.660 160.475 79.885 160.615 ;
        RECT 78.660 160.415 78.980 160.475 ;
        RECT 79.595 160.430 79.885 160.475 ;
        RECT 81.435 160.615 81.725 160.660 ;
        RECT 82.340 160.615 82.660 160.675 ;
        RECT 81.435 160.475 82.660 160.615 ;
        RECT 81.435 160.430 81.725 160.475 ;
        RECT 82.340 160.415 82.660 160.475 ;
        RECT 100.740 160.615 101.060 160.675 ;
        RECT 101.675 160.615 101.965 160.660 ;
        RECT 100.740 160.475 101.965 160.615 ;
        RECT 100.740 160.415 101.060 160.475 ;
        RECT 101.675 160.430 101.965 160.475 ;
        RECT 107.640 160.415 107.960 160.675 ;
        RECT 14.650 159.795 115.850 160.275 ;
        RECT 28.765 159.595 29.055 159.640 ;
        RECT 30.820 159.595 31.140 159.655 ;
        RECT 28.765 159.455 31.140 159.595 ;
        RECT 28.765 159.410 29.055 159.455 ;
        RECT 30.820 159.395 31.140 159.455 ;
        RECT 36.800 159.595 37.120 159.655 ;
        RECT 63.940 159.595 64.260 159.655 ;
        RECT 66.700 159.595 67.020 159.655 ;
        RECT 74.060 159.595 74.380 159.655 ;
        RECT 36.800 159.455 67.020 159.595 ;
        RECT 36.800 159.395 37.120 159.455 ;
        RECT 63.940 159.395 64.260 159.455 ;
        RECT 66.700 159.395 67.020 159.455 ;
        RECT 68.170 159.455 74.380 159.595 ;
        RECT 20.670 159.255 20.960 159.300 ;
        RECT 23.450 159.255 23.740 159.300 ;
        RECT 25.310 159.255 25.600 159.300 ;
        RECT 20.670 159.115 25.600 159.255 ;
        RECT 20.670 159.070 20.960 159.115 ;
        RECT 23.450 159.070 23.740 159.115 ;
        RECT 25.310 159.070 25.600 159.115 ;
        RECT 32.630 159.255 32.920 159.300 ;
        RECT 35.410 159.255 35.700 159.300 ;
        RECT 37.270 159.255 37.560 159.300 ;
        RECT 32.630 159.115 37.560 159.255 ;
        RECT 32.630 159.070 32.920 159.115 ;
        RECT 35.410 159.070 35.700 159.115 ;
        RECT 37.270 159.070 37.560 159.115 ;
        RECT 38.180 159.255 38.500 159.315 ;
        RECT 43.240 159.255 43.560 159.315 ;
        RECT 45.080 159.255 45.400 159.315 ;
        RECT 63.480 159.255 63.800 159.315 ;
        RECT 38.180 159.115 52.670 159.255 ;
        RECT 38.180 159.055 38.500 159.115 ;
        RECT 43.240 159.055 43.560 159.115 ;
        RECT 45.080 159.055 45.400 159.115 ;
        RECT 16.805 158.915 17.095 158.960 ;
        RECT 22.540 158.915 22.860 158.975 ;
        RECT 16.805 158.775 22.860 158.915 ;
        RECT 16.805 158.730 17.095 158.775 ;
        RECT 22.540 158.715 22.860 158.775 ;
        RECT 25.760 158.715 26.080 158.975 ;
        RECT 35.880 158.715 36.200 158.975 ;
        RECT 37.735 158.915 38.025 158.960 ;
        RECT 39.100 158.915 39.420 158.975 ;
        RECT 37.735 158.775 39.420 158.915 ;
        RECT 37.735 158.730 38.025 158.775 ;
        RECT 39.100 158.715 39.420 158.775 ;
        RECT 46.460 158.915 46.780 158.975 ;
        RECT 46.460 158.775 47.610 158.915 ;
        RECT 46.460 158.715 46.780 158.775 ;
        RECT 20.670 158.575 20.960 158.620 ;
        RECT 20.670 158.435 23.205 158.575 ;
        RECT 20.670 158.390 20.960 158.435 ;
        RECT 18.860 158.280 19.180 158.295 ;
        RECT 22.990 158.280 23.205 158.435 ;
        RECT 23.920 158.375 24.240 158.635 ;
        RECT 27.140 158.375 27.460 158.635 ;
        RECT 32.630 158.575 32.920 158.620 ;
        RECT 32.630 158.435 35.165 158.575 ;
        RECT 32.630 158.390 32.920 158.435 ;
        RECT 34.950 158.280 35.165 158.435 ;
        RECT 43.240 158.375 43.560 158.635 ;
        RECT 43.715 158.390 44.005 158.620 ;
        RECT 18.810 158.235 19.180 158.280 ;
        RECT 22.070 158.235 22.360 158.280 ;
        RECT 18.810 158.095 22.360 158.235 ;
        RECT 18.810 158.050 19.180 158.095 ;
        RECT 22.070 158.050 22.360 158.095 ;
        RECT 22.990 158.235 23.280 158.280 ;
        RECT 24.850 158.235 25.140 158.280 ;
        RECT 22.990 158.095 25.140 158.235 ;
        RECT 22.990 158.050 23.280 158.095 ;
        RECT 24.850 158.050 25.140 158.095 ;
        RECT 27.615 158.235 27.905 158.280 ;
        RECT 30.770 158.235 31.060 158.280 ;
        RECT 34.030 158.235 34.320 158.280 ;
        RECT 27.615 158.095 34.320 158.235 ;
        RECT 27.615 158.050 27.905 158.095 ;
        RECT 30.770 158.050 31.060 158.095 ;
        RECT 34.030 158.050 34.320 158.095 ;
        RECT 34.950 158.235 35.240 158.280 ;
        RECT 36.810 158.235 37.100 158.280 ;
        RECT 43.790 158.235 43.930 158.390 ;
        RECT 44.160 158.375 44.480 158.635 ;
        RECT 45.080 158.375 45.400 158.635 ;
        RECT 45.540 158.575 45.860 158.635 ;
        RECT 47.470 158.620 47.610 158.775 ;
        RECT 46.935 158.575 47.225 158.620 ;
        RECT 45.540 158.435 47.225 158.575 ;
        RECT 45.540 158.375 45.860 158.435 ;
        RECT 46.935 158.390 47.225 158.435 ;
        RECT 47.395 158.390 47.685 158.620 ;
        RECT 47.855 158.560 48.145 158.605 ;
        RECT 48.300 158.560 48.620 158.635 ;
        RECT 48.850 158.620 48.990 159.115 ;
        RECT 49.680 158.915 50.000 158.975 ;
        RECT 49.680 158.775 51.290 158.915 ;
        RECT 49.680 158.715 50.000 158.775 ;
        RECT 47.855 158.420 48.620 158.560 ;
        RECT 46.460 158.235 46.780 158.295 ;
        RECT 34.950 158.095 37.100 158.235 ;
        RECT 34.950 158.050 35.240 158.095 ;
        RECT 36.810 158.050 37.100 158.095 ;
        RECT 41.030 158.095 46.780 158.235 ;
        RECT 47.010 158.235 47.150 158.390 ;
        RECT 47.855 158.375 48.145 158.420 ;
        RECT 48.300 158.375 48.620 158.420 ;
        RECT 48.775 158.390 49.065 158.620 ;
        RECT 50.600 158.575 50.920 158.635 ;
        RECT 51.150 158.620 51.290 158.775 ;
        RECT 50.230 158.435 50.920 158.575 ;
        RECT 50.230 158.235 50.370 158.435 ;
        RECT 50.600 158.375 50.920 158.435 ;
        RECT 51.060 158.390 51.350 158.620 ;
        RECT 51.535 158.575 51.825 158.620 ;
        RECT 51.980 158.575 52.300 158.635 ;
        RECT 52.530 158.620 52.670 159.115 ;
        RECT 63.480 159.115 65.550 159.255 ;
        RECT 63.480 159.055 63.800 159.115 ;
        RECT 54.740 158.715 55.060 158.975 ;
        RECT 65.410 158.620 65.550 159.115 ;
        RECT 51.535 158.435 52.300 158.575 ;
        RECT 51.535 158.390 51.825 158.435 ;
        RECT 51.980 158.375 52.300 158.435 ;
        RECT 52.455 158.575 52.745 158.620 ;
        RECT 52.455 158.435 65.090 158.575 ;
        RECT 52.455 158.390 52.745 158.435 ;
        RECT 47.010 158.095 50.370 158.235 ;
        RECT 18.860 158.035 19.180 158.050 ;
        RECT 41.030 157.955 41.170 158.095 ;
        RECT 46.460 158.035 46.780 158.095 ;
        RECT 63.480 158.035 63.800 158.295 ;
        RECT 64.950 158.235 65.090 158.435 ;
        RECT 65.335 158.390 65.625 158.620 ;
        RECT 67.160 158.375 67.480 158.635 ;
        RECT 68.170 158.620 68.310 159.455 ;
        RECT 74.060 159.395 74.380 159.455 ;
        RECT 75.440 159.595 75.760 159.655 ;
        RECT 86.020 159.595 86.340 159.655 ;
        RECT 86.495 159.595 86.785 159.640 ;
        RECT 75.440 159.455 84.410 159.595 ;
        RECT 75.440 159.395 75.760 159.455 ;
        RECT 70.395 159.255 70.685 159.300 ;
        RECT 72.220 159.255 72.540 159.315 ;
        RECT 70.395 159.115 72.540 159.255 ;
        RECT 70.395 159.070 70.685 159.115 ;
        RECT 72.220 159.055 72.540 159.115 ;
        RECT 79.090 159.255 79.380 159.300 ;
        RECT 81.870 159.255 82.160 159.300 ;
        RECT 83.730 159.255 84.020 159.300 ;
        RECT 79.090 159.115 84.020 159.255 ;
        RECT 84.270 159.255 84.410 159.455 ;
        RECT 86.020 159.455 86.785 159.595 ;
        RECT 86.020 159.395 86.340 159.455 ;
        RECT 86.495 159.410 86.785 159.455 ;
        RECT 89.240 159.395 89.560 159.655 ;
        RECT 91.540 159.595 91.860 159.655 ;
        RECT 92.015 159.595 92.305 159.640 ;
        RECT 108.100 159.595 108.420 159.655 ;
        RECT 91.540 159.455 92.305 159.595 ;
        RECT 91.540 159.395 91.860 159.455 ;
        RECT 92.015 159.410 92.305 159.455 ;
        RECT 107.500 159.455 108.420 159.595 ;
        RECT 107.500 159.255 107.640 159.455 ;
        RECT 108.100 159.395 108.420 159.455 ;
        RECT 108.560 159.395 108.880 159.655 ;
        RECT 84.270 159.115 107.640 159.255 ;
        RECT 79.090 159.070 79.380 159.115 ;
        RECT 81.870 159.070 82.160 159.115 ;
        RECT 83.730 159.070 84.020 159.115 ;
        RECT 69.460 158.915 69.780 158.975 ;
        RECT 70.855 158.915 71.145 158.960 ;
        RECT 69.460 158.775 71.145 158.915 ;
        RECT 69.460 158.715 69.780 158.775 ;
        RECT 70.855 158.730 71.145 158.775 ;
        RECT 71.760 158.915 72.080 158.975 ;
        RECT 77.740 158.915 78.060 158.975 ;
        RECT 71.760 158.775 73.830 158.915 ;
        RECT 71.760 158.715 72.080 158.775 ;
        RECT 73.690 158.635 73.830 158.775 ;
        RECT 77.740 158.775 82.110 158.915 ;
        RECT 77.740 158.715 78.060 158.775 ;
        RECT 68.095 158.390 68.385 158.620 ;
        RECT 68.555 158.390 68.845 158.620 ;
        RECT 69.015 158.575 69.305 158.620 ;
        RECT 70.380 158.575 70.700 158.635 ;
        RECT 72.235 158.575 72.525 158.620 ;
        RECT 69.015 158.435 72.525 158.575 ;
        RECT 69.015 158.390 69.305 158.435 ;
        RECT 67.250 158.235 67.390 158.375 ;
        RECT 64.950 158.095 67.390 158.235 ;
        RECT 68.630 158.235 68.770 158.390 ;
        RECT 70.380 158.375 70.700 158.435 ;
        RECT 72.235 158.390 72.525 158.435 ;
        RECT 72.695 158.390 72.985 158.620 ;
        RECT 73.155 158.390 73.445 158.620 ;
        RECT 73.600 158.575 73.920 158.635 ;
        RECT 74.075 158.575 74.365 158.620 ;
        RECT 73.600 158.435 74.365 158.575 ;
        RECT 71.300 158.235 71.620 158.295 ;
        RECT 72.770 158.235 72.910 158.390 ;
        RECT 68.630 158.095 72.910 158.235 ;
        RECT 73.230 158.235 73.370 158.390 ;
        RECT 73.600 158.375 73.920 158.435 ;
        RECT 74.075 158.390 74.365 158.435 ;
        RECT 79.090 158.575 79.380 158.620 ;
        RECT 81.970 158.575 82.110 158.775 ;
        RECT 82.340 158.715 82.660 158.975 ;
        RECT 84.195 158.915 84.485 158.960 ;
        RECT 86.480 158.915 86.800 158.975 ;
        RECT 84.195 158.775 86.800 158.915 ;
        RECT 84.195 158.730 84.485 158.775 ;
        RECT 86.480 158.715 86.800 158.775 ;
        RECT 92.920 158.715 93.240 158.975 ;
        RECT 99.360 158.915 99.680 158.975 ;
        RECT 93.470 158.775 100.510 158.915 ;
        RECT 86.035 158.575 86.325 158.620 ;
        RECT 86.940 158.575 87.260 158.635 ;
        RECT 79.090 158.435 81.625 158.575 ;
        RECT 81.970 158.435 87.260 158.575 ;
        RECT 79.090 158.390 79.380 158.435 ;
        RECT 74.520 158.235 74.840 158.295 ;
        RECT 75.225 158.235 75.515 158.280 ;
        RECT 73.230 158.095 75.515 158.235 ;
        RECT 71.300 158.035 71.620 158.095 ;
        RECT 74.520 158.035 74.840 158.095 ;
        RECT 75.225 158.050 75.515 158.095 ;
        RECT 77.230 158.235 77.520 158.280 ;
        RECT 78.660 158.235 78.980 158.295 ;
        RECT 81.410 158.280 81.625 158.435 ;
        RECT 86.035 158.390 86.325 158.435 ;
        RECT 86.940 158.375 87.260 158.435 ;
        RECT 88.335 158.575 88.625 158.620 ;
        RECT 91.080 158.575 91.400 158.635 ;
        RECT 88.335 158.435 91.400 158.575 ;
        RECT 88.335 158.390 88.625 158.435 ;
        RECT 91.080 158.375 91.400 158.435 ;
        RECT 92.000 158.375 92.320 158.635 ;
        RECT 93.470 158.575 93.610 158.775 ;
        RECT 93.010 158.435 93.610 158.575 ;
        RECT 93.840 158.575 94.160 158.635 ;
        RECT 96.690 158.620 96.830 158.775 ;
        RECT 99.360 158.715 99.680 158.775 ;
        RECT 96.155 158.575 96.445 158.620 ;
        RECT 93.840 158.435 96.445 158.575 ;
        RECT 93.010 158.295 93.150 158.435 ;
        RECT 93.840 158.375 94.160 158.435 ;
        RECT 96.155 158.390 96.445 158.435 ;
        RECT 96.615 158.390 96.905 158.620 ;
        RECT 97.075 158.575 97.365 158.620 ;
        RECT 97.520 158.575 97.840 158.635 ;
        RECT 97.075 158.435 97.840 158.575 ;
        RECT 97.075 158.390 97.365 158.435 ;
        RECT 80.490 158.235 80.780 158.280 ;
        RECT 77.230 158.095 80.780 158.235 ;
        RECT 77.230 158.050 77.520 158.095 ;
        RECT 78.660 158.035 78.980 158.095 ;
        RECT 80.490 158.050 80.780 158.095 ;
        RECT 81.410 158.235 81.700 158.280 ;
        RECT 83.270 158.235 83.560 158.280 ;
        RECT 92.920 158.235 93.240 158.295 ;
        RECT 81.410 158.095 83.560 158.235 ;
        RECT 81.410 158.050 81.700 158.095 ;
        RECT 83.270 158.050 83.560 158.095 ;
        RECT 90.710 158.095 93.240 158.235 ;
        RECT 90.710 157.955 90.850 158.095 ;
        RECT 92.920 158.035 93.240 158.095 ;
        RECT 93.380 158.035 93.700 158.295 ;
        RECT 96.230 158.235 96.370 158.390 ;
        RECT 97.520 158.375 97.840 158.435 ;
        RECT 97.995 158.575 98.285 158.620 ;
        RECT 98.440 158.575 98.760 158.635 ;
        RECT 98.915 158.575 99.205 158.620 ;
        RECT 97.995 158.435 99.205 158.575 ;
        RECT 97.995 158.390 98.285 158.435 ;
        RECT 98.440 158.375 98.760 158.435 ;
        RECT 98.915 158.390 99.205 158.435 ;
        RECT 99.820 158.375 100.140 158.635 ;
        RECT 100.370 158.620 100.510 158.775 ;
        RECT 102.670 158.620 102.810 159.115 ;
        RECT 105.815 158.915 106.105 158.960 ;
        RECT 107.640 158.915 107.960 158.975 ;
        RECT 105.815 158.775 107.960 158.915 ;
        RECT 105.815 158.730 106.105 158.775 ;
        RECT 107.640 158.715 107.960 158.775 ;
        RECT 100.295 158.390 100.585 158.620 ;
        RECT 100.755 158.390 101.045 158.620 ;
        RECT 102.595 158.390 102.885 158.620 ;
        RECT 100.830 158.235 100.970 158.390 ;
        RECT 93.930 158.095 95.910 158.235 ;
        RECT 96.230 158.095 100.970 158.235 ;
        RECT 32.660 157.895 32.980 157.955 ;
        RECT 37.260 157.895 37.580 157.955 ;
        RECT 32.660 157.755 37.580 157.895 ;
        RECT 32.660 157.695 32.980 157.755 ;
        RECT 37.260 157.695 37.580 157.755 ;
        RECT 39.100 157.895 39.420 157.955 ;
        RECT 40.940 157.895 41.260 157.955 ;
        RECT 39.100 157.755 41.260 157.895 ;
        RECT 39.100 157.695 39.420 157.755 ;
        RECT 40.940 157.695 41.260 157.755 ;
        RECT 41.400 157.895 41.720 157.955 ;
        RECT 41.875 157.895 42.165 157.940 ;
        RECT 41.400 157.755 42.165 157.895 ;
        RECT 41.400 157.695 41.720 157.755 ;
        RECT 41.875 157.710 42.165 157.755 ;
        RECT 42.780 157.895 43.100 157.955 ;
        RECT 45.555 157.895 45.845 157.940 ;
        RECT 42.780 157.755 45.845 157.895 ;
        RECT 42.780 157.695 43.100 157.755 ;
        RECT 45.555 157.710 45.845 157.755 ;
        RECT 46.000 157.895 46.320 157.955 ;
        RECT 49.235 157.895 49.525 157.940 ;
        RECT 46.000 157.755 49.525 157.895 ;
        RECT 46.000 157.695 46.320 157.755 ;
        RECT 49.235 157.710 49.525 157.755 ;
        RECT 58.880 157.895 59.200 157.955 ;
        RECT 66.255 157.895 66.545 157.940 ;
        RECT 58.880 157.755 66.545 157.895 ;
        RECT 58.880 157.695 59.200 157.755 ;
        RECT 66.255 157.710 66.545 157.755 ;
        RECT 66.700 157.895 67.020 157.955 ;
        RECT 90.620 157.895 90.940 157.955 ;
        RECT 66.700 157.755 90.940 157.895 ;
        RECT 66.700 157.695 67.020 157.755 ;
        RECT 90.620 157.695 90.940 157.755 ;
        RECT 91.095 157.895 91.385 157.940 ;
        RECT 93.930 157.895 94.070 158.095 ;
        RECT 91.095 157.755 94.070 157.895 ;
        RECT 94.300 157.895 94.620 157.955 ;
        RECT 94.775 157.895 95.065 157.940 ;
        RECT 94.300 157.755 95.065 157.895 ;
        RECT 95.770 157.895 95.910 158.095 ;
        RECT 100.370 157.955 100.510 158.095 ;
        RECT 103.960 158.035 104.280 158.295 ;
        RECT 99.820 157.895 100.140 157.955 ;
        RECT 95.770 157.755 100.140 157.895 ;
        RECT 91.095 157.710 91.385 157.755 ;
        RECT 94.300 157.695 94.620 157.755 ;
        RECT 94.775 157.710 95.065 157.755 ;
        RECT 99.820 157.695 100.140 157.755 ;
        RECT 100.280 157.695 100.600 157.955 ;
        RECT 101.200 157.895 101.520 157.955 ;
        RECT 102.135 157.895 102.425 157.940 ;
        RECT 101.200 157.755 102.425 157.895 ;
        RECT 101.200 157.695 101.520 157.755 ;
        RECT 102.135 157.710 102.425 157.755 ;
        RECT 14.650 157.075 115.850 157.555 ;
        RECT 17.940 156.875 18.260 156.935 ;
        RECT 18.875 156.875 19.165 156.920 ;
        RECT 17.940 156.735 19.165 156.875 ;
        RECT 17.940 156.675 18.260 156.735 ;
        RECT 18.875 156.690 19.165 156.735 ;
        RECT 23.000 156.875 23.320 156.935 ;
        RECT 70.380 156.875 70.700 156.935 ;
        RECT 92.000 156.875 92.320 156.935 ;
        RECT 93.855 156.875 94.145 156.920 ;
        RECT 98.440 156.875 98.760 156.935 ;
        RECT 23.000 156.735 40.250 156.875 ;
        RECT 23.000 156.675 23.320 156.735 ;
        RECT 29.900 156.535 30.220 156.595 ;
        RECT 33.120 156.535 33.440 156.595 ;
        RECT 39.100 156.535 39.420 156.595 ;
        RECT 29.900 156.395 32.890 156.535 ;
        RECT 29.900 156.335 30.220 156.395 ;
        RECT 19.320 156.195 19.640 156.255 ;
        RECT 19.795 156.195 20.085 156.240 ;
        RECT 19.320 156.055 20.085 156.195 ;
        RECT 19.320 155.995 19.640 156.055 ;
        RECT 19.795 156.010 20.085 156.055 ;
        RECT 22.095 156.195 22.385 156.240 ;
        RECT 23.000 156.195 23.320 156.255 ;
        RECT 22.095 156.055 23.320 156.195 ;
        RECT 22.095 156.010 22.385 156.055 ;
        RECT 23.000 155.995 23.320 156.055 ;
        RECT 31.740 155.995 32.060 156.255 ;
        RECT 32.200 155.995 32.520 156.255 ;
        RECT 32.750 156.240 32.890 156.395 ;
        RECT 33.120 156.395 36.110 156.535 ;
        RECT 33.120 156.335 33.440 156.395 ;
        RECT 32.675 156.010 32.965 156.240 ;
        RECT 33.580 155.995 33.900 156.255 ;
        RECT 35.970 156.240 36.110 156.395 ;
        RECT 37.350 156.395 39.420 156.535 ;
        RECT 37.350 156.240 37.490 156.395 ;
        RECT 39.100 156.335 39.420 156.395 ;
        RECT 35.895 156.010 36.185 156.240 ;
        RECT 36.815 156.010 37.105 156.240 ;
        RECT 37.275 156.010 37.565 156.240 ;
        RECT 37.735 156.010 38.025 156.240 ;
        RECT 38.180 156.195 38.500 156.255 ;
        RECT 39.575 156.195 39.865 156.240 ;
        RECT 38.180 156.055 39.865 156.195 ;
        RECT 40.110 156.195 40.250 156.735 ;
        RECT 70.380 156.735 73.830 156.875 ;
        RECT 70.380 156.675 70.700 156.735 ;
        RECT 57.450 156.535 57.740 156.580 ;
        RECT 58.420 156.535 58.740 156.595 ;
        RECT 60.710 156.535 61.000 156.580 ;
        RECT 57.450 156.395 61.000 156.535 ;
        RECT 57.450 156.350 57.740 156.395 ;
        RECT 58.420 156.335 58.740 156.395 ;
        RECT 60.710 156.350 61.000 156.395 ;
        RECT 61.630 156.535 61.920 156.580 ;
        RECT 63.490 156.535 63.780 156.580 ;
        RECT 61.630 156.395 63.780 156.535 ;
        RECT 61.630 156.350 61.920 156.395 ;
        RECT 63.490 156.350 63.780 156.395 ;
        RECT 67.620 156.535 67.940 156.595 ;
        RECT 71.300 156.535 71.620 156.595 ;
        RECT 67.620 156.395 69.230 156.535 ;
        RECT 40.495 156.195 40.785 156.240 ;
        RECT 40.110 156.055 40.785 156.195 ;
        RECT 21.175 155.670 21.465 155.900 ;
        RECT 21.635 155.855 21.925 155.900 ;
        RECT 22.540 155.855 22.860 155.915 ;
        RECT 36.890 155.855 37.030 156.010 ;
        RECT 21.635 155.715 37.030 155.855 ;
        RECT 37.810 155.855 37.950 156.010 ;
        RECT 38.180 155.995 38.500 156.055 ;
        RECT 39.575 156.010 39.865 156.055 ;
        RECT 40.495 156.010 40.785 156.055 ;
        RECT 40.940 155.995 41.260 156.255 ;
        RECT 41.415 156.195 41.705 156.240 ;
        RECT 43.240 156.195 43.560 156.255 ;
        RECT 45.540 156.195 45.860 156.255 ;
        RECT 41.415 156.055 45.860 156.195 ;
        RECT 41.415 156.010 41.705 156.055 ;
        RECT 41.490 155.855 41.630 156.010 ;
        RECT 43.240 155.995 43.560 156.055 ;
        RECT 45.540 155.995 45.860 156.055 ;
        RECT 46.015 156.195 46.305 156.240 ;
        RECT 46.920 156.195 47.240 156.255 ;
        RECT 46.015 156.055 47.240 156.195 ;
        RECT 46.015 156.010 46.305 156.055 ;
        RECT 46.920 155.995 47.240 156.055 ;
        RECT 47.840 156.195 48.160 156.255 ;
        RECT 49.695 156.195 49.985 156.240 ;
        RECT 47.840 156.055 49.985 156.195 ;
        RECT 47.840 155.995 48.160 156.055 ;
        RECT 49.695 156.010 49.985 156.055 ;
        RECT 53.820 155.995 54.140 156.255 ;
        RECT 59.310 156.195 59.600 156.240 ;
        RECT 61.630 156.195 61.845 156.350 ;
        RECT 67.620 156.335 67.940 156.395 ;
        RECT 59.310 156.055 61.845 156.195 ;
        RECT 62.575 156.195 62.865 156.240 ;
        RECT 63.020 156.195 63.340 156.255 ;
        RECT 62.575 156.055 63.340 156.195 ;
        RECT 59.310 156.010 59.600 156.055 ;
        RECT 62.575 156.010 62.865 156.055 ;
        RECT 63.020 155.995 63.340 156.055 ;
        RECT 63.940 156.195 64.260 156.255 ;
        RECT 66.255 156.195 66.545 156.240 ;
        RECT 68.095 156.195 68.385 156.240 ;
        RECT 63.940 156.055 68.385 156.195 ;
        RECT 63.940 155.995 64.260 156.055 ;
        RECT 66.255 156.010 66.545 156.055 ;
        RECT 68.095 156.010 68.385 156.055 ;
        RECT 68.540 155.995 68.860 156.255 ;
        RECT 69.090 156.195 69.230 156.395 ;
        RECT 71.300 156.395 73.370 156.535 ;
        RECT 71.300 156.335 71.620 156.395 ;
        RECT 69.475 156.195 69.765 156.240 ;
        RECT 69.090 156.055 69.765 156.195 ;
        RECT 69.475 156.010 69.765 156.055 ;
        RECT 69.935 156.195 70.225 156.240 ;
        RECT 70.380 156.195 70.700 156.255 ;
        RECT 69.935 156.055 70.700 156.195 ;
        RECT 69.935 156.010 70.225 156.055 ;
        RECT 70.380 155.995 70.700 156.055 ;
        RECT 71.760 155.995 72.080 156.255 ;
        RECT 72.680 155.995 73.000 156.255 ;
        RECT 73.230 156.240 73.370 156.395 ;
        RECT 73.690 156.240 73.830 156.735 ;
        RECT 92.000 156.735 94.145 156.875 ;
        RECT 92.000 156.675 92.320 156.735 ;
        RECT 93.855 156.690 94.145 156.735 ;
        RECT 97.150 156.735 98.760 156.875 ;
        RECT 78.200 156.535 78.520 156.595 ;
        RECT 92.920 156.535 93.240 156.595 ;
        RECT 78.200 156.395 92.690 156.535 ;
        RECT 78.200 156.335 78.520 156.395 ;
        RECT 73.155 156.010 73.445 156.240 ;
        RECT 73.615 156.010 73.905 156.240 ;
        RECT 74.060 156.195 74.380 156.255 ;
        RECT 90.635 156.195 90.925 156.240 ;
        RECT 74.060 156.055 90.925 156.195 ;
        RECT 74.060 155.995 74.380 156.055 ;
        RECT 90.635 156.010 90.925 156.055 ;
        RECT 57.500 155.855 57.820 155.915 ;
        RECT 59.800 155.855 60.120 155.915 ;
        RECT 64.415 155.855 64.705 155.900 ;
        RECT 37.810 155.715 41.630 155.855 ;
        RECT 41.950 155.715 59.110 155.855 ;
        RECT 21.635 155.670 21.925 155.715 ;
        RECT 21.250 155.515 21.390 155.670 ;
        RECT 22.540 155.655 22.860 155.715 ;
        RECT 28.520 155.515 28.840 155.575 ;
        RECT 21.250 155.375 28.840 155.515 ;
        RECT 28.520 155.315 28.840 155.375 ;
        RECT 30.820 155.315 31.140 155.575 ;
        RECT 35.420 155.515 35.740 155.575 ;
        RECT 33.210 155.375 35.740 155.515 ;
        RECT 23.935 155.175 24.225 155.220 ;
        RECT 24.380 155.175 24.700 155.235 ;
        RECT 23.935 155.035 24.700 155.175 ;
        RECT 23.935 154.990 24.225 155.035 ;
        RECT 24.380 154.975 24.700 155.035 ;
        RECT 28.980 155.175 29.300 155.235 ;
        RECT 30.375 155.175 30.665 155.220 ;
        RECT 28.980 155.035 30.665 155.175 ;
        RECT 30.910 155.175 31.050 155.315 ;
        RECT 33.210 155.175 33.350 155.375 ;
        RECT 35.420 155.315 35.740 155.375 ;
        RECT 36.340 155.515 36.660 155.575 ;
        RECT 41.950 155.515 42.090 155.715 ;
        RECT 57.500 155.655 57.820 155.715 ;
        RECT 36.340 155.375 42.090 155.515 ;
        RECT 54.280 155.515 54.600 155.575 ;
        RECT 55.445 155.515 55.735 155.560 ;
        RECT 58.420 155.515 58.740 155.575 ;
        RECT 54.280 155.375 58.740 155.515 ;
        RECT 36.340 155.315 36.660 155.375 ;
        RECT 54.280 155.315 54.600 155.375 ;
        RECT 55.445 155.330 55.735 155.375 ;
        RECT 58.420 155.315 58.740 155.375 ;
        RECT 30.910 155.035 33.350 155.175 ;
        RECT 28.980 154.975 29.300 155.035 ;
        RECT 30.375 154.990 30.665 155.035 ;
        RECT 39.100 154.975 39.420 155.235 ;
        RECT 40.480 155.175 40.800 155.235 ;
        RECT 42.795 155.175 43.085 155.220 ;
        RECT 40.480 155.035 43.085 155.175 ;
        RECT 40.480 154.975 40.800 155.035 ;
        RECT 42.795 154.990 43.085 155.035 ;
        RECT 46.460 154.975 46.780 155.235 ;
        RECT 54.740 154.975 55.060 155.235 ;
        RECT 58.970 155.175 59.110 155.715 ;
        RECT 59.800 155.715 64.705 155.855 ;
        RECT 59.800 155.655 60.120 155.715 ;
        RECT 64.415 155.670 64.705 155.715 ;
        RECT 67.250 155.715 73.140 155.855 ;
        RECT 67.250 155.560 67.390 155.715 ;
        RECT 59.310 155.515 59.600 155.560 ;
        RECT 62.090 155.515 62.380 155.560 ;
        RECT 63.950 155.515 64.240 155.560 ;
        RECT 59.310 155.375 64.240 155.515 ;
        RECT 59.310 155.330 59.600 155.375 ;
        RECT 62.090 155.330 62.380 155.375 ;
        RECT 63.950 155.330 64.240 155.375 ;
        RECT 67.175 155.330 67.465 155.560 ;
        RECT 73.000 155.515 73.140 155.715 ;
        RECT 74.520 155.515 74.840 155.575 ;
        RECT 73.000 155.375 74.840 155.515 ;
        RECT 74.520 155.315 74.840 155.375 ;
        RECT 66.700 155.175 67.020 155.235 ;
        RECT 58.970 155.035 67.020 155.175 ;
        RECT 66.700 154.975 67.020 155.035 ;
        RECT 70.395 155.175 70.685 155.220 ;
        RECT 71.300 155.175 71.620 155.235 ;
        RECT 70.395 155.035 71.620 155.175 ;
        RECT 70.395 154.990 70.685 155.035 ;
        RECT 71.300 154.975 71.620 155.035 ;
        RECT 73.140 155.175 73.460 155.235 ;
        RECT 74.995 155.175 75.285 155.220 ;
        RECT 73.140 155.035 75.285 155.175 ;
        RECT 73.140 154.975 73.460 155.035 ;
        RECT 74.995 154.990 75.285 155.035 ;
        RECT 89.255 155.175 89.545 155.220 ;
        RECT 89.700 155.175 90.020 155.235 ;
        RECT 89.255 155.035 90.020 155.175 ;
        RECT 90.710 155.175 90.850 156.010 ;
        RECT 91.080 155.995 91.400 156.255 ;
        RECT 91.555 156.195 91.845 156.240 ;
        RECT 92.000 156.195 92.320 156.255 ;
        RECT 92.550 156.240 92.690 156.395 ;
        RECT 92.920 156.395 95.910 156.535 ;
        RECT 92.920 156.335 93.240 156.395 ;
        RECT 95.770 156.255 95.910 156.395 ;
        RECT 91.555 156.055 92.320 156.195 ;
        RECT 91.555 156.010 91.845 156.055 ;
        RECT 92.000 155.995 92.320 156.055 ;
        RECT 92.475 156.010 92.765 156.240 ;
        RECT 93.840 156.195 94.160 156.255 ;
        RECT 95.235 156.195 95.525 156.240 ;
        RECT 93.840 156.055 95.525 156.195 ;
        RECT 92.550 155.515 92.690 156.010 ;
        RECT 93.840 155.995 94.160 156.055 ;
        RECT 95.235 156.010 95.525 156.055 ;
        RECT 95.680 155.995 96.000 156.255 ;
        RECT 96.155 156.195 96.445 156.240 ;
        RECT 96.600 156.195 96.920 156.255 ;
        RECT 97.150 156.240 97.290 156.735 ;
        RECT 98.440 156.675 98.760 156.735 ;
        RECT 102.135 156.875 102.425 156.920 ;
        RECT 107.180 156.875 107.500 156.935 ;
        RECT 102.135 156.735 107.500 156.875 ;
        RECT 102.135 156.690 102.425 156.735 ;
        RECT 107.180 156.675 107.500 156.735 ;
        RECT 96.155 156.055 96.920 156.195 ;
        RECT 96.155 156.010 96.445 156.055 ;
        RECT 96.600 155.995 96.920 156.055 ;
        RECT 97.075 156.010 97.365 156.240 ;
        RECT 97.535 156.010 97.825 156.240 ;
        RECT 97.150 155.855 97.290 156.010 ;
        RECT 95.770 155.715 97.290 155.855 ;
        RECT 97.610 155.855 97.750 156.010 ;
        RECT 98.440 155.995 98.760 156.255 ;
        RECT 98.900 155.995 99.220 156.255 ;
        RECT 99.375 156.195 99.665 156.240 ;
        RECT 100.280 156.195 100.600 156.255 ;
        RECT 99.375 156.055 100.600 156.195 ;
        RECT 99.375 156.010 99.665 156.055 ;
        RECT 100.280 155.995 100.600 156.055 ;
        RECT 101.215 156.195 101.505 156.240 ;
        RECT 102.120 156.195 102.440 156.255 ;
        RECT 101.215 156.055 102.440 156.195 ;
        RECT 101.215 156.010 101.505 156.055 ;
        RECT 102.120 155.995 102.440 156.055 ;
        RECT 109.020 155.995 109.340 156.255 ;
        RECT 110.415 156.010 110.705 156.240 ;
        RECT 97.610 155.715 99.590 155.855 ;
        RECT 95.770 155.575 95.910 155.715 ;
        RECT 99.450 155.575 99.590 155.715 ;
        RECT 99.820 155.655 100.140 155.915 ;
        RECT 104.880 155.855 105.200 155.915 ;
        RECT 110.490 155.855 110.630 156.010 ;
        RECT 104.880 155.715 110.630 155.855 ;
        RECT 104.880 155.655 105.200 155.715 ;
        RECT 95.680 155.515 96.000 155.575 ;
        RECT 92.550 155.375 96.000 155.515 ;
        RECT 95.680 155.315 96.000 155.375 ;
        RECT 99.360 155.315 99.680 155.575 ;
        RECT 99.910 155.515 100.050 155.655 ;
        RECT 108.100 155.515 108.420 155.575 ;
        RECT 99.910 155.375 108.420 155.515 ;
        RECT 108.100 155.315 108.420 155.375 ;
        RECT 93.840 155.175 94.160 155.235 ;
        RECT 90.710 155.035 94.160 155.175 ;
        RECT 89.255 154.990 89.545 155.035 ;
        RECT 89.700 154.975 90.020 155.035 ;
        RECT 93.840 154.975 94.160 155.035 ;
        RECT 99.820 155.175 100.140 155.235 ;
        RECT 100.755 155.175 101.045 155.220 ;
        RECT 99.820 155.035 101.045 155.175 ;
        RECT 99.820 154.975 100.140 155.035 ;
        RECT 100.755 154.990 101.045 155.035 ;
        RECT 107.180 155.175 107.500 155.235 ;
        RECT 108.575 155.175 108.865 155.220 ;
        RECT 107.180 155.035 108.865 155.175 ;
        RECT 107.180 154.975 107.500 155.035 ;
        RECT 108.575 154.990 108.865 155.035 ;
        RECT 111.335 155.175 111.625 155.220 ;
        RECT 112.700 155.175 113.020 155.235 ;
        RECT 111.335 155.035 113.020 155.175 ;
        RECT 111.335 154.990 111.625 155.035 ;
        RECT 112.700 154.975 113.020 155.035 ;
        RECT 14.650 154.355 115.850 154.835 ;
        RECT 23.920 154.155 24.240 154.215 ;
        RECT 25.775 154.155 26.065 154.200 ;
        RECT 23.920 154.015 26.065 154.155 ;
        RECT 23.920 153.955 24.240 154.015 ;
        RECT 25.775 153.970 26.065 154.015 ;
        RECT 30.360 153.955 30.680 154.215 ;
        RECT 31.740 154.155 32.060 154.215 ;
        RECT 34.500 154.155 34.820 154.215 ;
        RECT 36.340 154.155 36.660 154.215 ;
        RECT 31.740 154.015 36.660 154.155 ;
        RECT 31.740 153.955 32.060 154.015 ;
        RECT 20.210 153.815 20.500 153.860 ;
        RECT 22.990 153.815 23.280 153.860 ;
        RECT 24.850 153.815 25.140 153.860 ;
        RECT 20.210 153.675 25.140 153.815 ;
        RECT 20.210 153.630 20.500 153.675 ;
        RECT 22.990 153.630 23.280 153.675 ;
        RECT 24.850 153.630 25.140 153.675 ;
        RECT 24.380 153.275 24.700 153.535 ;
        RECT 25.315 153.475 25.605 153.520 ;
        RECT 25.760 153.475 26.080 153.535 ;
        RECT 25.315 153.335 26.080 153.475 ;
        RECT 25.315 153.290 25.605 153.335 ;
        RECT 25.760 153.275 26.080 153.335 ;
        RECT 29.440 153.275 29.760 153.535 ;
        RECT 20.210 153.135 20.500 153.180 ;
        RECT 20.210 152.995 22.745 153.135 ;
        RECT 20.210 152.950 20.500 152.995 ;
        RECT 18.350 152.795 18.640 152.840 ;
        RECT 19.320 152.795 19.640 152.855 ;
        RECT 22.530 152.840 22.745 152.995 ;
        RECT 23.460 152.935 23.780 153.195 ;
        RECT 24.470 153.135 24.610 153.275 ;
        RECT 26.695 153.135 26.985 153.180 ;
        RECT 24.470 152.995 26.985 153.135 ;
        RECT 26.695 152.950 26.985 152.995 ;
        RECT 28.980 152.935 29.300 153.195 ;
        RECT 32.290 153.180 32.430 154.015 ;
        RECT 34.500 153.955 34.820 154.015 ;
        RECT 36.340 153.955 36.660 154.015 ;
        RECT 37.720 154.155 38.040 154.215 ;
        RECT 38.655 154.155 38.945 154.200 ;
        RECT 37.720 154.015 38.945 154.155 ;
        RECT 37.720 153.955 38.040 154.015 ;
        RECT 38.655 153.970 38.945 154.015 ;
        RECT 44.175 154.155 44.465 154.200 ;
        RECT 45.080 154.155 45.400 154.215 ;
        RECT 57.515 154.155 57.805 154.200 ;
        RECT 44.175 154.015 45.400 154.155 ;
        RECT 44.175 153.970 44.465 154.015 ;
        RECT 45.080 153.955 45.400 154.015 ;
        RECT 48.850 154.015 57.805 154.155 ;
        RECT 36.800 153.815 37.120 153.875 ;
        RECT 40.955 153.815 41.245 153.860 ;
        RECT 36.800 153.675 41.245 153.815 ;
        RECT 36.800 153.615 37.120 153.675 ;
        RECT 40.955 153.630 41.245 153.675 ;
        RECT 43.240 153.815 43.560 153.875 ;
        RECT 44.620 153.815 44.940 153.875 ;
        RECT 48.315 153.815 48.605 153.860 ;
        RECT 43.240 153.675 44.940 153.815 ;
        RECT 43.240 153.615 43.560 153.675 ;
        RECT 44.620 153.615 44.940 153.675 ;
        RECT 45.170 153.675 48.605 153.815 ;
        RECT 38.180 153.475 38.500 153.535 ;
        RECT 34.590 153.335 38.500 153.475 ;
        RECT 32.215 152.950 32.505 153.180 ;
        RECT 32.660 152.935 32.980 153.195 ;
        RECT 33.120 152.935 33.440 153.195 ;
        RECT 33.580 153.135 33.900 153.195 ;
        RECT 34.590 153.180 34.730 153.335 ;
        RECT 38.180 153.275 38.500 153.335 ;
        RECT 39.100 153.275 39.420 153.535 ;
        RECT 43.700 153.275 44.020 153.535 ;
        RECT 44.160 153.475 44.480 153.535 ;
        RECT 45.170 153.520 45.310 153.675 ;
        RECT 48.315 153.630 48.605 153.675 ;
        RECT 45.095 153.475 45.385 153.520 ;
        RECT 48.850 153.475 48.990 154.015 ;
        RECT 57.515 153.970 57.805 154.015 ;
        RECT 63.020 154.155 63.340 154.215 ;
        RECT 68.095 154.155 68.385 154.200 ;
        RECT 63.020 154.015 68.385 154.155 ;
        RECT 63.020 153.955 63.340 154.015 ;
        RECT 68.095 153.970 68.385 154.015 ;
        RECT 68.540 154.155 68.860 154.215 ;
        RECT 70.380 154.155 70.700 154.215 ;
        RECT 93.380 154.155 93.700 154.215 ;
        RECT 96.155 154.155 96.445 154.200 ;
        RECT 68.540 154.015 71.530 154.155 ;
        RECT 68.540 153.955 68.860 154.015 ;
        RECT 70.380 153.955 70.700 154.015 ;
        RECT 51.175 153.815 51.465 153.860 ;
        RECT 54.295 153.815 54.585 153.860 ;
        RECT 56.185 153.815 56.475 153.860 ;
        RECT 59.800 153.815 60.120 153.875 ;
        RECT 51.175 153.675 56.475 153.815 ;
        RECT 51.175 153.630 51.465 153.675 ;
        RECT 54.295 153.630 54.585 153.675 ;
        RECT 56.185 153.630 56.475 153.675 ;
        RECT 57.130 153.675 60.120 153.815 ;
        RECT 44.160 153.335 45.385 153.475 ;
        RECT 44.160 153.275 44.480 153.335 ;
        RECT 45.095 153.290 45.385 153.335 ;
        RECT 45.630 153.335 48.990 153.475 ;
        RECT 34.055 153.135 34.345 153.180 ;
        RECT 33.580 152.995 34.345 153.135 ;
        RECT 33.580 152.935 33.900 152.995 ;
        RECT 34.055 152.950 34.345 152.995 ;
        RECT 34.515 152.950 34.805 153.180 ;
        RECT 35.420 152.935 35.740 153.195 ;
        RECT 35.880 152.935 36.200 153.195 ;
        RECT 36.340 152.935 36.660 153.195 ;
        RECT 37.260 153.135 37.580 153.195 ;
        RECT 38.655 153.135 38.945 153.180 ;
        RECT 37.260 152.995 38.945 153.135 ;
        RECT 37.260 152.935 37.580 152.995 ;
        RECT 38.655 152.950 38.945 152.995 ;
        RECT 40.035 153.135 40.325 153.180 ;
        RECT 40.940 153.135 41.260 153.195 ;
        RECT 40.035 152.995 41.260 153.135 ;
        RECT 40.035 152.950 40.325 152.995 ;
        RECT 40.940 152.935 41.260 152.995 ;
        RECT 42.780 152.935 43.100 153.195 ;
        RECT 45.630 153.135 45.770 153.335 ;
        RECT 55.660 153.275 55.980 153.535 ;
        RECT 43.790 152.995 45.770 153.135 ;
        RECT 47.855 153.135 48.145 153.180 ;
        RECT 48.300 153.135 48.620 153.195 ;
        RECT 57.130 153.180 57.270 153.675 ;
        RECT 59.800 153.615 60.120 153.675 ;
        RECT 60.720 153.815 61.040 153.875 ;
        RECT 62.115 153.815 62.405 153.860 ;
        RECT 60.720 153.675 70.150 153.815 ;
        RECT 60.720 153.615 61.040 153.675 ;
        RECT 62.115 153.630 62.405 153.675 ;
        RECT 58.420 153.475 58.740 153.535 ;
        RECT 64.415 153.475 64.705 153.520 ;
        RECT 58.420 153.335 64.705 153.475 ;
        RECT 58.420 153.275 58.740 153.335 ;
        RECT 47.855 152.995 48.620 153.135 ;
        RECT 21.610 152.795 21.900 152.840 ;
        RECT 18.350 152.655 21.900 152.795 ;
        RECT 18.350 152.610 18.640 152.655 ;
        RECT 19.320 152.595 19.640 152.655 ;
        RECT 21.610 152.610 21.900 152.655 ;
        RECT 22.530 152.795 22.820 152.840 ;
        RECT 24.390 152.795 24.680 152.840 ;
        RECT 22.530 152.655 24.680 152.795 ;
        RECT 22.530 152.610 22.820 152.655 ;
        RECT 24.390 152.610 24.680 152.655 ;
        RECT 30.375 152.795 30.665 152.840 ;
        RECT 43.790 152.795 43.930 152.995 ;
        RECT 47.855 152.950 48.145 152.995 ;
        RECT 48.300 152.935 48.620 152.995 ;
        RECT 30.375 152.655 43.930 152.795 ;
        RECT 44.175 152.795 44.465 152.840 ;
        RECT 44.620 152.795 44.940 152.855 ;
        RECT 44.175 152.655 44.940 152.795 ;
        RECT 30.375 152.610 30.665 152.655 ;
        RECT 44.175 152.610 44.465 152.655 ;
        RECT 44.620 152.595 44.940 152.655 ;
        RECT 46.460 152.795 46.780 152.855 ;
        RECT 50.095 152.840 50.385 153.155 ;
        RECT 51.175 153.135 51.465 153.180 ;
        RECT 54.755 153.135 55.045 153.180 ;
        RECT 56.590 153.135 56.880 153.180 ;
        RECT 51.175 152.995 56.880 153.135 ;
        RECT 51.175 152.950 51.465 152.995 ;
        RECT 54.755 152.950 55.045 152.995 ;
        RECT 56.590 152.950 56.880 152.995 ;
        RECT 57.055 152.950 57.345 153.180 ;
        RECT 58.895 152.950 59.185 153.180 ;
        RECT 49.795 152.795 50.385 152.840 ;
        RECT 53.035 152.795 53.685 152.840 ;
        RECT 57.130 152.795 57.270 152.950 ;
        RECT 46.460 152.655 53.685 152.795 ;
        RECT 46.460 152.595 46.780 152.655 ;
        RECT 49.795 152.610 50.085 152.655 ;
        RECT 53.035 152.610 53.685 152.655 ;
        RECT 56.670 152.655 57.270 152.795 ;
        RECT 58.420 152.795 58.740 152.855 ;
        RECT 58.970 152.795 59.110 152.950 ;
        RECT 59.340 152.935 59.660 153.195 ;
        RECT 59.890 153.180 60.030 153.335 ;
        RECT 64.415 153.290 64.705 153.335 ;
        RECT 67.160 153.475 67.480 153.535 ;
        RECT 67.160 153.335 69.690 153.475 ;
        RECT 67.160 153.275 67.480 153.335 ;
        RECT 59.815 152.950 60.105 153.180 ;
        RECT 60.260 153.135 60.580 153.195 ;
        RECT 60.735 153.135 61.025 153.180 ;
        RECT 60.260 152.995 61.025 153.135 ;
        RECT 60.260 152.935 60.580 152.995 ;
        RECT 60.735 152.950 61.025 152.995 ;
        RECT 61.180 153.135 61.500 153.195 ;
        RECT 69.550 153.180 69.690 153.335 ;
        RECT 70.010 153.180 70.150 153.675 ;
        RECT 69.015 153.135 69.305 153.180 ;
        RECT 61.180 152.995 69.305 153.135 ;
        RECT 61.180 152.935 61.500 152.995 ;
        RECT 69.015 152.950 69.305 152.995 ;
        RECT 69.475 152.950 69.765 153.180 ;
        RECT 69.935 152.950 70.225 153.180 ;
        RECT 70.855 152.950 71.145 153.180 ;
        RECT 71.390 153.135 71.530 154.015 ;
        RECT 93.380 154.015 96.445 154.155 ;
        RECT 93.380 153.955 93.700 154.015 ;
        RECT 96.155 153.970 96.445 154.015 ;
        RECT 97.060 154.155 97.380 154.215 ;
        RECT 100.280 154.155 100.600 154.215 ;
        RECT 97.060 154.015 100.600 154.155 ;
        RECT 97.060 153.955 97.380 154.015 ;
        RECT 100.280 153.955 100.600 154.015 ;
        RECT 104.880 153.955 105.200 154.215 ;
        RECT 98.440 153.815 98.760 153.875 ;
        RECT 105.340 153.815 105.660 153.875 ;
        RECT 78.750 153.675 98.210 153.815 ;
        RECT 73.155 153.475 73.445 153.520 ;
        RECT 76.360 153.475 76.680 153.535 ;
        RECT 78.750 153.520 78.890 153.675 ;
        RECT 85.190 153.520 85.330 153.675 ;
        RECT 78.675 153.475 78.965 153.520 ;
        RECT 73.155 153.335 78.965 153.475 ;
        RECT 73.155 153.290 73.445 153.335 ;
        RECT 76.360 153.275 76.680 153.335 ;
        RECT 78.675 153.290 78.965 153.335 ;
        RECT 79.135 153.475 79.425 153.520 ;
        RECT 79.135 153.335 83.030 153.475 ;
        RECT 79.135 153.290 79.425 153.335 ;
        RECT 74.075 153.135 74.365 153.180 ;
        RECT 71.390 152.995 74.365 153.135 ;
        RECT 74.075 152.950 74.365 152.995 ;
        RECT 77.295 152.950 77.585 153.180 ;
        RECT 78.200 153.135 78.520 153.195 ;
        RECT 79.210 153.135 79.350 153.290 ;
        RECT 82.355 153.135 82.645 153.180 ;
        RECT 78.200 152.995 79.350 153.135 ;
        RECT 81.510 152.995 82.645 153.135 ;
        RECT 82.890 153.135 83.030 153.335 ;
        RECT 85.115 153.290 85.405 153.520 ;
        RECT 96.140 153.475 96.460 153.535 ;
        RECT 94.390 153.335 96.460 153.475 ;
        RECT 98.070 153.475 98.210 153.675 ;
        RECT 98.440 153.675 105.660 153.815 ;
        RECT 98.440 153.615 98.760 153.675 ;
        RECT 105.340 153.615 105.660 153.675 ;
        RECT 108.215 153.815 108.505 153.860 ;
        RECT 111.335 153.815 111.625 153.860 ;
        RECT 113.225 153.815 113.515 153.860 ;
        RECT 108.215 153.675 113.515 153.815 ;
        RECT 108.215 153.630 108.505 153.675 ;
        RECT 111.335 153.630 111.625 153.675 ;
        RECT 113.225 153.630 113.515 153.675 ;
        RECT 101.675 153.475 101.965 153.520 ;
        RECT 103.500 153.475 103.820 153.535 ;
        RECT 98.070 153.335 103.820 153.475 ;
        RECT 86.495 153.135 86.785 153.180 ;
        RECT 82.890 152.995 86.785 153.135 ;
        RECT 58.420 152.655 59.110 152.795 ;
        RECT 16.345 152.455 16.635 152.500 ;
        RECT 23.000 152.455 23.320 152.515 ;
        RECT 16.345 152.315 23.320 152.455 ;
        RECT 16.345 152.270 16.635 152.315 ;
        RECT 23.000 152.255 23.320 152.315 ;
        RECT 24.840 152.455 25.160 152.515 ;
        RECT 28.075 152.455 28.365 152.500 ;
        RECT 24.840 152.315 28.365 152.455 ;
        RECT 24.840 152.255 25.160 152.315 ;
        RECT 28.075 152.270 28.365 152.315 ;
        RECT 30.835 152.455 31.125 152.500 ;
        RECT 31.280 152.455 31.600 152.515 ;
        RECT 30.835 152.315 31.600 152.455 ;
        RECT 30.835 152.270 31.125 152.315 ;
        RECT 31.280 152.255 31.600 152.315 ;
        RECT 37.735 152.455 38.025 152.500 ;
        RECT 39.560 152.455 39.880 152.515 ;
        RECT 37.735 152.315 39.880 152.455 ;
        RECT 37.735 152.270 38.025 152.315 ;
        RECT 39.560 152.255 39.880 152.315 ;
        RECT 41.860 152.255 42.180 152.515 ;
        RECT 47.840 152.455 48.160 152.515 ;
        RECT 56.670 152.455 56.810 152.655 ;
        RECT 58.420 152.595 58.740 152.655 ;
        RECT 63.035 152.610 63.325 152.840 ;
        RECT 67.635 152.795 67.925 152.840 ;
        RECT 70.930 152.795 71.070 152.950 ;
        RECT 67.635 152.655 71.070 152.795 ;
        RECT 67.635 152.610 67.925 152.655 ;
        RECT 71.775 152.610 72.065 152.840 ;
        RECT 77.370 152.795 77.510 152.950 ;
        RECT 78.200 152.935 78.520 152.995 ;
        RECT 79.120 152.795 79.440 152.855 ;
        RECT 77.370 152.655 79.440 152.795 ;
        RECT 47.840 152.315 56.810 152.455 ;
        RECT 63.110 152.455 63.250 152.610 ;
        RECT 71.300 152.455 71.620 152.515 ;
        RECT 71.850 152.455 71.990 152.610 ;
        RECT 79.120 152.595 79.440 152.655 ;
        RECT 63.110 152.315 71.990 152.455 ;
        RECT 74.995 152.455 75.285 152.500 ;
        RECT 75.440 152.455 75.760 152.515 ;
        RECT 74.995 152.315 75.760 152.455 ;
        RECT 47.840 152.255 48.160 152.315 ;
        RECT 71.300 152.255 71.620 152.315 ;
        RECT 74.995 152.270 75.285 152.315 ;
        RECT 75.440 152.255 75.760 152.315 ;
        RECT 76.820 152.255 77.140 152.515 ;
        RECT 77.740 152.455 78.060 152.515 ;
        RECT 81.510 152.500 81.650 152.995 ;
        RECT 82.355 152.950 82.645 152.995 ;
        RECT 86.495 152.950 86.785 152.995 ;
        RECT 93.840 152.935 94.160 153.195 ;
        RECT 94.390 153.180 94.530 153.335 ;
        RECT 96.140 153.275 96.460 153.335 ;
        RECT 101.675 153.290 101.965 153.335 ;
        RECT 103.500 153.275 103.820 153.335 ;
        RECT 112.700 153.275 113.020 153.535 ;
        RECT 94.315 152.950 94.605 153.180 ;
        RECT 94.775 152.950 95.065 153.180 ;
        RECT 94.850 152.795 94.990 152.950 ;
        RECT 95.680 152.935 96.000 153.195 ;
        RECT 97.060 153.135 97.380 153.195 ;
        RECT 97.535 153.135 97.825 153.180 ;
        RECT 97.060 152.995 97.825 153.135 ;
        RECT 97.060 152.935 97.380 152.995 ;
        RECT 97.535 152.950 97.825 152.995 ;
        RECT 97.980 152.935 98.300 153.195 ;
        RECT 98.440 152.935 98.760 153.195 ;
        RECT 99.360 152.935 99.680 153.195 ;
        RECT 105.800 153.135 106.120 153.195 ;
        RECT 107.180 153.155 107.500 153.195 ;
        RECT 101.750 152.995 106.120 153.135 ;
        RECT 101.750 152.795 101.890 152.995 ;
        RECT 105.800 152.935 106.120 152.995 ;
        RECT 107.135 152.935 107.500 153.155 ;
        RECT 108.215 153.135 108.505 153.180 ;
        RECT 111.795 153.135 112.085 153.180 ;
        RECT 113.630 153.135 113.920 153.180 ;
        RECT 108.215 152.995 113.920 153.135 ;
        RECT 108.215 152.950 108.505 152.995 ;
        RECT 111.795 152.950 112.085 152.995 ;
        RECT 113.630 152.950 113.920 152.995 ;
        RECT 114.095 152.950 114.385 153.180 ;
        RECT 94.850 152.655 101.890 152.795 ;
        RECT 102.120 152.795 102.440 152.855 ;
        RECT 107.135 152.840 107.425 152.935 ;
        RECT 103.055 152.795 103.345 152.840 ;
        RECT 102.120 152.655 103.345 152.795 ;
        RECT 102.120 152.595 102.440 152.655 ;
        RECT 103.055 152.610 103.345 152.655 ;
        RECT 106.835 152.795 107.425 152.840 ;
        RECT 110.075 152.795 110.725 152.840 ;
        RECT 106.835 152.655 110.725 152.795 ;
        RECT 106.835 152.610 107.125 152.655 ;
        RECT 110.075 152.610 110.725 152.655 ;
        RECT 113.160 152.795 113.480 152.855 ;
        RECT 114.170 152.795 114.310 152.950 ;
        RECT 113.160 152.655 114.310 152.795 ;
        RECT 113.160 152.595 113.480 152.655 ;
        RECT 79.595 152.455 79.885 152.500 ;
        RECT 77.740 152.315 79.885 152.455 ;
        RECT 77.740 152.255 78.060 152.315 ;
        RECT 79.595 152.270 79.885 152.315 ;
        RECT 81.435 152.270 81.725 152.500 ;
        RECT 83.275 152.455 83.565 152.500 ;
        RECT 84.640 152.455 84.960 152.515 ;
        RECT 83.275 152.315 84.960 152.455 ;
        RECT 83.275 152.270 83.565 152.315 ;
        RECT 84.640 152.255 84.960 152.315 ;
        RECT 86.020 152.255 86.340 152.515 ;
        RECT 88.335 152.455 88.625 152.500 ;
        RECT 89.240 152.455 89.560 152.515 ;
        RECT 88.335 152.315 89.560 152.455 ;
        RECT 88.335 152.270 88.625 152.315 ;
        RECT 89.240 152.255 89.560 152.315 ;
        RECT 92.475 152.455 92.765 152.500 ;
        RECT 93.840 152.455 94.160 152.515 ;
        RECT 92.475 152.315 94.160 152.455 ;
        RECT 92.475 152.270 92.765 152.315 ;
        RECT 93.840 152.255 94.160 152.315 ;
        RECT 102.595 152.455 102.885 152.500 ;
        RECT 107.640 152.455 107.960 152.515 ;
        RECT 102.595 152.315 107.960 152.455 ;
        RECT 102.595 152.270 102.885 152.315 ;
        RECT 107.640 152.255 107.960 152.315 ;
        RECT 14.650 151.635 115.850 152.115 ;
        RECT 18.860 151.435 19.180 151.495 ;
        RECT 20.255 151.435 20.545 151.480 ;
        RECT 30.835 151.435 31.125 151.480 ;
        RECT 49.220 151.435 49.540 151.495 ;
        RECT 18.860 151.295 20.545 151.435 ;
        RECT 18.860 151.235 19.180 151.295 ;
        RECT 20.255 151.250 20.545 151.295 ;
        RECT 24.010 151.295 36.110 151.435 ;
        RECT 24.010 150.815 24.150 151.295 ;
        RECT 30.835 151.250 31.125 151.295 ;
        RECT 29.900 151.095 30.220 151.155 ;
        RECT 31.295 151.095 31.585 151.140 ;
        RECT 29.900 150.955 31.585 151.095 ;
        RECT 29.900 150.895 30.220 150.955 ;
        RECT 31.295 150.910 31.585 150.955 ;
        RECT 32.660 151.095 32.980 151.155 ;
        RECT 32.660 150.955 35.650 151.095 ;
        RECT 32.660 150.895 32.980 150.955 ;
        RECT 18.860 150.755 19.180 150.815 ;
        RECT 19.795 150.755 20.085 150.800 ;
        RECT 18.860 150.615 20.085 150.755 ;
        RECT 18.860 150.555 19.180 150.615 ;
        RECT 19.795 150.570 20.085 150.615 ;
        RECT 23.015 150.755 23.305 150.800 ;
        RECT 23.920 150.755 24.240 150.815 ;
        RECT 23.015 150.615 24.240 150.755 ;
        RECT 23.015 150.570 23.305 150.615 ;
        RECT 23.920 150.555 24.240 150.615 ;
        RECT 27.140 150.555 27.460 150.815 ;
        RECT 33.120 150.555 33.440 150.815 ;
        RECT 34.500 150.755 34.820 150.815 ;
        RECT 35.510 150.800 35.650 150.955 ;
        RECT 35.970 150.800 36.110 151.295 ;
        RECT 43.330 151.295 49.540 151.435 ;
        RECT 39.115 151.095 39.405 151.140 ;
        RECT 41.875 151.095 42.165 151.140 ;
        RECT 39.115 150.955 42.165 151.095 ;
        RECT 39.115 150.910 39.405 150.955 ;
        RECT 41.875 150.910 42.165 150.955 ;
        RECT 34.975 150.755 35.265 150.800 ;
        RECT 34.500 150.615 35.265 150.755 ;
        RECT 34.500 150.555 34.820 150.615 ;
        RECT 34.975 150.570 35.265 150.615 ;
        RECT 35.435 150.570 35.725 150.800 ;
        RECT 35.895 150.570 36.185 150.800 ;
        RECT 36.800 150.555 37.120 150.815 ;
        RECT 40.020 150.555 40.340 150.815 ;
        RECT 40.480 150.555 40.800 150.815 ;
        RECT 43.330 150.800 43.470 151.295 ;
        RECT 49.220 151.235 49.540 151.295 ;
        RECT 52.455 151.435 52.745 151.480 ;
        RECT 53.820 151.435 54.140 151.495 ;
        RECT 52.455 151.295 54.140 151.435 ;
        RECT 52.455 151.250 52.745 151.295 ;
        RECT 53.820 151.235 54.140 151.295 ;
        RECT 54.280 151.235 54.600 151.495 ;
        RECT 77.525 151.435 77.815 151.480 ;
        RECT 78.200 151.435 78.520 151.495 ;
        RECT 75.070 151.295 78.520 151.435 ;
        RECT 46.460 151.095 46.780 151.155 ;
        RECT 46.935 151.095 47.225 151.140 ;
        RECT 46.460 150.955 47.225 151.095 ;
        RECT 46.460 150.895 46.780 150.955 ;
        RECT 46.935 150.910 47.225 150.955 ;
        RECT 47.395 151.095 47.685 151.140 ;
        RECT 48.300 151.095 48.620 151.155 ;
        RECT 54.755 151.095 55.045 151.140 ;
        RECT 47.395 150.955 55.045 151.095 ;
        RECT 47.395 150.910 47.685 150.955 ;
        RECT 48.300 150.895 48.620 150.955 ;
        RECT 54.755 150.910 55.045 150.955 ;
        RECT 61.590 151.095 61.880 151.140 ;
        RECT 63.020 151.095 63.340 151.155 ;
        RECT 64.850 151.095 65.140 151.140 ;
        RECT 61.590 150.955 65.140 151.095 ;
        RECT 61.590 150.910 61.880 150.955 ;
        RECT 63.020 150.895 63.340 150.955 ;
        RECT 64.850 150.910 65.140 150.955 ;
        RECT 65.770 151.095 66.060 151.140 ;
        RECT 67.630 151.095 67.920 151.140 ;
        RECT 65.770 150.955 67.920 151.095 ;
        RECT 65.770 150.910 66.060 150.955 ;
        RECT 67.630 150.910 67.920 150.955 ;
        RECT 72.235 151.095 72.525 151.140 ;
        RECT 72.695 151.095 72.985 151.140 ;
        RECT 72.235 150.955 72.985 151.095 ;
        RECT 72.235 150.910 72.525 150.955 ;
        RECT 72.695 150.910 72.985 150.955 ;
        RECT 43.255 150.570 43.545 150.800 ;
        RECT 43.715 150.570 44.005 150.800 ;
        RECT 23.475 150.230 23.765 150.460 ;
        RECT 24.395 150.415 24.685 150.460 ;
        RECT 28.520 150.415 28.840 150.475 ;
        RECT 29.915 150.415 30.205 150.460 ;
        RECT 33.210 150.415 33.350 150.555 ;
        RECT 24.395 150.275 30.205 150.415 ;
        RECT 24.395 150.230 24.685 150.275 ;
        RECT 23.000 150.075 23.320 150.135 ;
        RECT 23.550 150.075 23.690 150.230 ;
        RECT 28.520 150.215 28.840 150.275 ;
        RECT 29.915 150.230 30.205 150.275 ;
        RECT 30.450 150.275 33.350 150.415 ;
        RECT 43.790 150.415 43.930 150.570 ;
        RECT 44.160 150.555 44.480 150.815 ;
        RECT 45.095 150.755 45.385 150.800 ;
        RECT 48.760 150.755 49.080 150.815 ;
        RECT 45.095 150.615 49.080 150.755 ;
        RECT 45.095 150.570 45.385 150.615 ;
        RECT 48.760 150.555 49.080 150.615 ;
        RECT 63.450 150.755 63.740 150.800 ;
        RECT 65.770 150.755 65.985 150.910 ;
        RECT 63.450 150.615 65.985 150.755 ;
        RECT 70.855 150.755 71.145 150.800 ;
        RECT 71.760 150.755 72.080 150.815 ;
        RECT 70.855 150.615 72.080 150.755 ;
        RECT 63.450 150.570 63.740 150.615 ;
        RECT 70.855 150.570 71.145 150.615 ;
        RECT 71.760 150.555 72.080 150.615 ;
        RECT 74.060 150.555 74.380 150.815 ;
        RECT 74.520 150.555 74.840 150.815 ;
        RECT 75.070 150.800 75.210 151.295 ;
        RECT 77.525 151.250 77.815 151.295 ;
        RECT 78.200 151.235 78.520 151.295 ;
        RECT 86.020 151.435 86.340 151.495 ;
        RECT 99.375 151.435 99.665 151.480 ;
        RECT 102.120 151.435 102.440 151.495 ;
        RECT 86.020 151.295 102.440 151.435 ;
        RECT 86.020 151.235 86.340 151.295 ;
        RECT 99.375 151.250 99.665 151.295 ;
        RECT 102.120 151.235 102.440 151.295 ;
        RECT 107.195 151.435 107.485 151.480 ;
        RECT 107.640 151.435 107.960 151.495 ;
        RECT 109.495 151.435 109.785 151.480 ;
        RECT 107.195 151.295 109.785 151.435 ;
        RECT 107.195 151.250 107.485 151.295 ;
        RECT 107.640 151.235 107.960 151.295 ;
        RECT 109.495 151.250 109.785 151.295 ;
        RECT 76.820 151.095 77.140 151.155 ;
        RECT 79.530 151.095 79.820 151.140 ;
        RECT 82.790 151.095 83.080 151.140 ;
        RECT 76.820 150.955 83.080 151.095 ;
        RECT 76.820 150.895 77.140 150.955 ;
        RECT 79.530 150.910 79.820 150.955 ;
        RECT 82.790 150.910 83.080 150.955 ;
        RECT 83.710 151.095 84.000 151.140 ;
        RECT 85.570 151.095 85.860 151.140 ;
        RECT 83.710 150.955 85.860 151.095 ;
        RECT 83.710 150.910 84.000 150.955 ;
        RECT 85.570 150.910 85.860 150.955 ;
        RECT 87.860 151.095 88.180 151.155 ;
        RECT 90.615 151.095 91.265 151.140 ;
        RECT 94.215 151.095 94.505 151.140 ;
        RECT 87.860 150.955 94.505 151.095 ;
        RECT 74.995 150.570 75.285 150.800 ;
        RECT 75.440 150.755 75.760 150.815 ;
        RECT 75.915 150.755 76.205 150.800 ;
        RECT 75.440 150.615 76.205 150.755 ;
        RECT 75.440 150.555 75.760 150.615 ;
        RECT 75.915 150.570 76.205 150.615 ;
        RECT 81.390 150.755 81.680 150.800 ;
        RECT 83.710 150.755 83.925 150.910 ;
        RECT 87.860 150.895 88.180 150.955 ;
        RECT 90.615 150.910 91.265 150.955 ;
        RECT 93.915 150.910 94.505 150.955 ;
        RECT 81.390 150.615 83.925 150.755 ;
        RECT 81.390 150.570 81.680 150.615 ;
        RECT 84.640 150.555 84.960 150.815 ;
        RECT 87.420 150.755 87.710 150.800 ;
        RECT 89.255 150.755 89.545 150.800 ;
        RECT 92.835 150.755 93.125 150.800 ;
        RECT 87.420 150.615 93.125 150.755 ;
        RECT 87.420 150.570 87.710 150.615 ;
        RECT 89.255 150.570 89.545 150.615 ;
        RECT 92.835 150.570 93.125 150.615 ;
        RECT 93.915 150.595 94.205 150.910 ;
        RECT 99.820 150.895 100.140 151.155 ;
        RECT 101.200 150.555 101.520 150.815 ;
        RECT 105.340 150.755 105.660 150.815 ;
        RECT 112.255 150.755 112.545 150.800 ;
        RECT 105.340 150.615 112.545 150.755 ;
        RECT 105.340 150.555 105.660 150.615 ;
        RECT 112.255 150.570 112.545 150.615 ;
        RECT 114.095 150.570 114.385 150.800 ;
        RECT 45.540 150.415 45.860 150.475 ;
        RECT 43.790 150.275 45.860 150.415 ;
        RECT 30.450 150.075 30.590 150.275 ;
        RECT 45.540 150.215 45.860 150.275 ;
        RECT 46.475 150.415 46.765 150.460 ;
        RECT 55.215 150.415 55.505 150.460 ;
        RECT 59.340 150.415 59.660 150.475 ;
        RECT 60.720 150.415 61.040 150.475 ;
        RECT 46.475 150.275 61.040 150.415 ;
        RECT 46.475 150.230 46.765 150.275 ;
        RECT 55.215 150.230 55.505 150.275 ;
        RECT 59.340 150.215 59.660 150.275 ;
        RECT 60.720 150.215 61.040 150.275 ;
        RECT 65.320 150.415 65.640 150.475 ;
        RECT 66.715 150.415 67.005 150.460 ;
        RECT 65.320 150.275 67.005 150.415 ;
        RECT 65.320 150.215 65.640 150.275 ;
        RECT 66.715 150.230 67.005 150.275 ;
        RECT 68.540 150.215 68.860 150.475 ;
        RECT 69.920 150.415 70.240 150.475 ;
        RECT 71.315 150.415 71.605 150.460 ;
        RECT 69.920 150.275 71.605 150.415 ;
        RECT 69.920 150.215 70.240 150.275 ;
        RECT 71.315 150.230 71.605 150.275 ;
        RECT 86.480 150.415 86.800 150.475 ;
        RECT 86.955 150.415 87.245 150.460 ;
        RECT 86.480 150.275 87.245 150.415 ;
        RECT 86.480 150.215 86.800 150.275 ;
        RECT 86.955 150.230 87.245 150.275 ;
        RECT 88.320 150.215 88.640 150.475 ;
        RECT 95.695 150.415 95.985 150.460 ;
        RECT 96.155 150.415 96.445 150.460 ;
        RECT 98.440 150.415 98.760 150.475 ;
        RECT 95.695 150.275 98.760 150.415 ;
        RECT 95.695 150.230 95.985 150.275 ;
        RECT 96.155 150.230 96.445 150.275 ;
        RECT 98.440 150.215 98.760 150.275 ;
        RECT 100.755 150.415 101.045 150.460 ;
        RECT 103.040 150.415 103.360 150.475 ;
        RECT 100.755 150.275 103.360 150.415 ;
        RECT 100.755 150.230 101.045 150.275 ;
        RECT 103.040 150.215 103.360 150.275 ;
        RECT 103.500 150.415 103.820 150.475 ;
        RECT 105.815 150.415 106.105 150.460 ;
        RECT 103.500 150.275 106.105 150.415 ;
        RECT 103.500 150.215 103.820 150.275 ;
        RECT 105.815 150.230 106.105 150.275 ;
        RECT 106.720 150.215 107.040 150.475 ;
        RECT 114.170 150.415 114.310 150.570 ;
        RECT 109.110 150.275 114.310 150.415 ;
        RECT 23.000 149.935 30.590 150.075 ;
        RECT 33.135 150.075 33.425 150.120 ;
        RECT 34.500 150.075 34.820 150.135 ;
        RECT 33.135 149.935 34.820 150.075 ;
        RECT 23.000 149.875 23.320 149.935 ;
        RECT 33.135 149.890 33.425 149.935 ;
        RECT 34.500 149.875 34.820 149.935 ;
        RECT 41.415 150.075 41.705 150.120 ;
        RECT 62.100 150.075 62.420 150.135 ;
        RECT 109.110 150.120 109.250 150.275 ;
        RECT 41.415 149.935 62.420 150.075 ;
        RECT 41.415 149.890 41.705 149.935 ;
        RECT 62.100 149.875 62.420 149.935 ;
        RECT 63.450 150.075 63.740 150.120 ;
        RECT 66.230 150.075 66.520 150.120 ;
        RECT 68.090 150.075 68.380 150.120 ;
        RECT 63.450 149.935 68.380 150.075 ;
        RECT 63.450 149.890 63.740 149.935 ;
        RECT 66.230 149.890 66.520 149.935 ;
        RECT 68.090 149.890 68.380 149.935 ;
        RECT 81.390 150.075 81.680 150.120 ;
        RECT 84.170 150.075 84.460 150.120 ;
        RECT 86.030 150.075 86.320 150.120 ;
        RECT 81.390 149.935 86.320 150.075 ;
        RECT 81.390 149.890 81.680 149.935 ;
        RECT 84.170 149.890 84.460 149.935 ;
        RECT 86.030 149.890 86.320 149.935 ;
        RECT 87.825 150.075 88.115 150.120 ;
        RECT 89.715 150.075 90.005 150.120 ;
        RECT 92.835 150.075 93.125 150.120 ;
        RECT 87.825 149.935 93.125 150.075 ;
        RECT 87.825 149.890 88.115 149.935 ;
        RECT 89.715 149.890 90.005 149.935 ;
        RECT 92.835 149.890 93.125 149.935 ;
        RECT 109.035 149.890 109.325 150.120 ;
        RECT 21.175 149.735 21.465 149.780 ;
        RECT 22.540 149.735 22.860 149.795 ;
        RECT 21.175 149.595 22.860 149.735 ;
        RECT 21.175 149.550 21.465 149.595 ;
        RECT 22.540 149.535 22.860 149.595 ;
        RECT 27.600 149.535 27.920 149.795 ;
        RECT 33.580 149.535 33.900 149.795 ;
        RECT 38.180 149.735 38.500 149.795 ;
        RECT 39.115 149.735 39.405 149.780 ;
        RECT 38.180 149.595 39.405 149.735 ;
        RECT 38.180 149.535 38.500 149.595 ;
        RECT 39.115 149.550 39.405 149.595 ;
        RECT 40.480 149.735 40.800 149.795 ;
        RECT 46.920 149.735 47.240 149.795 ;
        RECT 40.480 149.595 47.240 149.735 ;
        RECT 40.480 149.535 40.800 149.595 ;
        RECT 46.920 149.535 47.240 149.595 ;
        RECT 49.235 149.735 49.525 149.780 ;
        RECT 51.980 149.735 52.300 149.795 ;
        RECT 49.235 149.595 52.300 149.735 ;
        RECT 49.235 149.550 49.525 149.595 ;
        RECT 51.980 149.535 52.300 149.595 ;
        RECT 58.880 149.735 59.200 149.795 ;
        RECT 59.585 149.735 59.875 149.780 ;
        RECT 58.880 149.595 59.875 149.735 ;
        RECT 58.880 149.535 59.200 149.595 ;
        RECT 59.585 149.550 59.875 149.595 ;
        RECT 69.920 149.535 70.240 149.795 ;
        RECT 72.220 149.535 72.540 149.795 ;
        RECT 99.820 149.535 100.140 149.795 ;
        RECT 102.135 149.735 102.425 149.780 ;
        RECT 108.560 149.735 108.880 149.795 ;
        RECT 102.135 149.595 108.880 149.735 ;
        RECT 102.135 149.550 102.425 149.595 ;
        RECT 108.560 149.535 108.880 149.595 ;
        RECT 112.240 149.735 112.560 149.795 ;
        RECT 113.175 149.735 113.465 149.780 ;
        RECT 112.240 149.595 113.465 149.735 ;
        RECT 112.240 149.535 112.560 149.595 ;
        RECT 113.175 149.550 113.465 149.595 ;
        RECT 14.650 148.915 115.850 149.395 ;
        RECT 23.460 148.515 23.780 148.775 ;
        RECT 23.920 148.760 24.240 148.775 ;
        RECT 23.920 148.530 24.455 148.760 ;
        RECT 40.940 148.715 41.260 148.775 ;
        RECT 61.180 148.715 61.500 148.775 ;
        RECT 40.940 148.575 61.500 148.715 ;
        RECT 23.920 148.515 24.240 148.530 ;
        RECT 40.940 148.515 41.260 148.575 ;
        RECT 61.180 148.515 61.500 148.575 ;
        RECT 63.020 148.515 63.340 148.775 ;
        RECT 65.320 148.515 65.640 148.775 ;
        RECT 69.935 148.715 70.225 148.760 ;
        RECT 69.935 148.575 71.070 148.715 ;
        RECT 69.935 148.530 70.225 148.575 ;
        RECT 28.030 148.375 28.320 148.420 ;
        RECT 30.810 148.375 31.100 148.420 ;
        RECT 32.670 148.375 32.960 148.420 ;
        RECT 28.030 148.235 32.960 148.375 ;
        RECT 28.030 148.190 28.320 148.235 ;
        RECT 30.810 148.190 31.100 148.235 ;
        RECT 32.670 148.190 32.960 148.235 ;
        RECT 33.595 148.190 33.885 148.420 ;
        RECT 42.750 148.375 43.040 148.420 ;
        RECT 45.530 148.375 45.820 148.420 ;
        RECT 47.390 148.375 47.680 148.420 ;
        RECT 48.300 148.375 48.620 148.435 ;
        RECT 42.750 148.235 47.680 148.375 ;
        RECT 42.750 148.190 43.040 148.235 ;
        RECT 45.530 148.190 45.820 148.235 ;
        RECT 47.390 148.190 47.680 148.235 ;
        RECT 47.930 148.235 48.620 148.375 ;
        RECT 19.320 148.035 19.640 148.095 ;
        RECT 20.255 148.035 20.545 148.080 ;
        RECT 19.320 147.895 20.545 148.035 ;
        RECT 19.320 147.835 19.640 147.895 ;
        RECT 20.255 147.850 20.545 147.895 ;
        RECT 25.760 148.035 26.080 148.095 ;
        RECT 31.295 148.035 31.585 148.080 ;
        RECT 33.670 148.035 33.810 148.190 ;
        RECT 25.760 147.895 31.050 148.035 ;
        RECT 25.760 147.835 26.080 147.895 ;
        RECT 18.860 147.695 19.180 147.755 ;
        RECT 20.715 147.695 21.005 147.740 ;
        RECT 18.860 147.555 22.310 147.695 ;
        RECT 18.860 147.495 19.180 147.555 ;
        RECT 20.715 147.510 21.005 147.555 ;
        RECT 22.170 147.015 22.310 147.555 ;
        RECT 22.540 147.495 22.860 147.755 ;
        RECT 28.030 147.695 28.320 147.740 ;
        RECT 30.910 147.695 31.050 147.895 ;
        RECT 31.295 147.895 33.810 148.035 ;
        RECT 38.885 148.035 39.175 148.080 ;
        RECT 42.320 148.035 42.640 148.095 ;
        RECT 46.460 148.035 46.780 148.095 ;
        RECT 47.930 148.080 48.070 148.235 ;
        RECT 48.300 148.175 48.620 148.235 ;
        RECT 57.500 148.375 57.820 148.435 ;
        RECT 59.800 148.375 60.120 148.435 ;
        RECT 57.500 148.235 60.120 148.375 ;
        RECT 57.500 148.175 57.820 148.235 ;
        RECT 59.800 148.175 60.120 148.235 ;
        RECT 66.700 148.175 67.020 148.435 ;
        RECT 38.885 147.895 46.780 148.035 ;
        RECT 31.295 147.850 31.585 147.895 ;
        RECT 38.885 147.850 39.175 147.895 ;
        RECT 42.320 147.835 42.640 147.895 ;
        RECT 46.460 147.835 46.780 147.895 ;
        RECT 47.820 147.850 48.110 148.080 ;
        RECT 58.420 148.035 58.740 148.095 ;
        RECT 59.890 148.035 60.030 148.175 ;
        RECT 57.590 147.895 58.740 148.035 ;
        RECT 33.135 147.695 33.425 147.740 ;
        RECT 28.030 147.555 30.565 147.695 ;
        RECT 30.910 147.555 33.425 147.695 ;
        RECT 28.030 147.510 28.320 147.555 ;
        RECT 26.170 147.355 26.460 147.400 ;
        RECT 27.600 147.355 27.920 147.415 ;
        RECT 30.350 147.400 30.565 147.555 ;
        RECT 33.135 147.510 33.425 147.555 ;
        RECT 34.500 147.495 34.820 147.755 ;
        RECT 36.815 147.695 37.105 147.740 ;
        RECT 40.020 147.695 40.340 147.755 ;
        RECT 36.815 147.555 40.340 147.695 ;
        RECT 36.815 147.510 37.105 147.555 ;
        RECT 29.430 147.355 29.720 147.400 ;
        RECT 26.170 147.215 29.720 147.355 ;
        RECT 26.170 147.170 26.460 147.215 ;
        RECT 27.600 147.155 27.920 147.215 ;
        RECT 29.430 147.170 29.720 147.215 ;
        RECT 30.350 147.355 30.640 147.400 ;
        RECT 32.210 147.355 32.500 147.400 ;
        RECT 30.350 147.215 32.500 147.355 ;
        RECT 30.350 147.170 30.640 147.215 ;
        RECT 32.210 147.170 32.500 147.215 ;
        RECT 27.140 147.015 27.460 147.075 ;
        RECT 36.890 147.015 37.030 147.510 ;
        RECT 40.020 147.495 40.340 147.555 ;
        RECT 42.750 147.695 43.040 147.740 ;
        RECT 46.015 147.695 46.305 147.740 ;
        RECT 49.220 147.695 49.540 147.755 ;
        RECT 49.695 147.695 49.985 147.740 ;
        RECT 42.750 147.555 45.285 147.695 ;
        RECT 42.750 147.510 43.040 147.555 ;
        RECT 45.070 147.400 45.285 147.555 ;
        RECT 46.015 147.555 48.990 147.695 ;
        RECT 46.015 147.510 46.305 147.555 ;
        RECT 37.275 147.355 37.565 147.400 ;
        RECT 40.890 147.355 41.180 147.400 ;
        RECT 44.150 147.355 44.440 147.400 ;
        RECT 37.275 147.215 44.440 147.355 ;
        RECT 37.275 147.170 37.565 147.215 ;
        RECT 40.890 147.170 41.180 147.215 ;
        RECT 44.150 147.170 44.440 147.215 ;
        RECT 45.070 147.355 45.360 147.400 ;
        RECT 46.930 147.355 47.220 147.400 ;
        RECT 45.070 147.215 47.220 147.355 ;
        RECT 48.850 147.355 48.990 147.555 ;
        RECT 49.220 147.555 49.985 147.695 ;
        RECT 49.220 147.495 49.540 147.555 ;
        RECT 49.695 147.510 49.985 147.555 ;
        RECT 50.140 147.495 50.460 147.755 ;
        RECT 50.600 147.495 50.920 147.755 ;
        RECT 51.520 147.495 51.840 147.755 ;
        RECT 52.440 147.695 52.760 147.755 ;
        RECT 52.915 147.695 53.205 147.740 ;
        RECT 52.440 147.555 53.205 147.695 ;
        RECT 52.440 147.495 52.760 147.555 ;
        RECT 52.915 147.510 53.205 147.555 ;
        RECT 57.590 147.355 57.730 147.895 ;
        RECT 58.420 147.835 58.740 147.895 ;
        RECT 59.430 147.895 60.030 148.035 ;
        RECT 57.960 147.495 58.280 147.755 ;
        RECT 58.880 147.680 59.200 147.765 ;
        RECT 59.430 147.740 59.570 147.895 ;
        RECT 61.180 147.835 61.500 148.095 ;
        RECT 68.080 148.035 68.400 148.095 ;
        RECT 70.380 148.035 70.700 148.095 ;
        RECT 65.870 147.895 68.400 148.035 ;
        RECT 58.710 147.540 59.200 147.680 ;
        RECT 58.880 147.505 59.200 147.540 ;
        RECT 59.355 147.510 59.645 147.740 ;
        RECT 59.915 147.695 60.205 147.740 ;
        RECT 61.640 147.695 61.960 147.755 ;
        RECT 62.575 147.695 62.865 147.740 ;
        RECT 59.915 147.555 60.490 147.695 ;
        RECT 59.915 147.510 60.205 147.555 ;
        RECT 58.895 147.495 59.185 147.505 ;
        RECT 60.350 147.355 60.490 147.555 ;
        RECT 61.640 147.555 62.865 147.695 ;
        RECT 61.640 147.495 61.960 147.555 ;
        RECT 62.575 147.510 62.865 147.555 ;
        RECT 64.400 147.495 64.720 147.755 ;
        RECT 65.870 147.740 66.010 147.895 ;
        RECT 68.080 147.835 68.400 147.895 ;
        RECT 68.630 147.895 70.700 148.035 ;
        RECT 70.930 148.035 71.070 148.575 ;
        RECT 71.300 148.515 71.620 148.775 ;
        RECT 87.415 148.715 87.705 148.760 ;
        RECT 87.860 148.715 88.180 148.775 ;
        RECT 87.415 148.575 88.180 148.715 ;
        RECT 87.415 148.530 87.705 148.575 ;
        RECT 87.860 148.515 88.180 148.575 ;
        RECT 88.320 148.515 88.640 148.775 ;
        RECT 95.235 148.715 95.525 148.760 ;
        RECT 97.060 148.715 97.380 148.775 ;
        RECT 95.235 148.575 97.380 148.715 ;
        RECT 95.235 148.530 95.525 148.575 ;
        RECT 97.060 148.515 97.380 148.575 ;
        RECT 98.440 148.715 98.760 148.775 ;
        RECT 103.040 148.715 103.360 148.775 ;
        RECT 105.125 148.715 105.415 148.760 ;
        RECT 106.720 148.715 107.040 148.775 ;
        RECT 98.440 148.575 107.040 148.715 ;
        RECT 98.440 148.515 98.760 148.575 ;
        RECT 103.040 148.515 103.360 148.575 ;
        RECT 105.125 148.530 105.415 148.575 ;
        RECT 106.720 148.515 107.040 148.575 ;
        RECT 74.060 148.375 74.380 148.435 ;
        RECT 74.980 148.375 75.300 148.435 ;
        RECT 101.200 148.375 101.520 148.435 ;
        RECT 74.060 148.235 75.300 148.375 ;
        RECT 74.060 148.175 74.380 148.235 ;
        RECT 74.980 148.175 75.300 148.235 ;
        RECT 97.150 148.235 101.520 148.375 ;
        RECT 70.930 147.895 71.530 148.035 ;
        RECT 65.795 147.510 66.085 147.740 ;
        RECT 67.635 147.695 67.925 147.740 ;
        RECT 68.630 147.695 68.770 147.895 ;
        RECT 70.380 147.835 70.700 147.895 ;
        RECT 67.635 147.555 68.770 147.695 ;
        RECT 69.000 147.695 69.320 147.755 ;
        RECT 70.855 147.695 71.145 147.740 ;
        RECT 69.000 147.555 71.145 147.695 ;
        RECT 71.390 147.695 71.530 147.895 ;
        RECT 71.760 147.835 72.080 148.095 ;
        RECT 73.600 147.695 73.920 147.755 ;
        RECT 74.150 147.740 74.290 148.175 ;
        RECT 77.740 148.035 78.060 148.095 ;
        RECT 75.070 147.895 78.060 148.035 ;
        RECT 71.390 147.555 73.920 147.695 ;
        RECT 67.635 147.510 67.925 147.555 ;
        RECT 69.000 147.495 69.320 147.555 ;
        RECT 70.855 147.510 71.145 147.555 ;
        RECT 73.600 147.495 73.920 147.555 ;
        RECT 74.075 147.510 74.365 147.740 ;
        RECT 74.520 147.495 74.840 147.755 ;
        RECT 75.070 147.740 75.210 147.895 ;
        RECT 77.740 147.835 78.060 147.895 ;
        RECT 94.760 147.835 95.080 148.095 ;
        RECT 74.995 147.510 75.285 147.740 ;
        RECT 75.440 147.695 75.760 147.755 ;
        RECT 75.915 147.695 76.205 147.740 ;
        RECT 75.440 147.555 76.205 147.695 ;
        RECT 75.440 147.495 75.760 147.555 ;
        RECT 75.915 147.510 76.205 147.555 ;
        RECT 79.120 147.695 79.440 147.755 ;
        RECT 79.595 147.695 79.885 147.740 ;
        RECT 79.120 147.555 79.885 147.695 ;
        RECT 79.120 147.495 79.440 147.555 ;
        RECT 79.595 147.510 79.885 147.555 ;
        RECT 80.975 147.695 81.265 147.740 ;
        RECT 81.880 147.695 82.200 147.755 ;
        RECT 80.975 147.555 82.200 147.695 ;
        RECT 80.975 147.510 81.265 147.555 ;
        RECT 81.880 147.495 82.200 147.555 ;
        RECT 86.940 147.495 87.260 147.755 ;
        RECT 89.240 147.495 89.560 147.755 ;
        RECT 93.840 147.495 94.160 147.755 ;
        RECT 96.600 147.695 96.920 147.755 ;
        RECT 97.150 147.740 97.290 148.235 ;
        RECT 101.200 148.175 101.520 148.235 ;
        RECT 108.990 148.375 109.280 148.420 ;
        RECT 111.770 148.375 112.060 148.420 ;
        RECT 113.630 148.375 113.920 148.420 ;
        RECT 108.990 148.235 113.920 148.375 ;
        RECT 108.990 148.190 109.280 148.235 ;
        RECT 111.770 148.190 112.060 148.235 ;
        RECT 113.630 148.190 113.920 148.235 ;
        RECT 97.610 147.895 100.970 148.035 ;
        RECT 97.610 147.740 97.750 147.895 ;
        RECT 97.075 147.695 97.365 147.740 ;
        RECT 94.390 147.555 97.365 147.695 ;
        RECT 48.850 147.215 52.210 147.355 ;
        RECT 57.590 147.215 60.490 147.355 ;
        RECT 66.700 147.355 67.020 147.415 ;
        RECT 68.080 147.355 68.400 147.415 ;
        RECT 66.700 147.215 68.400 147.355 ;
        RECT 45.070 147.170 45.360 147.215 ;
        RECT 46.930 147.170 47.220 147.215 ;
        RECT 22.170 146.875 37.030 147.015 ;
        RECT 38.640 147.015 38.960 147.075 ;
        RECT 40.020 147.015 40.340 147.075 ;
        RECT 38.640 146.875 40.340 147.015 ;
        RECT 27.140 146.815 27.460 146.875 ;
        RECT 38.640 146.815 38.960 146.875 ;
        RECT 40.020 146.815 40.340 146.875 ;
        RECT 44.620 147.015 44.940 147.075 ;
        RECT 52.070 147.060 52.210 147.215 ;
        RECT 66.700 147.155 67.020 147.215 ;
        RECT 68.080 147.155 68.400 147.215 ;
        RECT 72.235 147.355 72.525 147.400 ;
        RECT 72.695 147.355 72.985 147.400 ;
        RECT 74.610 147.355 74.750 147.495 ;
        RECT 72.235 147.215 72.985 147.355 ;
        RECT 72.235 147.170 72.525 147.215 ;
        RECT 72.695 147.170 72.985 147.215 ;
        RECT 74.150 147.215 74.750 147.355 ;
        RECT 93.380 147.355 93.700 147.415 ;
        RECT 94.390 147.355 94.530 147.555 ;
        RECT 96.600 147.495 96.920 147.555 ;
        RECT 97.075 147.510 97.365 147.555 ;
        RECT 97.535 147.510 97.825 147.740 ;
        RECT 97.995 147.695 98.285 147.740 ;
        RECT 98.440 147.695 98.760 147.755 ;
        RECT 97.995 147.555 98.760 147.695 ;
        RECT 97.995 147.510 98.285 147.555 ;
        RECT 93.380 147.215 94.530 147.355 ;
        RECT 95.235 147.355 95.525 147.400 ;
        RECT 95.695 147.355 95.985 147.400 ;
        RECT 95.235 147.215 95.985 147.355 ;
        RECT 97.610 147.355 97.750 147.510 ;
        RECT 98.440 147.495 98.760 147.555 ;
        RECT 98.900 147.740 99.220 147.755 ;
        RECT 100.280 147.740 100.600 147.755 ;
        RECT 100.830 147.740 100.970 147.895 ;
        RECT 112.240 147.835 112.560 148.095 ;
        RECT 98.900 147.675 99.265 147.740 ;
        RECT 99.495 147.695 99.785 147.740 ;
        RECT 100.270 147.695 100.600 147.740 ;
        RECT 99.450 147.675 99.785 147.695 ;
        RECT 98.900 147.535 99.785 147.675 ;
        RECT 100.085 147.555 100.600 147.695 ;
        RECT 98.900 147.510 99.265 147.535 ;
        RECT 99.495 147.510 99.785 147.535 ;
        RECT 100.270 147.510 100.600 147.555 ;
        RECT 100.755 147.510 101.045 147.740 ;
        RECT 98.900 147.495 99.220 147.510 ;
        RECT 100.280 147.495 100.600 147.510 ;
        RECT 101.200 147.495 101.520 147.755 ;
        RECT 108.990 147.695 109.280 147.740 ;
        RECT 108.990 147.555 111.525 147.695 ;
        RECT 108.990 147.510 109.280 147.555 ;
        RECT 107.130 147.355 107.420 147.400 ;
        RECT 107.640 147.355 107.960 147.415 ;
        RECT 111.310 147.400 111.525 147.555 ;
        RECT 114.080 147.495 114.400 147.755 ;
        RECT 110.390 147.355 110.680 147.400 ;
        RECT 97.610 147.215 98.210 147.355 ;
        RECT 48.315 147.015 48.605 147.060 ;
        RECT 44.620 146.875 48.605 147.015 ;
        RECT 44.620 146.815 44.940 146.875 ;
        RECT 48.315 146.830 48.605 146.875 ;
        RECT 51.995 146.830 52.285 147.060 ;
        RECT 52.440 147.015 52.760 147.075 ;
        RECT 68.555 147.015 68.845 147.060 ;
        RECT 74.150 147.015 74.290 147.215 ;
        RECT 93.380 147.155 93.700 147.215 ;
        RECT 95.235 147.170 95.525 147.215 ;
        RECT 95.695 147.170 95.985 147.215 ;
        RECT 98.070 147.075 98.210 147.215 ;
        RECT 107.130 147.215 110.680 147.355 ;
        RECT 107.130 147.170 107.420 147.215 ;
        RECT 107.640 147.155 107.960 147.215 ;
        RECT 110.390 147.170 110.680 147.215 ;
        RECT 111.310 147.355 111.600 147.400 ;
        RECT 113.170 147.355 113.460 147.400 ;
        RECT 111.310 147.215 113.460 147.355 ;
        RECT 111.310 147.170 111.600 147.215 ;
        RECT 113.170 147.170 113.460 147.215 ;
        RECT 52.440 146.875 74.290 147.015 ;
        RECT 52.440 146.815 52.760 146.875 ;
        RECT 68.555 146.830 68.845 146.875 ;
        RECT 80.040 146.815 80.360 147.075 ;
        RECT 81.895 147.015 82.185 147.060 ;
        RECT 84.640 147.015 84.960 147.075 ;
        RECT 81.895 146.875 84.960 147.015 ;
        RECT 81.895 146.830 82.185 146.875 ;
        RECT 84.640 146.815 84.960 146.875 ;
        RECT 92.920 146.815 93.240 147.075 ;
        RECT 97.980 146.815 98.300 147.075 ;
        RECT 102.120 147.015 102.440 147.075 ;
        RECT 102.595 147.015 102.885 147.060 ;
        RECT 102.120 146.875 102.885 147.015 ;
        RECT 102.120 146.815 102.440 146.875 ;
        RECT 102.595 146.830 102.885 146.875 ;
        RECT 14.650 146.195 115.850 146.675 ;
        RECT 45.540 145.995 45.860 146.055 ;
        RECT 47.840 145.995 48.160 146.055 ;
        RECT 50.140 145.995 50.460 146.055 ;
        RECT 52.440 145.995 52.760 146.055 ;
        RECT 45.540 145.855 52.760 145.995 ;
        RECT 45.540 145.795 45.860 145.855 ;
        RECT 47.840 145.795 48.160 145.855 ;
        RECT 50.140 145.795 50.460 145.855 ;
        RECT 52.440 145.795 52.760 145.855 ;
        RECT 57.975 145.995 58.265 146.040 ;
        RECT 58.880 145.995 59.200 146.055 ;
        RECT 57.975 145.855 59.200 145.995 ;
        RECT 57.975 145.810 58.265 145.855 ;
        RECT 58.880 145.795 59.200 145.855 ;
        RECT 60.275 145.995 60.565 146.040 ;
        RECT 64.400 145.995 64.720 146.055 ;
        RECT 60.275 145.855 64.720 145.995 ;
        RECT 60.275 145.810 60.565 145.855 ;
        RECT 64.400 145.795 64.720 145.855 ;
        RECT 68.080 145.995 68.400 146.055 ;
        RECT 75.440 145.995 75.760 146.055 ;
        RECT 77.740 146.040 78.060 146.055 ;
        RECT 68.080 145.855 75.760 145.995 ;
        RECT 68.080 145.795 68.400 145.855 ;
        RECT 75.440 145.795 75.760 145.855 ;
        RECT 77.525 145.810 78.060 146.040 ;
        RECT 77.740 145.795 78.060 145.810 ;
        RECT 86.940 145.995 87.260 146.055 ;
        RECT 86.940 145.855 106.030 145.995 ;
        RECT 86.940 145.795 87.260 145.855 ;
        RECT 38.640 145.700 38.960 145.715 ;
        RECT 35.900 145.655 36.190 145.700 ;
        RECT 37.760 145.655 38.050 145.700 ;
        RECT 35.900 145.515 38.050 145.655 ;
        RECT 35.900 145.470 36.190 145.515 ;
        RECT 37.760 145.470 38.050 145.515 ;
        RECT 37.835 145.315 38.050 145.470 ;
        RECT 38.640 145.655 38.970 145.700 ;
        RECT 41.940 145.655 42.230 145.700 ;
        RECT 38.640 145.515 42.230 145.655 ;
        RECT 38.640 145.470 38.970 145.515 ;
        RECT 41.940 145.470 42.230 145.515 ;
        RECT 46.935 145.655 47.225 145.700 ;
        RECT 47.395 145.655 47.685 145.700 ;
        RECT 50.230 145.655 50.370 145.795 ;
        RECT 46.935 145.515 47.685 145.655 ;
        RECT 46.935 145.470 47.225 145.515 ;
        RECT 47.395 145.470 47.685 145.515 ;
        RECT 49.310 145.515 50.370 145.655 ;
        RECT 62.970 145.655 63.260 145.700 ;
        RECT 65.320 145.655 65.640 145.715 ;
        RECT 66.230 145.655 66.520 145.700 ;
        RECT 62.970 145.515 66.520 145.655 ;
        RECT 38.640 145.455 38.960 145.470 ;
        RECT 40.080 145.315 40.370 145.360 ;
        RECT 37.835 145.175 40.370 145.315 ;
        RECT 40.080 145.130 40.370 145.175 ;
        RECT 45.555 145.315 45.845 145.360 ;
        RECT 46.000 145.315 46.320 145.375 ;
        RECT 45.555 145.175 46.320 145.315 ;
        RECT 45.555 145.130 45.845 145.175 ;
        RECT 46.000 145.115 46.320 145.175 ;
        RECT 48.300 145.315 48.620 145.375 ;
        RECT 49.310 145.360 49.450 145.515 ;
        RECT 62.970 145.470 63.260 145.515 ;
        RECT 65.320 145.455 65.640 145.515 ;
        RECT 66.230 145.470 66.520 145.515 ;
        RECT 67.150 145.655 67.440 145.700 ;
        RECT 69.010 145.655 69.300 145.700 ;
        RECT 67.150 145.515 69.300 145.655 ;
        RECT 67.150 145.470 67.440 145.515 ;
        RECT 69.010 145.470 69.300 145.515 ;
        RECT 79.530 145.655 79.820 145.700 ;
        RECT 80.040 145.655 80.360 145.715 ;
        RECT 82.790 145.655 83.080 145.700 ;
        RECT 79.530 145.515 83.080 145.655 ;
        RECT 79.530 145.470 79.820 145.515 ;
        RECT 48.775 145.315 49.065 145.360 ;
        RECT 48.300 145.175 49.065 145.315 ;
        RECT 48.300 145.115 48.620 145.175 ;
        RECT 48.775 145.130 49.065 145.175 ;
        RECT 49.235 145.130 49.525 145.360 ;
        RECT 49.680 145.115 50.000 145.375 ;
        RECT 50.615 145.315 50.905 145.360 ;
        RECT 51.520 145.315 51.840 145.375 ;
        RECT 50.615 145.175 51.840 145.315 ;
        RECT 50.615 145.130 50.905 145.175 ;
        RECT 51.520 145.115 51.840 145.175 ;
        RECT 58.435 145.315 58.725 145.360 ;
        RECT 59.800 145.315 60.120 145.375 ;
        RECT 60.965 145.315 61.255 145.360 ;
        RECT 58.435 145.175 61.255 145.315 ;
        RECT 58.435 145.130 58.725 145.175 ;
        RECT 59.800 145.115 60.120 145.175 ;
        RECT 60.965 145.130 61.255 145.175 ;
        RECT 64.830 145.315 65.120 145.360 ;
        RECT 67.150 145.315 67.365 145.470 ;
        RECT 80.040 145.455 80.360 145.515 ;
        RECT 82.790 145.470 83.080 145.515 ;
        RECT 83.710 145.655 84.000 145.700 ;
        RECT 85.570 145.655 85.860 145.700 ;
        RECT 83.710 145.515 85.860 145.655 ;
        RECT 83.710 145.470 84.000 145.515 ;
        RECT 85.570 145.470 85.860 145.515 ;
        RECT 95.695 145.655 95.985 145.700 ;
        RECT 96.155 145.655 96.445 145.700 ;
        RECT 98.900 145.655 99.220 145.715 ;
        RECT 95.695 145.515 96.445 145.655 ;
        RECT 95.695 145.470 95.985 145.515 ;
        RECT 96.155 145.470 96.445 145.515 ;
        RECT 98.070 145.515 99.220 145.655 ;
        RECT 64.830 145.175 67.365 145.315 ;
        RECT 68.540 145.315 68.860 145.375 ;
        RECT 69.935 145.315 70.225 145.360 ;
        RECT 68.540 145.175 70.225 145.315 ;
        RECT 64.830 145.130 65.120 145.175 ;
        RECT 68.540 145.115 68.860 145.175 ;
        RECT 69.935 145.130 70.225 145.175 ;
        RECT 81.390 145.315 81.680 145.360 ;
        RECT 83.710 145.315 83.925 145.470 ;
        RECT 81.390 145.175 83.925 145.315 ;
        RECT 81.390 145.130 81.680 145.175 ;
        RECT 25.300 144.975 25.620 145.035 ;
        RECT 34.975 144.975 35.265 145.020 ;
        RECT 25.300 144.835 35.265 144.975 ;
        RECT 25.300 144.775 25.620 144.835 ;
        RECT 34.975 144.790 35.265 144.835 ;
        RECT 36.815 144.975 37.105 145.020 ;
        RECT 37.720 144.975 38.040 145.035 ;
        RECT 36.815 144.835 38.040 144.975 ;
        RECT 36.815 144.790 37.105 144.835 ;
        RECT 37.720 144.775 38.040 144.835 ;
        RECT 46.475 144.975 46.765 145.020 ;
        RECT 47.380 144.975 47.700 145.035 ;
        RECT 46.475 144.835 47.700 144.975 ;
        RECT 46.475 144.790 46.765 144.835 ;
        RECT 47.380 144.775 47.700 144.835 ;
        RECT 57.515 144.975 57.805 145.020 ;
        RECT 59.340 144.975 59.660 145.035 ;
        RECT 57.515 144.835 59.660 144.975 ;
        RECT 57.515 144.790 57.805 144.835 ;
        RECT 59.340 144.775 59.660 144.835 ;
        RECT 68.080 144.775 68.400 145.035 ;
        RECT 70.010 144.975 70.150 145.130 ;
        RECT 84.640 145.115 84.960 145.375 ;
        RECT 94.300 145.115 94.620 145.375 ;
        RECT 98.070 145.360 98.210 145.515 ;
        RECT 98.900 145.455 99.220 145.515 ;
        RECT 97.535 145.315 97.825 145.360 ;
        RECT 94.850 145.175 97.825 145.315 ;
        RECT 86.480 144.975 86.800 145.035 ;
        RECT 70.010 144.835 86.800 144.975 ;
        RECT 86.480 144.775 86.800 144.835 ;
        RECT 91.080 144.975 91.400 145.035 ;
        RECT 93.380 144.975 93.700 145.035 ;
        RECT 94.850 144.975 94.990 145.175 ;
        RECT 97.535 145.130 97.825 145.175 ;
        RECT 97.995 145.130 98.285 145.360 ;
        RECT 98.440 145.115 98.760 145.375 ;
        RECT 99.360 145.115 99.680 145.375 ;
        RECT 105.890 145.360 106.030 145.855 ;
        RECT 107.640 145.795 107.960 146.055 ;
        RECT 105.815 145.315 106.105 145.360 ;
        RECT 107.195 145.315 107.485 145.360 ;
        RECT 109.020 145.315 109.340 145.375 ;
        RECT 109.495 145.315 109.785 145.360 ;
        RECT 105.815 145.175 109.785 145.315 ;
        RECT 105.815 145.130 106.105 145.175 ;
        RECT 107.195 145.130 107.485 145.175 ;
        RECT 109.020 145.115 109.340 145.175 ;
        RECT 109.495 145.130 109.785 145.175 ;
        RECT 91.080 144.835 94.990 144.975 ;
        RECT 95.235 144.975 95.525 145.020 ;
        RECT 95.235 144.835 97.750 144.975 ;
        RECT 91.080 144.775 91.400 144.835 ;
        RECT 93.380 144.775 93.700 144.835 ;
        RECT 95.235 144.790 95.525 144.835 ;
        RECT 97.610 144.695 97.750 144.835 ;
        RECT 35.440 144.635 35.730 144.680 ;
        RECT 37.300 144.635 37.590 144.680 ;
        RECT 40.080 144.635 40.370 144.680 ;
        RECT 35.440 144.495 40.370 144.635 ;
        RECT 35.440 144.450 35.730 144.495 ;
        RECT 37.300 144.450 37.590 144.495 ;
        RECT 40.080 144.450 40.370 144.495 ;
        RECT 44.635 144.635 44.925 144.680 ;
        RECT 52.440 144.635 52.760 144.695 ;
        RECT 44.635 144.495 52.760 144.635 ;
        RECT 44.635 144.450 44.925 144.495 ;
        RECT 52.440 144.435 52.760 144.495 ;
        RECT 64.830 144.635 65.120 144.680 ;
        RECT 67.610 144.635 67.900 144.680 ;
        RECT 69.470 144.635 69.760 144.680 ;
        RECT 64.830 144.495 69.760 144.635 ;
        RECT 64.830 144.450 65.120 144.495 ;
        RECT 67.610 144.450 67.900 144.495 ;
        RECT 69.470 144.450 69.760 144.495 ;
        RECT 81.390 144.635 81.680 144.680 ;
        RECT 84.170 144.635 84.460 144.680 ;
        RECT 86.030 144.635 86.320 144.680 ;
        RECT 81.390 144.495 86.320 144.635 ;
        RECT 81.390 144.450 81.680 144.495 ;
        RECT 84.170 144.450 84.460 144.495 ;
        RECT 86.030 144.450 86.320 144.495 ;
        RECT 97.520 144.435 97.840 144.695 ;
        RECT 43.945 144.295 44.235 144.340 ;
        RECT 45.540 144.295 45.860 144.355 ;
        RECT 43.945 144.155 45.860 144.295 ;
        RECT 43.945 144.110 44.235 144.155 ;
        RECT 45.540 144.095 45.860 144.155 ;
        RECT 46.935 144.295 47.225 144.340 ;
        RECT 47.380 144.295 47.700 144.355 ;
        RECT 46.935 144.155 47.700 144.295 ;
        RECT 46.935 144.110 47.225 144.155 ;
        RECT 47.380 144.095 47.700 144.155 ;
        RECT 93.380 144.095 93.700 144.355 ;
        RECT 93.840 144.295 94.160 144.355 ;
        RECT 94.315 144.295 94.605 144.340 ;
        RECT 93.840 144.155 94.605 144.295 ;
        RECT 93.840 144.095 94.160 144.155 ;
        RECT 94.315 144.110 94.605 144.155 ;
        RECT 106.260 144.095 106.580 144.355 ;
        RECT 109.035 144.295 109.325 144.340 ;
        RECT 109.480 144.295 109.800 144.355 ;
        RECT 109.035 144.155 109.800 144.295 ;
        RECT 109.035 144.110 109.325 144.155 ;
        RECT 109.480 144.095 109.800 144.155 ;
        RECT 14.650 143.475 115.850 143.955 ;
        RECT 22.080 143.275 22.400 143.335 ;
        RECT 22.080 143.135 27.370 143.275 ;
        RECT 22.080 143.075 22.400 143.135 ;
        RECT 20.210 142.935 20.500 142.980 ;
        RECT 22.990 142.935 23.280 142.980 ;
        RECT 24.850 142.935 25.140 142.980 ;
        RECT 20.210 142.795 25.140 142.935 ;
        RECT 20.210 142.750 20.500 142.795 ;
        RECT 22.990 142.750 23.280 142.795 ;
        RECT 24.850 142.750 25.140 142.795 ;
        RECT 25.300 142.395 25.620 142.655 ;
        RECT 27.230 142.595 27.370 143.135 ;
        RECT 31.740 143.075 32.060 143.335 ;
        RECT 33.120 143.275 33.440 143.335 ;
        RECT 33.595 143.275 33.885 143.320 ;
        RECT 33.120 143.135 33.885 143.275 ;
        RECT 33.120 143.075 33.440 143.135 ;
        RECT 33.595 143.090 33.885 143.135 ;
        RECT 37.720 143.275 38.040 143.335 ;
        RECT 40.035 143.275 40.325 143.320 ;
        RECT 57.515 143.275 57.805 143.320 ;
        RECT 37.720 143.135 40.325 143.275 ;
        RECT 37.720 143.075 38.040 143.135 ;
        RECT 40.035 143.090 40.325 143.135 ;
        RECT 40.570 143.135 57.805 143.275 ;
        RECT 37.275 142.935 37.565 142.980 ;
        RECT 38.640 142.935 38.960 142.995 ;
        RECT 37.275 142.795 38.960 142.935 ;
        RECT 37.275 142.750 37.565 142.795 ;
        RECT 38.640 142.735 38.960 142.795 ;
        RECT 31.755 142.595 32.045 142.640 ;
        RECT 27.230 142.455 32.045 142.595 ;
        RECT 31.755 142.410 32.045 142.455 ;
        RECT 34.040 142.395 34.360 142.655 ;
        RECT 40.570 142.595 40.710 143.135 ;
        RECT 57.515 143.090 57.805 143.135 ;
        RECT 64.875 143.275 65.165 143.320 ;
        RECT 65.320 143.275 65.640 143.335 ;
        RECT 64.875 143.135 65.640 143.275 ;
        RECT 64.875 143.090 65.165 143.135 ;
        RECT 65.320 143.075 65.640 143.135 ;
        RECT 66.715 143.275 67.005 143.320 ;
        RECT 68.080 143.275 68.400 143.335 ;
        RECT 66.715 143.135 68.400 143.275 ;
        RECT 66.715 143.090 67.005 143.135 ;
        RECT 68.080 143.075 68.400 143.135 ;
        RECT 80.055 143.275 80.345 143.320 ;
        RECT 81.880 143.275 82.200 143.335 ;
        RECT 80.055 143.135 82.200 143.275 ;
        RECT 80.055 143.090 80.345 143.135 ;
        RECT 81.880 143.075 82.200 143.135 ;
        RECT 89.255 143.275 89.545 143.320 ;
        RECT 90.160 143.275 90.480 143.335 ;
        RECT 89.255 143.135 90.480 143.275 ;
        RECT 89.255 143.090 89.545 143.135 ;
        RECT 90.160 143.075 90.480 143.135 ;
        RECT 51.950 142.935 52.240 142.980 ;
        RECT 54.730 142.935 55.020 142.980 ;
        RECT 56.590 142.935 56.880 142.980 ;
        RECT 51.950 142.795 56.880 142.935 ;
        RECT 51.950 142.750 52.240 142.795 ;
        RECT 54.730 142.750 55.020 142.795 ;
        RECT 56.590 142.750 56.880 142.795 ;
        RECT 61.180 142.935 61.500 142.995 ;
        RECT 99.360 142.935 99.680 142.995 ;
        RECT 61.180 142.795 99.680 142.935 ;
        RECT 61.180 142.735 61.500 142.795 ;
        RECT 36.430 142.455 40.710 142.595 ;
        RECT 44.635 142.595 44.925 142.640 ;
        RECT 46.920 142.595 47.240 142.655 ;
        RECT 44.635 142.455 47.240 142.595 ;
        RECT 20.210 142.255 20.500 142.300 ;
        RECT 20.210 142.115 22.745 142.255 ;
        RECT 20.210 142.070 20.500 142.115 ;
        RECT 18.400 141.960 18.720 141.975 ;
        RECT 22.530 141.960 22.745 142.115 ;
        RECT 23.460 142.055 23.780 142.315 ;
        RECT 30.835 142.255 31.125 142.300 ;
        RECT 31.280 142.255 31.600 142.315 ;
        RECT 30.835 142.115 31.600 142.255 ;
        RECT 30.835 142.070 31.125 142.115 ;
        RECT 31.280 142.055 31.600 142.115 ;
        RECT 33.580 142.055 33.900 142.315 ;
        RECT 36.430 142.255 36.570 142.455 ;
        RECT 44.635 142.410 44.925 142.455 ;
        RECT 46.920 142.395 47.240 142.455 ;
        RECT 57.055 142.595 57.345 142.640 ;
        RECT 60.260 142.595 60.580 142.655 ;
        RECT 57.055 142.455 60.580 142.595 ;
        RECT 57.055 142.410 57.345 142.455 ;
        RECT 60.260 142.395 60.580 142.455 ;
        RECT 76.360 142.595 76.680 142.655 ;
        RECT 76.835 142.595 77.125 142.640 ;
        RECT 76.360 142.455 77.125 142.595 ;
        RECT 76.360 142.395 76.680 142.455 ;
        RECT 76.835 142.410 77.125 142.455 ;
        RECT 77.740 142.395 78.060 142.655 ;
        RECT 88.780 142.395 89.100 142.655 ;
        RECT 34.655 142.115 36.570 142.255 ;
        RECT 36.815 142.255 37.105 142.300 ;
        RECT 40.480 142.255 40.800 142.315 ;
        RECT 36.815 142.115 40.800 142.255 ;
        RECT 18.350 141.915 18.720 141.960 ;
        RECT 21.610 141.915 21.900 141.960 ;
        RECT 18.350 141.775 21.900 141.915 ;
        RECT 18.350 141.730 18.720 141.775 ;
        RECT 21.610 141.730 21.900 141.775 ;
        RECT 22.530 141.915 22.820 141.960 ;
        RECT 24.390 141.915 24.680 141.960 ;
        RECT 22.530 141.775 24.680 141.915 ;
        RECT 22.530 141.730 22.820 141.775 ;
        RECT 24.390 141.730 24.680 141.775 ;
        RECT 32.215 141.915 32.505 141.960 ;
        RECT 34.655 141.915 34.795 142.115 ;
        RECT 36.815 142.070 37.105 142.115 ;
        RECT 40.480 142.055 40.800 142.115 ;
        RECT 40.955 142.255 41.245 142.300 ;
        RECT 42.320 142.255 42.640 142.315 ;
        RECT 43.255 142.255 43.545 142.300 ;
        RECT 40.955 142.115 41.630 142.255 ;
        RECT 40.955 142.070 41.245 142.115 ;
        RECT 32.215 141.775 34.795 141.915 ;
        RECT 34.975 141.915 35.265 141.960 ;
        RECT 37.260 141.915 37.580 141.975 ;
        RECT 34.975 141.775 37.580 141.915 ;
        RECT 32.215 141.730 32.505 141.775 ;
        RECT 34.975 141.730 35.265 141.775 ;
        RECT 18.400 141.715 18.720 141.730 ;
        RECT 37.260 141.715 37.580 141.775 ;
        RECT 16.345 141.575 16.635 141.620 ;
        RECT 19.320 141.575 19.640 141.635 ;
        RECT 16.345 141.435 19.640 141.575 ;
        RECT 16.345 141.390 16.635 141.435 ;
        RECT 19.320 141.375 19.640 141.435 ;
        RECT 29.915 141.575 30.205 141.620 ;
        RECT 31.280 141.575 31.600 141.635 ;
        RECT 29.915 141.435 31.600 141.575 ;
        RECT 29.915 141.390 30.205 141.435 ;
        RECT 31.280 141.375 31.600 141.435 ;
        RECT 32.660 141.375 32.980 141.635 ;
        RECT 41.490 141.620 41.630 142.115 ;
        RECT 42.320 142.115 43.545 142.255 ;
        RECT 42.320 142.055 42.640 142.115 ;
        RECT 43.255 142.070 43.545 142.115 ;
        RECT 43.715 142.255 44.005 142.300 ;
        RECT 45.540 142.255 45.860 142.315 ;
        RECT 49.220 142.255 49.540 142.315 ;
        RECT 43.715 142.115 49.540 142.255 ;
        RECT 43.715 142.070 44.005 142.115 ;
        RECT 45.540 142.055 45.860 142.115 ;
        RECT 49.220 142.055 49.540 142.115 ;
        RECT 51.950 142.255 52.240 142.300 ;
        RECT 51.950 142.115 54.485 142.255 ;
        RECT 51.950 142.070 52.240 142.115 ;
        RECT 50.090 141.915 50.380 141.960 ;
        RECT 51.520 141.915 51.840 141.975 ;
        RECT 54.270 141.960 54.485 142.115 ;
        RECT 55.200 142.055 55.520 142.315 ;
        RECT 58.880 142.055 59.200 142.315 ;
        RECT 59.355 142.070 59.645 142.300 ;
        RECT 53.350 141.915 53.640 141.960 ;
        RECT 50.090 141.775 53.640 141.915 ;
        RECT 50.090 141.730 50.380 141.775 ;
        RECT 51.520 141.715 51.840 141.775 ;
        RECT 53.350 141.730 53.640 141.775 ;
        RECT 54.270 141.915 54.560 141.960 ;
        RECT 56.130 141.915 56.420 141.960 ;
        RECT 54.270 141.775 56.420 141.915 ;
        RECT 54.270 141.730 54.560 141.775 ;
        RECT 56.130 141.730 56.420 141.775 ;
        RECT 57.500 141.915 57.820 141.975 ;
        RECT 59.430 141.915 59.570 142.070 ;
        RECT 59.800 142.055 60.120 142.315 ;
        RECT 60.720 142.055 61.040 142.315 ;
        RECT 61.640 142.255 61.960 142.315 ;
        RECT 63.480 142.255 63.800 142.315 ;
        RECT 65.335 142.255 65.625 142.300 ;
        RECT 61.640 142.115 65.625 142.255 ;
        RECT 61.640 142.055 61.960 142.115 ;
        RECT 63.480 142.055 63.800 142.115 ;
        RECT 65.335 142.070 65.625 142.115 ;
        RECT 65.795 142.070 66.085 142.300 ;
        RECT 87.875 142.255 88.165 142.300 ;
        RECT 89.700 142.255 90.020 142.315 ;
        RECT 87.875 142.115 90.020 142.255 ;
        RECT 87.875 142.070 88.165 142.115 ;
        RECT 57.500 141.775 59.570 141.915 ;
        RECT 64.400 141.915 64.720 141.975 ;
        RECT 65.870 141.915 66.010 142.070 ;
        RECT 89.700 142.055 90.020 142.115 ;
        RECT 91.080 142.255 91.400 142.315 ;
        RECT 91.555 142.255 91.845 142.300 ;
        RECT 91.080 142.115 91.845 142.255 ;
        RECT 91.080 142.055 91.400 142.115 ;
        RECT 91.555 142.070 91.845 142.115 ;
        RECT 92.000 142.055 92.320 142.315 ;
        RECT 92.460 142.055 92.780 142.315 ;
        RECT 93.010 142.255 93.150 142.795 ;
        RECT 99.360 142.735 99.680 142.795 ;
        RECT 108.990 142.935 109.280 142.980 ;
        RECT 111.770 142.935 112.060 142.980 ;
        RECT 113.630 142.935 113.920 142.980 ;
        RECT 108.990 142.795 113.920 142.935 ;
        RECT 108.990 142.750 109.280 142.795 ;
        RECT 111.770 142.750 112.060 142.795 ;
        RECT 113.630 142.750 113.920 142.795 ;
        RECT 97.075 142.595 97.365 142.640 ;
        RECT 101.675 142.595 101.965 142.640 ;
        RECT 103.500 142.595 103.820 142.655 ;
        RECT 97.075 142.455 103.820 142.595 ;
        RECT 97.075 142.410 97.365 142.455 ;
        RECT 101.675 142.410 101.965 142.455 ;
        RECT 103.500 142.395 103.820 142.455 ;
        RECT 114.080 142.395 114.400 142.655 ;
        RECT 93.395 142.255 93.685 142.300 ;
        RECT 93.010 142.115 93.685 142.255 ;
        RECT 93.395 142.070 93.685 142.115 ;
        RECT 102.595 142.255 102.885 142.300 ;
        RECT 103.040 142.255 103.360 142.315 ;
        RECT 102.595 142.115 103.360 142.255 ;
        RECT 102.595 142.070 102.885 142.115 ;
        RECT 103.040 142.055 103.360 142.115 ;
        RECT 108.990 142.255 109.280 142.300 ;
        RECT 112.255 142.255 112.545 142.300 ;
        RECT 112.700 142.255 113.020 142.315 ;
        RECT 108.990 142.115 111.525 142.255 ;
        RECT 108.990 142.070 109.280 142.115 ;
        RECT 89.255 141.915 89.545 141.960 ;
        RECT 90.175 141.915 90.465 141.960 ;
        RECT 64.400 141.775 66.010 141.915 ;
        RECT 66.330 141.775 89.010 141.915 ;
        RECT 57.500 141.715 57.820 141.775 ;
        RECT 64.400 141.715 64.720 141.775 ;
        RECT 41.415 141.390 41.705 141.620 ;
        RECT 48.085 141.575 48.375 141.620 ;
        RECT 48.760 141.575 49.080 141.635 ;
        RECT 48.085 141.435 49.080 141.575 ;
        RECT 48.085 141.390 48.375 141.435 ;
        RECT 48.760 141.375 49.080 141.435 ;
        RECT 58.880 141.575 59.200 141.635 ;
        RECT 66.330 141.575 66.470 141.775 ;
        RECT 58.880 141.435 66.470 141.575 ;
        RECT 77.740 141.575 78.060 141.635 ;
        RECT 78.215 141.575 78.505 141.620 ;
        RECT 77.740 141.435 78.505 141.575 ;
        RECT 58.880 141.375 59.200 141.435 ;
        RECT 77.740 141.375 78.060 141.435 ;
        RECT 78.215 141.390 78.505 141.435 ;
        RECT 86.940 141.375 87.260 141.635 ;
        RECT 88.870 141.575 89.010 141.775 ;
        RECT 89.255 141.775 90.465 141.915 ;
        RECT 89.255 141.730 89.545 141.775 ;
        RECT 90.175 141.730 90.465 141.775 ;
        RECT 91.170 141.575 91.310 142.055 ;
        RECT 92.550 141.915 92.690 142.055 ;
        RECT 96.155 141.915 96.445 141.960 ;
        RECT 92.550 141.775 96.445 141.915 ;
        RECT 96.155 141.730 96.445 141.775 ;
        RECT 100.280 141.915 100.600 141.975 ;
        RECT 105.125 141.915 105.415 141.960 ;
        RECT 100.280 141.775 105.415 141.915 ;
        RECT 100.280 141.715 100.600 141.775 ;
        RECT 102.210 141.635 102.350 141.775 ;
        RECT 105.125 141.730 105.415 141.775 ;
        RECT 107.130 141.915 107.420 141.960 ;
        RECT 109.480 141.915 109.800 141.975 ;
        RECT 111.310 141.960 111.525 142.115 ;
        RECT 112.255 142.115 113.020 142.255 ;
        RECT 112.255 142.070 112.545 142.115 ;
        RECT 112.700 142.055 113.020 142.115 ;
        RECT 110.390 141.915 110.680 141.960 ;
        RECT 107.130 141.775 110.680 141.915 ;
        RECT 107.130 141.730 107.420 141.775 ;
        RECT 109.480 141.715 109.800 141.775 ;
        RECT 110.390 141.730 110.680 141.775 ;
        RECT 111.310 141.915 111.600 141.960 ;
        RECT 113.170 141.915 113.460 141.960 ;
        RECT 111.310 141.775 113.460 141.915 ;
        RECT 111.310 141.730 111.600 141.775 ;
        RECT 113.170 141.730 113.460 141.775 ;
        RECT 88.870 141.435 91.310 141.575 ;
        RECT 93.855 141.575 94.145 141.620 ;
        RECT 94.300 141.575 94.620 141.635 ;
        RECT 93.855 141.435 94.620 141.575 ;
        RECT 93.855 141.390 94.145 141.435 ;
        RECT 94.300 141.375 94.620 141.435 ;
        RECT 95.695 141.575 95.985 141.620 ;
        RECT 97.980 141.575 98.300 141.635 ;
        RECT 95.695 141.435 98.300 141.575 ;
        RECT 95.695 141.390 95.985 141.435 ;
        RECT 97.980 141.375 98.300 141.435 ;
        RECT 102.120 141.375 102.440 141.635 ;
        RECT 104.420 141.375 104.740 141.635 ;
        RECT 14.650 140.755 115.850 141.235 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 23.460 140.355 23.780 140.615 ;
        RECT 31.740 140.355 32.060 140.615 ;
        RECT 48.775 140.555 49.065 140.600 ;
        RECT 49.220 140.555 49.540 140.615 ;
        RECT 48.775 140.415 49.540 140.555 ;
        RECT 48.775 140.370 49.065 140.415 ;
        RECT 49.220 140.355 49.540 140.415 ;
        RECT 51.520 140.555 51.840 140.615 ;
        RECT 51.995 140.555 52.285 140.600 ;
        RECT 51.520 140.415 52.285 140.555 ;
        RECT 51.520 140.355 51.840 140.415 ;
        RECT 51.995 140.370 52.285 140.415 ;
        RECT 54.295 140.555 54.585 140.600 ;
        RECT 55.200 140.555 55.520 140.615 ;
        RECT 54.295 140.415 55.520 140.555 ;
        RECT 54.295 140.370 54.585 140.415 ;
        RECT 55.200 140.355 55.520 140.415 ;
        RECT 59.800 140.555 60.120 140.615 ;
        RECT 62.115 140.555 62.405 140.600 ;
        RECT 59.800 140.415 62.405 140.555 ;
        RECT 59.800 140.355 60.120 140.415 ;
        RECT 62.115 140.370 62.405 140.415 ;
        RECT 64.400 140.355 64.720 140.615 ;
        RECT 89.945 140.555 90.235 140.600 ;
        RECT 92.460 140.555 92.780 140.615 ;
        RECT 89.945 140.415 92.780 140.555 ;
        RECT 89.945 140.370 90.235 140.415 ;
        RECT 92.460 140.355 92.780 140.415 ;
        RECT 104.420 140.555 104.740 140.615 ;
        RECT 104.420 140.415 112.010 140.555 ;
        RECT 104.420 140.355 104.740 140.415 ;
        RECT 37.260 140.215 37.580 140.275 ;
        RECT 56.595 140.215 56.885 140.260 ;
        RECT 37.260 140.075 56.885 140.215 ;
        RECT 37.260 140.015 37.580 140.075 ;
        RECT 56.595 140.030 56.885 140.075 ;
        RECT 57.500 140.215 57.820 140.275 ;
        RECT 61.180 140.215 61.500 140.275 ;
        RECT 75.440 140.215 75.760 140.275 ;
        RECT 57.500 140.075 58.650 140.215 ;
        RECT 57.500 140.015 57.820 140.075 ;
        RECT 21.175 139.690 21.465 139.920 ;
        RECT 21.250 139.535 21.390 139.690 ;
        RECT 22.540 139.675 22.860 139.935 ;
        RECT 26.220 139.875 26.540 139.935 ;
        RECT 28.075 139.875 28.365 139.920 ;
        RECT 26.220 139.735 28.365 139.875 ;
        RECT 26.220 139.675 26.540 139.735 ;
        RECT 28.075 139.690 28.365 139.735 ;
        RECT 30.820 139.675 31.140 139.935 ;
        RECT 40.480 139.875 40.800 139.935 ;
        RECT 52.455 139.875 52.745 139.920 ;
        RECT 52.900 139.875 53.220 139.935 ;
        RECT 40.480 139.735 53.220 139.875 ;
        RECT 40.480 139.675 40.800 139.735 ;
        RECT 52.455 139.690 52.745 139.735 ;
        RECT 52.900 139.675 53.220 139.735 ;
        RECT 53.375 139.690 53.665 139.920 ;
        RECT 24.840 139.535 25.160 139.595 ;
        RECT 21.250 139.395 25.160 139.535 ;
        RECT 24.840 139.335 25.160 139.395 ;
        RECT 29.900 139.335 30.220 139.595 ;
        RECT 46.920 139.535 47.240 139.595 ;
        RECT 47.395 139.535 47.685 139.580 ;
        RECT 46.920 139.395 47.685 139.535 ;
        RECT 46.920 139.335 47.240 139.395 ;
        RECT 47.395 139.350 47.685 139.395 ;
        RECT 48.315 139.535 48.605 139.580 ;
        RECT 48.760 139.535 49.080 139.595 ;
        RECT 53.450 139.535 53.590 139.690 ;
        RECT 57.960 139.675 58.280 139.935 ;
        RECT 58.510 139.920 58.650 140.075 ;
        RECT 59.890 140.075 61.500 140.215 ;
        RECT 59.890 139.920 60.030 140.075 ;
        RECT 61.180 140.015 61.500 140.075 ;
        RECT 73.230 140.075 75.760 140.215 ;
        RECT 58.435 139.690 58.725 139.920 ;
        RECT 58.895 139.690 59.185 139.920 ;
        RECT 59.815 139.690 60.105 139.920 ;
        RECT 60.720 139.875 61.040 139.935 ;
        RECT 73.230 139.920 73.370 140.075 ;
        RECT 75.440 140.015 75.760 140.075 ;
        RECT 82.290 140.215 82.580 140.260 ;
        RECT 84.640 140.215 84.960 140.275 ;
        RECT 92.000 140.260 92.320 140.275 ;
        RECT 85.550 140.215 85.840 140.260 ;
        RECT 82.290 140.075 85.840 140.215 ;
        RECT 82.290 140.030 82.580 140.075 ;
        RECT 84.640 140.015 84.960 140.075 ;
        RECT 85.550 140.030 85.840 140.075 ;
        RECT 86.470 140.215 86.760 140.260 ;
        RECT 88.330 140.215 88.620 140.260 ;
        RECT 86.470 140.075 88.620 140.215 ;
        RECT 86.470 140.030 86.760 140.075 ;
        RECT 88.330 140.030 88.620 140.075 ;
        RECT 91.950 140.215 92.320 140.260 ;
        RECT 95.210 140.215 95.500 140.260 ;
        RECT 91.950 140.075 95.500 140.215 ;
        RECT 91.950 140.030 92.320 140.075 ;
        RECT 95.210 140.030 95.500 140.075 ;
        RECT 96.130 140.215 96.420 140.260 ;
        RECT 97.990 140.215 98.280 140.260 ;
        RECT 96.130 140.075 98.280 140.215 ;
        RECT 96.130 140.030 96.420 140.075 ;
        RECT 97.990 140.030 98.280 140.075 ;
        RECT 62.575 139.875 62.865 139.920 ;
        RECT 60.350 139.735 62.865 139.875 ;
        RECT 48.315 139.395 49.080 139.535 ;
        RECT 48.315 139.350 48.605 139.395 ;
        RECT 48.760 139.335 49.080 139.395 ;
        RECT 50.690 139.395 53.590 139.535 ;
        RECT 58.970 139.535 59.110 139.690 ;
        RECT 60.350 139.535 60.490 139.735 ;
        RECT 60.720 139.675 61.040 139.735 ;
        RECT 62.575 139.690 62.865 139.735 ;
        RECT 73.155 139.690 73.445 139.920 ;
        RECT 74.075 139.690 74.365 139.920 ;
        RECT 58.970 139.395 60.490 139.535 ;
        RECT 50.690 139.240 50.830 139.395 ;
        RECT 61.195 139.350 61.485 139.580 ;
        RECT 74.150 139.535 74.290 139.690 ;
        RECT 74.520 139.675 74.840 139.935 ;
        RECT 74.980 139.675 75.300 139.935 ;
        RECT 77.280 139.675 77.600 139.935 ;
        RECT 79.120 139.875 79.440 139.935 ;
        RECT 79.595 139.875 79.885 139.920 ;
        RECT 79.120 139.735 79.885 139.875 ;
        RECT 79.120 139.675 79.440 139.735 ;
        RECT 79.595 139.690 79.885 139.735 ;
        RECT 84.150 139.875 84.440 139.920 ;
        RECT 86.470 139.875 86.685 140.030 ;
        RECT 92.000 140.015 92.320 140.030 ;
        RECT 84.150 139.735 86.685 139.875 ;
        RECT 84.150 139.690 84.440 139.735 ;
        RECT 87.400 139.675 87.720 139.935 ;
        RECT 93.810 139.875 94.100 139.920 ;
        RECT 96.130 139.875 96.345 140.030 ;
        RECT 101.660 140.015 101.980 140.275 ;
        RECT 105.290 140.215 105.580 140.260 ;
        RECT 106.260 140.215 106.580 140.275 ;
        RECT 108.550 140.215 108.840 140.260 ;
        RECT 105.290 140.075 108.840 140.215 ;
        RECT 105.290 140.030 105.580 140.075 ;
        RECT 106.260 140.015 106.580 140.075 ;
        RECT 108.550 140.030 108.840 140.075 ;
        RECT 109.470 140.215 109.760 140.260 ;
        RECT 111.330 140.215 111.620 140.260 ;
        RECT 109.470 140.075 111.620 140.215 ;
        RECT 111.870 140.215 112.010 140.415 ;
        RECT 112.700 140.355 113.020 140.615 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 111.870 140.075 113.850 140.215 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 109.470 140.030 109.760 140.075 ;
        RECT 111.330 140.030 111.620 140.075 ;
        RECT 93.810 139.735 96.345 139.875 ;
        RECT 100.295 139.875 100.585 139.920 ;
        RECT 100.740 139.875 101.060 139.935 ;
        RECT 102.580 139.875 102.900 139.935 ;
        RECT 100.295 139.735 101.060 139.875 ;
        RECT 93.810 139.690 94.100 139.735 ;
        RECT 100.295 139.690 100.585 139.735 ;
        RECT 100.740 139.675 101.060 139.735 ;
        RECT 101.290 139.735 102.900 139.875 ;
        RECT 86.480 139.535 86.800 139.595 ;
        RECT 89.255 139.535 89.545 139.580 ;
        RECT 74.150 139.395 79.810 139.535 ;
        RECT 50.615 139.010 50.905 139.240 ;
        RECT 59.340 139.195 59.660 139.255 ;
        RECT 61.270 139.195 61.410 139.350 ;
        RECT 59.340 139.055 61.410 139.195 ;
        RECT 59.340 138.995 59.660 139.055 ;
        RECT 21.635 138.855 21.925 138.900 ;
        RECT 22.080 138.855 22.400 138.915 ;
        RECT 21.635 138.715 22.400 138.855 ;
        RECT 21.635 138.670 21.925 138.715 ;
        RECT 22.080 138.655 22.400 138.715 ;
        RECT 27.140 138.655 27.460 138.915 ;
        RECT 76.360 138.655 76.680 138.915 ;
        RECT 78.200 138.655 78.520 138.915 ;
        RECT 78.660 138.855 78.980 138.915 ;
        RECT 79.135 138.855 79.425 138.900 ;
        RECT 78.660 138.715 79.425 138.855 ;
        RECT 79.670 138.855 79.810 139.395 ;
        RECT 86.480 139.395 89.545 139.535 ;
        RECT 86.480 139.335 86.800 139.395 ;
        RECT 89.255 139.350 89.545 139.395 ;
        RECT 95.220 139.535 95.540 139.595 ;
        RECT 97.075 139.535 97.365 139.580 ;
        RECT 95.220 139.395 97.365 139.535 ;
        RECT 95.220 139.335 95.540 139.395 ;
        RECT 97.075 139.350 97.365 139.395 ;
        RECT 97.520 139.535 97.840 139.595 ;
        RECT 101.290 139.580 101.430 139.735 ;
        RECT 102.580 139.675 102.900 139.735 ;
        RECT 107.150 139.875 107.440 139.920 ;
        RECT 109.470 139.875 109.685 140.030 ;
        RECT 107.150 139.735 109.685 139.875 ;
        RECT 110.415 139.875 110.705 139.920 ;
        RECT 112.700 139.875 113.020 139.935 ;
        RECT 113.710 139.920 113.850 140.075 ;
        RECT 110.415 139.735 113.020 139.875 ;
        RECT 107.150 139.690 107.440 139.735 ;
        RECT 110.415 139.690 110.705 139.735 ;
        RECT 112.700 139.675 113.020 139.735 ;
        RECT 113.635 139.690 113.925 139.920 ;
        RECT 98.915 139.535 99.205 139.580 ;
        RECT 97.520 139.395 99.590 139.535 ;
        RECT 97.520 139.335 97.840 139.395 ;
        RECT 98.915 139.350 99.205 139.395 ;
        RECT 84.150 139.195 84.440 139.240 ;
        RECT 86.930 139.195 87.220 139.240 ;
        RECT 88.790 139.195 89.080 139.240 ;
        RECT 84.150 139.055 89.080 139.195 ;
        RECT 84.150 139.010 84.440 139.055 ;
        RECT 86.930 139.010 87.220 139.055 ;
        RECT 88.790 139.010 89.080 139.055 ;
        RECT 93.810 139.195 94.100 139.240 ;
        RECT 96.590 139.195 96.880 139.240 ;
        RECT 98.450 139.195 98.740 139.240 ;
        RECT 93.810 139.055 98.740 139.195 ;
        RECT 99.450 139.195 99.590 139.395 ;
        RECT 101.215 139.350 101.505 139.580 ;
        RECT 112.255 139.535 112.545 139.580 ;
        RECT 114.080 139.535 114.400 139.595 ;
        RECT 101.750 139.395 114.400 139.535 ;
        RECT 101.750 139.195 101.890 139.395 ;
        RECT 112.255 139.350 112.545 139.395 ;
        RECT 114.080 139.335 114.400 139.395 ;
        RECT 99.450 139.055 101.890 139.195 ;
        RECT 107.150 139.195 107.440 139.240 ;
        RECT 109.930 139.195 110.220 139.240 ;
        RECT 111.790 139.195 112.080 139.240 ;
        RECT 107.150 139.055 112.080 139.195 ;
        RECT 93.810 139.010 94.100 139.055 ;
        RECT 96.590 139.010 96.880 139.055 ;
        RECT 98.450 139.010 98.740 139.055 ;
        RECT 107.150 139.010 107.440 139.055 ;
        RECT 109.930 139.010 110.220 139.055 ;
        RECT 111.790 139.010 112.080 139.055 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 80.285 138.855 80.575 138.900 ;
        RECT 86.020 138.855 86.340 138.915 ;
        RECT 79.670 138.715 86.340 138.855 ;
        RECT 78.660 138.655 78.980 138.715 ;
        RECT 79.135 138.670 79.425 138.715 ;
        RECT 80.285 138.670 80.575 138.715 ;
        RECT 86.020 138.655 86.340 138.715 ;
        RECT 99.360 138.655 99.680 138.915 ;
        RECT 100.280 138.855 100.600 138.915 ;
        RECT 100.755 138.855 101.045 138.900 ;
        RECT 100.280 138.715 101.045 138.855 ;
        RECT 100.280 138.655 100.600 138.715 ;
        RECT 100.755 138.670 101.045 138.715 ;
        RECT 103.285 138.855 103.575 138.900 ;
        RECT 104.420 138.855 104.740 138.915 ;
        RECT 103.285 138.715 104.740 138.855 ;
        RECT 103.285 138.670 103.575 138.715 ;
        RECT 104.420 138.655 104.740 138.715 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 14.650 138.035 115.850 138.515 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 17.955 137.835 18.245 137.880 ;
        RECT 18.400 137.835 18.720 137.895 ;
        RECT 17.955 137.695 18.720 137.835 ;
        RECT 17.955 137.650 18.245 137.695 ;
        RECT 18.400 137.635 18.720 137.695 ;
        RECT 23.460 137.835 23.780 137.895 ;
        RECT 23.460 137.695 28.750 137.835 ;
        RECT 23.460 137.635 23.780 137.695 ;
        RECT 22.970 137.495 23.260 137.540 ;
        RECT 25.750 137.495 26.040 137.540 ;
        RECT 27.610 137.495 27.900 137.540 ;
        RECT 22.970 137.355 27.900 137.495 ;
        RECT 22.970 137.310 23.260 137.355 ;
        RECT 25.750 137.310 26.040 137.355 ;
        RECT 27.610 137.310 27.900 137.355 ;
        RECT 24.840 137.155 25.160 137.215 ;
        RECT 17.570 137.015 25.160 137.155 ;
        RECT 17.570 136.860 17.710 137.015 ;
        RECT 24.840 136.955 25.160 137.015 ;
        RECT 25.300 137.155 25.620 137.215 ;
        RECT 26.235 137.155 26.525 137.200 ;
        RECT 27.140 137.155 27.460 137.215 ;
        RECT 28.610 137.200 28.750 137.695 ;
        RECT 30.360 137.635 30.680 137.895 ;
        RECT 32.675 137.835 32.965 137.880 ;
        RECT 33.120 137.835 33.440 137.895 ;
        RECT 32.675 137.695 33.440 137.835 ;
        RECT 32.675 137.650 32.965 137.695 ;
        RECT 33.120 137.635 33.440 137.695 ;
        RECT 34.975 137.835 35.265 137.880 ;
        RECT 37.260 137.835 37.580 137.895 ;
        RECT 34.975 137.695 37.580 137.835 ;
        RECT 34.975 137.650 35.265 137.695 ;
        RECT 37.260 137.635 37.580 137.695 ;
        RECT 37.735 137.835 38.025 137.880 ;
        RECT 38.180 137.835 38.500 137.895 ;
        RECT 37.735 137.695 38.500 137.835 ;
        RECT 37.735 137.650 38.025 137.695 ;
        RECT 38.180 137.635 38.500 137.695 ;
        RECT 40.480 137.635 40.800 137.895 ;
        RECT 48.300 137.835 48.620 137.895 ;
        RECT 48.300 137.695 66.470 137.835 ;
        RECT 48.300 137.635 48.620 137.695 ;
        RECT 30.820 137.495 31.140 137.555 ;
        RECT 64.400 137.495 64.720 137.555 ;
        RECT 65.795 137.495 66.085 137.540 ;
        RECT 30.820 137.355 66.085 137.495 ;
        RECT 66.330 137.495 66.470 137.695 ;
        RECT 70.380 137.635 70.700 137.895 ;
        RECT 74.980 137.835 75.300 137.895 ;
        RECT 73.000 137.695 75.300 137.835 ;
        RECT 73.000 137.495 73.140 137.695 ;
        RECT 74.980 137.635 75.300 137.695 ;
        RECT 76.820 137.835 77.140 137.895 ;
        RECT 76.820 137.695 85.330 137.835 ;
        RECT 76.820 137.635 77.140 137.695 ;
        RECT 66.330 137.355 73.140 137.495 ;
        RECT 30.820 137.295 31.140 137.355 ;
        RECT 25.300 137.015 25.990 137.155 ;
        RECT 25.300 136.955 25.620 137.015 ;
        RECT 17.495 136.630 17.785 136.860 ;
        RECT 22.970 136.815 23.260 136.860 ;
        RECT 25.850 136.815 25.990 137.015 ;
        RECT 26.235 137.015 27.460 137.155 ;
        RECT 26.235 136.970 26.525 137.015 ;
        RECT 27.140 136.955 27.460 137.015 ;
        RECT 28.535 136.970 28.825 137.200 ;
        RECT 31.830 137.155 31.970 137.355 ;
        RECT 33.135 137.155 33.425 137.200 ;
        RECT 29.530 137.015 31.970 137.155 ;
        RECT 29.530 136.860 29.670 137.015 ;
        RECT 31.830 136.860 31.970 137.015 ;
        RECT 32.290 137.015 33.425 137.155 ;
        RECT 28.075 136.815 28.365 136.860 ;
        RECT 22.970 136.675 25.505 136.815 ;
        RECT 25.850 136.675 28.365 136.815 ;
        RECT 22.970 136.630 23.260 136.675 ;
        RECT 21.110 136.475 21.400 136.520 ;
        RECT 22.080 136.475 22.400 136.535 ;
        RECT 25.290 136.520 25.505 136.675 ;
        RECT 28.075 136.630 28.365 136.675 ;
        RECT 29.455 136.630 29.745 136.860 ;
        RECT 30.835 136.630 31.125 136.860 ;
        RECT 31.755 136.630 32.045 136.860 ;
        RECT 24.370 136.475 24.660 136.520 ;
        RECT 21.110 136.335 24.660 136.475 ;
        RECT 21.110 136.290 21.400 136.335 ;
        RECT 22.080 136.275 22.400 136.335 ;
        RECT 24.370 136.290 24.660 136.335 ;
        RECT 25.290 136.475 25.580 136.520 ;
        RECT 27.150 136.475 27.440 136.520 ;
        RECT 25.290 136.335 27.440 136.475 ;
        RECT 25.290 136.290 25.580 136.335 ;
        RECT 27.150 136.290 27.440 136.335 ;
        RECT 28.520 136.475 28.840 136.535 ;
        RECT 30.910 136.475 31.050 136.630 ;
        RECT 28.520 136.335 31.050 136.475 ;
        RECT 28.520 136.275 28.840 136.335 ;
        RECT 19.105 136.135 19.395 136.180 ;
        RECT 21.620 136.135 21.940 136.195 ;
        RECT 19.105 135.995 21.940 136.135 ;
        RECT 19.105 135.950 19.395 135.995 ;
        RECT 21.620 135.935 21.940 135.995 ;
        RECT 23.000 136.135 23.320 136.195 ;
        RECT 32.290 136.135 32.430 137.015 ;
        RECT 33.135 136.970 33.425 137.015 ;
        RECT 34.130 136.860 34.270 137.355 ;
        RECT 64.400 137.295 64.720 137.355 ;
        RECT 65.795 137.310 66.085 137.355 ;
        RECT 40.020 136.955 40.340 137.215 ;
        RECT 46.460 137.155 46.780 137.215 ;
        RECT 51.980 137.155 52.300 137.215 ;
        RECT 46.460 137.015 52.300 137.155 ;
        RECT 46.460 136.955 46.780 137.015 ;
        RECT 34.055 136.630 34.345 136.860 ;
        RECT 35.895 136.630 36.185 136.860 ;
        RECT 36.815 136.630 37.105 136.860 ;
        RECT 33.580 136.475 33.900 136.535 ;
        RECT 35.970 136.475 36.110 136.630 ;
        RECT 33.580 136.335 36.110 136.475 ;
        RECT 36.890 136.475 37.030 136.630 ;
        RECT 39.560 136.615 39.880 136.875 ;
        RECT 44.620 136.815 44.940 136.875 ;
        RECT 48.300 136.815 48.620 136.875 ;
        RECT 50.230 136.860 50.370 137.015 ;
        RECT 51.980 136.955 52.300 137.015 ;
        RECT 70.395 137.155 70.685 137.200 ;
        RECT 71.760 137.155 72.080 137.215 ;
        RECT 70.395 137.015 72.080 137.155 ;
        RECT 70.395 136.970 70.685 137.015 ;
        RECT 71.760 136.955 72.080 137.015 ;
        RECT 44.620 136.675 48.620 136.815 ;
        RECT 44.620 136.615 44.940 136.675 ;
        RECT 48.300 136.615 48.620 136.675 ;
        RECT 48.775 136.630 49.065 136.860 ;
        RECT 49.235 136.630 49.525 136.860 ;
        RECT 50.155 136.630 50.445 136.860 ;
        RECT 51.535 136.815 51.825 136.860 ;
        RECT 52.900 136.815 53.220 136.875 ;
        RECT 51.535 136.675 53.220 136.815 ;
        RECT 51.535 136.630 51.825 136.675 ;
        RECT 40.955 136.475 41.245 136.520 ;
        RECT 46.935 136.475 47.225 136.520 ;
        RECT 36.890 136.335 39.790 136.475 ;
        RECT 33.580 136.275 33.900 136.335 ;
        RECT 39.650 136.195 39.790 136.335 ;
        RECT 40.955 136.335 47.225 136.475 ;
        RECT 40.955 136.290 41.245 136.335 ;
        RECT 46.935 136.290 47.225 136.335 ;
        RECT 47.840 136.475 48.160 136.535 ;
        RECT 48.850 136.475 48.990 136.630 ;
        RECT 47.840 136.335 48.990 136.475 ;
        RECT 49.310 136.475 49.450 136.630 ;
        RECT 52.900 136.615 53.220 136.675 ;
        RECT 58.880 136.815 59.200 136.875 ;
        RECT 63.480 136.815 63.800 136.875 ;
        RECT 58.880 136.675 63.800 136.815 ;
        RECT 58.880 136.615 59.200 136.675 ;
        RECT 63.480 136.615 63.800 136.675 ;
        RECT 66.715 136.815 67.005 136.860 ;
        RECT 67.620 136.815 67.940 136.875 ;
        RECT 66.715 136.675 67.940 136.815 ;
        RECT 66.715 136.630 67.005 136.675 ;
        RECT 67.620 136.615 67.940 136.675 ;
        RECT 69.460 136.615 69.780 136.875 ;
        RECT 72.770 136.860 72.910 137.355 ;
        RECT 74.520 137.295 74.840 137.555 ;
        RECT 79.090 137.495 79.380 137.540 ;
        RECT 81.870 137.495 82.160 137.540 ;
        RECT 83.730 137.495 84.020 137.540 ;
        RECT 79.090 137.355 84.020 137.495 ;
        RECT 79.090 137.310 79.380 137.355 ;
        RECT 81.870 137.310 82.160 137.355 ;
        RECT 83.730 137.310 84.020 137.355 ;
        RECT 74.610 137.155 74.750 137.295 ;
        RECT 73.230 137.015 74.750 137.155 ;
        RECT 78.200 137.155 78.520 137.215 ;
        RECT 85.190 137.200 85.330 137.695 ;
        RECT 92.000 137.635 92.320 137.895 ;
        RECT 95.220 137.635 95.540 137.895 ;
        RECT 95.695 137.835 95.985 137.880 ;
        RECT 97.060 137.835 97.380 137.895 ;
        RECT 95.695 137.695 97.380 137.835 ;
        RECT 95.695 137.650 95.985 137.695 ;
        RECT 97.060 137.635 97.380 137.695 ;
        RECT 108.575 137.835 108.865 137.880 ;
        RECT 112.700 137.835 113.020 137.895 ;
        RECT 108.575 137.695 113.020 137.835 ;
        RECT 108.575 137.650 108.865 137.695 ;
        RECT 112.700 137.635 113.020 137.695 ;
        RECT 97.980 137.495 98.300 137.555 ;
        RECT 97.980 137.355 104.650 137.495 ;
        RECT 97.980 137.295 98.300 137.355 ;
        RECT 104.510 137.215 104.650 137.355 ;
        RECT 106.735 137.310 107.025 137.540 ;
        RECT 82.355 137.155 82.645 137.200 ;
        RECT 78.200 137.015 82.645 137.155 ;
        RECT 73.230 136.860 73.370 137.015 ;
        RECT 78.200 136.955 78.520 137.015 ;
        RECT 82.355 136.970 82.645 137.015 ;
        RECT 85.115 136.970 85.405 137.200 ;
        RECT 86.020 136.955 86.340 137.215 ;
        RECT 86.480 136.955 86.800 137.215 ;
        RECT 103.500 136.955 103.820 137.215 ;
        RECT 104.420 136.955 104.740 137.215 ;
        RECT 106.810 137.155 106.950 137.310 ;
        RECT 106.810 137.015 107.870 137.155 ;
        RECT 72.695 136.630 72.985 136.860 ;
        RECT 73.155 136.630 73.445 136.860 ;
        RECT 73.615 136.630 73.905 136.860 ;
        RECT 74.535 136.815 74.825 136.860 ;
        RECT 75.440 136.815 75.760 136.875 ;
        RECT 74.535 136.675 75.760 136.815 ;
        RECT 74.535 136.630 74.825 136.675 ;
        RECT 54.740 136.475 55.060 136.535 ;
        RECT 49.310 136.335 55.060 136.475 ;
        RECT 47.840 136.275 48.160 136.335 ;
        RECT 54.740 136.275 55.060 136.335 ;
        RECT 70.855 136.475 71.145 136.520 ;
        RECT 71.315 136.475 71.605 136.520 ;
        RECT 70.855 136.335 71.605 136.475 ;
        RECT 70.855 136.290 71.145 136.335 ;
        RECT 71.315 136.290 71.605 136.335 ;
        RECT 23.000 135.995 32.430 136.135 ;
        RECT 38.655 136.135 38.945 136.180 ;
        RECT 39.100 136.135 39.420 136.195 ;
        RECT 38.655 135.995 39.420 136.135 ;
        RECT 23.000 135.935 23.320 135.995 ;
        RECT 38.655 135.950 38.945 135.995 ;
        RECT 39.100 135.935 39.420 135.995 ;
        RECT 39.560 135.935 39.880 136.195 ;
        RECT 51.980 135.935 52.300 136.195 ;
        RECT 63.035 136.135 63.325 136.180 ;
        RECT 63.480 136.135 63.800 136.195 ;
        RECT 63.035 135.995 63.800 136.135 ;
        RECT 63.035 135.950 63.325 135.995 ;
        RECT 63.480 135.935 63.800 135.995 ;
        RECT 68.555 136.135 68.845 136.180 ;
        RECT 71.760 136.135 72.080 136.195 ;
        RECT 68.555 135.995 72.080 136.135 ;
        RECT 73.690 136.135 73.830 136.630 ;
        RECT 75.440 136.615 75.760 136.675 ;
        RECT 79.090 136.815 79.380 136.860 ;
        RECT 84.180 136.815 84.500 136.875 ;
        RECT 86.570 136.815 86.710 136.955 ;
        RECT 79.090 136.675 81.625 136.815 ;
        RECT 79.090 136.630 79.380 136.675 ;
        RECT 77.230 136.475 77.520 136.520 ;
        RECT 78.660 136.475 78.980 136.535 ;
        RECT 81.410 136.520 81.625 136.675 ;
        RECT 84.180 136.675 86.710 136.815 ;
        RECT 91.080 136.815 91.400 136.875 ;
        RECT 91.555 136.815 91.845 136.860 ;
        RECT 91.080 136.675 91.845 136.815 ;
        RECT 84.180 136.615 84.500 136.675 ;
        RECT 91.080 136.615 91.400 136.675 ;
        RECT 91.555 136.630 91.845 136.675 ;
        RECT 94.300 136.615 94.620 136.875 ;
        RECT 96.615 136.630 96.905 136.860 ;
        RECT 80.490 136.475 80.780 136.520 ;
        RECT 77.230 136.335 80.780 136.475 ;
        RECT 77.230 136.290 77.520 136.335 ;
        RECT 78.660 136.275 78.980 136.335 ;
        RECT 80.490 136.290 80.780 136.335 ;
        RECT 81.410 136.475 81.700 136.520 ;
        RECT 83.270 136.475 83.560 136.520 ;
        RECT 81.410 136.335 83.560 136.475 ;
        RECT 81.410 136.290 81.700 136.335 ;
        RECT 83.270 136.290 83.560 136.335 ;
        RECT 86.495 136.475 86.785 136.520 ;
        RECT 92.460 136.475 92.780 136.535 ;
        RECT 96.690 136.475 96.830 136.630 ;
        RECT 97.060 136.615 97.380 136.875 ;
        RECT 102.120 136.815 102.440 136.875 ;
        RECT 107.730 136.860 107.870 137.015 ;
        RECT 104.895 136.815 105.185 136.860 ;
        RECT 102.120 136.675 105.185 136.815 ;
        RECT 102.120 136.615 102.440 136.675 ;
        RECT 104.895 136.630 105.185 136.675 ;
        RECT 107.695 136.630 107.985 136.860 ;
        RECT 86.495 136.335 92.780 136.475 ;
        RECT 86.495 136.290 86.785 136.335 ;
        RECT 92.460 136.275 92.780 136.335 ;
        RECT 94.390 136.335 96.830 136.475 ;
        RECT 94.390 136.195 94.530 136.335 ;
        RECT 75.225 136.135 75.515 136.180 ;
        RECT 77.740 136.135 78.060 136.195 ;
        RECT 79.580 136.135 79.900 136.195 ;
        RECT 73.690 135.995 79.900 136.135 ;
        RECT 68.555 135.950 68.845 135.995 ;
        RECT 71.760 135.935 72.080 135.995 ;
        RECT 75.225 135.950 75.515 135.995 ;
        RECT 77.740 135.935 78.060 135.995 ;
        RECT 79.580 135.935 79.900 135.995 ;
        RECT 88.320 135.935 88.640 136.195 ;
        RECT 94.300 135.935 94.620 136.195 ;
        RECT 14.650 135.315 115.850 135.795 ;
        RECT 19.320 135.115 19.640 135.175 ;
        RECT 22.080 135.115 22.400 135.175 ;
        RECT 19.320 134.975 22.400 135.115 ;
        RECT 19.320 134.915 19.640 134.975 ;
        RECT 22.080 134.915 22.400 134.975 ;
        RECT 22.540 135.115 22.860 135.175 ;
        RECT 23.935 135.115 24.225 135.160 ;
        RECT 22.540 134.975 24.225 135.115 ;
        RECT 22.540 134.915 22.860 134.975 ;
        RECT 23.935 134.930 24.225 134.975 ;
        RECT 26.220 134.915 26.540 135.175 ;
        RECT 28.075 135.115 28.365 135.160 ;
        RECT 29.900 135.115 30.220 135.175 ;
        RECT 28.075 134.975 30.220 135.115 ;
        RECT 28.075 134.930 28.365 134.975 ;
        RECT 21.620 134.775 21.940 134.835 ;
        RECT 28.150 134.775 28.290 134.930 ;
        RECT 29.900 134.915 30.220 134.975 ;
        RECT 37.720 134.915 38.040 135.175 ;
        RECT 40.495 135.115 40.785 135.160 ;
        RECT 44.160 135.115 44.480 135.175 ;
        RECT 47.840 135.115 48.160 135.175 ;
        RECT 40.495 134.975 44.480 135.115 ;
        RECT 40.495 134.930 40.785 134.975 ;
        RECT 44.160 134.915 44.480 134.975 ;
        RECT 45.170 134.975 48.160 135.115 ;
        RECT 21.620 134.635 28.290 134.775 ;
        RECT 28.520 134.775 28.840 134.835 ;
        RECT 33.595 134.775 33.885 134.820 ;
        RECT 28.520 134.635 33.885 134.775 ;
        RECT 21.620 134.575 21.940 134.635 ;
        RECT 28.520 134.575 28.840 134.635 ;
        RECT 33.595 134.590 33.885 134.635 ;
        RECT 42.795 134.775 43.085 134.820 ;
        RECT 43.255 134.775 43.545 134.820 ;
        RECT 42.795 134.635 43.545 134.775 ;
        RECT 42.795 134.590 43.085 134.635 ;
        RECT 43.255 134.590 43.545 134.635 ;
        RECT 24.840 134.435 25.160 134.495 ;
        RECT 28.980 134.435 29.300 134.495 ;
        RECT 30.375 134.435 30.665 134.480 ;
        RECT 24.840 134.295 30.665 134.435 ;
        RECT 24.840 134.235 25.160 134.295 ;
        RECT 28.980 134.235 29.300 134.295 ;
        RECT 30.375 134.250 30.665 134.295 ;
        RECT 30.820 134.235 31.140 134.495 ;
        RECT 38.640 134.235 38.960 134.495 ;
        RECT 40.035 134.435 40.325 134.480 ;
        RECT 40.940 134.435 41.260 134.495 ;
        RECT 40.035 134.295 41.260 134.435 ;
        RECT 40.035 134.250 40.325 134.295 ;
        RECT 40.940 134.235 41.260 134.295 ;
        RECT 41.400 134.235 41.720 134.495 ;
        RECT 44.620 134.235 44.940 134.495 ;
        RECT 45.170 134.480 45.310 134.975 ;
        RECT 47.840 134.915 48.160 134.975 ;
        RECT 50.615 134.930 50.905 135.160 ;
        RECT 57.055 135.115 57.345 135.160 ;
        RECT 58.420 135.115 58.740 135.175 ;
        RECT 57.055 134.975 58.740 135.115 ;
        RECT 57.055 134.930 57.345 134.975 ;
        RECT 48.760 134.775 49.080 134.835 ;
        RECT 45.630 134.635 49.080 134.775 ;
        RECT 45.630 134.480 45.770 134.635 ;
        RECT 48.760 134.575 49.080 134.635 ;
        RECT 45.095 134.250 45.385 134.480 ;
        RECT 45.555 134.250 45.845 134.480 ;
        RECT 46.460 134.235 46.780 134.495 ;
        RECT 46.920 134.435 47.240 134.495 ;
        RECT 50.690 134.435 50.830 134.930 ;
        RECT 58.420 134.915 58.740 134.975 ;
        RECT 72.235 135.115 72.525 135.160 ;
        RECT 72.680 135.115 73.000 135.175 ;
        RECT 72.235 134.975 73.000 135.115 ;
        RECT 72.235 134.930 72.525 134.975 ;
        RECT 72.680 134.915 73.000 134.975 ;
        RECT 77.280 134.915 77.600 135.175 ;
        RECT 79.580 134.915 79.900 135.175 ;
        RECT 84.195 135.115 84.485 135.160 ;
        RECT 84.640 135.115 84.960 135.175 ;
        RECT 84.195 134.975 84.960 135.115 ;
        RECT 84.195 134.930 84.485 134.975 ;
        RECT 84.640 134.915 84.960 134.975 ;
        RECT 87.400 134.915 87.720 135.175 ;
        RECT 94.300 135.115 94.620 135.175 ;
        RECT 93.930 134.975 99.590 135.115 ;
        RECT 61.130 134.775 61.420 134.820 ;
        RECT 63.480 134.775 63.800 134.835 ;
        RECT 64.390 134.775 64.680 134.820 ;
        RECT 61.130 134.635 64.680 134.775 ;
        RECT 61.130 134.590 61.420 134.635 ;
        RECT 63.480 134.575 63.800 134.635 ;
        RECT 64.390 134.590 64.680 134.635 ;
        RECT 65.310 134.775 65.600 134.820 ;
        RECT 67.170 134.775 67.460 134.820 ;
        RECT 65.310 134.635 67.460 134.775 ;
        RECT 65.310 134.590 65.600 134.635 ;
        RECT 67.170 134.590 67.460 134.635 ;
        RECT 74.535 134.775 74.825 134.820 ;
        RECT 76.360 134.775 76.680 134.835 ;
        RECT 74.535 134.635 76.680 134.775 ;
        RECT 74.535 134.590 74.825 134.635 ;
        RECT 51.995 134.435 52.285 134.480 ;
        RECT 55.215 134.435 55.505 134.480 ;
        RECT 46.920 134.295 47.610 134.435 ;
        RECT 50.690 134.295 52.285 134.435 ;
        RECT 46.920 134.235 47.240 134.295 ;
        RECT 21.175 133.910 21.465 134.140 ;
        RECT 21.250 133.755 21.390 133.910 ;
        RECT 28.520 133.895 28.840 134.155 ;
        RECT 29.455 133.910 29.745 134.140 ;
        RECT 32.215 133.910 32.505 134.140 ;
        RECT 33.135 134.095 33.425 134.140 ;
        RECT 38.180 134.095 38.500 134.155 ;
        RECT 33.135 133.955 38.500 134.095 ;
        RECT 33.135 133.910 33.425 133.955 ;
        RECT 29.530 133.755 29.670 133.910 ;
        RECT 30.360 133.755 30.680 133.815 ;
        RECT 32.290 133.755 32.430 133.910 ;
        RECT 38.180 133.895 38.500 133.955 ;
        RECT 39.575 134.095 39.865 134.140 ;
        RECT 41.860 134.095 42.180 134.155 ;
        RECT 39.575 133.955 42.180 134.095 ;
        RECT 39.575 133.910 39.865 133.955 ;
        RECT 41.860 133.895 42.180 133.955 ;
        RECT 42.335 134.095 42.625 134.140 ;
        RECT 43.240 134.095 43.560 134.155 ;
        RECT 47.470 134.140 47.610 134.295 ;
        RECT 51.995 134.250 52.285 134.295 ;
        RECT 52.530 134.295 55.505 134.435 ;
        RECT 47.395 134.095 47.685 134.140 ;
        RECT 42.335 133.955 43.560 134.095 ;
        RECT 42.335 133.910 42.625 133.955 ;
        RECT 43.240 133.895 43.560 133.955 ;
        RECT 46.550 133.955 47.685 134.095 ;
        RECT 21.250 133.615 32.430 133.755 ;
        RECT 30.360 133.555 30.680 133.615 ;
        RECT 35.435 133.415 35.725 133.460 ;
        RECT 37.260 133.415 37.580 133.475 ;
        RECT 35.435 133.275 37.580 133.415 ;
        RECT 35.435 133.230 35.725 133.275 ;
        RECT 37.260 133.215 37.580 133.275 ;
        RECT 40.020 133.215 40.340 133.475 ;
        RECT 42.320 133.215 42.640 133.475 ;
        RECT 46.550 133.415 46.690 133.955 ;
        RECT 47.395 133.910 47.685 133.955 ;
        RECT 48.315 134.095 48.605 134.140 ;
        RECT 52.530 134.095 52.670 134.295 ;
        RECT 55.215 134.250 55.505 134.295 ;
        RECT 62.990 134.435 63.280 134.480 ;
        RECT 65.310 134.435 65.525 134.590 ;
        RECT 76.360 134.575 76.680 134.635 ;
        RECT 79.135 134.775 79.425 134.820 ;
        RECT 86.020 134.775 86.340 134.835 ;
        RECT 79.135 134.635 86.340 134.775 ;
        RECT 79.135 134.590 79.425 134.635 ;
        RECT 86.020 134.575 86.340 134.635 ;
        RECT 62.990 134.295 65.525 134.435 ;
        RECT 62.990 134.250 63.280 134.295 ;
        RECT 66.240 134.235 66.560 134.495 ;
        RECT 73.140 134.235 73.460 134.495 ;
        RECT 79.580 134.435 79.900 134.495 ;
        RECT 84.655 134.435 84.945 134.480 ;
        RECT 79.580 134.295 84.945 134.435 ;
        RECT 79.580 134.235 79.900 134.295 ;
        RECT 84.655 134.250 84.945 134.295 ;
        RECT 85.100 134.435 85.420 134.495 ;
        RECT 86.955 134.435 87.245 134.480 ;
        RECT 85.100 134.295 87.245 134.435 ;
        RECT 48.315 133.955 52.670 134.095 ;
        RECT 48.315 133.910 48.605 133.955 ;
        RECT 53.835 133.910 54.125 134.140 ;
        RECT 46.920 133.755 47.240 133.815 ;
        RECT 48.390 133.755 48.530 133.910 ;
        RECT 53.910 133.755 54.050 133.910 ;
        RECT 54.740 133.895 55.060 134.155 ;
        RECT 59.340 134.095 59.660 134.155 ;
        RECT 59.200 133.895 59.660 134.095 ;
        RECT 60.260 134.095 60.580 134.155 ;
        RECT 68.095 134.095 68.385 134.140 ;
        RECT 60.260 133.955 68.385 134.095 ;
        RECT 60.260 133.895 60.580 133.955 ;
        RECT 68.095 133.910 68.385 133.955 ;
        RECT 74.075 134.095 74.365 134.140 ;
        RECT 75.900 134.095 76.220 134.155 ;
        RECT 74.075 133.955 76.220 134.095 ;
        RECT 74.075 133.910 74.365 133.955 ;
        RECT 75.900 133.895 76.220 133.955 ;
        RECT 76.820 134.095 77.140 134.155 ;
        RECT 80.055 134.095 80.345 134.140 ;
        RECT 76.820 133.955 80.345 134.095 ;
        RECT 84.730 134.095 84.870 134.250 ;
        RECT 85.100 134.235 85.420 134.295 ;
        RECT 86.955 134.250 87.245 134.295 ;
        RECT 88.320 134.235 88.640 134.495 ;
        RECT 90.620 134.435 90.940 134.495 ;
        RECT 88.870 134.295 90.940 134.435 ;
        RECT 88.870 134.095 89.010 134.295 ;
        RECT 90.620 134.235 90.940 134.295 ;
        RECT 91.095 134.435 91.385 134.480 ;
        RECT 93.395 134.435 93.685 134.480 ;
        RECT 93.930 134.435 94.070 134.975 ;
        RECT 94.300 134.915 94.620 134.975 ;
        RECT 97.520 134.575 97.840 134.835 ;
        RECT 91.095 134.295 94.070 134.435 ;
        RECT 91.095 134.250 91.385 134.295 ;
        RECT 93.395 134.250 93.685 134.295 ;
        RECT 84.730 133.955 89.010 134.095 ;
        RECT 76.820 133.895 77.140 133.955 ;
        RECT 80.055 133.910 80.345 133.955 ;
        RECT 90.160 133.895 90.480 134.155 ;
        RECT 59.200 133.755 59.340 133.895 ;
        RECT 46.920 133.615 48.530 133.755 ;
        RECT 52.530 133.615 59.340 133.755 ;
        RECT 62.990 133.755 63.280 133.800 ;
        RECT 65.770 133.755 66.060 133.800 ;
        RECT 67.630 133.755 67.920 133.800 ;
        RECT 91.170 133.755 91.310 134.250 ;
        RECT 94.300 134.235 94.620 134.495 ;
        RECT 99.450 134.480 99.590 134.975 ;
        RECT 100.280 134.915 100.600 135.175 ;
        RECT 99.375 134.435 99.665 134.480 ;
        RECT 100.280 134.435 100.600 134.495 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 99.375 134.295 100.600 134.435 ;
        RECT 99.375 134.250 99.665 134.295 ;
        RECT 100.280 134.235 100.600 134.295 ;
        RECT 92.000 133.895 92.320 134.155 ;
        RECT 97.980 134.095 98.300 134.155 ;
        RECT 98.455 134.095 98.745 134.140 ;
        RECT 97.980 133.955 98.745 134.095 ;
        RECT 97.980 133.895 98.300 133.955 ;
        RECT 98.455 133.910 98.745 133.955 ;
        RECT 62.990 133.615 67.920 133.755 ;
        RECT 46.920 133.555 47.240 133.615 ;
        RECT 52.530 133.415 52.670 133.615 ;
        RECT 62.990 133.570 63.280 133.615 ;
        RECT 65.770 133.570 66.060 133.615 ;
        RECT 67.630 133.570 67.920 133.615 ;
        RECT 74.150 133.615 91.310 133.755 ;
        RECT 46.550 133.275 52.670 133.415 ;
        RECT 52.915 133.415 53.205 133.460 ;
        RECT 55.660 133.415 55.980 133.475 ;
        RECT 52.915 133.275 55.980 133.415 ;
        RECT 52.915 133.230 53.205 133.275 ;
        RECT 55.660 133.215 55.980 133.275 ;
        RECT 59.125 133.415 59.415 133.460 ;
        RECT 60.720 133.415 61.040 133.475 ;
        RECT 59.125 133.275 61.040 133.415 ;
        RECT 59.125 133.230 59.415 133.275 ;
        RECT 60.720 133.215 61.040 133.275 ;
        RECT 64.400 133.415 64.720 133.475 ;
        RECT 74.150 133.415 74.290 133.615 ;
        RECT 64.400 133.275 74.290 133.415 ;
        RECT 74.535 133.415 74.825 133.460 ;
        RECT 77.280 133.415 77.600 133.475 ;
        RECT 74.535 133.275 77.600 133.415 ;
        RECT 64.400 133.215 64.720 133.275 ;
        RECT 74.535 133.230 74.825 133.275 ;
        RECT 77.280 133.215 77.600 133.275 ;
        RECT 85.560 133.415 85.880 133.475 ;
        RECT 86.035 133.415 86.325 133.460 ;
        RECT 85.560 133.275 86.325 133.415 ;
        RECT 85.560 133.215 85.880 133.275 ;
        RECT 86.035 133.230 86.325 133.275 ;
        RECT 91.540 133.415 91.860 133.475 ;
        RECT 92.475 133.415 92.765 133.460 ;
        RECT 91.540 133.275 92.765 133.415 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 91.540 133.215 91.860 133.275 ;
        RECT 92.475 133.230 92.765 133.275 ;
        RECT 14.650 132.595 115.850 133.075 ;
        RECT 16.805 132.395 17.095 132.440 ;
        RECT 23.000 132.395 23.320 132.455 ;
        RECT 16.805 132.255 23.320 132.395 ;
        RECT 16.805 132.210 17.095 132.255 ;
        RECT 23.000 132.195 23.320 132.255 ;
        RECT 27.845 132.395 28.135 132.440 ;
        RECT 28.520 132.395 28.840 132.455 ;
        RECT 27.845 132.255 28.840 132.395 ;
        RECT 27.845 132.210 28.135 132.255 ;
        RECT 28.520 132.195 28.840 132.255 ;
        RECT 40.480 132.195 40.800 132.455 ;
        RECT 42.320 132.195 42.640 132.455 ;
        RECT 72.220 132.195 72.540 132.455 ;
        RECT 78.215 132.395 78.505 132.440 ;
        RECT 84.180 132.395 84.500 132.455 ;
        RECT 78.215 132.255 84.500 132.395 ;
        RECT 78.215 132.210 78.505 132.255 ;
        RECT 84.180 132.195 84.500 132.255 ;
        RECT 85.100 132.195 85.420 132.455 ;
        RECT 92.460 132.395 92.780 132.455 ;
        RECT 97.520 132.395 97.840 132.455 ;
        RECT 92.460 132.255 97.840 132.395 ;
        RECT 92.460 132.195 92.780 132.255 ;
        RECT 97.520 132.195 97.840 132.255 ;
        RECT 99.820 132.395 100.140 132.455 ;
        RECT 101.215 132.395 101.505 132.440 ;
        RECT 99.820 132.255 101.505 132.395 ;
        RECT 99.820 132.195 100.140 132.255 ;
        RECT 101.215 132.210 101.505 132.255 ;
        RECT 20.670 132.055 20.960 132.100 ;
        RECT 23.450 132.055 23.740 132.100 ;
        RECT 25.310 132.055 25.600 132.100 ;
        RECT 20.670 131.915 25.600 132.055 ;
        RECT 20.670 131.870 20.960 131.915 ;
        RECT 23.450 131.870 23.740 131.915 ;
        RECT 25.310 131.870 25.600 131.915 ;
        RECT 31.710 132.055 32.000 132.100 ;
        RECT 34.490 132.055 34.780 132.100 ;
        RECT 36.350 132.055 36.640 132.100 ;
        RECT 31.710 131.915 36.640 132.055 ;
        RECT 31.710 131.870 32.000 131.915 ;
        RECT 34.490 131.870 34.780 131.915 ;
        RECT 36.350 131.870 36.640 131.915 ;
        RECT 40.940 132.055 41.260 132.115 ;
        RECT 44.635 132.055 44.925 132.100 ;
        RECT 47.840 132.055 48.160 132.115 ;
        RECT 40.940 131.915 44.925 132.055 ;
        RECT 40.940 131.855 41.260 131.915 ;
        RECT 44.635 131.870 44.925 131.915 ;
        RECT 46.550 131.915 48.160 132.055 ;
        RECT 22.080 131.715 22.400 131.775 ;
        RECT 23.935 131.715 24.225 131.760 ;
        RECT 22.080 131.575 24.225 131.715 ;
        RECT 22.080 131.515 22.400 131.575 ;
        RECT 23.935 131.530 24.225 131.575 ;
        RECT 25.850 131.575 34.730 131.715 ;
        RECT 20.670 131.375 20.960 131.420 ;
        RECT 25.300 131.375 25.620 131.435 ;
        RECT 25.850 131.420 25.990 131.575 ;
        RECT 25.775 131.375 26.065 131.420 ;
        RECT 20.670 131.235 23.205 131.375 ;
        RECT 20.670 131.190 20.960 131.235 ;
        RECT 17.020 131.035 17.340 131.095 ;
        RECT 22.990 131.080 23.205 131.235 ;
        RECT 25.300 131.235 26.065 131.375 ;
        RECT 25.300 131.175 25.620 131.235 ;
        RECT 25.775 131.190 26.065 131.235 ;
        RECT 26.235 131.375 26.525 131.420 ;
        RECT 28.980 131.375 29.300 131.435 ;
        RECT 26.235 131.235 29.300 131.375 ;
        RECT 26.235 131.190 26.525 131.235 ;
        RECT 28.980 131.175 29.300 131.235 ;
        RECT 31.710 131.375 32.000 131.420 ;
        RECT 34.590 131.375 34.730 131.575 ;
        RECT 34.960 131.515 35.280 131.775 ;
        RECT 38.180 131.715 38.500 131.775 ;
        RECT 38.655 131.715 38.945 131.760 ;
        RECT 38.180 131.575 38.945 131.715 ;
        RECT 38.180 131.515 38.500 131.575 ;
        RECT 38.655 131.530 38.945 131.575 ;
        RECT 36.815 131.375 37.105 131.420 ;
        RECT 31.710 131.235 34.245 131.375 ;
        RECT 34.590 131.235 37.105 131.375 ;
        RECT 31.710 131.190 32.000 131.235 ;
        RECT 18.810 131.035 19.100 131.080 ;
        RECT 22.070 131.035 22.360 131.080 ;
        RECT 17.020 130.895 22.360 131.035 ;
        RECT 17.020 130.835 17.340 130.895 ;
        RECT 18.810 130.850 19.100 130.895 ;
        RECT 22.070 130.850 22.360 130.895 ;
        RECT 22.990 131.035 23.280 131.080 ;
        RECT 24.850 131.035 25.140 131.080 ;
        RECT 22.990 130.895 25.140 131.035 ;
        RECT 22.990 130.850 23.280 130.895 ;
        RECT 24.850 130.850 25.140 130.895 ;
        RECT 29.850 131.035 30.140 131.080 ;
        RECT 30.820 131.035 31.140 131.095 ;
        RECT 34.030 131.080 34.245 131.235 ;
        RECT 36.815 131.190 37.105 131.235 ;
        RECT 39.560 131.375 39.880 131.435 ;
        RECT 42.780 131.375 43.100 131.435 ;
        RECT 43.255 131.375 43.545 131.420 ;
        RECT 39.560 131.235 43.545 131.375 ;
        RECT 39.560 131.175 39.880 131.235 ;
        RECT 42.780 131.175 43.100 131.235 ;
        RECT 43.255 131.190 43.545 131.235 ;
        RECT 43.700 131.175 44.020 131.435 ;
        RECT 44.620 131.375 44.940 131.435 ;
        RECT 46.550 131.420 46.690 131.915 ;
        RECT 47.840 131.855 48.160 131.915 ;
        RECT 52.410 132.055 52.700 132.100 ;
        RECT 55.190 132.055 55.480 132.100 ;
        RECT 57.050 132.055 57.340 132.100 ;
        RECT 52.410 131.915 57.340 132.055 ;
        RECT 52.410 131.870 52.700 131.915 ;
        RECT 55.190 131.870 55.480 131.915 ;
        RECT 57.050 131.870 57.340 131.915 ;
        RECT 66.240 132.055 66.560 132.115 ;
        RECT 69.475 132.055 69.765 132.100 ;
        RECT 66.240 131.915 69.765 132.055 ;
        RECT 66.240 131.855 66.560 131.915 ;
        RECT 69.475 131.870 69.765 131.915 ;
        RECT 105.355 132.055 105.645 132.100 ;
        RECT 105.355 131.915 107.640 132.055 ;
        RECT 105.355 131.870 105.645 131.915 ;
        RECT 48.545 131.715 48.835 131.760 ;
        RECT 47.010 131.575 48.835 131.715 ;
        RECT 47.010 131.435 47.150 131.575 ;
        RECT 48.545 131.530 48.835 131.575 ;
        RECT 55.660 131.515 55.980 131.775 ;
        RECT 59.340 131.515 59.660 131.775 ;
        RECT 60.275 131.715 60.565 131.760 ;
        RECT 60.720 131.715 61.040 131.775 ;
        RECT 60.275 131.575 61.040 131.715 ;
        RECT 60.275 131.530 60.565 131.575 ;
        RECT 60.720 131.515 61.040 131.575 ;
        RECT 67.160 131.515 67.480 131.775 ;
        RECT 74.075 131.715 74.365 131.760 ;
        RECT 74.520 131.715 74.840 131.775 ;
        RECT 87.415 131.715 87.705 131.760 ;
        RECT 74.075 131.575 87.705 131.715 ;
        RECT 74.075 131.530 74.365 131.575 ;
        RECT 74.520 131.515 74.840 131.575 ;
        RECT 87.415 131.530 87.705 131.575 ;
        RECT 88.335 131.715 88.625 131.760 ;
        RECT 98.440 131.715 98.760 131.775 ;
        RECT 102.135 131.715 102.425 131.760 ;
        RECT 88.335 131.575 102.425 131.715 ;
        RECT 107.500 131.715 107.640 131.915 ;
        RECT 107.500 131.575 109.710 131.715 ;
        RECT 88.335 131.530 88.625 131.575 ;
        RECT 98.440 131.515 98.760 131.575 ;
        RECT 102.135 131.530 102.425 131.575 ;
        RECT 46.015 131.375 46.305 131.420 ;
        RECT 44.620 131.235 46.305 131.375 ;
        RECT 44.620 131.175 44.940 131.235 ;
        RECT 46.015 131.190 46.305 131.235 ;
        RECT 46.475 131.190 46.765 131.420 ;
        RECT 46.920 131.175 47.240 131.435 ;
        RECT 47.855 131.190 48.145 131.420 ;
        RECT 52.410 131.375 52.700 131.420 ;
        RECT 57.515 131.375 57.805 131.420 ;
        RECT 66.255 131.375 66.545 131.420 ;
        RECT 67.620 131.375 67.940 131.435 ;
        RECT 68.095 131.375 68.385 131.420 ;
        RECT 52.410 131.235 54.945 131.375 ;
        RECT 52.410 131.190 52.700 131.235 ;
        RECT 33.110 131.035 33.400 131.080 ;
        RECT 29.850 130.895 33.400 131.035 ;
        RECT 29.850 130.850 30.140 130.895 ;
        RECT 30.820 130.835 31.140 130.895 ;
        RECT 33.110 130.850 33.400 130.895 ;
        RECT 34.030 131.035 34.320 131.080 ;
        RECT 35.890 131.035 36.180 131.080 ;
        RECT 47.930 131.035 48.070 131.190 ;
        RECT 34.030 130.895 36.180 131.035 ;
        RECT 34.030 130.850 34.320 130.895 ;
        RECT 35.890 130.850 36.180 130.895 ;
        RECT 46.550 130.895 48.070 131.035 ;
        RECT 50.550 131.035 50.840 131.080 ;
        RECT 51.980 131.035 52.300 131.095 ;
        RECT 54.730 131.080 54.945 131.235 ;
        RECT 57.515 131.235 59.340 131.375 ;
        RECT 57.515 131.190 57.805 131.235 ;
        RECT 53.810 131.035 54.100 131.080 ;
        RECT 50.550 130.895 54.100 131.035 ;
        RECT 46.550 130.755 46.690 130.895 ;
        RECT 50.550 130.850 50.840 130.895 ;
        RECT 51.980 130.835 52.300 130.895 ;
        RECT 53.810 130.850 54.100 130.895 ;
        RECT 54.730 131.035 55.020 131.080 ;
        RECT 56.590 131.035 56.880 131.080 ;
        RECT 54.730 130.895 56.880 131.035 ;
        RECT 59.200 131.035 59.340 131.235 ;
        RECT 66.255 131.235 68.385 131.375 ;
        RECT 66.255 131.190 66.545 131.235 ;
        RECT 67.620 131.175 67.940 131.235 ;
        RECT 68.095 131.190 68.385 131.235 ;
        RECT 70.395 131.190 70.685 131.420 ;
        RECT 73.155 131.375 73.445 131.420 ;
        RECT 70.930 131.235 73.445 131.375 ;
        RECT 60.260 131.035 60.580 131.095 ;
        RECT 70.470 131.035 70.610 131.190 ;
        RECT 59.200 130.895 60.580 131.035 ;
        RECT 54.730 130.850 55.020 130.895 ;
        RECT 56.590 130.850 56.880 130.895 ;
        RECT 60.260 130.835 60.580 130.895 ;
        RECT 62.650 130.895 70.610 131.035 ;
        RECT 26.680 130.495 27.000 130.755 ;
        RECT 46.460 130.495 46.780 130.755 ;
        RECT 55.200 130.695 55.520 130.755 ;
        RECT 62.650 130.740 62.790 130.895 ;
        RECT 60.735 130.695 61.025 130.740 ;
        RECT 55.200 130.555 61.025 130.695 ;
        RECT 55.200 130.495 55.520 130.555 ;
        RECT 60.735 130.510 61.025 130.555 ;
        RECT 62.575 130.510 62.865 130.740 ;
        RECT 64.400 130.695 64.720 130.755 ;
        RECT 65.335 130.695 65.625 130.740 ;
        RECT 64.400 130.555 65.625 130.695 ;
        RECT 64.400 130.495 64.720 130.555 ;
        RECT 65.335 130.510 65.625 130.555 ;
        RECT 68.540 130.695 68.860 130.755 ;
        RECT 70.930 130.695 71.070 131.235 ;
        RECT 73.155 131.190 73.445 131.235 ;
        RECT 84.640 131.175 84.960 131.435 ;
        RECT 86.955 131.375 87.245 131.420 ;
        RECT 94.300 131.375 94.620 131.435 ;
        RECT 86.955 131.235 94.620 131.375 ;
        RECT 86.955 131.190 87.245 131.235 ;
        RECT 94.300 131.175 94.620 131.235 ;
        RECT 98.900 131.175 99.220 131.435 ;
        RECT 99.820 131.175 100.140 131.435 ;
        RECT 100.280 131.175 100.600 131.435 ;
        RECT 103.960 131.375 104.280 131.435 ;
        RECT 109.570 131.420 109.710 131.575 ;
        RECT 107.655 131.375 107.945 131.420 ;
        RECT 103.960 131.235 107.945 131.375 ;
        RECT 103.960 131.175 104.280 131.235 ;
        RECT 107.655 131.190 107.945 131.235 ;
        RECT 109.495 131.190 109.785 131.420 ;
        RECT 99.910 131.035 100.050 131.175 ;
        RECT 103.055 131.035 103.345 131.080 ;
        RECT 99.910 130.895 103.345 131.035 ;
        RECT 103.055 130.850 103.345 130.895 ;
        RECT 68.540 130.555 71.070 130.695 ;
        RECT 68.540 130.495 68.860 130.555 ;
        RECT 103.500 130.495 103.820 130.755 ;
        RECT 108.100 130.495 108.420 130.755 ;
        RECT 110.415 130.695 110.705 130.740 ;
        RECT 112.240 130.695 112.560 130.755 ;
        RECT 110.415 130.555 112.560 130.695 ;
        RECT 110.415 130.510 110.705 130.555 ;
        RECT 112.240 130.495 112.560 130.555 ;
        RECT 14.650 129.875 115.850 130.355 ;
        RECT 20.255 129.490 20.545 129.720 ;
        RECT 18.875 128.995 19.165 129.040 ;
        RECT 20.330 128.995 20.470 129.490 ;
        RECT 22.540 129.475 22.860 129.735 ;
        RECT 34.500 129.675 34.820 129.735 ;
        RECT 35.895 129.675 36.185 129.720 ;
        RECT 34.500 129.535 36.185 129.675 ;
        RECT 34.500 129.475 34.820 129.535 ;
        RECT 35.895 129.490 36.185 129.535 ;
        RECT 38.655 129.675 38.945 129.720 ;
        RECT 43.700 129.675 44.020 129.735 ;
        RECT 38.655 129.535 44.020 129.675 ;
        RECT 38.655 129.490 38.945 129.535 ;
        RECT 43.700 129.475 44.020 129.535 ;
        RECT 53.605 129.675 53.895 129.720 ;
        RECT 54.740 129.675 55.060 129.735 ;
        RECT 53.605 129.535 55.060 129.675 ;
        RECT 53.605 129.490 53.895 129.535 ;
        RECT 54.740 129.475 55.060 129.535 ;
        RECT 70.380 129.475 70.700 129.735 ;
        RECT 74.520 129.475 74.840 129.735 ;
        RECT 77.280 129.475 77.600 129.735 ;
        RECT 93.840 129.675 94.160 129.735 ;
        RECT 94.775 129.675 95.065 129.720 ;
        RECT 93.840 129.535 95.065 129.675 ;
        RECT 93.840 129.475 94.160 129.535 ;
        RECT 94.775 129.490 95.065 129.535 ;
        RECT 22.095 129.335 22.385 129.380 ;
        RECT 23.460 129.335 23.780 129.395 ;
        RECT 22.095 129.195 23.780 129.335 ;
        RECT 22.095 129.150 22.385 129.195 ;
        RECT 23.460 129.135 23.780 129.195 ;
        RECT 25.300 129.335 25.620 129.395 ;
        RECT 26.695 129.335 26.985 129.380 ;
        RECT 25.300 129.195 26.985 129.335 ;
        RECT 25.300 129.135 25.620 129.195 ;
        RECT 26.695 129.150 26.985 129.195 ;
        RECT 35.435 129.335 35.725 129.380 ;
        RECT 41.400 129.335 41.720 129.395 ;
        RECT 35.435 129.195 41.720 129.335 ;
        RECT 35.435 129.150 35.725 129.195 ;
        RECT 41.400 129.135 41.720 129.195 ;
        RECT 55.610 129.335 55.900 129.380 ;
        RECT 57.960 129.335 58.280 129.395 ;
        RECT 58.870 129.335 59.160 129.380 ;
        RECT 55.610 129.195 59.160 129.335 ;
        RECT 55.610 129.150 55.900 129.195 ;
        RECT 57.960 129.135 58.280 129.195 ;
        RECT 58.870 129.150 59.160 129.195 ;
        RECT 59.790 129.335 60.080 129.380 ;
        RECT 61.650 129.335 61.940 129.380 ;
        RECT 59.790 129.195 61.940 129.335 ;
        RECT 59.790 129.150 60.080 129.195 ;
        RECT 61.650 129.150 61.940 129.195 ;
        RECT 84.200 129.335 84.490 129.380 ;
        RECT 86.060 129.335 86.350 129.380 ;
        RECT 84.200 129.195 86.350 129.335 ;
        RECT 84.200 129.150 84.490 129.195 ;
        RECT 86.060 129.150 86.350 129.195 ;
        RECT 86.980 129.335 87.270 129.380 ;
        RECT 87.860 129.335 88.180 129.395 ;
        RECT 90.240 129.335 90.530 129.380 ;
        RECT 86.980 129.195 90.530 129.335 ;
        RECT 86.980 129.150 87.270 129.195 ;
        RECT 18.875 128.855 20.470 128.995 ;
        RECT 36.815 128.995 37.105 129.040 ;
        RECT 37.260 128.995 37.580 129.055 ;
        RECT 36.815 128.855 37.580 128.995 ;
        RECT 18.875 128.810 19.165 128.855 ;
        RECT 36.815 128.810 37.105 128.855 ;
        RECT 37.260 128.795 37.580 128.855 ;
        RECT 38.640 128.995 38.960 129.055 ;
        RECT 39.115 128.995 39.405 129.040 ;
        RECT 38.640 128.855 39.405 128.995 ;
        RECT 38.640 128.795 38.960 128.855 ;
        RECT 39.115 128.810 39.405 128.855 ;
        RECT 57.470 128.995 57.760 129.040 ;
        RECT 59.790 128.995 60.005 129.150 ;
        RECT 57.470 128.855 60.005 128.995 ;
        RECT 57.470 128.810 57.760 128.855 ;
        RECT 60.260 128.795 60.580 129.055 ;
        RECT 60.720 128.795 61.040 129.055 ;
        RECT 64.400 128.995 64.720 129.055 ;
        RECT 64.875 128.995 65.165 129.040 ;
        RECT 66.255 128.995 66.545 129.040 ;
        RECT 64.400 128.855 66.545 128.995 ;
        RECT 64.400 128.795 64.720 128.855 ;
        RECT 64.875 128.810 65.165 128.855 ;
        RECT 66.255 128.810 66.545 128.855 ;
        RECT 68.540 128.995 68.860 129.055 ;
        RECT 71.315 128.995 71.605 129.040 ;
        RECT 78.215 128.995 78.505 129.040 ;
        RECT 68.540 128.855 78.505 128.995 ;
        RECT 68.540 128.795 68.860 128.855 ;
        RECT 71.315 128.810 71.605 128.855 ;
        RECT 78.215 128.810 78.505 128.855 ;
        RECT 85.115 128.995 85.405 129.040 ;
        RECT 85.560 128.995 85.880 129.055 ;
        RECT 85.115 128.855 85.880 128.995 ;
        RECT 86.135 128.995 86.350 129.150 ;
        RECT 87.860 129.135 88.180 129.195 ;
        RECT 90.240 129.150 90.530 129.195 ;
        RECT 92.245 129.335 92.535 129.380 ;
        RECT 94.300 129.335 94.620 129.395 ;
        RECT 99.835 129.335 100.125 129.380 ;
        RECT 92.245 129.195 100.125 129.335 ;
        RECT 92.245 129.150 92.535 129.195 ;
        RECT 94.300 129.135 94.620 129.195 ;
        RECT 99.835 129.150 100.125 129.195 ;
        RECT 107.130 129.335 107.420 129.380 ;
        RECT 108.100 129.335 108.420 129.395 ;
        RECT 110.390 129.335 110.680 129.380 ;
        RECT 107.130 129.195 110.680 129.335 ;
        RECT 107.130 129.150 107.420 129.195 ;
        RECT 108.100 129.135 108.420 129.195 ;
        RECT 110.390 129.150 110.680 129.195 ;
        RECT 111.310 129.335 111.600 129.380 ;
        RECT 113.170 129.335 113.460 129.380 ;
        RECT 111.310 129.195 113.460 129.335 ;
        RECT 111.310 129.150 111.600 129.195 ;
        RECT 113.170 129.150 113.460 129.195 ;
        RECT 88.380 128.995 88.670 129.040 ;
        RECT 86.135 128.855 88.670 128.995 ;
        RECT 85.115 128.810 85.405 128.855 ;
        RECT 85.560 128.795 85.880 128.855 ;
        RECT 88.380 128.810 88.670 128.855 ;
        RECT 95.695 128.995 95.985 129.040 ;
        RECT 95.695 128.855 99.590 128.995 ;
        RECT 95.695 128.810 95.985 128.855 ;
        RECT 23.475 128.655 23.765 128.700 ;
        RECT 30.820 128.655 31.140 128.715 ;
        RECT 23.475 128.515 31.140 128.655 ;
        RECT 23.475 128.470 23.765 128.515 ;
        RECT 30.820 128.455 31.140 128.515 ;
        RECT 38.195 128.655 38.485 128.700 ;
        RECT 60.350 128.655 60.490 128.795 ;
        RECT 62.575 128.655 62.865 128.700 ;
        RECT 38.195 128.515 52.210 128.655 ;
        RECT 60.350 128.515 62.865 128.655 ;
        RECT 38.195 128.470 38.485 128.515 ;
        RECT 52.070 128.035 52.210 128.515 ;
        RECT 62.575 128.470 62.865 128.515 ;
        RECT 69.460 128.655 69.780 128.715 ;
        RECT 72.235 128.655 72.525 128.700 ;
        RECT 69.460 128.515 72.525 128.655 ;
        RECT 69.460 128.455 69.780 128.515 ;
        RECT 72.235 128.470 72.525 128.515 ;
        RECT 73.155 128.470 73.445 128.700 ;
        RECT 57.470 128.315 57.760 128.360 ;
        RECT 60.250 128.315 60.540 128.360 ;
        RECT 62.110 128.315 62.400 128.360 ;
        RECT 73.230 128.315 73.370 128.470 ;
        RECT 74.060 128.455 74.380 128.715 ;
        RECT 79.120 128.455 79.440 128.715 ;
        RECT 83.275 128.655 83.565 128.700 ;
        RECT 84.180 128.655 84.500 128.715 ;
        RECT 83.275 128.515 84.500 128.655 ;
        RECT 83.275 128.470 83.565 128.515 ;
        RECT 84.180 128.455 84.500 128.515 ;
        RECT 96.615 128.655 96.905 128.700 ;
        RECT 97.520 128.655 97.840 128.715 ;
        RECT 96.615 128.515 97.840 128.655 ;
        RECT 96.615 128.470 96.905 128.515 ;
        RECT 97.520 128.455 97.840 128.515 ;
        RECT 98.440 128.655 98.760 128.715 ;
        RECT 98.915 128.655 99.205 128.700 ;
        RECT 98.440 128.515 99.205 128.655 ;
        RECT 99.450 128.655 99.590 128.855 ;
        RECT 100.280 128.795 100.600 129.055 ;
        RECT 103.960 128.995 104.280 129.055 ;
        RECT 104.435 128.995 104.725 129.040 ;
        RECT 103.960 128.855 104.725 128.995 ;
        RECT 103.960 128.795 104.280 128.855 ;
        RECT 104.435 128.810 104.725 128.855 ;
        RECT 108.990 128.995 109.280 129.040 ;
        RECT 111.310 128.995 111.525 129.150 ;
        RECT 108.990 128.855 111.525 128.995 ;
        RECT 108.990 128.810 109.280 128.855 ;
        RECT 112.240 128.795 112.560 129.055 ;
        RECT 114.080 128.795 114.400 129.055 ;
        RECT 100.740 128.655 101.060 128.715 ;
        RECT 99.450 128.515 101.060 128.655 ;
        RECT 98.440 128.455 98.760 128.515 ;
        RECT 98.915 128.470 99.205 128.515 ;
        RECT 100.740 128.455 101.060 128.515 ;
        RECT 57.470 128.175 62.400 128.315 ;
        RECT 57.470 128.130 57.760 128.175 ;
        RECT 60.250 128.130 60.540 128.175 ;
        RECT 62.110 128.130 62.400 128.175 ;
        RECT 72.310 128.175 73.370 128.315 ;
        RECT 83.740 128.315 84.030 128.360 ;
        RECT 85.600 128.315 85.890 128.360 ;
        RECT 88.380 128.315 88.670 128.360 ;
        RECT 83.740 128.175 88.670 128.315 ;
        RECT 72.310 128.035 72.450 128.175 ;
        RECT 83.740 128.130 84.030 128.175 ;
        RECT 85.600 128.130 85.890 128.175 ;
        RECT 88.380 128.130 88.670 128.175 ;
        RECT 97.060 128.315 97.380 128.375 ;
        RECT 103.500 128.315 103.820 128.375 ;
        RECT 105.125 128.315 105.415 128.360 ;
        RECT 97.060 128.175 105.415 128.315 ;
        RECT 97.060 128.115 97.380 128.175 ;
        RECT 103.500 128.115 103.820 128.175 ;
        RECT 105.125 128.130 105.415 128.175 ;
        RECT 108.990 128.315 109.280 128.360 ;
        RECT 111.770 128.315 112.060 128.360 ;
        RECT 113.630 128.315 113.920 128.360 ;
        RECT 108.990 128.175 113.920 128.315 ;
        RECT 108.990 128.130 109.280 128.175 ;
        RECT 111.770 128.130 112.060 128.175 ;
        RECT 113.630 128.130 113.920 128.175 ;
        RECT 19.795 127.975 20.085 128.020 ;
        RECT 23.920 127.975 24.240 128.035 ;
        RECT 19.795 127.835 24.240 127.975 ;
        RECT 19.795 127.790 20.085 127.835 ;
        RECT 23.920 127.775 24.240 127.835 ;
        RECT 39.560 127.975 39.880 128.035 ;
        RECT 40.955 127.975 41.245 128.020 ;
        RECT 39.560 127.835 41.245 127.975 ;
        RECT 39.560 127.775 39.880 127.835 ;
        RECT 40.955 127.790 41.245 127.835 ;
        RECT 48.760 127.775 49.080 128.035 ;
        RECT 51.980 127.975 52.300 128.035 ;
        RECT 63.495 127.975 63.785 128.020 ;
        RECT 51.980 127.835 63.785 127.975 ;
        RECT 51.980 127.775 52.300 127.835 ;
        RECT 63.495 127.790 63.785 127.835 ;
        RECT 67.635 127.975 67.925 128.020 ;
        RECT 72.220 127.975 72.540 128.035 ;
        RECT 67.635 127.835 72.540 127.975 ;
        RECT 67.635 127.790 67.925 127.835 ;
        RECT 72.220 127.775 72.540 127.835 ;
        RECT 76.360 127.775 76.680 128.035 ;
        RECT 101.200 127.975 101.520 128.035 ;
        RECT 102.135 127.975 102.425 128.020 ;
        RECT 101.200 127.835 102.425 127.975 ;
        RECT 101.200 127.775 101.520 127.835 ;
        RECT 102.135 127.790 102.425 127.835 ;
        RECT 103.975 127.975 104.265 128.020 ;
        RECT 104.420 127.975 104.740 128.035 ;
        RECT 103.975 127.835 104.740 127.975 ;
        RECT 103.975 127.790 104.265 127.835 ;
        RECT 104.420 127.775 104.740 127.835 ;
        RECT 14.650 127.155 115.850 127.635 ;
        RECT 37.260 127.000 37.580 127.015 ;
        RECT 37.260 126.955 37.795 127.000 ;
        RECT 38.180 126.955 38.500 127.015 ;
        RECT 37.260 126.815 38.500 126.955 ;
        RECT 37.260 126.770 37.795 126.815 ;
        RECT 37.260 126.755 37.580 126.770 ;
        RECT 38.180 126.755 38.500 126.815 ;
        RECT 47.380 126.955 47.700 127.015 ;
        RECT 50.615 126.955 50.905 127.000 ;
        RECT 47.380 126.815 50.905 126.955 ;
        RECT 47.380 126.755 47.700 126.815 ;
        RECT 50.615 126.770 50.905 126.815 ;
        RECT 57.515 126.955 57.805 127.000 ;
        RECT 57.960 126.955 58.280 127.015 ;
        RECT 57.515 126.815 58.280 126.955 ;
        RECT 57.515 126.770 57.805 126.815 ;
        RECT 57.960 126.755 58.280 126.815 ;
        RECT 59.355 126.955 59.645 127.000 ;
        RECT 60.720 126.955 61.040 127.015 ;
        RECT 59.355 126.815 61.040 126.955 ;
        RECT 59.355 126.770 59.645 126.815 ;
        RECT 60.720 126.755 61.040 126.815 ;
        RECT 71.300 126.755 71.620 127.015 ;
        RECT 73.845 126.955 74.135 127.000 ;
        RECT 74.520 126.955 74.840 127.015 ;
        RECT 73.845 126.815 74.840 126.955 ;
        RECT 73.845 126.770 74.135 126.815 ;
        RECT 74.520 126.755 74.840 126.815 ;
        RECT 76.360 126.955 76.680 127.015 ;
        RECT 87.415 126.955 87.705 127.000 ;
        RECT 87.860 126.955 88.180 127.015 ;
        RECT 100.280 127.000 100.600 127.015 ;
        RECT 76.360 126.815 84.870 126.955 ;
        RECT 76.360 126.755 76.680 126.815 ;
        RECT 20.670 126.615 20.960 126.660 ;
        RECT 23.450 126.615 23.740 126.660 ;
        RECT 25.310 126.615 25.600 126.660 ;
        RECT 20.670 126.475 25.600 126.615 ;
        RECT 20.670 126.430 20.960 126.475 ;
        RECT 23.450 126.430 23.740 126.475 ;
        RECT 25.310 126.430 25.600 126.475 ;
        RECT 29.000 126.615 29.290 126.660 ;
        RECT 30.860 126.615 31.150 126.660 ;
        RECT 33.640 126.615 33.930 126.660 ;
        RECT 68.540 126.615 68.860 126.675 ;
        RECT 72.220 126.615 72.540 126.675 ;
        RECT 29.000 126.475 33.930 126.615 ;
        RECT 29.000 126.430 29.290 126.475 ;
        RECT 30.860 126.430 31.150 126.475 ;
        RECT 33.640 126.430 33.930 126.475 ;
        RECT 51.610 126.475 68.860 126.615 ;
        RECT 23.920 126.075 24.240 126.335 ;
        RECT 28.535 126.275 28.825 126.320 ;
        RECT 29.900 126.275 30.220 126.335 ;
        RECT 25.850 126.135 30.220 126.275 ;
        RECT 20.670 125.935 20.960 125.980 ;
        RECT 25.300 125.935 25.620 125.995 ;
        RECT 25.850 125.980 25.990 126.135 ;
        RECT 28.535 126.090 28.825 126.135 ;
        RECT 29.900 126.075 30.220 126.135 ;
        RECT 42.780 126.275 43.100 126.335 ;
        RECT 51.610 126.275 51.750 126.475 ;
        RECT 68.540 126.415 68.860 126.475 ;
        RECT 70.470 126.475 72.540 126.615 ;
        RECT 58.880 126.275 59.200 126.335 ;
        RECT 42.780 126.135 51.750 126.275 ;
        RECT 42.780 126.075 43.100 126.135 ;
        RECT 25.775 125.935 26.065 125.980 ;
        RECT 20.670 125.795 23.205 125.935 ;
        RECT 20.670 125.750 20.960 125.795 ;
        RECT 18.860 125.640 19.180 125.655 ;
        RECT 22.990 125.640 23.205 125.795 ;
        RECT 25.300 125.795 26.065 125.935 ;
        RECT 25.300 125.735 25.620 125.795 ;
        RECT 25.775 125.750 26.065 125.795 ;
        RECT 28.060 125.735 28.380 125.995 ;
        RECT 30.360 125.735 30.680 125.995 ;
        RECT 33.640 125.935 33.930 125.980 ;
        RECT 31.395 125.795 33.930 125.935 ;
        RECT 31.395 125.640 31.610 125.795 ;
        RECT 33.640 125.750 33.930 125.795 ;
        RECT 48.760 125.935 49.080 125.995 ;
        RECT 51.610 125.980 51.750 126.135 ;
        RECT 58.050 126.135 59.200 126.275 ;
        RECT 58.050 125.980 58.190 126.135 ;
        RECT 58.880 126.075 59.200 126.135 ;
        RECT 49.235 125.935 49.525 125.980 ;
        RECT 48.760 125.795 49.525 125.935 ;
        RECT 48.760 125.735 49.080 125.795 ;
        RECT 49.235 125.750 49.525 125.795 ;
        RECT 51.535 125.750 51.825 125.980 ;
        RECT 51.995 125.750 52.285 125.980 ;
        RECT 57.975 125.750 58.265 125.980 ;
        RECT 18.810 125.595 19.180 125.640 ;
        RECT 22.070 125.595 22.360 125.640 ;
        RECT 18.810 125.455 22.360 125.595 ;
        RECT 18.810 125.410 19.180 125.455 ;
        RECT 22.070 125.410 22.360 125.455 ;
        RECT 22.990 125.595 23.280 125.640 ;
        RECT 24.850 125.595 25.140 125.640 ;
        RECT 22.990 125.455 25.140 125.595 ;
        RECT 22.990 125.410 23.280 125.455 ;
        RECT 24.850 125.410 25.140 125.455 ;
        RECT 29.460 125.595 29.750 125.640 ;
        RECT 31.320 125.595 31.610 125.640 ;
        RECT 29.460 125.455 31.610 125.595 ;
        RECT 29.460 125.410 29.750 125.455 ;
        RECT 31.320 125.410 31.610 125.455 ;
        RECT 32.200 125.640 32.520 125.655 ;
        RECT 32.200 125.595 32.530 125.640 ;
        RECT 35.500 125.595 35.790 125.640 ;
        RECT 52.070 125.595 52.210 125.750 ;
        RECT 58.420 125.735 58.740 125.995 ;
        RECT 32.200 125.455 35.790 125.595 ;
        RECT 32.200 125.410 32.530 125.455 ;
        RECT 35.500 125.410 35.790 125.455 ;
        RECT 49.310 125.455 52.210 125.595 ;
        RECT 68.630 125.595 68.770 126.415 ;
        RECT 70.470 126.320 70.610 126.475 ;
        RECT 72.220 126.415 72.540 126.475 ;
        RECT 77.710 126.615 78.000 126.660 ;
        RECT 80.490 126.615 80.780 126.660 ;
        RECT 82.350 126.615 82.640 126.660 ;
        RECT 77.710 126.475 82.640 126.615 ;
        RECT 77.710 126.430 78.000 126.475 ;
        RECT 80.490 126.430 80.780 126.475 ;
        RECT 82.350 126.430 82.640 126.475 ;
        RECT 84.180 126.415 84.500 126.675 ;
        RECT 70.395 126.090 70.685 126.320 ;
        RECT 73.155 126.275 73.445 126.320 ;
        RECT 74.060 126.275 74.380 126.335 ;
        RECT 71.850 126.135 74.380 126.275 ;
        RECT 69.015 125.935 69.305 125.980 ;
        RECT 71.850 125.935 71.990 126.135 ;
        RECT 73.155 126.090 73.445 126.135 ;
        RECT 74.060 126.075 74.380 126.135 ;
        RECT 82.815 126.275 83.105 126.320 ;
        RECT 84.270 126.275 84.410 126.415 ;
        RECT 82.815 126.135 84.410 126.275 ;
        RECT 82.815 126.090 83.105 126.135 ;
        RECT 69.015 125.795 71.990 125.935 ;
        RECT 69.015 125.750 69.305 125.795 ;
        RECT 72.235 125.750 72.525 125.980 ;
        RECT 77.710 125.935 78.000 125.980 ;
        RECT 80.975 125.935 81.265 125.980 ;
        RECT 84.195 125.935 84.485 125.980 ;
        RECT 84.730 125.935 84.870 126.815 ;
        RECT 87.415 126.815 88.180 126.955 ;
        RECT 87.415 126.770 87.705 126.815 ;
        RECT 87.860 126.755 88.180 126.815 ;
        RECT 100.065 126.770 100.600 127.000 ;
        RECT 100.280 126.755 100.600 126.770 ;
        RECT 98.440 126.615 98.760 126.675 ;
        RECT 96.690 126.475 98.760 126.615 ;
        RECT 96.690 126.320 96.830 126.475 ;
        RECT 98.440 126.415 98.760 126.475 ;
        RECT 103.930 126.615 104.220 126.660 ;
        RECT 106.710 126.615 107.000 126.660 ;
        RECT 108.570 126.615 108.860 126.660 ;
        RECT 103.930 126.475 108.860 126.615 ;
        RECT 103.930 126.430 104.220 126.475 ;
        RECT 106.710 126.430 107.000 126.475 ;
        RECT 108.570 126.430 108.860 126.475 ;
        RECT 93.395 126.275 93.685 126.320 ;
        RECT 96.615 126.275 96.905 126.320 ;
        RECT 93.395 126.135 96.905 126.275 ;
        RECT 93.395 126.090 93.685 126.135 ;
        RECT 96.615 126.090 96.905 126.135 ;
        RECT 97.060 126.075 97.380 126.335 ;
        RECT 102.120 126.275 102.440 126.335 ;
        RECT 107.195 126.275 107.485 126.320 ;
        RECT 102.120 126.135 107.485 126.275 ;
        RECT 102.120 126.075 102.440 126.135 ;
        RECT 107.195 126.090 107.485 126.135 ;
        RECT 109.020 126.275 109.340 126.335 ;
        RECT 114.080 126.275 114.400 126.335 ;
        RECT 109.020 126.135 114.400 126.275 ;
        RECT 109.020 126.075 109.340 126.135 ;
        RECT 114.080 126.075 114.400 126.135 ;
        RECT 77.710 125.795 80.245 125.935 ;
        RECT 77.710 125.750 78.000 125.795 ;
        RECT 72.310 125.595 72.450 125.750 ;
        RECT 68.630 125.455 72.450 125.595 ;
        RECT 75.850 125.595 76.140 125.640 ;
        RECT 78.200 125.595 78.520 125.655 ;
        RECT 80.030 125.640 80.245 125.795 ;
        RECT 80.975 125.795 83.490 125.935 ;
        RECT 80.975 125.750 81.265 125.795 ;
        RECT 79.110 125.595 79.400 125.640 ;
        RECT 75.850 125.455 79.400 125.595 ;
        RECT 18.860 125.395 19.180 125.410 ;
        RECT 32.200 125.395 32.520 125.410 ;
        RECT 49.310 125.315 49.450 125.455 ;
        RECT 75.850 125.410 76.140 125.455 ;
        RECT 78.200 125.395 78.520 125.455 ;
        RECT 79.110 125.410 79.400 125.455 ;
        RECT 80.030 125.595 80.320 125.640 ;
        RECT 81.890 125.595 82.180 125.640 ;
        RECT 80.030 125.455 82.180 125.595 ;
        RECT 80.030 125.410 80.320 125.455 ;
        RECT 81.890 125.410 82.180 125.455 ;
        RECT 16.805 125.255 17.095 125.300 ;
        RECT 23.460 125.255 23.780 125.315 ;
        RECT 16.805 125.115 23.780 125.255 ;
        RECT 16.805 125.070 17.095 125.115 ;
        RECT 23.460 125.055 23.780 125.115 ;
        RECT 27.140 125.055 27.460 125.315 ;
        RECT 49.220 125.055 49.540 125.315 ;
        RECT 67.175 125.255 67.465 125.300 ;
        RECT 68.540 125.255 68.860 125.315 ;
        RECT 67.175 125.115 68.860 125.255 ;
        RECT 67.175 125.070 67.465 125.115 ;
        RECT 68.540 125.055 68.860 125.115 ;
        RECT 69.460 125.055 69.780 125.315 ;
        RECT 83.350 125.300 83.490 125.795 ;
        RECT 84.195 125.795 84.870 125.935 ;
        RECT 86.955 125.935 87.245 125.980 ;
        RECT 91.080 125.935 91.400 125.995 ;
        RECT 86.955 125.795 91.400 125.935 ;
        RECT 84.195 125.750 84.485 125.795 ;
        RECT 86.955 125.750 87.245 125.795 ;
        RECT 91.080 125.735 91.400 125.795 ;
        RECT 92.000 125.735 92.320 125.995 ;
        RECT 103.930 125.935 104.220 125.980 ;
        RECT 109.495 125.935 109.785 125.980 ;
        RECT 103.930 125.795 106.465 125.935 ;
        RECT 103.930 125.750 104.220 125.795 ;
        RECT 102.070 125.595 102.360 125.640 ;
        RECT 104.420 125.595 104.740 125.655 ;
        RECT 106.250 125.640 106.465 125.795 ;
        RECT 108.650 125.795 109.785 125.935 ;
        RECT 105.330 125.595 105.620 125.640 ;
        RECT 102.070 125.455 105.620 125.595 ;
        RECT 102.070 125.410 102.360 125.455 ;
        RECT 104.420 125.395 104.740 125.455 ;
        RECT 105.330 125.410 105.620 125.455 ;
        RECT 106.250 125.595 106.540 125.640 ;
        RECT 108.110 125.595 108.400 125.640 ;
        RECT 106.250 125.455 108.400 125.595 ;
        RECT 106.250 125.410 106.540 125.455 ;
        RECT 108.110 125.410 108.400 125.455 ;
        RECT 83.275 125.070 83.565 125.300 ;
        RECT 90.175 125.255 90.465 125.300 ;
        RECT 90.620 125.255 90.940 125.315 ;
        RECT 90.175 125.115 90.940 125.255 ;
        RECT 90.175 125.070 90.465 125.115 ;
        RECT 90.620 125.055 90.940 125.115 ;
        RECT 92.000 125.255 92.320 125.315 ;
        RECT 92.475 125.255 92.765 125.300 ;
        RECT 92.000 125.115 92.765 125.255 ;
        RECT 92.000 125.055 92.320 125.115 ;
        RECT 92.475 125.070 92.765 125.115 ;
        RECT 97.535 125.255 97.825 125.300 ;
        RECT 97.980 125.255 98.300 125.315 ;
        RECT 97.535 125.115 98.300 125.255 ;
        RECT 97.535 125.070 97.825 125.115 ;
        RECT 97.980 125.055 98.300 125.115 ;
        RECT 99.375 125.255 99.665 125.300 ;
        RECT 108.650 125.255 108.790 125.795 ;
        RECT 109.495 125.750 109.785 125.795 ;
        RECT 99.375 125.115 108.790 125.255 ;
        RECT 99.375 125.070 99.665 125.115 ;
        RECT 110.400 125.055 110.720 125.315 ;
        RECT 14.650 124.435 115.850 124.915 ;
        RECT 17.020 124.035 17.340 124.295 ;
        RECT 18.415 124.235 18.705 124.280 ;
        RECT 18.860 124.235 19.180 124.295 ;
        RECT 18.415 124.095 19.180 124.235 ;
        RECT 18.415 124.050 18.705 124.095 ;
        RECT 18.860 124.035 19.180 124.095 ;
        RECT 20.255 124.235 20.545 124.280 ;
        RECT 22.080 124.235 22.400 124.295 ;
        RECT 20.255 124.095 22.400 124.235 ;
        RECT 20.255 124.050 20.545 124.095 ;
        RECT 22.080 124.035 22.400 124.095 ;
        RECT 23.015 124.235 23.305 124.280 ;
        RECT 23.460 124.235 23.780 124.295 ;
        RECT 23.015 124.095 23.780 124.235 ;
        RECT 23.015 124.050 23.305 124.095 ;
        RECT 23.460 124.035 23.780 124.095 ;
        RECT 26.695 124.235 26.985 124.280 ;
        RECT 28.060 124.235 28.380 124.295 ;
        RECT 26.695 124.095 28.380 124.235 ;
        RECT 26.695 124.050 26.985 124.095 ;
        RECT 28.060 124.035 28.380 124.095 ;
        RECT 30.360 124.235 30.680 124.295 ;
        RECT 31.755 124.235 32.045 124.280 ;
        RECT 30.360 124.095 32.045 124.235 ;
        RECT 30.360 124.035 30.680 124.095 ;
        RECT 31.755 124.050 32.045 124.095 ;
        RECT 35.205 124.235 35.495 124.280 ;
        RECT 38.180 124.235 38.500 124.295 ;
        RECT 35.205 124.095 38.500 124.235 ;
        RECT 35.205 124.050 35.495 124.095 ;
        RECT 38.180 124.035 38.500 124.095 ;
        RECT 44.635 124.235 44.925 124.280 ;
        RECT 45.080 124.235 45.400 124.295 ;
        RECT 44.635 124.095 45.400 124.235 ;
        RECT 44.635 124.050 44.925 124.095 ;
        RECT 45.080 124.035 45.400 124.095 ;
        RECT 77.755 124.235 78.045 124.280 ;
        RECT 78.200 124.235 78.520 124.295 ;
        RECT 77.755 124.095 78.520 124.235 ;
        RECT 77.755 124.050 78.045 124.095 ;
        RECT 78.200 124.035 78.520 124.095 ;
        RECT 80.975 124.235 81.265 124.280 ;
        RECT 83.965 124.235 84.255 124.280 ;
        RECT 91.540 124.235 91.860 124.295 ;
        RECT 80.975 124.095 91.860 124.235 ;
        RECT 80.975 124.050 81.265 124.095 ;
        RECT 83.965 124.050 84.255 124.095 ;
        RECT 91.540 124.035 91.860 124.095 ;
        RECT 97.535 124.235 97.825 124.280 ;
        RECT 97.980 124.235 98.300 124.295 ;
        RECT 97.535 124.095 98.300 124.235 ;
        RECT 97.535 124.050 97.825 124.095 ;
        RECT 28.980 123.895 29.300 123.955 ;
        RECT 18.030 123.755 29.300 123.895 ;
        RECT 18.030 123.600 18.170 123.755 ;
        RECT 28.980 123.695 29.300 123.755 ;
        RECT 29.900 123.895 30.220 123.955 ;
        RECT 37.210 123.895 37.500 123.940 ;
        RECT 38.640 123.895 38.960 123.955 ;
        RECT 65.320 123.940 65.640 123.955 ;
        RECT 40.470 123.895 40.760 123.940 ;
        RECT 29.900 123.755 33.810 123.895 ;
        RECT 29.900 123.695 30.220 123.755 ;
        RECT 17.495 123.555 17.785 123.600 ;
        RECT 17.955 123.555 18.245 123.600 ;
        RECT 17.495 123.415 18.245 123.555 ;
        RECT 17.495 123.370 17.785 123.415 ;
        RECT 17.955 123.370 18.245 123.415 ;
        RECT 19.335 123.555 19.625 123.600 ;
        RECT 22.555 123.555 22.845 123.600 ;
        RECT 23.000 123.555 23.320 123.615 ;
        RECT 28.535 123.555 28.825 123.600 ;
        RECT 31.740 123.555 32.060 123.615 ;
        RECT 19.335 123.415 20.930 123.555 ;
        RECT 19.335 123.370 19.625 123.415 ;
        RECT 20.790 122.920 20.930 123.415 ;
        RECT 22.555 123.415 26.450 123.555 ;
        RECT 22.555 123.370 22.845 123.415 ;
        RECT 23.000 123.355 23.320 123.415 ;
        RECT 23.935 123.215 24.225 123.260 ;
        RECT 26.310 123.215 26.450 123.415 ;
        RECT 28.535 123.415 32.060 123.555 ;
        RECT 28.535 123.370 28.825 123.415 ;
        RECT 31.740 123.355 32.060 123.415 ;
        RECT 32.675 123.555 32.965 123.600 ;
        RECT 33.120 123.555 33.440 123.615 ;
        RECT 33.670 123.600 33.810 123.755 ;
        RECT 37.210 123.755 40.760 123.895 ;
        RECT 37.210 123.710 37.500 123.755 ;
        RECT 38.640 123.695 38.960 123.755 ;
        RECT 40.470 123.710 40.760 123.755 ;
        RECT 41.390 123.895 41.680 123.940 ;
        RECT 43.250 123.895 43.540 123.940 ;
        RECT 62.580 123.895 62.870 123.940 ;
        RECT 64.440 123.895 64.730 123.940 ;
        RECT 41.390 123.755 43.540 123.895 ;
        RECT 41.390 123.710 41.680 123.755 ;
        RECT 43.250 123.710 43.540 123.755 ;
        RECT 46.090 123.755 54.050 123.895 ;
        RECT 32.675 123.415 33.440 123.555 ;
        RECT 32.675 123.370 32.965 123.415 ;
        RECT 33.120 123.355 33.440 123.415 ;
        RECT 33.595 123.370 33.885 123.600 ;
        RECT 39.070 123.555 39.360 123.600 ;
        RECT 41.390 123.555 41.605 123.710 ;
        RECT 39.070 123.415 41.605 123.555 ;
        RECT 42.780 123.555 43.100 123.615 ;
        RECT 45.555 123.555 45.845 123.600 ;
        RECT 42.780 123.415 45.845 123.555 ;
        RECT 39.070 123.370 39.360 123.415 ;
        RECT 42.780 123.355 43.100 123.415 ;
        RECT 45.555 123.370 45.845 123.415 ;
        RECT 28.995 123.215 29.285 123.260 ;
        RECT 23.935 123.075 25.990 123.215 ;
        RECT 26.310 123.075 29.285 123.215 ;
        RECT 23.935 123.030 24.225 123.075 ;
        RECT 20.715 122.690 21.005 122.920 ;
        RECT 25.850 122.535 25.990 123.075 ;
        RECT 28.995 123.030 29.285 123.075 ;
        RECT 29.900 123.215 30.220 123.275 ;
        RECT 30.820 123.215 31.140 123.275 ;
        RECT 29.900 123.075 31.140 123.215 ;
        RECT 29.070 122.875 29.210 123.030 ;
        RECT 29.900 123.015 30.220 123.075 ;
        RECT 30.820 123.015 31.140 123.075 ;
        RECT 40.480 123.215 40.800 123.275 ;
        RECT 42.335 123.215 42.625 123.260 ;
        RECT 40.480 123.075 42.625 123.215 ;
        RECT 40.480 123.015 40.800 123.075 ;
        RECT 42.335 123.030 42.625 123.075 ;
        RECT 44.175 123.030 44.465 123.260 ;
        RECT 45.080 123.215 45.400 123.275 ;
        RECT 46.090 123.215 46.230 123.755 ;
        RECT 48.315 123.555 48.605 123.600 ;
        RECT 46.550 123.415 48.605 123.555 ;
        RECT 46.550 123.275 46.690 123.415 ;
        RECT 48.315 123.370 48.605 123.415 ;
        RECT 48.775 123.555 49.065 123.600 ;
        RECT 49.220 123.555 49.540 123.615 ;
        RECT 53.910 123.600 54.050 123.755 ;
        RECT 62.580 123.755 64.730 123.895 ;
        RECT 62.580 123.710 62.870 123.755 ;
        RECT 64.440 123.710 64.730 123.755 ;
        RECT 48.775 123.415 49.540 123.555 ;
        RECT 48.775 123.370 49.065 123.415 ;
        RECT 49.220 123.355 49.540 123.415 ;
        RECT 53.835 123.555 54.125 123.600 ;
        RECT 56.135 123.555 56.425 123.600 ;
        RECT 53.835 123.415 56.425 123.555 ;
        RECT 53.835 123.370 54.125 123.415 ;
        RECT 56.135 123.370 56.425 123.415 ;
        RECT 57.515 123.555 57.805 123.600 ;
        RECT 58.880 123.555 59.200 123.615 ;
        RECT 57.515 123.415 59.200 123.555 ;
        RECT 57.515 123.370 57.805 123.415 ;
        RECT 58.880 123.355 59.200 123.415 ;
        RECT 60.260 123.555 60.580 123.615 ;
        RECT 61.655 123.555 61.945 123.600 ;
        RECT 60.260 123.415 61.945 123.555 ;
        RECT 64.515 123.555 64.730 123.710 ;
        RECT 65.320 123.895 65.650 123.940 ;
        RECT 68.620 123.895 68.910 123.940 ;
        RECT 65.320 123.755 68.910 123.895 ;
        RECT 65.320 123.710 65.650 123.755 ;
        RECT 68.620 123.710 68.910 123.755 ;
        RECT 70.625 123.895 70.915 123.940 ;
        RECT 74.060 123.895 74.380 123.955 ;
        RECT 86.020 123.940 86.340 123.955 ;
        RECT 70.625 123.755 74.380 123.895 ;
        RECT 70.625 123.710 70.915 123.755 ;
        RECT 65.320 123.695 65.640 123.710 ;
        RECT 74.060 123.695 74.380 123.755 ;
        RECT 85.970 123.895 86.340 123.940 ;
        RECT 89.230 123.895 89.520 123.940 ;
        RECT 85.970 123.755 89.520 123.895 ;
        RECT 85.970 123.710 86.340 123.755 ;
        RECT 89.230 123.710 89.520 123.755 ;
        RECT 90.150 123.895 90.440 123.940 ;
        RECT 92.010 123.895 92.300 123.940 ;
        RECT 90.150 123.755 92.300 123.895 ;
        RECT 97.610 123.895 97.750 124.050 ;
        RECT 97.980 124.035 98.300 124.095 ;
        RECT 102.120 124.035 102.440 124.295 ;
        RECT 103.285 123.895 103.575 123.940 ;
        RECT 97.610 123.755 103.575 123.895 ;
        RECT 90.150 123.710 90.440 123.755 ;
        RECT 92.010 123.710 92.300 123.755 ;
        RECT 103.285 123.710 103.575 123.755 ;
        RECT 105.290 123.895 105.580 123.940 ;
        RECT 106.260 123.895 106.580 123.955 ;
        RECT 108.550 123.895 108.840 123.940 ;
        RECT 105.290 123.755 108.840 123.895 ;
        RECT 105.290 123.710 105.580 123.755 ;
        RECT 86.020 123.695 86.340 123.710 ;
        RECT 66.760 123.555 67.050 123.600 ;
        RECT 64.515 123.415 67.050 123.555 ;
        RECT 60.260 123.355 60.580 123.415 ;
        RECT 61.655 123.370 61.945 123.415 ;
        RECT 66.760 123.370 67.050 123.415 ;
        RECT 69.460 123.555 69.780 123.615 ;
        RECT 73.155 123.555 73.445 123.600 ;
        RECT 69.460 123.415 73.445 123.555 ;
        RECT 69.460 123.355 69.780 123.415 ;
        RECT 73.155 123.370 73.445 123.415 ;
        RECT 78.200 123.355 78.520 123.615 ;
        RECT 81.435 123.555 81.725 123.600 ;
        RECT 80.130 123.415 81.725 123.555 ;
        RECT 45.080 123.075 46.230 123.215 ;
        RECT 33.580 122.875 33.900 122.935 ;
        RECT 29.070 122.735 33.900 122.875 ;
        RECT 33.580 122.675 33.900 122.735 ;
        RECT 39.070 122.875 39.360 122.920 ;
        RECT 41.850 122.875 42.140 122.920 ;
        RECT 43.710 122.875 44.000 122.920 ;
        RECT 39.070 122.735 44.000 122.875 ;
        RECT 44.250 122.875 44.390 123.030 ;
        RECT 45.080 123.015 45.400 123.075 ;
        RECT 46.460 123.015 46.780 123.275 ;
        RECT 47.840 123.215 48.160 123.275 ;
        RECT 51.980 123.215 52.300 123.275 ;
        RECT 47.840 123.075 52.300 123.215 ;
        RECT 47.840 123.015 48.160 123.075 ;
        RECT 51.980 123.015 52.300 123.075 ;
        RECT 63.480 123.015 63.800 123.275 ;
        RECT 72.220 123.015 72.540 123.275 ;
        RECT 72.695 123.215 72.985 123.260 ;
        RECT 79.120 123.215 79.440 123.275 ;
        RECT 80.130 123.215 80.270 123.415 ;
        RECT 81.435 123.370 81.725 123.415 ;
        RECT 87.830 123.555 88.120 123.600 ;
        RECT 90.150 123.555 90.365 123.710 ;
        RECT 106.260 123.695 106.580 123.755 ;
        RECT 108.550 123.710 108.840 123.755 ;
        RECT 109.470 123.895 109.760 123.940 ;
        RECT 111.330 123.895 111.620 123.940 ;
        RECT 109.470 123.755 111.620 123.895 ;
        RECT 109.470 123.710 109.760 123.755 ;
        RECT 111.330 123.710 111.620 123.755 ;
        RECT 87.830 123.415 90.365 123.555 ;
        RECT 92.460 123.555 92.780 123.615 ;
        RECT 92.935 123.555 93.225 123.600 ;
        RECT 92.460 123.415 93.225 123.555 ;
        RECT 87.830 123.370 88.120 123.415 ;
        RECT 92.460 123.355 92.780 123.415 ;
        RECT 92.935 123.370 93.225 123.415 ;
        RECT 94.760 123.355 95.080 123.615 ;
        RECT 97.520 123.555 97.840 123.615 ;
        RECT 97.995 123.555 98.285 123.600 ;
        RECT 95.310 123.415 98.285 123.555 ;
        RECT 72.695 123.075 80.270 123.215 ;
        RECT 80.515 123.215 80.805 123.260 ;
        RECT 91.095 123.215 91.385 123.260 ;
        RECT 91.540 123.215 91.860 123.275 ;
        RECT 80.515 123.075 87.170 123.215 ;
        RECT 72.695 123.030 72.985 123.075 ;
        RECT 79.120 123.015 79.440 123.075 ;
        RECT 80.515 123.030 80.805 123.075 ;
        RECT 48.760 122.875 49.080 122.935 ;
        RECT 44.250 122.735 49.080 122.875 ;
        RECT 39.070 122.690 39.360 122.735 ;
        RECT 41.850 122.690 42.140 122.735 ;
        RECT 43.710 122.690 44.000 122.735 ;
        RECT 48.760 122.675 49.080 122.735 ;
        RECT 62.120 122.875 62.410 122.920 ;
        RECT 63.980 122.875 64.270 122.920 ;
        RECT 66.760 122.875 67.050 122.920 ;
        RECT 62.120 122.735 67.050 122.875 ;
        RECT 72.310 122.875 72.450 123.015 ;
        RECT 80.590 122.875 80.730 123.030 ;
        RECT 72.310 122.735 80.730 122.875 ;
        RECT 62.120 122.690 62.410 122.735 ;
        RECT 63.980 122.690 64.270 122.735 ;
        RECT 66.760 122.690 67.050 122.735 ;
        RECT 29.900 122.535 30.220 122.595 ;
        RECT 25.850 122.395 30.220 122.535 ;
        RECT 29.900 122.335 30.220 122.395 ;
        RECT 31.740 122.535 32.060 122.595 ;
        RECT 46.460 122.535 46.780 122.595 ;
        RECT 31.740 122.395 46.780 122.535 ;
        RECT 31.740 122.335 32.060 122.395 ;
        RECT 46.460 122.335 46.780 122.395 ;
        RECT 50.615 122.535 50.905 122.580 ;
        RECT 51.980 122.535 52.300 122.595 ;
        RECT 50.615 122.395 52.300 122.535 ;
        RECT 50.615 122.350 50.905 122.395 ;
        RECT 51.980 122.335 52.300 122.395 ;
        RECT 54.280 122.335 54.600 122.595 ;
        RECT 74.995 122.535 75.285 122.580 ;
        RECT 76.360 122.535 76.680 122.595 ;
        RECT 74.995 122.395 76.680 122.535 ;
        RECT 74.995 122.350 75.285 122.395 ;
        RECT 76.360 122.335 76.680 122.395 ;
        RECT 83.275 122.535 83.565 122.580 ;
        RECT 86.480 122.535 86.800 122.595 ;
        RECT 83.275 122.395 86.800 122.535 ;
        RECT 87.030 122.535 87.170 123.075 ;
        RECT 91.095 123.075 91.860 123.215 ;
        RECT 91.095 123.030 91.385 123.075 ;
        RECT 91.540 123.015 91.860 123.075 ;
        RECT 92.000 123.215 92.320 123.275 ;
        RECT 95.310 123.215 95.450 123.415 ;
        RECT 97.520 123.355 97.840 123.415 ;
        RECT 97.995 123.370 98.285 123.415 ;
        RECT 101.200 123.355 101.520 123.615 ;
        RECT 107.150 123.555 107.440 123.600 ;
        RECT 109.470 123.555 109.685 123.710 ;
        RECT 107.150 123.415 109.685 123.555 ;
        RECT 107.150 123.370 107.440 123.415 ;
        RECT 110.400 123.355 110.720 123.615 ;
        RECT 112.255 123.555 112.545 123.600 ;
        RECT 114.080 123.555 114.400 123.615 ;
        RECT 112.255 123.415 114.400 123.555 ;
        RECT 112.255 123.370 112.545 123.415 ;
        RECT 114.080 123.355 114.400 123.415 ;
        RECT 92.000 123.075 95.450 123.215 ;
        RECT 97.075 123.215 97.365 123.260 ;
        RECT 98.440 123.215 98.760 123.275 ;
        RECT 97.075 123.075 98.760 123.215 ;
        RECT 92.000 123.015 92.320 123.075 ;
        RECT 97.075 123.030 97.365 123.075 ;
        RECT 87.830 122.875 88.120 122.920 ;
        RECT 90.610 122.875 90.900 122.920 ;
        RECT 92.470 122.875 92.760 122.920 ;
        RECT 97.150 122.875 97.290 123.030 ;
        RECT 98.440 123.015 98.760 123.075 ;
        RECT 87.830 122.735 92.760 122.875 ;
        RECT 87.830 122.690 88.120 122.735 ;
        RECT 90.610 122.690 90.900 122.735 ;
        RECT 92.470 122.690 92.760 122.735 ;
        RECT 93.010 122.735 97.290 122.875 ;
        RECT 107.150 122.875 107.440 122.920 ;
        RECT 109.930 122.875 110.220 122.920 ;
        RECT 111.790 122.875 112.080 122.920 ;
        RECT 107.150 122.735 112.080 122.875 ;
        RECT 93.010 122.535 93.150 122.735 ;
        RECT 107.150 122.690 107.440 122.735 ;
        RECT 109.930 122.690 110.220 122.735 ;
        RECT 111.790 122.690 112.080 122.735 ;
        RECT 87.030 122.395 93.150 122.535 ;
        RECT 83.275 122.350 83.565 122.395 ;
        RECT 86.480 122.335 86.800 122.395 ;
        RECT 95.220 122.335 95.540 122.595 ;
        RECT 99.820 122.335 100.140 122.595 ;
        RECT 14.650 121.715 115.850 122.195 ;
        RECT 33.120 121.515 33.440 121.575 ;
        RECT 34.055 121.515 34.345 121.560 ;
        RECT 47.380 121.515 47.700 121.575 ;
        RECT 33.120 121.375 34.345 121.515 ;
        RECT 33.120 121.315 33.440 121.375 ;
        RECT 34.055 121.330 34.345 121.375 ;
        RECT 37.810 121.375 47.700 121.515 ;
        RECT 23.940 121.175 24.230 121.220 ;
        RECT 25.800 121.175 26.090 121.220 ;
        RECT 28.580 121.175 28.870 121.220 ;
        RECT 23.940 121.035 28.870 121.175 ;
        RECT 23.940 120.990 24.230 121.035 ;
        RECT 25.800 120.990 26.090 121.035 ;
        RECT 28.580 120.990 28.870 121.035 ;
        RECT 25.315 120.835 25.605 120.880 ;
        RECT 27.140 120.835 27.460 120.895 ;
        RECT 25.315 120.695 27.460 120.835 ;
        RECT 25.315 120.650 25.605 120.695 ;
        RECT 27.140 120.635 27.460 120.695 ;
        RECT 29.900 120.835 30.220 120.895 ;
        RECT 37.275 120.835 37.565 120.880 ;
        RECT 37.810 120.835 37.950 121.375 ;
        RECT 47.380 121.315 47.700 121.375 ;
        RECT 49.220 121.515 49.540 121.575 ;
        RECT 50.845 121.515 51.135 121.560 ;
        RECT 49.220 121.375 51.135 121.515 ;
        RECT 49.220 121.315 49.540 121.375 ;
        RECT 50.845 121.330 51.135 121.375 ;
        RECT 64.875 121.515 65.165 121.560 ;
        RECT 65.320 121.515 65.640 121.575 ;
        RECT 64.875 121.375 65.640 121.515 ;
        RECT 64.875 121.330 65.165 121.375 ;
        RECT 65.320 121.315 65.640 121.375 ;
        RECT 66.025 121.515 66.315 121.560 ;
        RECT 69.460 121.515 69.780 121.575 ;
        RECT 66.025 121.375 69.780 121.515 ;
        RECT 66.025 121.330 66.315 121.375 ;
        RECT 69.460 121.315 69.780 121.375 ;
        RECT 77.065 121.515 77.355 121.560 ;
        RECT 79.120 121.515 79.440 121.575 ;
        RECT 77.065 121.375 79.440 121.515 ;
        RECT 77.065 121.330 77.355 121.375 ;
        RECT 79.120 121.315 79.440 121.375 ;
        RECT 91.540 121.315 91.860 121.575 ;
        RECT 92.000 121.560 92.320 121.575 ;
        RECT 92.000 121.330 92.535 121.560 ;
        RECT 94.760 121.515 95.080 121.575 ;
        RECT 103.960 121.515 104.280 121.575 ;
        RECT 94.760 121.375 104.280 121.515 ;
        RECT 92.000 121.315 92.320 121.330 ;
        RECT 94.760 121.315 95.080 121.375 ;
        RECT 103.960 121.315 104.280 121.375 ;
        RECT 106.260 121.315 106.580 121.575 ;
        RECT 45.050 121.175 45.340 121.220 ;
        RECT 47.830 121.175 48.120 121.220 ;
        RECT 49.690 121.175 49.980 121.220 ;
        RECT 45.050 121.035 49.980 121.175 ;
        RECT 45.050 120.990 45.340 121.035 ;
        RECT 47.830 120.990 48.120 121.035 ;
        RECT 49.690 120.990 49.980 121.035 ;
        RECT 54.710 121.175 55.000 121.220 ;
        RECT 57.490 121.175 57.780 121.220 ;
        RECT 59.350 121.175 59.640 121.220 ;
        RECT 54.710 121.035 59.640 121.175 ;
        RECT 54.710 120.990 55.000 121.035 ;
        RECT 57.490 120.990 57.780 121.035 ;
        RECT 59.350 120.990 59.640 121.035 ;
        RECT 69.890 121.175 70.180 121.220 ;
        RECT 72.670 121.175 72.960 121.220 ;
        RECT 74.530 121.175 74.820 121.220 ;
        RECT 69.890 121.035 74.820 121.175 ;
        RECT 69.890 120.990 70.180 121.035 ;
        RECT 72.670 120.990 72.960 121.035 ;
        RECT 74.530 120.990 74.820 121.035 ;
        RECT 75.455 120.990 75.745 121.220 ;
        RECT 80.930 121.175 81.220 121.220 ;
        RECT 83.710 121.175 84.000 121.220 ;
        RECT 85.570 121.175 85.860 121.220 ;
        RECT 80.930 121.035 85.860 121.175 ;
        RECT 80.930 120.990 81.220 121.035 ;
        RECT 83.710 120.990 84.000 121.035 ;
        RECT 85.570 120.990 85.860 121.035 ;
        RECT 91.080 121.175 91.400 121.235 ;
        RECT 94.850 121.175 94.990 121.315 ;
        RECT 91.080 121.035 94.990 121.175 ;
        RECT 96.110 121.175 96.400 121.220 ;
        RECT 98.890 121.175 99.180 121.220 ;
        RECT 100.750 121.175 101.040 121.220 ;
        RECT 96.110 121.035 101.040 121.175 ;
        RECT 29.900 120.695 37.950 120.835 ;
        RECT 38.180 120.835 38.500 120.895 ;
        RECT 38.655 120.835 38.945 120.880 ;
        RECT 42.780 120.835 43.100 120.895 ;
        RECT 38.180 120.695 38.945 120.835 ;
        RECT 29.900 120.635 30.220 120.695 ;
        RECT 37.275 120.650 37.565 120.695 ;
        RECT 38.180 120.635 38.500 120.695 ;
        RECT 38.655 120.650 38.945 120.695 ;
        RECT 39.650 120.695 43.100 120.835 ;
        RECT 23.475 120.495 23.765 120.540 ;
        RECT 24.840 120.495 25.160 120.555 ;
        RECT 28.580 120.495 28.870 120.540 ;
        RECT 23.475 120.355 25.160 120.495 ;
        RECT 23.475 120.310 23.765 120.355 ;
        RECT 24.840 120.295 25.160 120.355 ;
        RECT 26.335 120.355 28.870 120.495 ;
        RECT 26.335 120.200 26.550 120.355 ;
        RECT 28.580 120.310 28.870 120.355 ;
        RECT 31.740 120.495 32.060 120.555 ;
        RECT 32.445 120.495 32.735 120.540 ;
        RECT 31.740 120.355 32.735 120.495 ;
        RECT 31.740 120.295 32.060 120.355 ;
        RECT 32.445 120.310 32.735 120.355 ;
        RECT 36.355 120.495 36.645 120.540 ;
        RECT 38.270 120.495 38.410 120.635 ;
        RECT 39.650 120.540 39.790 120.695 ;
        RECT 42.780 120.635 43.100 120.695 ;
        RECT 50.230 120.695 57.730 120.835 ;
        RECT 36.355 120.355 38.410 120.495 ;
        RECT 36.355 120.310 36.645 120.355 ;
        RECT 39.575 120.310 39.865 120.540 ;
        RECT 40.020 120.495 40.340 120.555 ;
        RECT 40.495 120.495 40.785 120.540 ;
        RECT 40.020 120.355 40.785 120.495 ;
        RECT 40.020 120.295 40.340 120.355 ;
        RECT 40.495 120.310 40.785 120.355 ;
        RECT 41.185 120.495 41.475 120.540 ;
        RECT 43.700 120.495 44.020 120.555 ;
        RECT 41.185 120.355 44.020 120.495 ;
        RECT 41.185 120.310 41.475 120.355 ;
        RECT 43.700 120.295 44.020 120.355 ;
        RECT 45.050 120.495 45.340 120.540 ;
        RECT 45.050 120.355 47.585 120.495 ;
        RECT 45.050 120.310 45.340 120.355 ;
        RECT 24.400 120.155 24.690 120.200 ;
        RECT 26.260 120.155 26.550 120.200 ;
        RECT 24.400 120.015 26.550 120.155 ;
        RECT 24.400 119.970 24.690 120.015 ;
        RECT 26.260 119.970 26.550 120.015 ;
        RECT 27.140 120.200 27.460 120.215 ;
        RECT 27.140 120.155 27.470 120.200 ;
        RECT 30.440 120.155 30.730 120.200 ;
        RECT 27.140 120.015 30.730 120.155 ;
        RECT 27.140 119.970 27.470 120.015 ;
        RECT 30.440 119.970 30.730 120.015 ;
        RECT 35.895 120.155 36.185 120.200 ;
        RECT 37.260 120.155 37.580 120.215 ;
        RECT 35.895 120.015 37.580 120.155 ;
        RECT 35.895 119.970 36.185 120.015 ;
        RECT 27.140 119.955 27.460 119.970 ;
        RECT 37.260 119.955 37.580 120.015 ;
        RECT 43.190 120.155 43.480 120.200 ;
        RECT 44.620 120.155 44.940 120.215 ;
        RECT 47.370 120.200 47.585 120.355 ;
        RECT 48.300 120.295 48.620 120.555 ;
        RECT 48.760 120.495 49.080 120.555 ;
        RECT 50.230 120.540 50.370 120.695 ;
        RECT 50.155 120.495 50.445 120.540 ;
        RECT 48.760 120.355 50.445 120.495 ;
        RECT 48.760 120.295 49.080 120.355 ;
        RECT 50.155 120.310 50.445 120.355 ;
        RECT 54.710 120.495 55.000 120.540 ;
        RECT 57.590 120.495 57.730 120.695 ;
        RECT 57.960 120.635 58.280 120.895 ;
        RECT 59.815 120.835 60.105 120.880 ;
        RECT 60.260 120.835 60.580 120.895 ;
        RECT 75.530 120.835 75.670 120.990 ;
        RECT 91.080 120.975 91.400 121.035 ;
        RECT 96.110 120.990 96.400 121.035 ;
        RECT 98.890 120.990 99.180 121.035 ;
        RECT 100.750 120.990 101.040 121.035 ;
        RECT 81.880 120.835 82.200 120.895 ;
        RECT 84.640 120.835 84.960 120.895 ;
        RECT 86.035 120.835 86.325 120.880 ;
        RECT 59.200 120.695 60.580 120.835 ;
        RECT 59.200 120.495 59.340 120.695 ;
        RECT 59.815 120.650 60.105 120.695 ;
        RECT 60.260 120.635 60.580 120.695 ;
        RECT 74.610 120.695 75.670 120.835 ;
        RECT 80.590 120.695 86.325 120.835 ;
        RECT 54.710 120.355 57.245 120.495 ;
        RECT 57.590 120.355 59.340 120.495 ;
        RECT 62.560 120.495 62.880 120.555 ;
        RECT 64.415 120.495 64.705 120.540 ;
        RECT 62.560 120.355 64.705 120.495 ;
        RECT 54.710 120.310 55.000 120.355 ;
        RECT 46.450 120.155 46.740 120.200 ;
        RECT 43.190 120.015 46.740 120.155 ;
        RECT 43.190 119.970 43.480 120.015 ;
        RECT 44.620 119.955 44.940 120.015 ;
        RECT 46.450 119.970 46.740 120.015 ;
        RECT 47.370 120.155 47.660 120.200 ;
        RECT 49.230 120.155 49.520 120.200 ;
        RECT 47.370 120.015 49.520 120.155 ;
        RECT 47.370 119.970 47.660 120.015 ;
        RECT 49.230 119.970 49.520 120.015 ;
        RECT 52.850 120.155 53.140 120.200 ;
        RECT 54.280 120.155 54.600 120.215 ;
        RECT 57.030 120.200 57.245 120.355 ;
        RECT 62.560 120.295 62.880 120.355 ;
        RECT 64.415 120.310 64.705 120.355 ;
        RECT 69.890 120.495 70.180 120.540 ;
        RECT 73.155 120.495 73.445 120.540 ;
        RECT 74.610 120.495 74.750 120.695 ;
        RECT 69.890 120.355 72.425 120.495 ;
        RECT 69.890 120.310 70.180 120.355 ;
        RECT 56.110 120.155 56.400 120.200 ;
        RECT 52.850 120.015 56.400 120.155 ;
        RECT 52.850 119.970 53.140 120.015 ;
        RECT 54.280 119.955 54.600 120.015 ;
        RECT 56.110 119.970 56.400 120.015 ;
        RECT 57.030 120.155 57.320 120.200 ;
        RECT 58.890 120.155 59.180 120.200 ;
        RECT 57.030 120.015 59.180 120.155 ;
        RECT 57.030 119.970 57.320 120.015 ;
        RECT 58.890 119.970 59.180 120.015 ;
        RECT 68.030 120.155 68.320 120.200 ;
        RECT 69.460 120.155 69.780 120.215 ;
        RECT 72.210 120.200 72.425 120.355 ;
        RECT 73.155 120.355 74.750 120.495 ;
        RECT 73.155 120.310 73.445 120.355 ;
        RECT 74.995 120.310 75.285 120.540 ;
        RECT 71.290 120.155 71.580 120.200 ;
        RECT 68.030 120.015 71.580 120.155 ;
        RECT 68.030 119.970 68.320 120.015 ;
        RECT 69.460 119.955 69.780 120.015 ;
        RECT 71.290 119.970 71.580 120.015 ;
        RECT 72.210 120.155 72.500 120.200 ;
        RECT 74.070 120.155 74.360 120.200 ;
        RECT 72.210 120.015 74.360 120.155 ;
        RECT 75.070 120.155 75.210 120.310 ;
        RECT 76.360 120.295 76.680 120.555 ;
        RECT 80.590 120.495 80.730 120.695 ;
        RECT 81.880 120.635 82.200 120.695 ;
        RECT 84.640 120.635 84.960 120.695 ;
        RECT 86.035 120.650 86.325 120.695 ;
        RECT 86.480 120.835 86.800 120.895 ;
        RECT 86.480 120.695 87.170 120.835 ;
        RECT 86.480 120.635 86.800 120.695 ;
        RECT 76.910 120.355 80.730 120.495 ;
        RECT 80.930 120.495 81.220 120.540 ;
        RECT 84.195 120.495 84.485 120.540 ;
        RECT 87.030 120.495 87.170 120.695 ;
        RECT 87.415 120.495 87.705 120.540 ;
        RECT 80.930 120.355 83.465 120.495 ;
        RECT 76.910 120.155 77.050 120.355 ;
        RECT 80.930 120.310 81.220 120.355 ;
        RECT 75.070 120.015 77.050 120.155 ;
        RECT 79.070 120.155 79.360 120.200 ;
        RECT 81.420 120.155 81.740 120.215 ;
        RECT 83.250 120.200 83.465 120.355 ;
        RECT 84.195 120.355 86.710 120.495 ;
        RECT 87.030 120.355 87.705 120.495 ;
        RECT 84.195 120.310 84.485 120.355 ;
        RECT 82.330 120.155 82.620 120.200 ;
        RECT 79.070 120.015 82.620 120.155 ;
        RECT 72.210 119.970 72.500 120.015 ;
        RECT 74.070 119.970 74.360 120.015 ;
        RECT 79.070 119.970 79.360 120.015 ;
        RECT 81.420 119.955 81.740 120.015 ;
        RECT 82.330 119.970 82.620 120.015 ;
        RECT 83.250 120.155 83.540 120.200 ;
        RECT 85.110 120.155 85.400 120.200 ;
        RECT 83.250 120.015 85.400 120.155 ;
        RECT 83.250 119.970 83.540 120.015 ;
        RECT 85.110 119.970 85.400 120.015 ;
        RECT 86.570 119.860 86.710 120.355 ;
        RECT 87.415 120.310 87.705 120.355 ;
        RECT 90.620 120.295 90.940 120.555 ;
        RECT 96.110 120.495 96.400 120.540 ;
        RECT 96.110 120.355 98.645 120.495 ;
        RECT 96.110 120.310 96.400 120.355 ;
        RECT 94.250 120.155 94.540 120.200 ;
        RECT 95.220 120.155 95.540 120.215 ;
        RECT 98.430 120.200 98.645 120.355 ;
        RECT 99.360 120.295 99.680 120.555 ;
        RECT 101.215 120.310 101.505 120.540 ;
        RECT 103.960 120.495 104.280 120.555 ;
        RECT 105.815 120.495 106.105 120.540 ;
        RECT 103.960 120.355 106.105 120.495 ;
        RECT 97.510 120.155 97.800 120.200 ;
        RECT 94.250 120.015 97.800 120.155 ;
        RECT 94.250 119.970 94.540 120.015 ;
        RECT 95.220 119.955 95.540 120.015 ;
        RECT 97.510 119.970 97.800 120.015 ;
        RECT 98.430 120.155 98.720 120.200 ;
        RECT 100.290 120.155 100.580 120.200 ;
        RECT 98.430 120.015 100.580 120.155 ;
        RECT 101.290 120.155 101.430 120.310 ;
        RECT 103.960 120.295 104.280 120.355 ;
        RECT 105.815 120.310 106.105 120.355 ;
        RECT 109.020 120.155 109.340 120.215 ;
        RECT 101.290 120.015 109.340 120.155 ;
        RECT 98.430 119.970 98.720 120.015 ;
        RECT 100.290 119.970 100.580 120.015 ;
        RECT 109.020 119.955 109.340 120.015 ;
        RECT 86.495 119.630 86.785 119.860 ;
        RECT 14.650 118.995 115.850 119.475 ;
        RECT 32.200 118.795 32.520 118.855 ;
        RECT 32.675 118.795 32.965 118.840 ;
        RECT 32.200 118.655 32.965 118.795 ;
        RECT 32.200 118.595 32.520 118.655 ;
        RECT 32.675 118.610 32.965 118.655 ;
        RECT 38.640 118.595 38.960 118.855 ;
        RECT 40.480 118.595 40.800 118.855 ;
        RECT 44.620 118.595 44.940 118.855 ;
        RECT 46.475 118.795 46.765 118.840 ;
        RECT 48.300 118.795 48.620 118.855 ;
        RECT 46.475 118.655 48.620 118.795 ;
        RECT 46.475 118.610 46.765 118.655 ;
        RECT 48.300 118.595 48.620 118.655 ;
        RECT 49.220 118.595 49.540 118.855 ;
        RECT 56.595 118.795 56.885 118.840 ;
        RECT 57.960 118.795 58.280 118.855 ;
        RECT 56.595 118.655 58.280 118.795 ;
        RECT 56.595 118.610 56.885 118.655 ;
        RECT 57.960 118.595 58.280 118.655 ;
        RECT 63.480 118.795 63.800 118.855 ;
        RECT 67.635 118.795 67.925 118.840 ;
        RECT 63.480 118.655 67.925 118.795 ;
        RECT 63.480 118.595 63.800 118.655 ;
        RECT 67.635 118.610 67.925 118.655 ;
        RECT 69.460 118.595 69.780 118.855 ;
        RECT 80.975 118.795 81.265 118.840 ;
        RECT 81.420 118.795 81.740 118.855 ;
        RECT 80.975 118.655 81.740 118.795 ;
        RECT 80.975 118.610 81.265 118.655 ;
        RECT 81.420 118.595 81.740 118.655 ;
        RECT 84.195 118.795 84.485 118.840 ;
        RECT 86.020 118.795 86.340 118.855 ;
        RECT 84.195 118.655 86.340 118.795 ;
        RECT 84.195 118.610 84.485 118.655 ;
        RECT 86.020 118.595 86.340 118.655 ;
        RECT 98.915 118.795 99.205 118.840 ;
        RECT 99.360 118.795 99.680 118.855 ;
        RECT 98.915 118.655 99.680 118.795 ;
        RECT 98.915 118.610 99.205 118.655 ;
        RECT 99.360 118.595 99.680 118.655 ;
        RECT 105.800 118.795 106.120 118.855 ;
        RECT 109.495 118.795 109.785 118.840 ;
        RECT 105.800 118.655 109.785 118.795 ;
        RECT 105.800 118.595 106.120 118.655 ;
        RECT 109.495 118.610 109.785 118.655 ;
        RECT 43.700 118.455 44.020 118.515 ;
        RECT 48.775 118.455 49.065 118.500 ;
        RECT 43.700 118.315 49.065 118.455 ;
        RECT 43.700 118.255 44.020 118.315 ;
        RECT 48.775 118.270 49.065 118.315 ;
        RECT 62.560 118.455 62.880 118.515 ;
        RECT 78.200 118.455 78.520 118.515 ;
        RECT 62.560 118.315 78.520 118.455 ;
        RECT 62.560 118.255 62.880 118.315 ;
        RECT 28.980 118.115 29.300 118.175 ;
        RECT 33.135 118.115 33.425 118.160 ;
        RECT 38.195 118.115 38.485 118.160 ;
        RECT 28.980 117.975 38.485 118.115 ;
        RECT 28.980 117.915 29.300 117.975 ;
        RECT 33.135 117.930 33.425 117.975 ;
        RECT 38.195 117.930 38.485 117.975 ;
        RECT 38.270 117.775 38.410 117.930 ;
        RECT 39.560 117.915 39.880 118.175 ;
        RECT 44.175 118.115 44.465 118.160 ;
        RECT 45.080 118.115 45.400 118.175 ;
        RECT 44.175 117.975 45.400 118.115 ;
        RECT 44.175 117.930 44.465 117.975 ;
        RECT 44.250 117.775 44.390 117.930 ;
        RECT 45.080 117.915 45.400 117.975 ;
        RECT 45.555 118.115 45.845 118.160 ;
        RECT 51.980 118.115 52.300 118.175 ;
        RECT 55.675 118.115 55.965 118.160 ;
        RECT 45.555 117.975 47.150 118.115 ;
        RECT 45.555 117.930 45.845 117.975 ;
        RECT 38.270 117.635 44.390 117.775 ;
        RECT 47.010 117.480 47.150 117.975 ;
        RECT 51.980 117.975 55.965 118.115 ;
        RECT 51.980 117.915 52.300 117.975 ;
        RECT 55.675 117.930 55.965 117.975 ;
        RECT 68.540 117.915 68.860 118.175 ;
        RECT 69.090 118.160 69.230 118.315 ;
        RECT 78.200 118.255 78.520 118.315 ;
        RECT 107.640 118.455 107.960 118.515 ;
        RECT 107.640 118.315 112.010 118.455 ;
        RECT 107.640 118.255 107.960 118.315 ;
        RECT 69.015 117.930 69.305 118.160 ;
        RECT 78.290 118.115 78.430 118.255 ;
        RECT 81.435 118.115 81.725 118.160 ;
        RECT 83.735 118.115 84.025 118.160 ;
        RECT 78.290 117.975 84.025 118.115 ;
        RECT 81.435 117.930 81.725 117.975 ;
        RECT 83.735 117.930 84.025 117.975 ;
        RECT 99.820 117.915 100.140 118.175 ;
        RECT 108.100 117.915 108.420 118.175 ;
        RECT 108.560 118.115 108.880 118.175 ;
        RECT 111.870 118.160 112.010 118.315 ;
        RECT 110.415 118.115 110.705 118.160 ;
        RECT 108.560 117.975 110.705 118.115 ;
        RECT 108.560 117.915 108.880 117.975 ;
        RECT 110.415 117.930 110.705 117.975 ;
        RECT 111.795 117.930 112.085 118.160 ;
        RECT 114.080 117.915 114.400 118.175 ;
        RECT 47.840 117.775 48.160 117.835 ;
        RECT 49.695 117.775 49.985 117.820 ;
        RECT 47.840 117.635 49.985 117.775 ;
        RECT 47.840 117.575 48.160 117.635 ;
        RECT 49.695 117.590 49.985 117.635 ;
        RECT 72.220 117.775 72.540 117.835 ;
        RECT 72.220 117.635 113.390 117.775 ;
        RECT 72.220 117.575 72.540 117.635 ;
        RECT 46.935 117.250 47.225 117.480 ;
        RECT 105.340 117.435 105.660 117.495 ;
        RECT 113.250 117.480 113.390 117.635 ;
        RECT 110.875 117.435 111.165 117.480 ;
        RECT 105.340 117.295 111.165 117.435 ;
        RECT 105.340 117.235 105.660 117.295 ;
        RECT 110.875 117.250 111.165 117.295 ;
        RECT 113.175 117.250 113.465 117.480 ;
        RECT 108.560 116.895 108.880 117.155 ;
        RECT 14.650 116.275 115.850 116.755 ;
        RECT 24.840 116.075 25.160 116.135 ;
        RECT 67.160 116.075 67.480 116.135 ;
        RECT 71.775 116.075 72.065 116.120 ;
        RECT 109.020 116.075 109.340 116.135 ;
        RECT 24.840 115.935 26.910 116.075 ;
        RECT 24.840 115.875 25.160 115.935 ;
        RECT 21.275 115.735 21.565 115.780 ;
        RECT 24.395 115.735 24.685 115.780 ;
        RECT 26.285 115.735 26.575 115.780 ;
        RECT 21.275 115.595 26.575 115.735 ;
        RECT 21.275 115.550 21.565 115.595 ;
        RECT 24.395 115.550 24.685 115.595 ;
        RECT 26.285 115.550 26.575 115.595 ;
        RECT 26.770 115.395 26.910 115.935 ;
        RECT 67.160 115.935 72.065 116.075 ;
        RECT 67.160 115.875 67.480 115.935 ;
        RECT 71.775 115.890 72.065 115.935 ;
        RECT 104.050 115.935 109.340 116.075 ;
        RECT 72.680 115.735 73.000 115.795 ;
        RECT 99.835 115.735 100.125 115.780 ;
        RECT 101.660 115.735 101.980 115.795 ;
        RECT 72.680 115.595 86.710 115.735 ;
        RECT 72.680 115.535 73.000 115.595 ;
        RECT 27.140 115.395 27.460 115.455 ;
        RECT 26.770 115.255 27.460 115.395 ;
        RECT 27.140 115.195 27.460 115.255 ;
        RECT 58.420 115.195 58.740 115.455 ;
        RECT 66.330 115.255 73.830 115.395 ;
        RECT 17.035 114.715 17.325 114.760 ;
        RECT 17.940 114.715 18.260 114.775 ;
        RECT 20.195 114.760 20.485 115.075 ;
        RECT 21.275 115.055 21.565 115.100 ;
        RECT 24.855 115.055 25.145 115.100 ;
        RECT 26.690 115.055 26.980 115.100 ;
        RECT 21.275 114.915 26.980 115.055 ;
        RECT 21.275 114.870 21.565 114.915 ;
        RECT 24.855 114.870 25.145 114.915 ;
        RECT 26.690 114.870 26.980 114.915 ;
        RECT 28.060 114.855 28.380 115.115 ;
        RECT 29.440 115.055 29.760 115.115 ;
        RECT 30.375 115.055 30.665 115.100 ;
        RECT 29.440 114.915 30.665 115.055 ;
        RECT 29.440 114.855 29.760 114.915 ;
        RECT 30.375 114.870 30.665 114.915 ;
        RECT 31.280 115.055 31.600 115.115 ;
        RECT 32.215 115.055 32.505 115.100 ;
        RECT 31.280 114.915 32.505 115.055 ;
        RECT 31.280 114.855 31.600 114.915 ;
        RECT 32.215 114.870 32.505 114.915 ;
        RECT 32.660 115.055 32.980 115.115 ;
        RECT 33.135 115.055 33.425 115.100 ;
        RECT 32.660 114.915 33.425 115.055 ;
        RECT 32.660 114.855 32.980 114.915 ;
        RECT 33.135 114.870 33.425 114.915 ;
        RECT 44.160 115.055 44.480 115.115 ;
        RECT 47.395 115.055 47.685 115.100 ;
        RECT 44.160 114.915 47.685 115.055 ;
        RECT 44.160 114.855 44.480 114.915 ;
        RECT 47.395 114.870 47.685 114.915 ;
        RECT 57.515 115.055 57.805 115.100 ;
        RECT 58.880 115.055 59.200 115.115 ;
        RECT 66.330 115.055 66.470 115.255 ;
        RECT 57.515 114.915 66.470 115.055 ;
        RECT 57.515 114.870 57.805 114.915 ;
        RECT 58.880 114.855 59.200 114.915 ;
        RECT 69.475 114.870 69.765 115.100 ;
        RECT 17.035 114.575 18.260 114.715 ;
        RECT 17.035 114.530 17.325 114.575 ;
        RECT 17.940 114.515 18.260 114.575 ;
        RECT 19.895 114.715 20.485 114.760 ;
        RECT 22.080 114.715 22.400 114.775 ;
        RECT 23.135 114.715 23.785 114.760 ;
        RECT 19.895 114.575 23.785 114.715 ;
        RECT 19.895 114.530 20.185 114.575 ;
        RECT 22.080 114.515 22.400 114.575 ;
        RECT 23.135 114.530 23.785 114.575 ;
        RECT 25.775 114.530 26.065 114.760 ;
        RECT 25.850 114.375 25.990 114.530 ;
        RECT 28.520 114.515 28.840 114.775 ;
        RECT 69.550 114.715 69.690 114.870 ;
        RECT 69.920 114.855 70.240 115.115 ;
        RECT 72.220 114.855 72.540 115.115 ;
        RECT 73.690 115.100 73.830 115.255 ;
        RECT 86.570 115.100 86.710 115.595 ;
        RECT 99.835 115.595 101.980 115.735 ;
        RECT 99.835 115.550 100.125 115.595 ;
        RECT 101.660 115.535 101.980 115.595 ;
        RECT 92.920 115.395 93.240 115.455 ;
        RECT 103.040 115.395 103.360 115.455 ;
        RECT 104.050 115.440 104.190 115.935 ;
        RECT 109.020 115.875 109.340 115.935 ;
        RECT 104.845 115.735 105.135 115.780 ;
        RECT 106.735 115.735 107.025 115.780 ;
        RECT 109.855 115.735 110.145 115.780 ;
        RECT 104.845 115.595 110.145 115.735 ;
        RECT 104.845 115.550 105.135 115.595 ;
        RECT 106.735 115.550 107.025 115.595 ;
        RECT 109.855 115.550 110.145 115.595 ;
        RECT 103.975 115.395 104.265 115.440 ;
        RECT 92.920 115.255 100.510 115.395 ;
        RECT 92.920 115.195 93.240 115.255 ;
        RECT 73.615 114.870 73.905 115.100 ;
        RECT 86.495 114.870 86.785 115.100 ;
        RECT 86.940 115.055 87.260 115.115 ;
        RECT 92.015 115.055 92.305 115.100 ;
        RECT 86.940 114.915 92.305 115.055 ;
        RECT 86.940 114.855 87.260 114.915 ;
        RECT 92.015 114.870 92.305 114.915 ;
        RECT 93.380 115.055 93.700 115.115 ;
        RECT 97.075 115.055 97.365 115.100 ;
        RECT 93.380 114.915 97.365 115.055 ;
        RECT 93.380 114.855 93.700 114.915 ;
        RECT 97.075 114.870 97.365 114.915 ;
        RECT 98.900 114.855 99.220 115.115 ;
        RECT 100.370 115.100 100.510 115.255 ;
        RECT 103.040 115.255 104.265 115.395 ;
        RECT 103.040 115.195 103.360 115.255 ;
        RECT 103.975 115.210 104.265 115.255 ;
        RECT 105.340 115.195 105.660 115.455 ;
        RECT 100.295 114.870 100.585 115.100 ;
        RECT 104.440 115.055 104.730 115.100 ;
        RECT 106.275 115.055 106.565 115.100 ;
        RECT 109.855 115.055 110.145 115.100 ;
        RECT 104.440 114.915 110.145 115.055 ;
        RECT 104.440 114.870 104.730 114.915 ;
        RECT 106.275 114.870 106.565 114.915 ;
        RECT 109.855 114.870 110.145 114.915 ;
        RECT 74.995 114.715 75.285 114.760 ;
        RECT 78.200 114.715 78.520 114.775 ;
        RECT 69.550 114.575 78.520 114.715 ;
        RECT 74.995 114.530 75.285 114.575 ;
        RECT 78.200 114.515 78.520 114.575 ;
        RECT 107.635 114.715 108.285 114.760 ;
        RECT 108.560 114.715 108.880 114.775 ;
        RECT 110.935 114.760 111.225 115.075 ;
        RECT 110.935 114.715 111.525 114.760 ;
        RECT 107.635 114.575 111.525 114.715 ;
        RECT 107.635 114.530 108.285 114.575 ;
        RECT 108.560 114.515 108.880 114.575 ;
        RECT 111.235 114.530 111.525 114.575 ;
        RECT 114.095 114.715 114.385 114.760 ;
        RECT 117.300 114.715 117.620 114.775 ;
        RECT 114.095 114.575 117.620 114.715 ;
        RECT 114.095 114.530 114.385 114.575 ;
        RECT 117.300 114.515 117.620 114.575 ;
        RECT 29.455 114.375 29.745 114.420 ;
        RECT 25.850 114.235 29.745 114.375 ;
        RECT 29.455 114.190 29.745 114.235 ;
        RECT 29.900 114.375 30.220 114.435 ;
        RECT 31.295 114.375 31.585 114.420 ;
        RECT 29.900 114.235 31.585 114.375 ;
        RECT 29.900 114.175 30.220 114.235 ;
        RECT 31.295 114.190 31.585 114.235 ;
        RECT 34.055 114.375 34.345 114.420 ;
        RECT 34.500 114.375 34.820 114.435 ;
        RECT 34.055 114.235 34.820 114.375 ;
        RECT 34.055 114.190 34.345 114.235 ;
        RECT 34.500 114.175 34.820 114.235 ;
        RECT 48.315 114.375 48.605 114.420 ;
        RECT 49.220 114.375 49.540 114.435 ;
        RECT 48.315 114.235 49.540 114.375 ;
        RECT 48.315 114.190 48.605 114.235 ;
        RECT 49.220 114.175 49.540 114.235 ;
        RECT 69.000 114.175 69.320 114.435 ;
        RECT 70.840 114.175 71.160 114.435 ;
        RECT 87.415 114.375 87.705 114.420 ;
        RECT 89.700 114.375 90.020 114.435 ;
        RECT 87.415 114.235 90.020 114.375 ;
        RECT 87.415 114.190 87.705 114.235 ;
        RECT 89.700 114.175 90.020 114.235 ;
        RECT 92.920 114.175 93.240 114.435 ;
        RECT 97.995 114.375 98.285 114.420 ;
        RECT 100.280 114.375 100.600 114.435 ;
        RECT 97.995 114.235 100.600 114.375 ;
        RECT 97.995 114.190 98.285 114.235 ;
        RECT 100.280 114.175 100.600 114.235 ;
        RECT 101.215 114.375 101.505 114.420 ;
        RECT 104.420 114.375 104.740 114.435 ;
        RECT 101.215 114.235 104.740 114.375 ;
        RECT 101.215 114.190 101.505 114.235 ;
        RECT 104.420 114.175 104.740 114.235 ;
        RECT 14.650 113.555 115.850 114.035 ;
        RECT 21.635 113.355 21.925 113.400 ;
        RECT 22.080 113.355 22.400 113.415 ;
        RECT 21.635 113.215 22.400 113.355 ;
        RECT 21.635 113.170 21.925 113.215 ;
        RECT 22.080 113.155 22.400 113.215 ;
        RECT 62.100 113.355 62.420 113.415 ;
        RECT 70.840 113.355 71.160 113.415 ;
        RECT 62.100 113.215 64.630 113.355 ;
        RECT 62.100 113.155 62.420 113.215 ;
        RECT 28.060 113.015 28.380 113.075 ;
        RECT 23.550 112.875 28.380 113.015 ;
        RECT 23.550 112.720 23.690 112.875 ;
        RECT 28.060 112.815 28.380 112.875 ;
        RECT 28.520 113.015 28.840 113.075 ;
        RECT 29.095 113.015 29.385 113.060 ;
        RECT 32.335 113.015 32.985 113.060 ;
        RECT 28.520 112.875 32.985 113.015 ;
        RECT 28.520 112.815 28.840 112.875 ;
        RECT 29.095 112.830 29.685 112.875 ;
        RECT 32.335 112.830 32.985 112.875 ;
        RECT 34.500 113.015 34.820 113.075 ;
        RECT 34.975 113.015 35.265 113.060 ;
        RECT 34.500 112.875 35.265 113.015 ;
        RECT 20.715 112.675 21.005 112.720 ;
        RECT 22.095 112.675 22.385 112.720 ;
        RECT 23.475 112.675 23.765 112.720 ;
        RECT 20.715 112.535 23.765 112.675 ;
        RECT 20.715 112.490 21.005 112.535 ;
        RECT 22.095 112.490 22.385 112.535 ;
        RECT 23.475 112.490 23.765 112.535 ;
        RECT 23.935 112.675 24.225 112.720 ;
        RECT 24.380 112.675 24.700 112.735 ;
        RECT 23.935 112.535 24.700 112.675 ;
        RECT 23.935 112.490 24.225 112.535 ;
        RECT 24.380 112.475 24.700 112.535 ;
        RECT 29.395 112.515 29.685 112.830 ;
        RECT 34.500 112.815 34.820 112.875 ;
        RECT 34.975 112.830 35.265 112.875 ;
        RECT 37.720 113.015 38.040 113.075 ;
        RECT 46.920 113.060 47.240 113.075 ;
        RECT 43.355 113.015 43.645 113.060 ;
        RECT 46.595 113.015 47.245 113.060 ;
        RECT 37.720 112.875 39.330 113.015 ;
        RECT 37.720 112.815 38.040 112.875 ;
        RECT 30.475 112.675 30.765 112.720 ;
        RECT 34.055 112.675 34.345 112.720 ;
        RECT 35.890 112.675 36.180 112.720 ;
        RECT 30.475 112.535 36.180 112.675 ;
        RECT 30.475 112.490 30.765 112.535 ;
        RECT 34.055 112.490 34.345 112.535 ;
        RECT 35.890 112.490 36.180 112.535 ;
        RECT 38.640 112.475 38.960 112.735 ;
        RECT 39.190 112.720 39.330 112.875 ;
        RECT 43.355 112.875 47.245 113.015 ;
        RECT 43.355 112.830 43.945 112.875 ;
        RECT 46.595 112.830 47.245 112.875 ;
        RECT 39.115 112.490 39.405 112.720 ;
        RECT 43.655 112.515 43.945 112.830 ;
        RECT 46.920 112.815 47.240 112.830 ;
        RECT 49.220 112.815 49.540 113.075 ;
        RECT 56.695 113.015 56.985 113.060 ;
        RECT 58.880 113.015 59.200 113.075 ;
        RECT 59.935 113.015 60.585 113.060 ;
        RECT 56.695 112.875 60.585 113.015 ;
        RECT 56.695 112.830 57.285 112.875 ;
        RECT 44.735 112.675 45.025 112.720 ;
        RECT 48.315 112.675 48.605 112.720 ;
        RECT 50.150 112.675 50.440 112.720 ;
        RECT 44.735 112.535 50.440 112.675 ;
        RECT 44.735 112.490 45.025 112.535 ;
        RECT 48.315 112.490 48.605 112.535 ;
        RECT 50.150 112.490 50.440 112.535 ;
        RECT 52.440 112.475 52.760 112.735 ;
        RECT 56.995 112.515 57.285 112.830 ;
        RECT 58.880 112.815 59.200 112.875 ;
        RECT 59.935 112.830 60.585 112.875 ;
        RECT 61.180 113.015 61.500 113.075 ;
        RECT 62.575 113.015 62.865 113.060 ;
        RECT 61.180 112.875 62.865 113.015 ;
        RECT 61.180 112.815 61.500 112.875 ;
        RECT 62.575 112.830 62.865 112.875 ;
        RECT 64.490 112.720 64.630 113.215 ;
        RECT 70.840 113.215 74.750 113.355 ;
        RECT 70.840 113.155 71.160 113.215 ;
        RECT 74.610 113.060 74.750 113.215 ;
        RECT 68.655 113.015 68.945 113.060 ;
        RECT 71.895 113.015 72.545 113.060 ;
        RECT 68.655 112.875 72.545 113.015 ;
        RECT 68.655 112.830 69.245 112.875 ;
        RECT 71.895 112.830 72.545 112.875 ;
        RECT 74.535 112.830 74.825 113.060 ;
        RECT 74.980 113.015 75.300 113.075 ;
        RECT 81.880 113.015 82.200 113.075 ;
        RECT 86.940 113.060 87.260 113.075 ;
        RECT 74.980 112.875 78.430 113.015 ;
        RECT 68.955 112.735 69.245 112.830 ;
        RECT 74.980 112.815 75.300 112.875 ;
        RECT 58.075 112.675 58.365 112.720 ;
        RECT 61.655 112.675 61.945 112.720 ;
        RECT 63.490 112.675 63.780 112.720 ;
        RECT 58.075 112.535 63.780 112.675 ;
        RECT 58.075 112.490 58.365 112.535 ;
        RECT 61.655 112.490 61.945 112.535 ;
        RECT 63.490 112.490 63.780 112.535 ;
        RECT 64.415 112.490 64.705 112.720 ;
        RECT 68.955 112.515 69.320 112.735 ;
        RECT 78.290 112.720 78.430 112.875 ;
        RECT 79.210 112.875 82.200 113.015 ;
        RECT 69.000 112.475 69.320 112.515 ;
        RECT 70.035 112.675 70.325 112.720 ;
        RECT 73.615 112.675 73.905 112.720 ;
        RECT 75.450 112.675 75.740 112.720 ;
        RECT 70.035 112.535 75.740 112.675 ;
        RECT 70.035 112.490 70.325 112.535 ;
        RECT 73.615 112.490 73.905 112.535 ;
        RECT 75.450 112.490 75.740 112.535 ;
        RECT 78.215 112.490 78.505 112.720 ;
        RECT 26.235 112.150 26.525 112.380 ;
        RECT 27.140 112.335 27.460 112.395 ;
        RECT 36.355 112.335 36.645 112.380 ;
        RECT 37.720 112.335 38.040 112.395 ;
        RECT 27.140 112.195 38.040 112.335 ;
        RECT 26.310 111.995 26.450 112.150 ;
        RECT 27.140 112.135 27.460 112.195 ;
        RECT 36.355 112.150 36.645 112.195 ;
        RECT 37.720 112.135 38.040 112.195 ;
        RECT 40.495 112.335 40.785 112.380 ;
        RECT 45.540 112.335 45.860 112.395 ;
        RECT 40.495 112.195 45.860 112.335 ;
        RECT 40.495 112.150 40.785 112.195 ;
        RECT 45.540 112.135 45.860 112.195 ;
        RECT 48.760 112.335 49.080 112.395 ;
        RECT 50.615 112.335 50.905 112.380 ;
        RECT 48.760 112.195 50.905 112.335 ;
        RECT 48.760 112.135 49.080 112.195 ;
        RECT 50.615 112.150 50.905 112.195 ;
        RECT 53.835 112.335 54.125 112.380 ;
        RECT 56.580 112.335 56.900 112.395 ;
        RECT 53.835 112.195 56.900 112.335 ;
        RECT 53.835 112.150 54.125 112.195 ;
        RECT 56.580 112.135 56.900 112.195 ;
        RECT 60.260 112.335 60.580 112.395 ;
        RECT 63.955 112.335 64.245 112.380 ;
        RECT 60.260 112.195 64.245 112.335 ;
        RECT 60.260 112.135 60.580 112.195 ;
        RECT 63.955 112.150 64.245 112.195 ;
        RECT 65.795 112.335 66.085 112.380 ;
        RECT 67.620 112.335 67.940 112.395 ;
        RECT 65.795 112.195 67.940 112.335 ;
        RECT 65.795 112.150 66.085 112.195 ;
        RECT 67.620 112.135 67.940 112.195 ;
        RECT 74.520 112.335 74.840 112.395 ;
        RECT 75.915 112.335 76.205 112.380 ;
        RECT 79.210 112.335 79.350 112.875 ;
        RECT 81.880 112.815 82.200 112.875 ;
        RECT 83.835 113.015 84.125 113.060 ;
        RECT 86.940 113.015 87.725 113.060 ;
        RECT 83.835 112.875 87.725 113.015 ;
        RECT 83.835 112.830 84.425 112.875 ;
        RECT 79.595 112.490 79.885 112.720 ;
        RECT 80.975 112.675 81.265 112.720 ;
        RECT 83.260 112.675 83.580 112.735 ;
        RECT 80.975 112.535 83.580 112.675 ;
        RECT 80.975 112.490 81.265 112.535 ;
        RECT 74.520 112.195 79.350 112.335 ;
        RECT 74.520 112.135 74.840 112.195 ;
        RECT 75.915 112.150 76.205 112.195 ;
        RECT 28.980 111.995 29.300 112.055 ;
        RECT 26.310 111.855 29.300 111.995 ;
        RECT 28.980 111.795 29.300 111.855 ;
        RECT 30.475 111.995 30.765 112.040 ;
        RECT 33.595 111.995 33.885 112.040 ;
        RECT 35.485 111.995 35.775 112.040 ;
        RECT 30.475 111.855 35.775 111.995 ;
        RECT 30.475 111.810 30.765 111.855 ;
        RECT 33.595 111.810 33.885 111.855 ;
        RECT 35.485 111.810 35.775 111.855 ;
        RECT 44.735 111.995 45.025 112.040 ;
        RECT 47.855 111.995 48.145 112.040 ;
        RECT 49.745 111.995 50.035 112.040 ;
        RECT 44.735 111.855 50.035 111.995 ;
        RECT 44.735 111.810 45.025 111.855 ;
        RECT 47.855 111.810 48.145 111.855 ;
        RECT 49.745 111.810 50.035 111.855 ;
        RECT 58.075 111.995 58.365 112.040 ;
        RECT 61.195 111.995 61.485 112.040 ;
        RECT 63.085 111.995 63.375 112.040 ;
        RECT 58.075 111.855 63.375 111.995 ;
        RECT 58.075 111.810 58.365 111.855 ;
        RECT 61.195 111.810 61.485 111.855 ;
        RECT 63.085 111.810 63.375 111.855 ;
        RECT 70.035 111.995 70.325 112.040 ;
        RECT 73.155 111.995 73.445 112.040 ;
        RECT 75.045 111.995 75.335 112.040 ;
        RECT 79.670 111.995 79.810 112.490 ;
        RECT 83.260 112.475 83.580 112.535 ;
        RECT 84.135 112.515 84.425 112.830 ;
        RECT 86.940 112.830 87.725 112.875 ;
        RECT 86.940 112.815 87.260 112.830 ;
        RECT 89.700 112.815 90.020 113.075 ;
        RECT 94.415 113.015 94.705 113.060 ;
        RECT 97.060 113.015 97.380 113.075 ;
        RECT 97.655 113.015 98.305 113.060 ;
        RECT 94.415 112.875 98.305 113.015 ;
        RECT 94.415 112.830 95.005 112.875 ;
        RECT 85.215 112.675 85.505 112.720 ;
        RECT 88.795 112.675 89.085 112.720 ;
        RECT 90.630 112.675 90.920 112.720 ;
        RECT 85.215 112.535 90.920 112.675 ;
        RECT 85.215 112.490 85.505 112.535 ;
        RECT 88.795 112.490 89.085 112.535 ;
        RECT 90.630 112.490 90.920 112.535 ;
        RECT 94.715 112.515 95.005 112.830 ;
        RECT 97.060 112.815 97.380 112.875 ;
        RECT 97.655 112.830 98.305 112.875 ;
        RECT 100.280 112.815 100.600 113.075 ;
        RECT 104.420 112.815 104.740 113.075 ;
        RECT 106.715 113.015 107.365 113.060 ;
        RECT 110.315 113.015 110.605 113.060 ;
        RECT 112.240 113.015 112.560 113.075 ;
        RECT 106.715 112.875 112.560 113.015 ;
        RECT 106.715 112.830 107.365 112.875 ;
        RECT 110.015 112.830 110.605 112.875 ;
        RECT 95.795 112.675 96.085 112.720 ;
        RECT 99.375 112.675 99.665 112.720 ;
        RECT 101.210 112.675 101.500 112.720 ;
        RECT 95.795 112.535 101.500 112.675 ;
        RECT 95.795 112.490 96.085 112.535 ;
        RECT 99.375 112.490 99.665 112.535 ;
        RECT 101.210 112.490 101.500 112.535 ;
        RECT 101.675 112.675 101.965 112.720 ;
        RECT 103.040 112.675 103.360 112.735 ;
        RECT 101.675 112.535 103.360 112.675 ;
        RECT 101.675 112.490 101.965 112.535 ;
        RECT 103.040 112.475 103.360 112.535 ;
        RECT 103.520 112.675 103.810 112.720 ;
        RECT 105.355 112.675 105.645 112.720 ;
        RECT 108.935 112.675 109.225 112.720 ;
        RECT 103.520 112.535 109.225 112.675 ;
        RECT 103.520 112.490 103.810 112.535 ;
        RECT 105.355 112.490 105.645 112.535 ;
        RECT 108.935 112.490 109.225 112.535 ;
        RECT 110.015 112.515 110.305 112.830 ;
        RECT 112.240 112.815 112.560 112.875 ;
        RECT 81.880 112.335 82.200 112.395 ;
        RECT 86.020 112.335 86.340 112.395 ;
        RECT 91.095 112.335 91.385 112.380 ;
        RECT 81.880 112.195 91.385 112.335 ;
        RECT 81.880 112.135 82.200 112.195 ;
        RECT 86.020 112.135 86.340 112.195 ;
        RECT 91.095 112.150 91.385 112.195 ;
        RECT 91.555 112.335 91.845 112.380 ;
        RECT 94.300 112.335 94.620 112.395 ;
        RECT 91.555 112.195 94.620 112.335 ;
        RECT 91.555 112.150 91.845 112.195 ;
        RECT 94.300 112.135 94.620 112.195 ;
        RECT 106.260 112.335 106.580 112.395 ;
        RECT 113.175 112.335 113.465 112.380 ;
        RECT 106.260 112.195 113.465 112.335 ;
        RECT 106.260 112.135 106.580 112.195 ;
        RECT 113.175 112.150 113.465 112.195 ;
        RECT 70.035 111.855 75.335 111.995 ;
        RECT 70.035 111.810 70.325 111.855 ;
        RECT 73.155 111.810 73.445 111.855 ;
        RECT 75.045 111.810 75.335 111.855 ;
        RECT 75.530 111.855 79.810 111.995 ;
        RECT 85.215 111.995 85.505 112.040 ;
        RECT 88.335 111.995 88.625 112.040 ;
        RECT 90.225 111.995 90.515 112.040 ;
        RECT 85.215 111.855 90.515 111.995 ;
        RECT 20.255 111.655 20.545 111.700 ;
        RECT 22.080 111.655 22.400 111.715 ;
        RECT 20.255 111.515 22.400 111.655 ;
        RECT 20.255 111.470 20.545 111.515 ;
        RECT 22.080 111.455 22.400 111.515 ;
        RECT 23.000 111.455 23.320 111.715 ;
        RECT 24.840 111.455 25.160 111.715 ;
        RECT 36.340 111.655 36.660 111.715 ;
        RECT 37.735 111.655 38.025 111.700 ;
        RECT 36.340 111.515 38.025 111.655 ;
        RECT 36.340 111.455 36.660 111.515 ;
        RECT 37.735 111.470 38.025 111.515 ;
        RECT 40.035 111.655 40.325 111.700 ;
        RECT 40.480 111.655 40.800 111.715 ;
        RECT 40.035 111.515 40.800 111.655 ;
        RECT 40.035 111.470 40.325 111.515 ;
        RECT 40.480 111.455 40.800 111.515 ;
        RECT 53.360 111.455 53.680 111.715 ;
        RECT 65.320 111.455 65.640 111.715 ;
        RECT 71.760 111.655 72.080 111.715 ;
        RECT 75.530 111.655 75.670 111.855 ;
        RECT 85.215 111.810 85.505 111.855 ;
        RECT 88.335 111.810 88.625 111.855 ;
        RECT 90.225 111.810 90.515 111.855 ;
        RECT 95.795 111.995 96.085 112.040 ;
        RECT 98.915 111.995 99.205 112.040 ;
        RECT 100.805 111.995 101.095 112.040 ;
        RECT 95.795 111.855 101.095 111.995 ;
        RECT 95.795 111.810 96.085 111.855 ;
        RECT 98.915 111.810 99.205 111.855 ;
        RECT 100.805 111.810 101.095 111.855 ;
        RECT 103.925 111.995 104.215 112.040 ;
        RECT 105.815 111.995 106.105 112.040 ;
        RECT 108.935 111.995 109.225 112.040 ;
        RECT 103.925 111.855 109.225 111.995 ;
        RECT 103.925 111.810 104.215 111.855 ;
        RECT 105.815 111.810 106.105 111.855 ;
        RECT 108.935 111.810 109.225 111.855 ;
        RECT 71.760 111.515 75.670 111.655 ;
        RECT 71.760 111.455 72.080 111.515 ;
        RECT 77.280 111.455 77.600 111.715 ;
        RECT 80.515 111.655 80.805 111.700 ;
        RECT 84.640 111.655 84.960 111.715 ;
        RECT 80.515 111.515 84.960 111.655 ;
        RECT 80.515 111.470 80.805 111.515 ;
        RECT 84.640 111.455 84.960 111.515 ;
        RECT 14.650 110.835 115.850 111.315 ;
        RECT 28.060 110.635 28.380 110.695 ;
        RECT 46.920 110.635 47.240 110.695 ;
        RECT 47.395 110.635 47.685 110.680 ;
        RECT 28.060 110.495 39.790 110.635 ;
        RECT 28.060 110.435 28.380 110.495 ;
        RECT 21.275 110.295 21.565 110.340 ;
        RECT 24.395 110.295 24.685 110.340 ;
        RECT 26.285 110.295 26.575 110.340 ;
        RECT 21.275 110.155 26.575 110.295 ;
        RECT 21.275 110.110 21.565 110.155 ;
        RECT 24.395 110.110 24.685 110.155 ;
        RECT 26.285 110.110 26.575 110.155 ;
        RECT 31.855 110.295 32.145 110.340 ;
        RECT 34.975 110.295 35.265 110.340 ;
        RECT 36.865 110.295 37.155 110.340 ;
        RECT 31.855 110.155 37.155 110.295 ;
        RECT 31.855 110.110 32.145 110.155 ;
        RECT 34.975 110.110 35.265 110.155 ;
        RECT 36.865 110.110 37.155 110.155 ;
        RECT 17.035 109.955 17.325 110.000 ;
        RECT 23.460 109.955 23.780 110.015 ;
        RECT 17.035 109.815 23.780 109.955 ;
        RECT 17.035 109.770 17.325 109.815 ;
        RECT 23.460 109.755 23.780 109.815 ;
        RECT 27.140 109.755 27.460 110.015 ;
        RECT 27.615 109.955 27.905 110.000 ;
        RECT 34.500 109.955 34.820 110.015 ;
        RECT 27.615 109.815 34.820 109.955 ;
        RECT 27.615 109.770 27.905 109.815 ;
        RECT 34.500 109.755 34.820 109.815 ;
        RECT 36.340 109.755 36.660 110.015 ;
        RECT 37.720 109.755 38.040 110.015 ;
        RECT 39.650 109.660 39.790 110.495 ;
        RECT 46.920 110.495 47.685 110.635 ;
        RECT 46.920 110.435 47.240 110.495 ;
        RECT 47.395 110.450 47.685 110.495 ;
        RECT 60.735 110.635 61.025 110.680 ;
        RECT 61.180 110.635 61.500 110.695 ;
        RECT 60.735 110.495 61.500 110.635 ;
        RECT 60.735 110.450 61.025 110.495 ;
        RECT 61.180 110.435 61.500 110.495 ;
        RECT 86.940 110.435 87.260 110.695 ;
        RECT 109.020 110.635 109.340 110.695 ;
        RECT 111.795 110.635 112.085 110.680 ;
        RECT 112.240 110.635 112.560 110.695 ;
        RECT 109.020 110.495 110.630 110.635 ;
        RECT 109.020 110.435 109.340 110.495 ;
        RECT 52.555 110.295 52.845 110.340 ;
        RECT 55.675 110.295 55.965 110.340 ;
        RECT 57.565 110.295 57.855 110.340 ;
        RECT 52.555 110.155 57.855 110.295 ;
        RECT 52.555 110.110 52.845 110.155 ;
        RECT 55.675 110.110 55.965 110.155 ;
        RECT 57.565 110.110 57.855 110.155 ;
        RECT 68.655 110.295 68.945 110.340 ;
        RECT 71.775 110.295 72.065 110.340 ;
        RECT 73.665 110.295 73.955 110.340 ;
        RECT 68.655 110.155 73.955 110.295 ;
        RECT 68.655 110.110 68.945 110.155 ;
        RECT 71.775 110.110 72.065 110.155 ;
        RECT 73.665 110.110 73.955 110.155 ;
        RECT 80.155 110.295 80.445 110.340 ;
        RECT 83.275 110.295 83.565 110.340 ;
        RECT 85.165 110.295 85.455 110.340 ;
        RECT 80.155 110.155 85.455 110.295 ;
        RECT 80.155 110.110 80.445 110.155 ;
        RECT 83.275 110.110 83.565 110.155 ;
        RECT 85.165 110.110 85.455 110.155 ;
        RECT 94.415 110.295 94.705 110.340 ;
        RECT 97.535 110.295 97.825 110.340 ;
        RECT 99.425 110.295 99.715 110.340 ;
        RECT 103.040 110.295 103.360 110.355 ;
        RECT 94.415 110.155 99.715 110.295 ;
        RECT 94.415 110.110 94.705 110.155 ;
        RECT 97.535 110.110 97.825 110.155 ;
        RECT 99.425 110.110 99.715 110.155 ;
        RECT 100.370 110.155 103.360 110.295 ;
        RECT 53.360 109.955 53.680 110.015 ;
        RECT 57.055 109.955 57.345 110.000 ;
        RECT 53.360 109.815 57.345 109.955 ;
        RECT 53.360 109.755 53.680 109.815 ;
        RECT 57.055 109.770 57.345 109.815 ;
        RECT 58.435 109.955 58.725 110.000 ;
        RECT 60.260 109.955 60.580 110.015 ;
        RECT 58.435 109.815 60.580 109.955 ;
        RECT 58.435 109.770 58.725 109.815 ;
        RECT 60.260 109.755 60.580 109.815 ;
        RECT 65.320 109.955 65.640 110.015 ;
        RECT 73.155 109.955 73.445 110.000 ;
        RECT 65.320 109.815 73.445 109.955 ;
        RECT 65.320 109.755 65.640 109.815 ;
        RECT 73.155 109.770 73.445 109.815 ;
        RECT 74.520 109.755 74.840 110.015 ;
        RECT 75.915 109.955 76.205 110.000 ;
        RECT 78.660 109.955 78.980 110.015 ;
        RECT 75.915 109.815 78.980 109.955 ;
        RECT 75.915 109.770 76.205 109.815 ;
        RECT 78.660 109.755 78.980 109.815 ;
        RECT 84.640 109.755 84.960 110.015 ;
        RECT 86.020 109.755 86.340 110.015 ;
        RECT 92.920 109.955 93.240 110.015 ;
        RECT 100.370 110.000 100.510 110.155 ;
        RECT 103.040 110.095 103.360 110.155 ;
        RECT 104.995 110.295 105.285 110.340 ;
        RECT 108.115 110.295 108.405 110.340 ;
        RECT 110.005 110.295 110.295 110.340 ;
        RECT 104.995 110.155 110.295 110.295 ;
        RECT 104.995 110.110 105.285 110.155 ;
        RECT 108.115 110.110 108.405 110.155 ;
        RECT 110.005 110.110 110.295 110.155 ;
        RECT 98.915 109.955 99.205 110.000 ;
        RECT 92.920 109.815 99.205 109.955 ;
        RECT 92.920 109.755 93.240 109.815 ;
        RECT 98.915 109.770 99.205 109.815 ;
        RECT 100.295 109.770 100.585 110.000 ;
        RECT 100.755 109.955 101.045 110.000 ;
        RECT 101.200 109.955 101.520 110.015 ;
        RECT 100.755 109.815 101.520 109.955 ;
        RECT 100.755 109.770 101.045 109.815 ;
        RECT 101.200 109.755 101.520 109.815 ;
        RECT 101.660 109.955 101.980 110.015 ;
        RECT 109.495 109.955 109.785 110.000 ;
        RECT 101.660 109.815 109.785 109.955 ;
        RECT 110.490 109.955 110.630 110.495 ;
        RECT 111.795 110.495 112.560 110.635 ;
        RECT 111.795 110.450 112.085 110.495 ;
        RECT 112.240 110.435 112.560 110.495 ;
        RECT 110.875 109.955 111.165 110.000 ;
        RECT 110.490 109.815 111.165 109.955 ;
        RECT 101.660 109.755 101.980 109.815 ;
        RECT 109.495 109.770 109.785 109.815 ;
        RECT 110.875 109.770 111.165 109.815 ;
        RECT 20.195 109.320 20.485 109.635 ;
        RECT 21.275 109.615 21.565 109.660 ;
        RECT 24.855 109.615 25.145 109.660 ;
        RECT 26.690 109.615 26.980 109.660 ;
        RECT 21.275 109.475 26.980 109.615 ;
        RECT 21.275 109.430 21.565 109.475 ;
        RECT 24.855 109.430 25.145 109.475 ;
        RECT 26.690 109.430 26.980 109.475 ;
        RECT 19.895 109.275 20.485 109.320 ;
        RECT 23.000 109.320 23.320 109.335 ;
        RECT 23.000 109.275 23.785 109.320 ;
        RECT 19.895 109.135 23.785 109.275 ;
        RECT 19.895 109.090 20.185 109.135 ;
        RECT 23.000 109.090 23.785 109.135 ;
        RECT 25.775 109.275 26.065 109.320 ;
        RECT 29.900 109.275 30.220 109.335 ;
        RECT 30.775 109.320 31.065 109.635 ;
        RECT 31.855 109.615 32.145 109.660 ;
        RECT 35.435 109.615 35.725 109.660 ;
        RECT 37.270 109.615 37.560 109.660 ;
        RECT 31.855 109.475 37.560 109.615 ;
        RECT 31.855 109.430 32.145 109.475 ;
        RECT 35.435 109.430 35.725 109.475 ;
        RECT 37.270 109.430 37.560 109.475 ;
        RECT 39.575 109.615 39.865 109.660 ;
        RECT 40.955 109.615 41.245 109.660 ;
        RECT 47.855 109.615 48.145 109.660 ;
        RECT 39.575 109.475 48.145 109.615 ;
        RECT 39.575 109.430 39.865 109.475 ;
        RECT 40.955 109.430 41.245 109.475 ;
        RECT 47.855 109.430 48.145 109.475 ;
        RECT 25.775 109.135 30.220 109.275 ;
        RECT 25.775 109.090 26.065 109.135 ;
        RECT 23.000 109.075 23.320 109.090 ;
        RECT 29.900 109.075 30.220 109.135 ;
        RECT 30.475 109.275 31.065 109.320 ;
        RECT 33.715 109.275 34.365 109.320 ;
        RECT 39.115 109.275 39.405 109.320 ;
        RECT 30.475 109.135 39.405 109.275 ;
        RECT 30.475 109.090 30.765 109.135 ;
        RECT 33.715 109.090 34.365 109.135 ;
        RECT 39.115 109.090 39.405 109.135 ;
        RECT 41.415 108.935 41.705 108.980 ;
        RECT 41.860 108.935 42.180 108.995 ;
        RECT 41.415 108.795 42.180 108.935 ;
        RECT 47.930 108.935 48.070 109.430 ;
        RECT 48.300 109.075 48.620 109.335 ;
        RECT 51.475 109.320 51.765 109.635 ;
        RECT 52.555 109.615 52.845 109.660 ;
        RECT 56.135 109.615 56.425 109.660 ;
        RECT 57.970 109.615 58.260 109.660 ;
        RECT 52.555 109.475 58.260 109.615 ;
        RECT 52.555 109.430 52.845 109.475 ;
        RECT 56.135 109.430 56.425 109.475 ;
        RECT 57.970 109.430 58.260 109.475 ;
        RECT 59.800 109.415 60.120 109.675 ;
        RECT 61.195 109.430 61.485 109.660 ;
        RECT 61.655 109.615 61.945 109.660 ;
        RECT 67.575 109.615 67.865 109.635 ;
        RECT 61.655 109.475 67.865 109.615 ;
        RECT 61.655 109.430 61.945 109.475 ;
        RECT 51.175 109.275 51.765 109.320 ;
        RECT 53.360 109.275 53.680 109.335 ;
        RECT 54.415 109.275 55.065 109.320 ;
        RECT 51.175 109.135 55.065 109.275 ;
        RECT 51.175 109.090 51.465 109.135 ;
        RECT 53.360 109.075 53.680 109.135 ;
        RECT 54.415 109.090 55.065 109.135 ;
        RECT 58.420 109.275 58.740 109.335 ;
        RECT 61.270 109.275 61.410 109.430 ;
        RECT 58.420 109.135 61.410 109.275 ;
        RECT 62.100 109.275 62.420 109.335 ;
        RECT 67.575 109.320 67.865 109.475 ;
        RECT 68.655 109.615 68.945 109.660 ;
        RECT 72.235 109.615 72.525 109.660 ;
        RECT 74.070 109.615 74.360 109.660 ;
        RECT 68.655 109.475 74.360 109.615 ;
        RECT 68.655 109.430 68.945 109.475 ;
        RECT 72.235 109.430 72.525 109.475 ;
        RECT 74.070 109.430 74.360 109.475 ;
        RECT 79.075 109.320 79.365 109.635 ;
        RECT 80.155 109.615 80.445 109.660 ;
        RECT 83.735 109.615 84.025 109.660 ;
        RECT 85.570 109.615 85.860 109.660 ;
        RECT 80.155 109.475 85.860 109.615 ;
        RECT 80.155 109.430 80.445 109.475 ;
        RECT 83.735 109.430 84.025 109.475 ;
        RECT 85.570 109.430 85.860 109.475 ;
        RECT 87.415 109.615 87.705 109.660 ;
        RECT 88.335 109.615 88.625 109.660 ;
        RECT 87.415 109.475 88.625 109.615 ;
        RECT 87.415 109.430 87.705 109.475 ;
        RECT 88.335 109.430 88.625 109.475 ;
        RECT 88.795 109.615 89.085 109.660 ;
        RECT 93.335 109.615 93.625 109.635 ;
        RECT 88.795 109.475 93.625 109.615 ;
        RECT 88.795 109.430 89.085 109.475 ;
        RECT 64.415 109.275 64.705 109.320 ;
        RECT 62.100 109.135 64.705 109.275 ;
        RECT 58.420 109.075 58.740 109.135 ;
        RECT 62.100 109.075 62.420 109.135 ;
        RECT 64.415 109.090 64.705 109.135 ;
        RECT 67.275 109.275 67.865 109.320 ;
        RECT 70.515 109.275 71.165 109.320 ;
        RECT 67.275 109.135 71.165 109.275 ;
        RECT 67.275 109.090 67.565 109.135 ;
        RECT 70.515 109.090 71.165 109.135 ;
        RECT 78.775 109.275 79.365 109.320 ;
        RECT 80.960 109.275 81.280 109.335 ;
        RECT 82.015 109.275 82.665 109.320 ;
        RECT 78.775 109.135 82.665 109.275 ;
        RECT 78.775 109.090 79.065 109.135 ;
        RECT 80.960 109.075 81.280 109.135 ;
        RECT 82.015 109.090 82.665 109.135 ;
        RECT 53.820 108.935 54.140 108.995 ;
        RECT 47.930 108.795 54.140 108.935 ;
        RECT 41.415 108.750 41.705 108.795 ;
        RECT 41.860 108.735 42.180 108.795 ;
        RECT 53.820 108.735 54.140 108.795 ;
        RECT 78.200 108.935 78.520 108.995 ;
        RECT 87.490 108.935 87.630 109.430 ;
        RECT 89.700 109.275 90.020 109.335 ;
        RECT 93.335 109.320 93.625 109.475 ;
        RECT 94.415 109.615 94.705 109.660 ;
        RECT 97.995 109.615 98.285 109.660 ;
        RECT 99.830 109.615 100.120 109.660 ;
        RECT 94.415 109.475 100.120 109.615 ;
        RECT 94.415 109.430 94.705 109.475 ;
        RECT 97.995 109.430 98.285 109.475 ;
        RECT 99.830 109.430 100.120 109.475 ;
        RECT 90.175 109.275 90.465 109.320 ;
        RECT 89.700 109.135 90.465 109.275 ;
        RECT 89.700 109.075 90.020 109.135 ;
        RECT 90.175 109.090 90.465 109.135 ;
        RECT 93.035 109.275 93.625 109.320 ;
        RECT 96.275 109.275 96.925 109.320 ;
        RECT 93.035 109.135 96.925 109.275 ;
        RECT 93.035 109.090 93.325 109.135 ;
        RECT 96.275 109.090 96.925 109.135 ;
        RECT 100.740 109.275 101.060 109.335 ;
        RECT 103.915 109.320 104.205 109.635 ;
        RECT 104.995 109.615 105.285 109.660 ;
        RECT 108.575 109.615 108.865 109.660 ;
        RECT 110.410 109.615 110.700 109.660 ;
        RECT 104.995 109.475 110.700 109.615 ;
        RECT 104.995 109.430 105.285 109.475 ;
        RECT 108.575 109.430 108.865 109.475 ;
        RECT 110.410 109.430 110.700 109.475 ;
        RECT 112.240 109.615 112.560 109.675 ;
        RECT 112.715 109.615 113.005 109.660 ;
        RECT 112.240 109.475 113.005 109.615 ;
        RECT 112.240 109.415 112.560 109.475 ;
        RECT 112.715 109.430 113.005 109.475 ;
        RECT 103.615 109.275 104.205 109.320 ;
        RECT 106.855 109.275 107.505 109.320 ;
        RECT 100.740 109.135 107.505 109.275 ;
        RECT 100.740 109.075 101.060 109.135 ;
        RECT 103.615 109.090 103.905 109.135 ;
        RECT 106.855 109.090 107.505 109.135 ;
        RECT 78.200 108.795 87.630 108.935 ;
        RECT 78.200 108.735 78.520 108.795 ;
        RECT 113.160 108.735 113.480 108.995 ;
        RECT 14.650 108.115 115.850 108.595 ;
        RECT 53.360 107.715 53.680 107.975 ;
        RECT 58.435 107.915 58.725 107.960 ;
        RECT 58.880 107.915 59.200 107.975 ;
        RECT 77.755 107.915 78.045 107.960 ;
        RECT 58.435 107.775 59.200 107.915 ;
        RECT 58.435 107.730 58.725 107.775 ;
        RECT 58.880 107.715 59.200 107.775 ;
        RECT 74.610 107.775 78.045 107.915 ;
        RECT 22.080 107.575 22.400 107.635 ;
        RECT 28.635 107.575 28.925 107.620 ;
        RECT 31.875 107.575 32.525 107.620 ;
        RECT 22.080 107.435 32.525 107.575 ;
        RECT 22.080 107.375 22.400 107.435 ;
        RECT 28.635 107.390 29.225 107.435 ;
        RECT 31.875 107.390 32.525 107.435 ;
        RECT 41.515 107.575 41.805 107.620 ;
        RECT 44.755 107.575 45.405 107.620 ;
        RECT 41.515 107.435 45.405 107.575 ;
        RECT 41.515 107.390 42.105 107.435 ;
        RECT 44.755 107.390 45.405 107.435 ;
        RECT 69.115 107.575 69.405 107.620 ;
        RECT 72.355 107.575 73.005 107.620 ;
        RECT 74.610 107.575 74.750 107.775 ;
        RECT 77.755 107.730 78.045 107.775 ;
        RECT 80.515 107.915 80.805 107.960 ;
        RECT 80.960 107.915 81.280 107.975 ;
        RECT 80.515 107.775 81.280 107.915 ;
        RECT 80.515 107.730 80.805 107.775 ;
        RECT 80.960 107.715 81.280 107.775 ;
        RECT 96.155 107.915 96.445 107.960 ;
        RECT 97.060 107.915 97.380 107.975 ;
        RECT 96.155 107.775 97.380 107.915 ;
        RECT 96.155 107.730 96.445 107.775 ;
        RECT 97.060 107.715 97.380 107.775 ;
        RECT 100.740 107.715 101.060 107.975 ;
        RECT 108.560 107.915 108.880 107.975 ;
        RECT 112.240 107.915 112.560 107.975 ;
        RECT 101.290 107.775 112.560 107.915 ;
        RECT 69.115 107.435 74.750 107.575 ;
        RECT 74.995 107.575 75.285 107.620 ;
        RECT 77.280 107.575 77.600 107.635 ;
        RECT 101.290 107.575 101.430 107.775 ;
        RECT 108.560 107.715 108.880 107.775 ;
        RECT 112.240 107.715 112.560 107.775 ;
        RECT 74.995 107.435 77.600 107.575 ;
        RECT 69.115 107.390 69.705 107.435 ;
        RECT 72.355 107.390 73.005 107.435 ;
        RECT 74.995 107.390 75.285 107.435 ;
        RECT 28.935 107.075 29.225 107.390 ;
        RECT 41.815 107.295 42.105 107.390 ;
        RECT 30.015 107.235 30.305 107.280 ;
        RECT 33.595 107.235 33.885 107.280 ;
        RECT 35.430 107.235 35.720 107.280 ;
        RECT 30.015 107.095 35.720 107.235 ;
        RECT 30.015 107.050 30.305 107.095 ;
        RECT 33.595 107.050 33.885 107.095 ;
        RECT 35.430 107.050 35.720 107.095 ;
        RECT 35.895 107.235 36.185 107.280 ;
        RECT 37.720 107.235 38.040 107.295 ;
        RECT 35.895 107.095 38.040 107.235 ;
        RECT 35.895 107.050 36.185 107.095 ;
        RECT 37.720 107.035 38.040 107.095 ;
        RECT 41.815 107.075 42.180 107.295 ;
        RECT 41.860 107.035 42.180 107.075 ;
        RECT 42.895 107.235 43.185 107.280 ;
        RECT 46.475 107.235 46.765 107.280 ;
        RECT 48.310 107.235 48.600 107.280 ;
        RECT 42.895 107.095 48.600 107.235 ;
        RECT 42.895 107.050 43.185 107.095 ;
        RECT 46.475 107.050 46.765 107.095 ;
        RECT 48.310 107.050 48.600 107.095 ;
        RECT 48.760 107.035 49.080 107.295 ;
        RECT 53.820 107.235 54.140 107.295 ;
        RECT 58.420 107.235 58.740 107.295 ;
        RECT 58.895 107.235 59.185 107.280 ;
        RECT 53.820 107.095 59.185 107.235 ;
        RECT 53.820 107.035 54.140 107.095 ;
        RECT 58.420 107.035 58.740 107.095 ;
        RECT 58.895 107.050 59.185 107.095 ;
        RECT 69.415 107.075 69.705 107.390 ;
        RECT 77.280 107.375 77.600 107.435 ;
        RECT 100.370 107.435 101.430 107.575 ;
        RECT 105.355 107.575 105.645 107.620 ;
        RECT 105.800 107.575 106.120 107.635 ;
        RECT 105.355 107.435 106.120 107.575 ;
        RECT 70.495 107.235 70.785 107.280 ;
        RECT 74.075 107.235 74.365 107.280 ;
        RECT 75.910 107.235 76.200 107.280 ;
        RECT 70.495 107.095 76.200 107.235 ;
        RECT 70.495 107.050 70.785 107.095 ;
        RECT 74.075 107.050 74.365 107.095 ;
        RECT 75.910 107.050 76.200 107.095 ;
        RECT 78.200 107.235 78.520 107.295 ;
        RECT 100.370 107.280 100.510 107.435 ;
        RECT 105.355 107.390 105.645 107.435 ;
        RECT 105.800 107.375 106.120 107.435 ;
        RECT 107.635 107.575 108.285 107.620 ;
        RECT 111.235 107.575 111.525 107.620 ;
        RECT 113.160 107.575 113.480 107.635 ;
        RECT 107.635 107.435 113.480 107.575 ;
        RECT 107.635 107.390 108.285 107.435 ;
        RECT 110.935 107.390 111.525 107.435 ;
        RECT 80.975 107.235 81.265 107.280 ;
        RECT 96.615 107.235 96.905 107.280 ;
        RECT 100.295 107.235 100.585 107.280 ;
        RECT 78.200 107.095 100.585 107.235 ;
        RECT 78.200 107.035 78.520 107.095 ;
        RECT 80.975 107.050 81.265 107.095 ;
        RECT 96.615 107.050 96.905 107.095 ;
        RECT 100.295 107.050 100.585 107.095 ;
        RECT 103.040 107.235 103.360 107.295 ;
        RECT 103.975 107.235 104.265 107.280 ;
        RECT 103.040 107.095 104.265 107.235 ;
        RECT 103.040 107.035 103.360 107.095 ;
        RECT 103.975 107.050 104.265 107.095 ;
        RECT 104.440 107.235 104.730 107.280 ;
        RECT 106.275 107.235 106.565 107.280 ;
        RECT 109.855 107.235 110.145 107.280 ;
        RECT 104.440 107.095 110.145 107.235 ;
        RECT 104.440 107.050 104.730 107.095 ;
        RECT 106.275 107.050 106.565 107.095 ;
        RECT 109.855 107.050 110.145 107.095 ;
        RECT 110.935 107.075 111.225 107.390 ;
        RECT 113.160 107.375 113.480 107.435 ;
        RECT 12.420 106.895 12.740 106.955 ;
        RECT 25.775 106.895 26.065 106.940 ;
        RECT 12.420 106.755 26.065 106.895 ;
        RECT 12.420 106.695 12.740 106.755 ;
        RECT 25.775 106.710 26.065 106.755 ;
        RECT 38.655 106.895 38.945 106.940 ;
        RECT 40.020 106.895 40.340 106.955 ;
        RECT 38.655 106.755 40.340 106.895 ;
        RECT 38.655 106.710 38.945 106.755 ;
        RECT 40.020 106.695 40.340 106.755 ;
        RECT 40.480 106.895 40.800 106.955 ;
        RECT 47.395 106.895 47.685 106.940 ;
        RECT 40.480 106.755 47.685 106.895 ;
        RECT 40.480 106.695 40.800 106.755 ;
        RECT 47.395 106.710 47.685 106.755 ;
        RECT 66.255 106.895 66.545 106.940 ;
        RECT 73.140 106.895 73.460 106.955 ;
        RECT 66.255 106.755 73.460 106.895 ;
        RECT 66.255 106.710 66.545 106.755 ;
        RECT 73.140 106.695 73.460 106.755 ;
        RECT 74.520 106.895 74.840 106.955 ;
        RECT 76.375 106.895 76.665 106.940 ;
        RECT 74.520 106.755 76.665 106.895 ;
        RECT 74.520 106.695 74.840 106.755 ;
        RECT 76.375 106.710 76.665 106.755 ;
        RECT 112.240 106.895 112.560 106.955 ;
        RECT 114.095 106.895 114.385 106.940 ;
        RECT 112.240 106.755 114.385 106.895 ;
        RECT 112.240 106.695 112.560 106.755 ;
        RECT 114.095 106.710 114.385 106.755 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 30.015 106.555 30.305 106.600 ;
        RECT 33.135 106.555 33.425 106.600 ;
        RECT 35.025 106.555 35.315 106.600 ;
        RECT 30.015 106.415 35.315 106.555 ;
        RECT 30.015 106.370 30.305 106.415 ;
        RECT 33.135 106.370 33.425 106.415 ;
        RECT 35.025 106.370 35.315 106.415 ;
        RECT 42.895 106.555 43.185 106.600 ;
        RECT 46.015 106.555 46.305 106.600 ;
        RECT 47.905 106.555 48.195 106.600 ;
        RECT 42.895 106.415 48.195 106.555 ;
        RECT 42.895 106.370 43.185 106.415 ;
        RECT 46.015 106.370 46.305 106.415 ;
        RECT 47.905 106.370 48.195 106.415 ;
        RECT 70.495 106.555 70.785 106.600 ;
        RECT 73.615 106.555 73.905 106.600 ;
        RECT 75.505 106.555 75.795 106.600 ;
        RECT 70.495 106.415 75.795 106.555 ;
        RECT 70.495 106.370 70.785 106.415 ;
        RECT 73.615 106.370 73.905 106.415 ;
        RECT 75.505 106.370 75.795 106.415 ;
        RECT 104.845 106.555 105.135 106.600 ;
        RECT 106.735 106.555 107.025 106.600 ;
        RECT 109.855 106.555 110.145 106.600 ;
        RECT 104.845 106.415 110.145 106.555 ;
        RECT 104.845 106.370 105.135 106.415 ;
        RECT 106.735 106.370 107.025 106.415 ;
        RECT 109.855 106.370 110.145 106.415 ;
        RECT 24.840 106.215 25.160 106.275 ;
        RECT 34.580 106.215 34.870 106.260 ;
        RECT 24.840 106.075 34.870 106.215 ;
        RECT 24.840 106.015 25.160 106.075 ;
        RECT 34.580 106.030 34.870 106.075 ;
        RECT 14.650 105.395 115.850 105.875 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 34.910 206.090 36.790 206.460 ;
        RECT 64.910 206.090 66.790 206.460 ;
        RECT 94.910 206.090 96.790 206.460 ;
        RECT 19.910 203.370 21.790 203.740 ;
        RECT 49.910 203.370 51.790 203.740 ;
        RECT 79.910 203.370 81.790 203.740 ;
        RECT 109.910 203.370 111.790 203.740 ;
        RECT 72.250 202.885 72.510 203.205 ;
        RECT 63.510 202.545 63.770 202.865 ;
        RECT 58.910 201.865 59.170 202.185 ;
        RECT 34.910 200.650 36.790 201.020 ;
        RECT 58.970 199.805 59.110 201.865 ;
        RECT 59.370 201.525 59.630 201.845 ;
        RECT 58.910 199.485 59.170 199.805 ;
        RECT 58.450 198.465 58.710 198.785 ;
        RECT 19.910 197.930 21.790 198.300 ;
        RECT 49.910 197.930 51.790 198.300 ;
        RECT 53.390 196.425 53.650 196.745 ;
        RECT 34.910 195.210 36.790 195.580 ;
        RECT 42.810 193.705 43.070 194.025 ;
        RECT 46.490 193.705 46.750 194.025 ;
        RECT 19.910 192.490 21.790 192.860 ;
        RECT 31.770 191.325 32.030 191.645 ;
        RECT 30.850 190.985 31.110 191.305 ;
        RECT 27.630 188.605 27.890 188.925 ;
        RECT 25.790 187.585 26.050 187.905 ;
        RECT 19.910 187.050 21.790 187.420 ;
        RECT 25.850 186.205 25.990 187.585 ;
        RECT 27.690 186.885 27.830 188.605 ;
        RECT 27.630 186.565 27.890 186.885 ;
        RECT 30.910 186.545 31.050 190.985 ;
        RECT 30.850 186.225 31.110 186.545 ;
        RECT 25.790 185.885 26.050 186.205 ;
        RECT 26.250 185.885 26.510 186.205 ;
        RECT 21.650 185.545 21.910 185.865 ;
        RECT 24.410 185.605 24.670 185.865 ;
        RECT 24.410 185.545 25.070 185.605 ;
        RECT 21.710 184.165 21.850 185.545 ;
        RECT 24.470 185.465 25.070 185.545 ;
        RECT 24.930 185.185 25.070 185.465 ;
        RECT 23.950 184.865 24.210 185.185 ;
        RECT 24.870 184.865 25.130 185.185 ;
        RECT 21.650 183.845 21.910 184.165 ;
        RECT 22.570 182.825 22.830 183.145 ;
        RECT 19.910 181.610 21.790 181.980 ;
        RECT 22.630 179.745 22.770 182.825 ;
        RECT 24.010 182.465 24.150 184.865 ;
        RECT 26.310 184.245 26.450 185.885 ;
        RECT 30.850 184.865 31.110 185.185 ;
        RECT 25.850 184.105 26.450 184.245 ;
        RECT 25.850 183.485 25.990 184.105 ;
        RECT 25.790 183.165 26.050 183.485 ;
        RECT 26.710 183.165 26.970 183.485 ;
        RECT 24.410 182.825 24.670 183.145 ;
        RECT 23.950 182.145 24.210 182.465 ;
        RECT 24.470 180.085 24.610 182.825 ;
        RECT 26.770 182.465 26.910 183.165 ;
        RECT 30.910 182.805 31.050 184.865 ;
        RECT 31.830 183.145 31.970 191.325 ;
        RECT 37.290 190.985 37.550 191.305 ;
        RECT 33.150 190.305 33.410 190.625 ;
        RECT 34.070 190.305 34.330 190.625 ;
        RECT 33.210 189.265 33.350 190.305 ;
        RECT 33.150 188.945 33.410 189.265 ;
        RECT 34.130 187.905 34.270 190.305 ;
        RECT 34.910 189.770 36.790 190.140 ;
        RECT 34.070 187.585 34.330 187.905 ;
        RECT 33.610 186.225 33.870 186.545 ;
        RECT 33.150 185.205 33.410 185.525 ;
        RECT 32.230 184.865 32.490 185.185 ;
        RECT 31.770 182.825 32.030 183.145 ;
        RECT 30.850 182.485 31.110 182.805 ;
        RECT 26.710 182.145 26.970 182.465 ;
        RECT 24.410 179.765 24.670 180.085 ;
        RECT 21.650 179.425 21.910 179.745 ;
        RECT 22.570 179.425 22.830 179.745 ;
        RECT 26.250 179.425 26.510 179.745 ;
        RECT 21.710 178.385 21.850 179.425 ;
        RECT 21.650 178.065 21.910 178.385 ;
        RECT 22.630 177.705 22.770 179.425 ;
        RECT 26.310 178.725 26.450 179.425 ;
        RECT 26.250 178.405 26.510 178.725 ;
        RECT 26.770 178.045 26.910 182.145 ;
        RECT 30.910 180.765 31.050 182.485 ;
        RECT 30.850 180.445 31.110 180.765 ;
        RECT 26.710 177.725 26.970 178.045 ;
        RECT 30.390 177.725 30.650 178.045 ;
        RECT 22.570 177.385 22.830 177.705 ;
        RECT 19.910 176.170 21.790 176.540 ;
        RECT 22.630 175.665 22.770 177.385 ;
        RECT 22.570 175.345 22.830 175.665 ;
        RECT 20.730 174.665 20.990 174.985 ;
        RECT 20.790 172.945 20.930 174.665 ;
        RECT 24.410 174.325 24.670 174.645 ;
        RECT 22.110 173.985 22.370 174.305 ;
        RECT 20.730 172.625 20.990 172.945 ;
        RECT 18.890 171.265 19.150 171.585 ;
        RECT 18.950 169.545 19.090 171.265 ;
        RECT 19.910 170.730 21.790 171.100 ;
        RECT 18.890 169.225 19.150 169.545 ;
        RECT 17.050 168.885 17.310 169.205 ;
        RECT 17.110 167.845 17.250 168.885 ;
        RECT 17.970 168.545 18.230 168.865 ;
        RECT 17.050 167.525 17.310 167.845 ;
        RECT 18.030 167.505 18.170 168.545 ;
        RECT 17.970 167.185 18.230 167.505 ;
        RECT 16.130 166.505 16.390 166.825 ;
        RECT 16.190 164.105 16.330 166.505 ;
        RECT 19.910 165.290 21.790 165.660 ;
        RECT 17.970 164.125 18.230 164.445 ;
        RECT 16.130 163.785 16.390 164.105 ;
        RECT 18.030 156.965 18.170 164.125 ;
        RECT 19.810 163.445 20.070 163.765 ;
        RECT 19.870 162.405 20.010 163.445 ;
        RECT 19.810 162.085 20.070 162.405 ;
        RECT 18.430 161.405 18.690 161.725 ;
        RECT 17.970 156.645 18.230 156.965 ;
        RECT 18.490 150.925 18.630 161.405 ;
        RECT 19.350 160.385 19.610 160.705 ;
        RECT 18.890 158.005 19.150 158.325 ;
        RECT 18.950 151.525 19.090 158.005 ;
        RECT 19.410 156.285 19.550 160.385 ;
        RECT 19.910 159.850 21.790 160.220 ;
        RECT 19.350 155.965 19.610 156.285 ;
        RECT 19.910 154.410 21.790 154.780 ;
        RECT 19.350 152.565 19.610 152.885 ;
        RECT 18.890 151.205 19.150 151.525 ;
        RECT 18.490 150.845 19.090 150.925 ;
        RECT 18.490 150.785 19.150 150.845 ;
        RECT 18.890 150.525 19.150 150.785 ;
        RECT 18.950 147.785 19.090 150.525 ;
        RECT 19.410 148.125 19.550 152.565 ;
        RECT 19.910 148.970 21.790 149.340 ;
        RECT 19.350 147.805 19.610 148.125 ;
        RECT 18.890 147.465 19.150 147.785 ;
        RECT 19.910 143.530 21.790 143.900 ;
        RECT 22.170 143.365 22.310 173.985 ;
        RECT 24.470 172.265 24.610 174.325 ;
        RECT 26.770 172.605 26.910 177.725 ;
        RECT 27.630 176.705 27.890 177.025 ;
        RECT 27.690 174.645 27.830 176.705 ;
        RECT 30.450 175.665 30.590 177.725 ;
        RECT 30.390 175.345 30.650 175.665 ;
        RECT 27.630 174.325 27.890 174.645 ;
        RECT 26.710 172.285 26.970 172.605 ;
        RECT 27.630 172.285 27.890 172.605 ;
        RECT 23.490 171.945 23.750 172.265 ;
        RECT 24.410 171.945 24.670 172.265 ;
        RECT 26.770 172.005 26.910 172.285 ;
        RECT 23.030 169.905 23.290 170.225 ;
        RECT 22.570 161.745 22.830 162.065 ;
        RECT 22.630 159.005 22.770 161.745 ;
        RECT 22.570 158.685 22.830 159.005 ;
        RECT 22.630 155.945 22.770 158.685 ;
        RECT 23.090 156.965 23.230 169.905 ;
        RECT 23.550 166.485 23.690 171.945 ;
        RECT 26.770 171.865 27.370 172.005 ;
        RECT 27.690 171.925 27.830 172.285 ;
        RECT 26.710 171.265 26.970 171.585 ;
        RECT 24.410 169.565 24.670 169.885 ;
        RECT 24.470 167.165 24.610 169.565 ;
        RECT 26.770 169.205 26.910 171.265 ;
        RECT 27.230 170.565 27.370 171.865 ;
        RECT 27.630 171.605 27.890 171.925 ;
        RECT 29.470 171.265 29.730 171.585 ;
        RECT 27.170 170.245 27.430 170.565 ;
        RECT 26.710 168.885 26.970 169.205 ;
        RECT 24.410 166.845 24.670 167.165 ;
        RECT 23.490 166.165 23.750 166.485 ;
        RECT 24.470 162.405 24.610 166.845 ;
        RECT 29.010 166.505 29.270 166.825 ;
        RECT 29.070 164.445 29.210 166.505 ;
        RECT 25.790 164.125 26.050 164.445 ;
        RECT 29.010 164.125 29.270 164.445 ;
        RECT 24.410 162.085 24.670 162.405 ;
        RECT 25.850 159.005 25.990 164.125 ;
        RECT 29.070 161.385 29.210 164.125 ;
        RECT 29.010 161.125 29.270 161.385 ;
        RECT 28.610 161.065 29.270 161.125 ;
        RECT 28.610 160.985 29.210 161.065 ;
        RECT 25.790 158.685 26.050 159.005 ;
        RECT 23.950 158.345 24.210 158.665 ;
        RECT 23.030 156.645 23.290 156.965 ;
        RECT 23.030 155.965 23.290 156.285 ;
        RECT 22.570 155.625 22.830 155.945 ;
        RECT 23.090 152.545 23.230 155.965 ;
        RECT 24.010 154.245 24.150 158.345 ;
        RECT 24.410 154.945 24.670 155.265 ;
        RECT 23.950 153.925 24.210 154.245 ;
        RECT 24.470 153.565 24.610 154.945 ;
        RECT 25.850 153.565 25.990 158.685 ;
        RECT 27.170 158.345 27.430 158.665 ;
        RECT 24.410 153.245 24.670 153.565 ;
        RECT 25.790 153.245 26.050 153.565 ;
        RECT 23.490 152.905 23.750 153.225 ;
        RECT 23.030 152.225 23.290 152.545 ;
        RECT 23.090 150.165 23.230 152.225 ;
        RECT 23.030 149.845 23.290 150.165 ;
        RECT 22.570 149.505 22.830 149.825 ;
        RECT 22.630 147.785 22.770 149.505 ;
        RECT 23.550 148.805 23.690 152.905 ;
        RECT 24.870 152.285 25.130 152.545 ;
        RECT 24.470 152.225 25.130 152.285 ;
        RECT 24.470 152.145 25.070 152.225 ;
        RECT 23.950 150.525 24.210 150.845 ;
        RECT 24.010 148.805 24.150 150.525 ;
        RECT 23.490 148.485 23.750 148.805 ;
        RECT 23.950 148.485 24.210 148.805 ;
        RECT 22.570 147.465 22.830 147.785 ;
        RECT 22.110 143.045 22.370 143.365 ;
        RECT 23.490 142.025 23.750 142.345 ;
        RECT 18.430 141.685 18.690 142.005 ;
        RECT 18.490 137.925 18.630 141.685 ;
        RECT 19.350 141.345 19.610 141.665 ;
        RECT 18.430 137.605 18.690 137.925 ;
        RECT 19.410 135.205 19.550 141.345 ;
        RECT 23.550 140.645 23.690 142.025 ;
        RECT 23.490 140.325 23.750 140.645 ;
        RECT 22.570 139.645 22.830 139.965 ;
        RECT 22.110 138.625 22.370 138.945 ;
        RECT 19.910 138.090 21.790 138.460 ;
        RECT 22.170 136.565 22.310 138.625 ;
        RECT 22.110 136.245 22.370 136.565 ;
        RECT 21.650 135.905 21.910 136.225 ;
        RECT 19.350 134.885 19.610 135.205 ;
        RECT 21.710 134.865 21.850 135.905 ;
        RECT 22.630 135.205 22.770 139.645 ;
        RECT 23.490 137.605 23.750 137.925 ;
        RECT 23.030 135.905 23.290 136.225 ;
        RECT 22.110 134.885 22.370 135.205 ;
        RECT 22.570 134.885 22.830 135.205 ;
        RECT 21.650 134.545 21.910 134.865 ;
        RECT 22.170 134.605 22.310 134.885 ;
        RECT 23.090 134.605 23.230 135.905 ;
        RECT 22.170 134.465 23.230 134.605 ;
        RECT 19.910 132.650 21.790 133.020 ;
        RECT 22.110 131.485 22.370 131.805 ;
        RECT 17.050 130.805 17.310 131.125 ;
        RECT 17.110 124.325 17.250 130.805 ;
        RECT 19.910 127.210 21.790 127.580 ;
        RECT 18.890 125.365 19.150 125.685 ;
        RECT 18.950 124.325 19.090 125.365 ;
        RECT 22.170 124.325 22.310 131.485 ;
        RECT 22.630 129.765 22.770 134.465 ;
        RECT 23.030 132.165 23.290 132.485 ;
        RECT 22.570 129.445 22.830 129.765 ;
        RECT 17.050 124.005 17.310 124.325 ;
        RECT 18.890 124.005 19.150 124.325 ;
        RECT 22.110 124.005 22.370 124.325 ;
        RECT 23.090 123.645 23.230 132.165 ;
        RECT 23.550 129.425 23.690 137.605 ;
        RECT 23.490 129.105 23.750 129.425 ;
        RECT 23.550 125.345 23.690 129.105 ;
        RECT 23.950 127.745 24.210 128.065 ;
        RECT 24.010 126.365 24.150 127.745 ;
        RECT 23.950 126.045 24.210 126.365 ;
        RECT 23.490 125.025 23.750 125.345 ;
        RECT 23.550 124.325 23.690 125.025 ;
        RECT 23.490 124.005 23.750 124.325 ;
        RECT 23.030 123.325 23.290 123.645 ;
        RECT 19.910 121.770 21.790 122.140 ;
        RECT 19.910 116.330 21.790 116.700 ;
        RECT 17.970 114.485 18.230 114.805 ;
        RECT 22.110 114.485 22.370 114.805 ;
        RECT 12.450 106.665 12.710 106.985 ;
        RECT 12.510 95.885 12.650 106.665 ;
        RECT 18.030 95.885 18.170 114.485 ;
        RECT 22.170 113.445 22.310 114.485 ;
        RECT 22.110 113.125 22.370 113.445 ;
        RECT 24.470 112.765 24.610 152.145 ;
        RECT 25.850 148.125 25.990 153.245 ;
        RECT 27.230 150.845 27.370 158.345 ;
        RECT 28.610 155.605 28.750 160.985 ;
        RECT 28.550 155.285 28.810 155.605 ;
        RECT 27.170 150.525 27.430 150.845 ;
        RECT 25.790 147.805 26.050 148.125 ;
        RECT 27.230 147.105 27.370 150.525 ;
        RECT 28.610 150.505 28.750 155.285 ;
        RECT 29.010 154.945 29.270 155.265 ;
        RECT 29.070 153.225 29.210 154.945 ;
        RECT 29.530 153.565 29.670 171.265 ;
        RECT 30.910 169.205 31.050 180.445 ;
        RECT 31.830 177.705 31.970 182.825 ;
        RECT 32.290 178.125 32.430 184.865 ;
        RECT 33.210 182.465 33.350 185.205 ;
        RECT 33.670 184.165 33.810 186.225 ;
        RECT 33.610 183.845 33.870 184.165 ;
        RECT 33.150 182.145 33.410 182.465 ;
        RECT 33.210 181.105 33.350 182.145 ;
        RECT 33.150 180.785 33.410 181.105 ;
        RECT 33.150 180.105 33.410 180.425 ;
        RECT 32.290 177.985 32.890 178.125 ;
        RECT 31.770 177.385 32.030 177.705 ;
        RECT 32.750 175.325 32.890 177.985 ;
        RECT 32.690 175.005 32.950 175.325 ;
        RECT 31.770 173.985 32.030 174.305 ;
        RECT 31.830 172.605 31.970 173.985 ;
        RECT 31.310 172.285 31.570 172.605 ;
        RECT 31.770 172.285 32.030 172.605 ;
        RECT 32.220 172.430 32.500 172.800 ;
        RECT 32.750 172.605 32.890 175.005 ;
        RECT 32.230 172.285 32.490 172.430 ;
        RECT 32.690 172.285 32.950 172.605 ;
        RECT 31.370 171.925 31.510 172.285 ;
        RECT 31.310 171.605 31.570 171.925 ;
        RECT 29.930 168.885 30.190 169.205 ;
        RECT 30.850 168.885 31.110 169.205 ;
        RECT 29.990 167.845 30.130 168.885 ;
        RECT 29.930 167.525 30.190 167.845 ;
        RECT 30.390 166.845 30.650 167.165 ;
        RECT 29.930 163.105 30.190 163.425 ;
        RECT 29.990 161.725 30.130 163.105 ;
        RECT 30.450 162.405 30.590 166.845 ;
        RECT 30.910 164.105 31.050 168.885 ;
        RECT 31.370 168.865 31.510 171.605 ;
        RECT 32.750 169.885 32.890 172.285 ;
        RECT 33.210 170.225 33.350 180.105 ;
        RECT 33.670 172.945 33.810 183.845 ;
        RECT 34.130 173.285 34.270 187.585 ;
        RECT 34.530 186.225 34.790 186.545 ;
        RECT 34.590 185.865 34.730 186.225 ;
        RECT 34.530 185.545 34.790 185.865 ;
        RECT 35.910 185.720 36.170 185.865 ;
        RECT 35.900 185.350 36.180 185.720 ;
        RECT 36.370 185.545 36.630 185.865 ;
        RECT 36.430 185.185 36.570 185.545 ;
        RECT 36.370 184.865 36.630 185.185 ;
        RECT 34.910 184.330 36.790 184.700 ;
        RECT 34.530 183.505 34.790 183.825 ;
        RECT 37.350 183.565 37.490 190.985 ;
        RECT 42.870 190.625 43.010 193.705 ;
        RECT 44.190 193.025 44.450 193.345 ;
        RECT 39.130 190.305 39.390 190.625 ;
        RECT 42.810 190.305 43.070 190.625 ;
        RECT 39.190 188.925 39.330 190.305 ;
        RECT 39.130 188.605 39.390 188.925 ;
        RECT 39.590 188.605 39.850 188.925 ;
        RECT 38.210 188.265 38.470 188.585 ;
        RECT 38.270 186.885 38.410 188.265 ;
        RECT 39.650 187.905 39.790 188.605 ;
        RECT 42.350 187.925 42.610 188.245 ;
        RECT 39.590 187.585 39.850 187.905 ;
        RECT 40.970 187.585 41.230 187.905 ;
        RECT 38.210 186.565 38.470 186.885 ;
        RECT 39.120 185.350 39.400 185.720 ;
        RECT 38.210 184.925 38.470 185.185 ;
        RECT 38.210 184.865 38.870 184.925 ;
        RECT 38.270 184.785 38.870 184.865 ;
        RECT 34.590 181.445 34.730 183.505 ;
        RECT 36.890 183.425 37.490 183.565 ;
        RECT 34.530 181.125 34.790 181.445 ;
        RECT 36.890 180.425 37.030 183.425 ;
        RECT 37.290 182.825 37.550 183.145 ;
        RECT 36.830 180.105 37.090 180.425 ;
        RECT 34.910 178.890 36.790 179.260 ;
        RECT 37.350 175.325 37.490 182.825 ;
        RECT 37.750 176.705 38.010 177.025 ;
        RECT 37.290 175.005 37.550 175.325 ;
        RECT 37.810 174.985 37.950 176.705 ;
        RECT 37.750 174.665 38.010 174.985 ;
        RECT 34.910 173.450 36.790 173.820 ;
        RECT 34.070 172.965 34.330 173.285 ;
        RECT 33.610 172.625 33.870 172.945 ;
        RECT 34.530 172.285 34.790 172.605 ;
        RECT 34.070 171.265 34.330 171.585 ;
        RECT 33.150 169.905 33.410 170.225 ;
        RECT 32.690 169.565 32.950 169.885 ;
        RECT 33.610 168.885 33.870 169.205 ;
        RECT 31.310 168.545 31.570 168.865 ;
        RECT 33.150 168.545 33.410 168.865 ;
        RECT 30.850 163.785 31.110 164.105 ;
        RECT 30.390 162.085 30.650 162.405 ;
        RECT 30.850 161.745 31.110 162.065 ;
        RECT 29.930 161.405 30.190 161.725 ;
        RECT 29.990 156.625 30.130 161.405 ;
        RECT 30.910 159.685 31.050 161.745 ;
        RECT 30.850 159.365 31.110 159.685 ;
        RECT 29.930 156.305 30.190 156.625 ;
        RECT 30.910 155.685 31.050 159.365 ;
        RECT 32.690 157.665 32.950 157.985 ;
        RECT 32.750 156.365 32.890 157.665 ;
        RECT 33.210 156.625 33.350 168.545 ;
        RECT 33.670 167.165 33.810 168.885 ;
        RECT 33.610 166.845 33.870 167.165 ;
        RECT 32.290 156.285 32.890 156.365 ;
        RECT 33.150 156.305 33.410 156.625 ;
        RECT 31.770 155.965 32.030 156.285 ;
        RECT 32.230 156.225 32.890 156.285 ;
        RECT 32.230 155.965 32.490 156.225 ;
        RECT 30.450 155.605 31.050 155.685 ;
        RECT 30.450 155.545 31.110 155.605 ;
        RECT 30.450 155.125 30.590 155.545 ;
        RECT 30.850 155.285 31.110 155.545 ;
        RECT 29.990 154.985 30.590 155.125 ;
        RECT 29.470 153.245 29.730 153.565 ;
        RECT 29.010 152.905 29.270 153.225 ;
        RECT 29.460 152.710 29.740 153.080 ;
        RECT 28.550 150.185 28.810 150.505 ;
        RECT 27.630 149.505 27.890 149.825 ;
        RECT 27.690 147.445 27.830 149.505 ;
        RECT 27.630 147.125 27.890 147.445 ;
        RECT 27.170 146.785 27.430 147.105 ;
        RECT 25.330 144.745 25.590 145.065 ;
        RECT 25.390 142.685 25.530 144.745 ;
        RECT 25.330 142.365 25.590 142.685 ;
        RECT 24.870 139.305 25.130 139.625 ;
        RECT 24.930 137.245 25.070 139.305 ;
        RECT 25.390 137.245 25.530 142.365 ;
        RECT 26.250 139.645 26.510 139.965 ;
        RECT 24.870 136.925 25.130 137.245 ;
        RECT 25.330 136.925 25.590 137.245 ;
        RECT 24.930 134.525 25.070 136.925 ;
        RECT 24.870 134.205 25.130 134.525 ;
        RECT 25.390 131.465 25.530 136.925 ;
        RECT 26.310 135.205 26.450 139.645 ;
        RECT 27.170 138.625 27.430 138.945 ;
        RECT 27.230 137.245 27.370 138.625 ;
        RECT 27.170 136.925 27.430 137.245 ;
        RECT 28.550 136.245 28.810 136.565 ;
        RECT 26.250 134.885 26.510 135.205 ;
        RECT 28.610 134.865 28.750 136.245 ;
        RECT 28.550 134.545 28.810 134.865 ;
        RECT 28.610 134.185 28.750 134.545 ;
        RECT 29.010 134.205 29.270 134.525 ;
        RECT 28.550 133.865 28.810 134.185 ;
        RECT 28.610 132.485 28.750 133.865 ;
        RECT 28.550 132.165 28.810 132.485 ;
        RECT 29.070 131.465 29.210 134.205 ;
        RECT 25.330 131.145 25.590 131.465 ;
        RECT 29.010 131.145 29.270 131.465 ;
        RECT 25.390 129.425 25.530 131.145 ;
        RECT 26.710 130.465 26.970 130.785 ;
        RECT 25.330 129.105 25.590 129.425 ;
        RECT 25.390 126.025 25.530 129.105 ;
        RECT 25.330 125.705 25.590 126.025 ;
        RECT 25.390 121.005 25.530 125.705 ;
        RECT 24.930 120.865 25.530 121.005 ;
        RECT 24.930 120.585 25.070 120.865 ;
        RECT 24.870 120.265 25.130 120.585 ;
        RECT 26.770 120.325 26.910 130.465 ;
        RECT 28.090 125.705 28.350 126.025 ;
        RECT 27.170 125.025 27.430 125.345 ;
        RECT 27.230 120.925 27.370 125.025 ;
        RECT 28.150 124.325 28.290 125.705 ;
        RECT 28.090 124.005 28.350 124.325 ;
        RECT 29.070 123.985 29.210 131.145 ;
        RECT 29.010 123.665 29.270 123.985 ;
        RECT 27.170 120.605 27.430 120.925 ;
        RECT 24.930 116.165 25.070 120.265 ;
        RECT 26.770 120.245 27.370 120.325 ;
        RECT 26.770 120.185 27.430 120.245 ;
        RECT 27.170 119.925 27.430 120.185 ;
        RECT 29.070 118.205 29.210 123.665 ;
        RECT 29.010 117.885 29.270 118.205 ;
        RECT 24.870 115.845 25.130 116.165 ;
        RECT 27.170 115.165 27.430 115.485 ;
        RECT 24.410 112.445 24.670 112.765 ;
        RECT 27.230 112.425 27.370 115.165 ;
        RECT 29.530 115.145 29.670 152.710 ;
        RECT 29.990 151.185 30.130 154.985 ;
        RECT 31.830 154.245 31.970 155.965 ;
        RECT 30.390 153.925 30.650 154.245 ;
        RECT 31.770 153.925 32.030 154.245 ;
        RECT 29.930 150.865 30.190 151.185 ;
        RECT 29.930 139.305 30.190 139.625 ;
        RECT 29.990 135.205 30.130 139.305 ;
        RECT 30.450 137.925 30.590 153.925 ;
        RECT 32.750 153.225 32.890 156.225 ;
        RECT 33.610 155.965 33.870 156.285 ;
        RECT 33.670 153.225 33.810 155.965 ;
        RECT 32.690 152.905 32.950 153.225 ;
        RECT 33.150 152.905 33.410 153.225 ;
        RECT 33.610 152.905 33.870 153.225 ;
        RECT 31.310 152.225 31.570 152.545 ;
        RECT 31.370 142.345 31.510 152.225 ;
        RECT 32.750 151.185 32.890 152.905 ;
        RECT 32.690 150.865 32.950 151.185 ;
        RECT 33.210 150.845 33.350 152.905 ;
        RECT 33.670 151.040 33.810 152.905 ;
        RECT 33.150 150.525 33.410 150.845 ;
        RECT 33.600 150.670 33.880 151.040 ;
        RECT 33.610 149.505 33.870 149.825 ;
        RECT 31.770 143.045 32.030 143.365 ;
        RECT 33.150 143.045 33.410 143.365 ;
        RECT 31.310 142.025 31.570 142.345 ;
        RECT 31.310 141.345 31.570 141.665 ;
        RECT 30.850 139.645 31.110 139.965 ;
        RECT 30.390 137.605 30.650 137.925 ;
        RECT 30.910 137.585 31.050 139.645 ;
        RECT 30.850 137.265 31.110 137.585 ;
        RECT 29.930 134.885 30.190 135.205 ;
        RECT 30.850 134.205 31.110 134.525 ;
        RECT 30.390 133.525 30.650 133.845 ;
        RECT 30.450 130.525 30.590 133.525 ;
        RECT 30.910 131.125 31.050 134.205 ;
        RECT 30.850 130.805 31.110 131.125 ;
        RECT 30.450 130.385 31.050 130.525 ;
        RECT 30.910 128.745 31.050 130.385 ;
        RECT 30.850 128.425 31.110 128.745 ;
        RECT 29.930 126.045 30.190 126.365 ;
        RECT 29.990 123.985 30.130 126.045 ;
        RECT 30.390 125.705 30.650 126.025 ;
        RECT 30.450 124.325 30.590 125.705 ;
        RECT 30.390 124.005 30.650 124.325 ;
        RECT 29.930 123.665 30.190 123.985 ;
        RECT 30.910 123.305 31.050 128.425 ;
        RECT 29.930 122.985 30.190 123.305 ;
        RECT 30.850 122.985 31.110 123.305 ;
        RECT 29.990 122.625 30.130 122.985 ;
        RECT 29.930 122.305 30.190 122.625 ;
        RECT 29.990 120.925 30.130 122.305 ;
        RECT 29.930 120.605 30.190 120.925 ;
        RECT 31.370 115.145 31.510 141.345 ;
        RECT 31.830 140.645 31.970 143.045 ;
        RECT 32.690 141.345 32.950 141.665 ;
        RECT 31.770 140.325 32.030 140.645 ;
        RECT 32.230 125.365 32.490 125.685 ;
        RECT 31.770 123.325 32.030 123.645 ;
        RECT 31.830 122.625 31.970 123.325 ;
        RECT 31.770 122.305 32.030 122.625 ;
        RECT 31.830 120.585 31.970 122.305 ;
        RECT 31.770 120.265 32.030 120.585 ;
        RECT 32.290 118.885 32.430 125.365 ;
        RECT 32.230 118.565 32.490 118.885 ;
        RECT 32.750 115.145 32.890 141.345 ;
        RECT 33.210 137.925 33.350 143.045 ;
        RECT 33.670 142.345 33.810 149.505 ;
        RECT 34.130 142.685 34.270 171.265 ;
        RECT 34.590 170.565 34.730 172.285 ;
        RECT 34.990 171.945 35.250 172.265 ;
        RECT 34.530 170.245 34.790 170.565 ;
        RECT 35.050 169.965 35.190 171.945 ;
        RECT 38.210 171.265 38.470 171.585 ;
        RECT 34.590 169.825 35.190 169.965 ;
        RECT 34.590 167.845 34.730 169.825 ;
        RECT 37.290 169.225 37.550 169.545 ;
        RECT 34.910 168.010 36.790 168.380 ;
        RECT 34.530 167.525 34.790 167.845 ;
        RECT 37.350 164.785 37.490 169.225 ;
        RECT 37.750 168.885 38.010 169.205 ;
        RECT 36.820 164.270 37.100 164.640 ;
        RECT 37.290 164.465 37.550 164.785 ;
        RECT 36.890 164.105 37.030 164.270 ;
        RECT 37.810 164.105 37.950 168.885 ;
        RECT 36.830 163.785 37.090 164.105 ;
        RECT 37.290 163.785 37.550 164.105 ;
        RECT 37.750 163.785 38.010 164.105 ;
        RECT 34.910 162.570 36.790 162.940 ;
        RECT 37.350 161.385 37.490 163.785 ;
        RECT 38.270 163.165 38.410 171.265 ;
        RECT 37.810 163.025 38.410 163.165 ;
        RECT 37.290 161.065 37.550 161.385 ;
        RECT 35.910 160.385 36.170 160.705 ;
        RECT 35.970 159.005 36.110 160.385 ;
        RECT 36.830 159.365 37.090 159.685 ;
        RECT 35.910 158.685 36.170 159.005 ;
        RECT 36.890 158.405 37.030 159.365 ;
        RECT 36.890 158.265 37.490 158.405 ;
        RECT 37.350 157.985 37.490 158.265 ;
        RECT 37.290 157.665 37.550 157.985 ;
        RECT 34.910 157.130 36.790 157.500 ;
        RECT 37.350 156.365 37.490 157.665 ;
        RECT 35.970 156.225 37.490 156.365 ;
        RECT 35.450 155.285 35.710 155.605 ;
        RECT 34.530 153.925 34.790 154.245 ;
        RECT 34.590 150.845 34.730 153.925 ;
        RECT 35.510 153.225 35.650 155.285 ;
        RECT 35.970 153.225 36.110 156.225 ;
        RECT 36.370 155.285 36.630 155.605 ;
        RECT 36.430 154.245 36.570 155.285 ;
        RECT 37.810 155.125 37.950 163.025 ;
        RECT 38.210 159.025 38.470 159.345 ;
        RECT 38.270 156.285 38.410 159.025 ;
        RECT 38.210 155.965 38.470 156.285 ;
        RECT 37.350 154.985 37.950 155.125 ;
        RECT 36.370 153.925 36.630 154.245 ;
        RECT 36.430 153.225 36.570 153.925 ;
        RECT 36.830 153.585 37.090 153.905 ;
        RECT 35.450 152.905 35.710 153.225 ;
        RECT 35.910 152.905 36.170 153.225 ;
        RECT 36.370 152.905 36.630 153.225 ;
        RECT 36.890 153.080 37.030 153.585 ;
        RECT 37.350 153.225 37.490 154.985 ;
        RECT 37.750 153.925 38.010 154.245 ;
        RECT 36.820 152.710 37.100 153.080 ;
        RECT 37.290 152.905 37.550 153.225 ;
        RECT 37.810 152.285 37.950 153.925 ;
        RECT 38.270 153.565 38.410 155.965 ;
        RECT 38.210 153.245 38.470 153.565 ;
        RECT 37.350 152.145 37.950 152.285 ;
        RECT 34.910 151.690 36.790 152.060 ;
        RECT 34.530 150.525 34.790 150.845 ;
        RECT 36.820 150.670 37.100 151.040 ;
        RECT 36.830 150.525 37.090 150.670 ;
        RECT 34.530 149.845 34.790 150.165 ;
        RECT 34.590 147.785 34.730 149.845 ;
        RECT 34.530 147.465 34.790 147.785 ;
        RECT 34.910 146.250 36.790 146.620 ;
        RECT 37.350 142.765 37.490 152.145 ;
        RECT 38.210 149.505 38.470 149.825 ;
        RECT 37.750 144.745 38.010 145.065 ;
        RECT 37.810 143.365 37.950 144.745 ;
        RECT 37.750 143.045 38.010 143.365 ;
        RECT 34.070 142.365 34.330 142.685 ;
        RECT 37.350 142.625 37.950 142.765 ;
        RECT 33.610 142.025 33.870 142.345 ;
        RECT 37.290 141.685 37.550 142.005 ;
        RECT 34.910 140.810 36.790 141.180 ;
        RECT 37.350 140.305 37.490 141.685 ;
        RECT 37.290 139.985 37.550 140.305 ;
        RECT 37.810 139.535 37.950 142.625 ;
        RECT 37.350 139.395 37.950 139.535 ;
        RECT 37.350 137.925 37.490 139.395 ;
        RECT 38.270 137.925 38.410 149.505 ;
        RECT 38.730 147.105 38.870 184.785 ;
        RECT 39.190 172.800 39.330 185.350 ;
        RECT 41.030 183.825 41.170 187.585 ;
        RECT 40.970 183.505 41.230 183.825 ;
        RECT 42.410 183.485 42.550 187.925 ;
        RECT 42.350 183.165 42.610 183.485 ;
        RECT 40.970 180.105 41.230 180.425 ;
        RECT 41.030 178.045 41.170 180.105 ;
        RECT 41.430 179.425 41.690 179.745 ;
        RECT 42.350 179.425 42.610 179.745 ;
        RECT 40.970 177.725 41.230 178.045 ;
        RECT 40.050 176.705 40.310 177.025 ;
        RECT 39.120 172.430 39.400 172.800 ;
        RECT 39.590 168.545 39.850 168.865 ;
        RECT 39.650 167.845 39.790 168.545 ;
        RECT 39.590 167.525 39.850 167.845 ;
        RECT 39.130 166.505 39.390 166.825 ;
        RECT 39.190 165.125 39.330 166.505 ;
        RECT 39.130 164.805 39.390 165.125 ;
        RECT 39.120 164.270 39.400 164.640 ;
        RECT 39.190 159.005 39.330 164.270 ;
        RECT 39.590 160.385 39.850 160.705 ;
        RECT 39.130 158.685 39.390 159.005 ;
        RECT 39.130 157.665 39.390 157.985 ;
        RECT 39.190 156.625 39.330 157.665 ;
        RECT 39.130 156.305 39.390 156.625 ;
        RECT 39.130 154.945 39.390 155.265 ;
        RECT 39.190 153.565 39.330 154.945 ;
        RECT 39.130 153.245 39.390 153.565 ;
        RECT 39.650 152.965 39.790 160.385 ;
        RECT 39.190 152.825 39.790 152.965 ;
        RECT 38.670 146.785 38.930 147.105 ;
        RECT 38.670 145.425 38.930 145.745 ;
        RECT 38.730 143.025 38.870 145.425 ;
        RECT 38.670 142.705 38.930 143.025 ;
        RECT 39.190 142.255 39.330 152.825 ;
        RECT 39.590 152.225 39.850 152.545 ;
        RECT 38.730 142.115 39.330 142.255 ;
        RECT 33.150 137.605 33.410 137.925 ;
        RECT 37.290 137.605 37.550 137.925 ;
        RECT 38.210 137.605 38.470 137.925 ;
        RECT 33.610 136.245 33.870 136.565 ;
        RECT 33.150 123.325 33.410 123.645 ;
        RECT 33.210 121.605 33.350 123.325 ;
        RECT 33.670 122.965 33.810 136.245 ;
        RECT 34.910 135.370 36.790 135.740 ;
        RECT 37.750 134.885 38.010 135.205 ;
        RECT 37.290 133.185 37.550 133.505 ;
        RECT 34.990 131.715 35.250 131.805 ;
        RECT 34.590 131.575 35.250 131.715 ;
        RECT 34.590 129.765 34.730 131.575 ;
        RECT 34.990 131.485 35.250 131.575 ;
        RECT 34.910 129.930 36.790 130.300 ;
        RECT 34.530 129.445 34.790 129.765 ;
        RECT 37.350 129.085 37.490 133.185 ;
        RECT 37.290 128.765 37.550 129.085 ;
        RECT 37.290 126.725 37.550 127.045 ;
        RECT 34.910 124.490 36.790 124.860 ;
        RECT 33.610 122.645 33.870 122.965 ;
        RECT 33.150 121.285 33.410 121.605 ;
        RECT 37.350 120.245 37.490 126.725 ;
        RECT 37.290 119.925 37.550 120.245 ;
        RECT 34.910 119.050 36.790 119.420 ;
        RECT 28.090 114.825 28.350 115.145 ;
        RECT 29.470 114.825 29.730 115.145 ;
        RECT 31.310 114.825 31.570 115.145 ;
        RECT 32.690 114.825 32.950 115.145 ;
        RECT 28.150 113.105 28.290 114.825 ;
        RECT 28.550 114.485 28.810 114.805 ;
        RECT 28.610 113.105 28.750 114.485 ;
        RECT 29.930 114.145 30.190 114.465 ;
        RECT 34.530 114.145 34.790 114.465 ;
        RECT 28.090 112.785 28.350 113.105 ;
        RECT 28.550 112.785 28.810 113.105 ;
        RECT 27.170 112.105 27.430 112.425 ;
        RECT 22.110 111.425 22.370 111.745 ;
        RECT 23.030 111.425 23.290 111.745 ;
        RECT 24.870 111.425 25.130 111.745 ;
        RECT 19.910 110.890 21.790 111.260 ;
        RECT 22.170 107.665 22.310 111.425 ;
        RECT 23.090 109.365 23.230 111.425 ;
        RECT 23.490 109.725 23.750 110.045 ;
        RECT 23.030 109.045 23.290 109.365 ;
        RECT 22.110 107.345 22.370 107.665 ;
        RECT 19.910 105.450 21.790 105.820 ;
        RECT 23.550 95.885 23.690 109.725 ;
        RECT 24.930 106.305 25.070 111.425 ;
        RECT 27.230 110.045 27.370 112.105 ;
        RECT 28.150 110.725 28.290 112.785 ;
        RECT 29.010 111.765 29.270 112.085 ;
        RECT 28.090 110.405 28.350 110.725 ;
        RECT 27.170 109.725 27.430 110.045 ;
        RECT 24.870 105.985 25.130 106.305 ;
        RECT 29.070 95.885 29.210 111.765 ;
        RECT 29.990 109.365 30.130 114.145 ;
        RECT 34.590 113.105 34.730 114.145 ;
        RECT 34.910 113.610 36.790 113.980 ;
        RECT 37.810 113.105 37.950 134.885 ;
        RECT 38.730 134.525 38.870 142.115 ;
        RECT 39.650 136.905 39.790 152.225 ;
        RECT 40.110 150.845 40.250 176.705 ;
        RECT 40.510 171.265 40.770 171.585 ;
        RECT 40.570 163.425 40.710 171.265 ;
        RECT 40.970 166.845 41.230 167.165 ;
        RECT 41.030 166.680 41.170 166.845 ;
        RECT 40.960 166.310 41.240 166.680 ;
        RECT 41.030 163.765 41.170 166.310 ;
        RECT 40.970 163.445 41.230 163.765 ;
        RECT 40.510 163.105 40.770 163.425 ;
        RECT 40.570 162.065 40.710 163.105 ;
        RECT 40.510 161.745 40.770 162.065 ;
        RECT 41.490 161.805 41.630 179.425 ;
        RECT 42.410 178.045 42.550 179.425 ;
        RECT 42.870 178.045 43.010 190.305 ;
        RECT 44.250 189.265 44.390 193.025 ;
        RECT 46.030 192.005 46.290 192.325 ;
        RECT 44.190 188.945 44.450 189.265 ;
        RECT 43.270 186.225 43.530 186.545 ;
        RECT 43.330 179.745 43.470 186.225 ;
        RECT 43.730 185.205 43.990 185.525 ;
        RECT 43.790 184.165 43.930 185.205 ;
        RECT 44.190 185.095 44.450 185.185 ;
        RECT 44.190 184.955 44.850 185.095 ;
        RECT 44.190 184.865 44.450 184.955 ;
        RECT 43.730 183.845 43.990 184.165 ;
        RECT 43.730 182.825 43.990 183.145 ;
        RECT 43.270 179.425 43.530 179.745 ;
        RECT 43.330 178.045 43.470 179.425 ;
        RECT 41.890 177.725 42.150 178.045 ;
        RECT 42.350 177.725 42.610 178.045 ;
        RECT 42.810 177.725 43.070 178.045 ;
        RECT 43.270 177.725 43.530 178.045 ;
        RECT 41.950 174.895 42.090 177.725 ;
        RECT 42.410 175.405 42.550 177.725 ;
        RECT 43.330 175.665 43.470 177.725 ;
        RECT 42.410 175.265 43.010 175.405 ;
        RECT 43.270 175.345 43.530 175.665 ;
        RECT 42.350 174.895 42.610 174.985 ;
        RECT 41.950 174.755 42.610 174.895 ;
        RECT 42.350 174.665 42.610 174.755 ;
        RECT 42.870 174.645 43.010 175.265 ;
        RECT 42.810 174.325 43.070 174.645 ;
        RECT 42.870 172.945 43.010 174.325 ;
        RECT 43.330 173.285 43.470 175.345 ;
        RECT 43.790 175.325 43.930 182.825 ;
        RECT 44.710 182.465 44.850 184.955 ;
        RECT 45.570 184.865 45.830 185.185 ;
        RECT 45.630 184.165 45.770 184.865 ;
        RECT 45.570 183.845 45.830 184.165 ;
        RECT 46.090 183.145 46.230 192.005 ;
        RECT 46.550 189.605 46.690 193.705 ;
        RECT 48.330 193.025 48.590 193.345 ;
        RECT 49.250 193.025 49.510 193.345 ;
        RECT 48.390 190.965 48.530 193.025 ;
        RECT 49.310 191.985 49.450 193.025 ;
        RECT 49.910 192.490 51.790 192.860 ;
        RECT 49.250 191.665 49.510 191.985 ;
        RECT 53.450 191.645 53.590 196.425 ;
        RECT 58.510 196.405 58.650 198.465 ;
        RECT 58.450 196.085 58.710 196.405 ;
        RECT 53.850 194.385 54.110 194.705 ;
        RECT 52.010 191.325 52.270 191.645 ;
        RECT 53.390 191.325 53.650 191.645 ;
        RECT 51.550 190.985 51.810 191.305 ;
        RECT 48.330 190.645 48.590 190.965 ;
        RECT 51.610 189.605 51.750 190.985 ;
        RECT 46.490 189.285 46.750 189.605 ;
        RECT 51.550 189.285 51.810 189.605 ;
        RECT 47.410 188.265 47.670 188.585 ;
        RECT 48.790 188.265 49.050 188.585 ;
        RECT 47.470 186.205 47.610 188.265 ;
        RECT 47.410 185.885 47.670 186.205 ;
        RECT 46.030 182.825 46.290 183.145 ;
        RECT 46.950 182.485 47.210 182.805 ;
        RECT 44.650 182.145 44.910 182.465 ;
        RECT 44.710 180.425 44.850 182.145 ;
        RECT 47.010 181.445 47.150 182.485 ;
        RECT 45.110 181.125 45.370 181.445 ;
        RECT 46.950 181.125 47.210 181.445 ;
        RECT 45.170 180.425 45.310 181.125 ;
        RECT 47.470 180.845 47.610 185.885 ;
        RECT 48.850 184.165 48.990 188.265 ;
        RECT 49.910 187.050 51.790 187.420 ;
        RECT 52.070 185.865 52.210 191.325 ;
        RECT 53.910 188.925 54.050 194.385 ;
        RECT 58.970 191.305 59.110 199.485 ;
        RECT 59.430 198.785 59.570 201.525 ;
        RECT 61.210 201.185 61.470 201.505 ;
        RECT 63.050 201.185 63.310 201.505 ;
        RECT 61.270 199.805 61.410 201.185 ;
        RECT 61.210 199.485 61.470 199.805 ;
        RECT 59.370 198.465 59.630 198.785 ;
        RECT 59.430 195.045 59.570 198.465 ;
        RECT 63.110 197.085 63.250 201.185 ;
        RECT 63.570 197.425 63.710 202.545 ;
        RECT 67.190 201.865 67.450 202.185 ;
        RECT 64.910 200.650 66.790 201.020 ;
        RECT 63.510 197.105 63.770 197.425 ;
        RECT 63.050 196.765 63.310 197.085 ;
        RECT 59.370 194.725 59.630 195.045 ;
        RECT 63.570 194.705 63.710 197.105 ;
        RECT 67.250 197.085 67.390 201.865 ;
        RECT 69.030 201.525 69.290 201.845 ;
        RECT 68.110 201.185 68.370 201.505 ;
        RECT 68.170 199.465 68.310 201.185 ;
        RECT 68.110 199.145 68.370 199.465 ;
        RECT 67.190 196.765 67.450 197.085 ;
        RECT 63.970 196.425 64.230 196.745 ;
        RECT 63.510 194.385 63.770 194.705 ;
        RECT 62.130 194.045 62.390 194.365 ;
        RECT 62.590 194.045 62.850 194.365 ;
        RECT 60.750 192.005 61.010 192.325 ;
        RECT 60.810 191.305 60.950 192.005 ;
        RECT 62.190 191.645 62.330 194.045 ;
        RECT 62.130 191.325 62.390 191.645 ;
        RECT 62.650 191.305 62.790 194.045 ;
        RECT 58.910 190.985 59.170 191.305 ;
        RECT 60.750 190.985 61.010 191.305 ;
        RECT 62.590 190.985 62.850 191.305 ;
        RECT 55.690 190.645 55.950 190.965 ;
        RECT 55.750 189.605 55.890 190.645 ;
        RECT 55.690 189.285 55.950 189.605 ;
        RECT 53.850 188.605 54.110 188.925 ;
        RECT 52.010 185.545 52.270 185.865 ;
        RECT 48.790 183.845 49.050 184.165 ;
        RECT 47.010 180.765 47.610 180.845 ;
        RECT 48.330 180.785 48.590 181.105 ;
        RECT 46.950 180.705 47.610 180.765 ;
        RECT 46.950 180.445 47.210 180.705 ;
        RECT 44.650 180.105 44.910 180.425 ;
        RECT 45.110 180.105 45.370 180.425 ;
        RECT 47.010 177.705 47.150 180.445 ;
        RECT 48.390 178.805 48.530 180.785 ;
        RECT 47.930 178.725 48.530 178.805 ;
        RECT 47.930 178.665 48.590 178.725 ;
        RECT 46.950 177.385 47.210 177.705 ;
        RECT 47.010 175.325 47.150 177.385 ;
        RECT 43.730 175.005 43.990 175.325 ;
        RECT 46.950 175.005 47.210 175.325 ;
        RECT 46.490 174.665 46.750 174.985 ;
        RECT 45.570 174.325 45.830 174.645 ;
        RECT 43.730 173.985 43.990 174.305 ;
        RECT 43.270 172.965 43.530 173.285 ;
        RECT 42.810 172.625 43.070 172.945 ;
        RECT 41.890 168.545 42.150 168.865 ;
        RECT 41.950 164.105 42.090 168.545 ;
        RECT 42.350 167.185 42.610 167.505 ;
        RECT 41.890 163.785 42.150 164.105 ;
        RECT 41.950 162.405 42.090 163.785 ;
        RECT 41.890 162.085 42.150 162.405 ;
        RECT 41.490 161.665 42.090 161.805 ;
        RECT 42.410 161.725 42.550 167.185 ;
        RECT 42.810 166.505 43.070 166.825 ;
        RECT 42.870 164.640 43.010 166.505 ;
        RECT 42.800 164.270 43.080 164.640 ;
        RECT 40.970 157.665 41.230 157.985 ;
        RECT 41.430 157.665 41.690 157.985 ;
        RECT 41.030 156.285 41.170 157.665 ;
        RECT 40.970 155.965 41.230 156.285 ;
        RECT 40.510 154.945 40.770 155.265 ;
        RECT 40.570 150.845 40.710 154.945 ;
        RECT 40.970 152.905 41.230 153.225 ;
        RECT 40.050 150.525 40.310 150.845 ;
        RECT 40.510 150.525 40.770 150.845 ;
        RECT 40.510 149.505 40.770 149.825 ;
        RECT 40.050 147.695 40.310 147.785 ;
        RECT 40.570 147.695 40.710 149.505 ;
        RECT 41.030 148.805 41.170 152.905 ;
        RECT 40.970 148.485 41.230 148.805 ;
        RECT 40.050 147.555 40.710 147.695 ;
        RECT 40.050 147.465 40.310 147.555 ;
        RECT 40.050 146.785 40.310 147.105 ;
        RECT 40.110 137.245 40.250 146.785 ;
        RECT 40.570 142.345 40.710 147.555 ;
        RECT 40.510 142.025 40.770 142.345 ;
        RECT 40.570 139.965 40.710 142.025 ;
        RECT 40.510 139.645 40.770 139.965 ;
        RECT 40.510 137.605 40.770 137.925 ;
        RECT 40.050 136.925 40.310 137.245 ;
        RECT 39.590 136.585 39.850 136.905 ;
        RECT 39.130 135.905 39.390 136.225 ;
        RECT 39.590 135.905 39.850 136.225 ;
        RECT 38.670 134.205 38.930 134.525 ;
        RECT 38.210 133.865 38.470 134.185 ;
        RECT 38.270 131.805 38.410 133.865 ;
        RECT 38.210 131.485 38.470 131.805 ;
        RECT 38.270 127.045 38.410 131.485 ;
        RECT 38.670 128.765 38.930 129.085 ;
        RECT 38.210 126.725 38.470 127.045 ;
        RECT 38.730 124.405 38.870 128.765 ;
        RECT 38.270 124.325 38.870 124.405 ;
        RECT 38.210 124.265 38.870 124.325 ;
        RECT 38.210 124.005 38.470 124.265 ;
        RECT 38.270 120.925 38.410 124.005 ;
        RECT 38.670 123.665 38.930 123.985 ;
        RECT 38.210 120.605 38.470 120.925 ;
        RECT 38.730 118.885 38.870 123.665 ;
        RECT 38.670 118.565 38.930 118.885 ;
        RECT 39.190 118.285 39.330 135.905 ;
        RECT 39.650 131.465 39.790 135.905 ;
        RECT 40.050 133.185 40.310 133.505 ;
        RECT 39.590 131.145 39.850 131.465 ;
        RECT 39.590 127.745 39.850 128.065 ;
        RECT 38.730 118.145 39.330 118.285 ;
        RECT 39.650 118.205 39.790 127.745 ;
        RECT 40.110 120.585 40.250 133.185 ;
        RECT 40.570 132.485 40.710 137.605 ;
        RECT 41.490 134.525 41.630 157.665 ;
        RECT 41.950 152.965 42.090 161.665 ;
        RECT 42.350 161.405 42.610 161.725 ;
        RECT 43.270 161.405 43.530 161.725 ;
        RECT 42.810 160.385 43.070 160.705 ;
        RECT 42.870 158.575 43.010 160.385 ;
        RECT 43.330 159.345 43.470 161.405 ;
        RECT 43.270 159.025 43.530 159.345 ;
        RECT 43.270 158.575 43.530 158.665 ;
        RECT 42.870 158.435 43.530 158.575 ;
        RECT 43.270 158.345 43.530 158.435 ;
        RECT 42.810 157.665 43.070 157.985 ;
        RECT 42.870 153.225 43.010 157.665 ;
        RECT 43.330 156.285 43.470 158.345 ;
        RECT 43.270 155.965 43.530 156.285 ;
        RECT 43.270 153.585 43.530 153.905 ;
        RECT 41.950 152.825 42.550 152.965 ;
        RECT 42.810 152.905 43.070 153.225 ;
        RECT 41.890 152.400 42.150 152.545 ;
        RECT 41.880 152.030 42.160 152.400 ;
        RECT 42.410 148.715 42.550 152.825 ;
        RECT 41.950 148.575 42.550 148.715 ;
        RECT 40.970 134.205 41.230 134.525 ;
        RECT 41.430 134.205 41.690 134.525 ;
        RECT 40.510 132.165 40.770 132.485 ;
        RECT 41.030 132.145 41.170 134.205 ;
        RECT 41.950 134.185 42.090 148.575 ;
        RECT 42.350 147.805 42.610 148.125 ;
        RECT 42.410 142.345 42.550 147.805 ;
        RECT 42.350 142.025 42.610 142.345 ;
        RECT 43.330 134.185 43.470 153.585 ;
        RECT 43.790 153.565 43.930 173.985 ;
        RECT 45.630 172.605 45.770 174.325 ;
        RECT 45.570 172.285 45.830 172.605 ;
        RECT 46.550 172.265 46.690 174.665 ;
        RECT 46.950 172.965 47.210 173.285 ;
        RECT 47.010 172.605 47.150 172.965 ;
        RECT 47.930 172.945 48.070 178.665 ;
        RECT 48.330 178.405 48.590 178.665 ;
        RECT 48.330 177.725 48.590 178.045 ;
        RECT 48.390 174.985 48.530 177.725 ;
        RECT 48.330 174.665 48.590 174.985 ;
        RECT 48.850 174.645 48.990 183.845 ;
        RECT 49.250 182.825 49.510 183.145 ;
        RECT 49.310 180.425 49.450 182.825 ;
        RECT 49.910 181.610 51.790 181.980 ;
        RECT 52.070 180.765 52.210 185.545 ;
        RECT 53.910 183.485 54.050 188.605 ;
        RECT 53.850 183.165 54.110 183.485 ;
        RECT 56.150 183.165 56.410 183.485 ;
        RECT 52.010 180.445 52.270 180.765 ;
        RECT 49.250 180.105 49.510 180.425 ;
        RECT 49.910 176.170 51.790 176.540 ;
        RECT 50.630 175.685 50.890 176.005 ;
        RECT 49.710 175.345 49.970 175.665 ;
        RECT 48.790 174.325 49.050 174.645 ;
        RECT 49.240 174.470 49.520 174.840 ;
        RECT 47.870 172.625 48.130 172.945 ;
        RECT 49.310 172.605 49.450 174.470 ;
        RECT 49.770 172.605 49.910 175.345 ;
        RECT 50.170 175.005 50.430 175.325 ;
        RECT 50.230 172.945 50.370 175.005 ;
        RECT 50.690 173.285 50.830 175.685 ;
        RECT 55.690 174.325 55.950 174.645 ;
        RECT 51.550 173.985 51.810 174.305 ;
        RECT 50.630 172.965 50.890 173.285 ;
        RECT 51.610 172.945 51.750 173.985 ;
        RECT 55.750 173.285 55.890 174.325 ;
        RECT 55.690 172.965 55.950 173.285 ;
        RECT 50.170 172.625 50.430 172.945 ;
        RECT 51.550 172.625 51.810 172.945 ;
        RECT 56.210 172.605 56.350 183.165 ;
        RECT 57.990 182.145 58.250 182.465 ;
        RECT 58.050 180.425 58.190 182.145 ;
        RECT 58.970 180.765 59.110 190.985 ;
        RECT 59.370 190.305 59.630 190.625 ;
        RECT 59.430 189.265 59.570 190.305 ;
        RECT 59.370 188.945 59.630 189.265 ;
        RECT 60.810 187.905 60.950 190.985 ;
        RECT 63.510 190.305 63.770 190.625 ;
        RECT 63.570 188.585 63.710 190.305 ;
        RECT 63.510 188.265 63.770 188.585 ;
        RECT 60.750 187.585 61.010 187.905 ;
        RECT 62.590 187.585 62.850 187.905 ;
        RECT 58.910 180.445 59.170 180.765 ;
        RECT 61.210 180.445 61.470 180.765 ;
        RECT 57.990 180.165 58.250 180.425 ;
        RECT 57.990 180.105 58.650 180.165 ;
        RECT 58.050 180.025 58.650 180.105 ;
        RECT 57.990 179.425 58.250 179.745 ;
        RECT 58.050 178.725 58.190 179.425 ;
        RECT 57.990 178.405 58.250 178.725 ;
        RECT 46.950 172.285 47.210 172.605 ;
        RECT 49.250 172.285 49.510 172.605 ;
        RECT 49.710 172.285 49.970 172.605 ;
        RECT 56.150 172.285 56.410 172.605 ;
        RECT 46.490 171.945 46.750 172.265 ;
        RECT 46.550 171.585 46.690 171.945 ;
        RECT 57.990 171.605 58.250 171.925 ;
        RECT 44.650 171.265 44.910 171.585 ;
        RECT 46.490 171.265 46.750 171.585 ;
        RECT 47.410 171.265 47.670 171.585 ;
        RECT 44.190 170.080 44.450 170.225 ;
        RECT 44.180 169.710 44.460 170.080 ;
        RECT 44.190 161.405 44.450 161.725 ;
        RECT 44.250 158.665 44.390 161.405 ;
        RECT 44.190 158.345 44.450 158.665 ;
        RECT 44.710 153.905 44.850 171.265 ;
        RECT 46.950 163.105 47.210 163.425 ;
        RECT 47.010 162.405 47.150 163.105 ;
        RECT 46.950 162.085 47.210 162.405 ;
        RECT 46.950 161.065 47.210 161.385 ;
        RECT 46.490 160.385 46.750 160.705 ;
        RECT 45.110 159.025 45.370 159.345 ;
        RECT 45.170 158.665 45.310 159.025 ;
        RECT 46.550 159.005 46.690 160.385 ;
        RECT 46.490 158.685 46.750 159.005 ;
        RECT 45.110 158.345 45.370 158.665 ;
        RECT 45.570 158.345 45.830 158.665 ;
        RECT 45.630 156.285 45.770 158.345 ;
        RECT 46.550 158.325 46.690 158.685 ;
        RECT 46.490 158.005 46.750 158.325 ;
        RECT 46.030 157.665 46.290 157.985 ;
        RECT 45.570 155.965 45.830 156.285 ;
        RECT 45.110 153.925 45.370 154.245 ;
        RECT 44.650 153.585 44.910 153.905 ;
        RECT 43.730 153.245 43.990 153.565 ;
        RECT 44.190 153.245 44.450 153.565 ;
        RECT 44.250 150.845 44.390 153.245 ;
        RECT 44.650 152.565 44.910 152.885 ;
        RECT 44.190 150.525 44.450 150.845 ;
        RECT 44.710 147.105 44.850 152.565 ;
        RECT 44.650 146.785 44.910 147.105 ;
        RECT 44.650 136.585 44.910 136.905 ;
        RECT 44.190 134.885 44.450 135.205 ;
        RECT 41.890 133.865 42.150 134.185 ;
        RECT 43.270 133.865 43.530 134.185 ;
        RECT 42.350 133.185 42.610 133.505 ;
        RECT 42.410 132.485 42.550 133.185 ;
        RECT 42.350 132.165 42.610 132.485 ;
        RECT 40.970 131.825 41.230 132.145 ;
        RECT 42.810 131.145 43.070 131.465 ;
        RECT 43.730 131.145 43.990 131.465 ;
        RECT 41.420 129.590 41.700 129.960 ;
        RECT 41.490 129.425 41.630 129.590 ;
        RECT 41.430 129.105 41.690 129.425 ;
        RECT 42.870 126.365 43.010 131.145 ;
        RECT 43.790 129.765 43.930 131.145 ;
        RECT 43.730 129.445 43.990 129.765 ;
        RECT 42.810 126.045 43.070 126.365 ;
        RECT 42.870 123.645 43.010 126.045 ;
        RECT 42.810 123.325 43.070 123.645 ;
        RECT 40.510 122.985 40.770 123.305 ;
        RECT 40.050 120.265 40.310 120.585 ;
        RECT 40.570 118.885 40.710 122.985 ;
        RECT 42.870 120.925 43.010 123.325 ;
        RECT 42.810 120.605 43.070 120.925 ;
        RECT 43.790 120.585 43.930 129.445 ;
        RECT 43.730 120.265 43.990 120.585 ;
        RECT 40.510 118.565 40.770 118.885 ;
        RECT 43.790 118.545 43.930 120.265 ;
        RECT 43.730 118.225 43.990 118.545 ;
        RECT 34.530 112.785 34.790 113.105 ;
        RECT 37.750 112.785 38.010 113.105 ;
        RECT 38.730 112.765 38.870 118.145 ;
        RECT 39.590 117.885 39.850 118.205 ;
        RECT 44.250 115.145 44.390 134.885 ;
        RECT 44.710 134.525 44.850 136.585 ;
        RECT 44.650 134.205 44.910 134.525 ;
        RECT 44.710 131.465 44.850 134.205 ;
        RECT 44.650 131.145 44.910 131.465 ;
        RECT 45.170 124.325 45.310 153.925 ;
        RECT 45.570 150.185 45.830 150.505 ;
        RECT 45.630 146.085 45.770 150.185 ;
        RECT 45.570 145.765 45.830 146.085 ;
        RECT 46.090 145.405 46.230 157.665 ;
        RECT 47.010 156.285 47.150 161.065 ;
        RECT 46.950 155.965 47.210 156.285 ;
        RECT 46.490 154.945 46.750 155.265 ;
        RECT 46.550 152.885 46.690 154.945 ;
        RECT 46.490 152.565 46.750 152.885 ;
        RECT 46.490 150.865 46.750 151.185 ;
        RECT 46.550 148.320 46.690 150.865 ;
        RECT 47.010 149.825 47.150 155.965 ;
        RECT 46.950 149.505 47.210 149.825 ;
        RECT 46.480 147.950 46.760 148.320 ;
        RECT 46.490 147.805 46.750 147.950 ;
        RECT 46.030 145.085 46.290 145.405 ;
        RECT 47.470 145.065 47.610 171.265 ;
        RECT 49.910 170.730 51.790 171.100 ;
        RECT 58.050 170.225 58.190 171.605 ;
        RECT 51.080 169.710 51.360 170.080 ;
        RECT 57.990 169.905 58.250 170.225 ;
        RECT 51.150 169.545 51.290 169.710 ;
        RECT 50.630 169.225 50.890 169.545 ;
        RECT 51.090 169.225 51.350 169.545 ;
        RECT 49.250 168.885 49.510 169.205 ;
        RECT 48.790 166.165 49.050 166.485 ;
        RECT 47.870 165.825 48.130 166.145 ;
        RECT 47.930 156.285 48.070 165.825 ;
        RECT 48.850 163.765 48.990 166.165 ;
        RECT 49.310 165.125 49.450 168.885 ;
        RECT 50.690 166.145 50.830 169.225 ;
        RECT 53.390 168.885 53.650 169.205 ;
        RECT 52.010 168.545 52.270 168.865 ;
        RECT 52.070 167.845 52.210 168.545 ;
        RECT 52.010 167.525 52.270 167.845 ;
        RECT 52.470 167.525 52.730 167.845 ;
        RECT 52.010 166.165 52.270 166.485 ;
        RECT 50.630 165.825 50.890 166.145 ;
        RECT 49.910 165.290 51.790 165.660 ;
        RECT 49.250 164.805 49.510 165.125 ;
        RECT 52.070 163.845 52.210 166.165 ;
        RECT 52.530 164.445 52.670 167.525 ;
        RECT 53.450 167.165 53.590 168.885 ;
        RECT 58.510 167.505 58.650 180.025 ;
        RECT 60.750 179.765 61.010 180.085 ;
        RECT 60.810 175.325 60.950 179.765 ;
        RECT 60.750 175.005 61.010 175.325 ;
        RECT 59.370 174.325 59.630 174.645 ;
        RECT 59.430 173.285 59.570 174.325 ;
        RECT 59.370 172.965 59.630 173.285 ;
        RECT 60.290 170.245 60.550 170.565 ;
        RECT 58.450 167.185 58.710 167.505 ;
        RECT 53.390 166.845 53.650 167.165 ;
        RECT 57.070 166.505 57.330 166.825 ;
        RECT 57.130 165.125 57.270 166.505 ;
        RECT 57.070 164.805 57.330 165.125 ;
        RECT 52.470 164.125 52.730 164.445 ;
        RECT 58.510 164.105 58.650 167.185 ;
        RECT 48.790 163.445 49.050 163.765 ;
        RECT 51.610 163.705 52.210 163.845 ;
        RECT 48.330 163.105 48.590 163.425 ;
        RECT 48.390 162.405 48.530 163.105 ;
        RECT 48.330 162.085 48.590 162.405 ;
        RECT 48.850 159.765 48.990 163.445 ;
        RECT 51.610 161.725 51.750 163.705 ;
        RECT 54.760 163.590 55.040 163.960 ;
        RECT 56.150 163.785 56.410 164.105 ;
        RECT 58.450 163.785 58.710 164.105 ;
        RECT 52.010 163.105 52.270 163.425 ;
        RECT 52.070 161.725 52.210 163.105 ;
        RECT 51.550 161.405 51.810 161.725 ;
        RECT 52.010 161.405 52.270 161.725 ;
        RECT 51.610 161.125 51.750 161.405 ;
        RECT 51.610 160.985 52.210 161.125 ;
        RECT 49.250 160.385 49.510 160.705 ;
        RECT 48.390 159.625 48.990 159.765 ;
        RECT 48.390 158.665 48.530 159.625 ;
        RECT 49.310 158.915 49.450 160.385 ;
        RECT 49.910 159.850 51.790 160.220 ;
        RECT 49.710 158.915 49.970 159.005 ;
        RECT 49.310 158.775 49.970 158.915 ;
        RECT 49.710 158.685 49.970 158.775 ;
        RECT 52.070 158.665 52.210 160.985 ;
        RECT 54.830 159.200 54.970 163.590 ;
        RECT 56.210 162.405 56.350 163.785 ;
        RECT 58.450 163.105 58.710 163.425 ;
        RECT 59.830 163.105 60.090 163.425 ;
        RECT 56.150 162.085 56.410 162.405 ;
        RECT 57.530 161.745 57.790 162.065 ;
        RECT 54.760 158.830 55.040 159.200 ;
        RECT 54.770 158.685 55.030 158.830 ;
        RECT 48.330 158.345 48.590 158.665 ;
        RECT 50.630 158.520 50.890 158.665 ;
        RECT 50.620 158.150 50.900 158.520 ;
        RECT 52.010 158.345 52.270 158.665 ;
        RECT 47.870 155.965 48.130 156.285 ;
        RECT 53.850 155.965 54.110 156.285 ;
        RECT 47.930 152.545 48.070 155.965 ;
        RECT 49.910 154.410 51.790 154.780 ;
        RECT 48.330 152.905 48.590 153.225 ;
        RECT 47.870 152.225 48.130 152.545 ;
        RECT 47.930 150.415 48.070 152.225 ;
        RECT 48.390 151.185 48.530 152.905 ;
        RECT 53.910 151.525 54.050 155.965 ;
        RECT 57.590 155.945 57.730 161.745 ;
        RECT 57.990 160.725 58.250 161.045 ;
        RECT 57.530 155.625 57.790 155.945 ;
        RECT 54.310 155.285 54.570 155.605 ;
        RECT 54.370 151.525 54.510 155.285 ;
        RECT 54.770 155.125 55.030 155.265 ;
        RECT 54.770 154.985 55.890 155.125 ;
        RECT 54.770 154.945 55.030 154.985 ;
        RECT 55.750 153.565 55.890 154.985 ;
        RECT 55.690 153.245 55.950 153.565 ;
        RECT 49.250 151.205 49.510 151.525 ;
        RECT 53.850 151.205 54.110 151.525 ;
        RECT 54.310 151.205 54.570 151.525 ;
        RECT 48.330 150.865 48.590 151.185 ;
        RECT 48.790 150.525 49.050 150.845 ;
        RECT 47.930 150.275 48.530 150.415 ;
        RECT 48.390 148.465 48.530 150.275 ;
        RECT 48.330 148.145 48.590 148.465 ;
        RECT 48.850 147.640 48.990 150.525 ;
        RECT 49.310 147.785 49.450 151.205 ;
        RECT 58.050 151.040 58.190 160.725 ;
        RECT 58.510 156.625 58.650 163.105 ;
        RECT 59.890 161.725 60.030 163.105 ;
        RECT 59.830 161.405 60.090 161.725 ;
        RECT 59.830 160.560 60.090 160.705 ;
        RECT 59.820 160.190 60.100 160.560 ;
        RECT 58.910 157.665 59.170 157.985 ;
        RECT 58.450 156.305 58.710 156.625 ;
        RECT 58.450 155.285 58.710 155.605 ;
        RECT 58.510 153.565 58.650 155.285 ;
        RECT 58.450 153.245 58.710 153.565 ;
        RECT 58.450 152.795 58.710 152.885 ;
        RECT 58.970 152.795 59.110 157.665 ;
        RECT 59.830 155.625 60.090 155.945 ;
        RECT 59.890 153.905 60.030 155.625 ;
        RECT 59.830 153.585 60.090 153.905 ;
        RECT 60.350 153.225 60.490 170.245 ;
        RECT 60.810 166.485 60.950 175.005 ;
        RECT 61.270 174.985 61.410 180.445 ;
        RECT 62.650 178.045 62.790 187.585 ;
        RECT 64.030 183.565 64.170 196.425 ;
        RECT 64.430 195.745 64.690 196.065 ;
        RECT 64.490 194.615 64.630 195.745 ;
        RECT 64.910 195.210 66.790 195.580 ;
        RECT 64.890 194.615 65.150 194.705 ;
        RECT 64.490 194.475 65.150 194.615 ;
        RECT 64.890 194.385 65.150 194.475 ;
        RECT 66.730 193.935 66.990 194.025 ;
        RECT 67.250 193.935 67.390 196.765 ;
        RECT 67.650 194.385 67.910 194.705 ;
        RECT 66.730 193.795 67.390 193.935 ;
        RECT 66.730 193.705 66.990 193.795 ;
        RECT 67.190 193.255 67.450 193.345 ;
        RECT 67.710 193.255 67.850 194.385 ;
        RECT 67.190 193.115 67.850 193.255 ;
        RECT 67.190 193.025 67.450 193.115 ;
        RECT 67.650 190.645 67.910 190.965 ;
        RECT 64.910 189.770 66.790 190.140 ;
        RECT 64.910 184.330 66.790 184.700 ;
        RECT 63.570 183.425 64.170 183.565 ;
        RECT 67.710 183.485 67.850 190.645 ;
        RECT 68.170 188.925 68.310 199.145 ;
        RECT 69.090 195.045 69.230 201.525 ;
        RECT 72.310 199.805 72.450 202.885 ;
        RECT 80.530 202.205 80.790 202.525 ;
        RECT 75.470 201.525 75.730 201.845 ;
        RECT 76.390 201.525 76.650 201.845 ;
        RECT 75.530 200.145 75.670 201.525 ;
        RECT 76.450 200.485 76.590 201.525 ;
        RECT 76.390 200.165 76.650 200.485 ;
        RECT 72.710 199.825 72.970 200.145 ;
        RECT 75.470 199.825 75.730 200.145 ;
        RECT 78.690 199.885 78.950 200.145 ;
        RECT 76.910 199.825 78.950 199.885 ;
        RECT 71.330 199.485 71.590 199.805 ;
        RECT 72.250 199.715 72.510 199.805 ;
        RECT 71.850 199.575 72.510 199.715 ;
        RECT 69.950 197.105 70.210 197.425 ;
        RECT 69.490 196.425 69.750 196.745 ;
        RECT 69.030 194.725 69.290 195.045 ;
        RECT 69.550 193.685 69.690 196.425 ;
        RECT 70.010 193.685 70.150 197.105 ;
        RECT 71.390 197.085 71.530 199.485 ;
        RECT 71.850 197.085 71.990 199.575 ;
        RECT 72.250 199.485 72.510 199.575 ;
        RECT 72.770 199.125 72.910 199.825 ;
        RECT 76.910 199.745 78.890 199.825 ;
        RECT 80.590 199.805 80.730 202.205 ;
        RECT 81.910 201.185 82.170 201.505 ;
        RECT 76.910 199.465 77.050 199.745 ;
        RECT 80.530 199.485 80.790 199.805 ;
        RECT 80.990 199.485 81.250 199.805 ;
        RECT 72.710 198.805 72.970 199.125 ;
        RECT 76.380 198.950 76.660 199.320 ;
        RECT 76.850 199.145 77.110 199.465 ;
        RECT 78.230 199.145 78.490 199.465 ;
        RECT 81.050 199.320 81.190 199.485 ;
        RECT 76.390 198.805 76.650 198.950 ;
        RECT 71.330 196.765 71.590 197.085 ;
        RECT 71.790 196.765 72.050 197.085 ;
        RECT 72.250 196.765 72.510 197.085 ;
        RECT 69.490 193.365 69.750 193.685 ;
        RECT 69.950 193.365 70.210 193.685 ;
        RECT 68.570 191.325 68.830 191.645 ;
        RECT 68.110 188.605 68.370 188.925 ;
        RECT 68.630 188.325 68.770 191.325 ;
        RECT 69.550 191.305 69.690 193.365 ;
        RECT 69.490 190.985 69.750 191.305 ;
        RECT 68.170 188.185 68.770 188.325 ;
        RECT 68.170 183.485 68.310 188.185 ;
        RECT 68.570 183.505 68.830 183.825 ;
        RECT 62.590 177.725 62.850 178.045 ;
        RECT 62.650 177.560 62.790 177.725 ;
        RECT 62.580 177.190 62.860 177.560 ;
        RECT 61.210 174.665 61.470 174.985 ;
        RECT 63.050 172.965 63.310 173.285 ;
        RECT 63.110 172.800 63.250 172.965 ;
        RECT 63.040 172.430 63.320 172.800 ;
        RECT 62.130 171.945 62.390 172.265 ;
        RECT 60.750 166.165 61.010 166.485 ;
        RECT 62.190 164.445 62.330 171.945 ;
        RECT 62.590 168.545 62.850 168.865 ;
        RECT 62.650 167.505 62.790 168.545 ;
        RECT 62.590 167.185 62.850 167.505 ;
        RECT 62.130 164.125 62.390 164.445 ;
        RECT 61.670 163.445 61.930 163.765 ;
        RECT 60.750 153.585 61.010 153.905 ;
        RECT 59.370 153.080 59.630 153.225 ;
        RECT 58.450 152.655 59.110 152.795 ;
        RECT 59.360 152.965 59.640 153.080 ;
        RECT 59.360 152.825 60.030 152.965 ;
        RECT 60.290 152.905 60.550 153.225 ;
        RECT 59.360 152.710 59.640 152.825 ;
        RECT 58.450 152.565 58.710 152.655 ;
        RECT 57.980 150.670 58.260 151.040 ;
        RECT 52.010 149.505 52.270 149.825 ;
        RECT 49.910 148.970 51.790 149.340 ;
        RECT 50.620 147.950 50.900 148.320 ;
        RECT 50.690 147.785 50.830 147.950 ;
        RECT 48.780 147.270 49.060 147.640 ;
        RECT 49.250 147.465 49.510 147.785 ;
        RECT 50.170 147.465 50.430 147.785 ;
        RECT 50.630 147.465 50.890 147.785 ;
        RECT 51.550 147.640 51.810 147.785 ;
        RECT 52.070 147.695 52.210 149.505 ;
        RECT 57.530 148.145 57.790 148.465 ;
        RECT 52.470 147.695 52.730 147.785 ;
        RECT 47.870 145.765 48.130 146.085 ;
        RECT 47.410 144.745 47.670 145.065 ;
        RECT 45.570 144.065 45.830 144.385 ;
        RECT 47.410 144.065 47.670 144.385 ;
        RECT 45.630 142.345 45.770 144.065 ;
        RECT 46.950 142.365 47.210 142.685 ;
        RECT 45.570 142.025 45.830 142.345 ;
        RECT 47.010 139.625 47.150 142.365 ;
        RECT 46.950 139.305 47.210 139.625 ;
        RECT 46.490 136.925 46.750 137.245 ;
        RECT 46.550 134.525 46.690 136.925 ;
        RECT 47.010 134.525 47.150 139.305 ;
        RECT 46.490 134.205 46.750 134.525 ;
        RECT 46.950 134.205 47.210 134.525 ;
        RECT 46.550 130.785 46.690 134.205 ;
        RECT 46.950 133.525 47.210 133.845 ;
        RECT 47.010 131.465 47.150 133.525 ;
        RECT 46.950 131.145 47.210 131.465 ;
        RECT 46.490 130.465 46.750 130.785 ;
        RECT 47.470 127.045 47.610 144.065 ;
        RECT 47.930 136.565 48.070 145.765 ;
        RECT 48.330 145.315 48.590 145.405 ;
        RECT 49.310 145.315 49.450 147.465 ;
        RECT 50.230 146.085 50.370 147.465 ;
        RECT 51.540 147.270 51.820 147.640 ;
        RECT 52.070 147.555 52.730 147.695 ;
        RECT 52.470 147.465 52.730 147.555 ;
        RECT 50.170 145.765 50.430 146.085 ;
        RECT 51.610 145.405 51.750 147.270 ;
        RECT 52.470 146.785 52.730 147.105 ;
        RECT 52.530 146.085 52.670 146.785 ;
        RECT 52.470 145.765 52.730 146.085 ;
        RECT 48.330 145.175 49.450 145.315 ;
        RECT 48.330 145.085 48.590 145.175 ;
        RECT 49.710 145.085 49.970 145.405 ;
        RECT 51.550 145.315 51.810 145.405 ;
        RECT 51.550 145.175 52.210 145.315 ;
        RECT 51.550 145.085 51.810 145.175 ;
        RECT 48.390 137.925 48.530 145.085 ;
        RECT 49.770 144.295 49.910 145.085 ;
        RECT 49.310 144.155 49.910 144.295 ;
        RECT 49.310 142.345 49.450 144.155 ;
        RECT 49.910 143.530 51.790 143.900 ;
        RECT 49.250 142.025 49.510 142.345 ;
        RECT 48.790 141.345 49.050 141.665 ;
        RECT 48.850 139.625 48.990 141.345 ;
        RECT 49.310 140.645 49.450 142.025 ;
        RECT 51.550 141.685 51.810 142.005 ;
        RECT 51.610 140.645 51.750 141.685 ;
        RECT 49.250 140.325 49.510 140.645 ;
        RECT 51.550 140.325 51.810 140.645 ;
        RECT 48.790 139.305 49.050 139.625 ;
        RECT 48.330 137.605 48.590 137.925 ;
        RECT 48.390 136.905 48.530 137.605 ;
        RECT 48.330 136.585 48.590 136.905 ;
        RECT 47.870 136.245 48.130 136.565 ;
        RECT 47.930 135.205 48.070 136.245 ;
        RECT 47.870 134.885 48.130 135.205 ;
        RECT 47.930 132.145 48.070 134.885 ;
        RECT 48.850 134.865 48.990 139.305 ;
        RECT 49.910 138.090 51.790 138.460 ;
        RECT 52.070 137.245 52.210 145.175 ;
        RECT 52.470 144.405 52.730 144.725 ;
        RECT 52.010 136.925 52.270 137.245 ;
        RECT 52.010 135.905 52.270 136.225 ;
        RECT 48.790 134.545 49.050 134.865 ;
        RECT 49.910 132.650 51.790 133.020 ;
        RECT 47.870 131.825 48.130 132.145 ;
        RECT 52.070 131.125 52.210 135.905 ;
        RECT 52.010 130.805 52.270 131.125 ;
        RECT 48.790 127.745 49.050 128.065 ;
        RECT 52.010 127.745 52.270 128.065 ;
        RECT 47.410 126.725 47.670 127.045 ;
        RECT 48.850 126.025 48.990 127.745 ;
        RECT 49.910 127.210 51.790 127.580 ;
        RECT 48.790 125.705 49.050 126.025 ;
        RECT 45.110 124.005 45.370 124.325 ;
        RECT 45.110 122.985 45.370 123.305 ;
        RECT 46.490 122.985 46.750 123.305 ;
        RECT 47.870 122.985 48.130 123.305 ;
        RECT 44.650 119.925 44.910 120.245 ;
        RECT 44.710 118.885 44.850 119.925 ;
        RECT 44.650 118.565 44.910 118.885 ;
        RECT 45.170 118.205 45.310 122.985 ;
        RECT 46.550 122.625 46.690 122.985 ;
        RECT 46.490 122.305 46.750 122.625 ;
        RECT 47.930 121.685 48.070 122.985 ;
        RECT 48.850 122.965 48.990 125.705 ;
        RECT 49.250 125.025 49.510 125.345 ;
        RECT 49.310 123.645 49.450 125.025 ;
        RECT 49.250 123.325 49.510 123.645 ;
        RECT 48.790 122.645 49.050 122.965 ;
        RECT 47.470 121.605 48.070 121.685 ;
        RECT 47.410 121.545 48.070 121.605 ;
        RECT 47.410 121.285 47.670 121.545 ;
        RECT 45.110 117.885 45.370 118.205 ;
        RECT 47.930 117.865 48.070 121.545 ;
        RECT 48.850 120.585 48.990 122.645 ;
        RECT 49.310 121.605 49.450 123.325 ;
        RECT 52.070 123.305 52.210 127.745 ;
        RECT 52.010 122.985 52.270 123.305 ;
        RECT 52.010 122.305 52.270 122.625 ;
        RECT 49.910 121.770 51.790 122.140 ;
        RECT 49.250 121.285 49.510 121.605 ;
        RECT 48.330 120.265 48.590 120.585 ;
        RECT 48.790 120.265 49.050 120.585 ;
        RECT 48.390 118.885 48.530 120.265 ;
        RECT 48.330 118.565 48.590 118.885 ;
        RECT 47.870 117.545 48.130 117.865 ;
        RECT 44.190 114.825 44.450 115.145 ;
        RECT 46.950 112.785 47.210 113.105 ;
        RECT 38.670 112.445 38.930 112.765 ;
        RECT 37.750 112.105 38.010 112.425 ;
        RECT 45.570 112.105 45.830 112.425 ;
        RECT 36.370 111.425 36.630 111.745 ;
        RECT 36.430 110.045 36.570 111.425 ;
        RECT 37.810 110.045 37.950 112.105 ;
        RECT 40.510 111.425 40.770 111.745 ;
        RECT 34.530 109.725 34.790 110.045 ;
        RECT 36.370 109.725 36.630 110.045 ;
        RECT 37.750 109.725 38.010 110.045 ;
        RECT 29.930 109.045 30.190 109.365 ;
        RECT 34.590 95.885 34.730 109.725 ;
        RECT 34.910 108.170 36.790 108.540 ;
        RECT 37.810 107.325 37.950 109.725 ;
        RECT 37.750 107.005 38.010 107.325 ;
        RECT 40.570 106.985 40.710 111.425 ;
        RECT 41.890 108.705 42.150 109.025 ;
        RECT 41.950 107.325 42.090 108.705 ;
        RECT 41.890 107.005 42.150 107.325 ;
        RECT 40.050 106.665 40.310 106.985 ;
        RECT 40.510 106.665 40.770 106.985 ;
        RECT 40.110 95.885 40.250 106.665 ;
        RECT 45.630 95.885 45.770 112.105 ;
        RECT 47.010 110.725 47.150 112.785 ;
        RECT 48.850 112.425 48.990 120.265 ;
        RECT 49.310 118.885 49.450 121.285 ;
        RECT 49.250 118.565 49.510 118.885 ;
        RECT 52.070 118.205 52.210 122.305 ;
        RECT 52.010 117.885 52.270 118.205 ;
        RECT 49.910 116.330 51.790 116.700 ;
        RECT 49.250 114.145 49.510 114.465 ;
        RECT 49.310 113.105 49.450 114.145 ;
        RECT 49.250 112.785 49.510 113.105 ;
        RECT 52.530 112.765 52.670 144.405 ;
        RECT 55.230 142.025 55.490 142.345 ;
        RECT 55.290 140.645 55.430 142.025 ;
        RECT 57.590 142.005 57.730 148.145 ;
        RECT 58.050 147.785 58.190 150.670 ;
        RECT 58.510 148.125 58.650 152.565 ;
        RECT 59.370 150.185 59.630 150.505 ;
        RECT 58.910 149.505 59.170 149.825 ;
        RECT 58.450 147.805 58.710 148.125 ;
        RECT 57.990 147.465 58.250 147.785 ;
        RECT 57.530 141.685 57.790 142.005 ;
        RECT 55.230 140.325 55.490 140.645 ;
        RECT 57.590 140.305 57.730 141.685 ;
        RECT 58.510 141.575 58.650 147.805 ;
        RECT 58.970 147.795 59.110 149.505 ;
        RECT 58.910 147.475 59.170 147.795 ;
        RECT 58.970 146.085 59.110 147.475 ;
        RECT 58.910 145.765 59.170 146.085 ;
        RECT 59.430 145.065 59.570 150.185 ;
        RECT 59.890 148.465 60.030 152.825 ;
        RECT 59.830 148.145 60.090 148.465 ;
        RECT 60.350 148.205 60.490 152.905 ;
        RECT 60.810 150.505 60.950 153.585 ;
        RECT 61.210 152.905 61.470 153.225 ;
        RECT 60.750 150.185 61.010 150.505 ;
        RECT 61.270 148.805 61.410 152.905 ;
        RECT 61.210 148.485 61.470 148.805 ;
        RECT 60.350 148.065 60.950 148.205 ;
        RECT 61.270 148.125 61.410 148.485 ;
        RECT 59.830 145.085 60.090 145.405 ;
        RECT 59.370 144.745 59.630 145.065 ;
        RECT 58.910 142.025 59.170 142.345 ;
        RECT 58.970 141.665 59.110 142.025 ;
        RECT 58.910 141.575 59.170 141.665 ;
        RECT 58.050 141.435 59.170 141.575 ;
        RECT 57.530 139.985 57.790 140.305 ;
        RECT 58.050 139.965 58.190 141.435 ;
        RECT 58.910 141.345 59.170 141.435 ;
        RECT 52.930 139.645 53.190 139.965 ;
        RECT 57.990 139.645 58.250 139.965 ;
        RECT 52.990 136.905 53.130 139.645 ;
        RECT 59.430 139.285 59.570 144.745 ;
        RECT 59.890 142.345 60.030 145.085 ;
        RECT 60.290 142.365 60.550 142.685 ;
        RECT 59.830 142.025 60.090 142.345 ;
        RECT 59.890 140.645 60.030 142.025 ;
        RECT 59.830 140.325 60.090 140.645 ;
        RECT 59.370 138.965 59.630 139.285 ;
        RECT 52.930 136.585 53.190 136.905 ;
        RECT 58.910 136.585 59.170 136.905 ;
        RECT 54.770 136.245 55.030 136.565 ;
        RECT 54.830 134.185 54.970 136.245 ;
        RECT 58.450 134.885 58.710 135.205 ;
        RECT 54.770 133.865 55.030 134.185 ;
        RECT 54.830 130.525 54.970 133.865 ;
        RECT 55.690 133.185 55.950 133.505 ;
        RECT 55.750 131.805 55.890 133.185 ;
        RECT 55.690 131.485 55.950 131.805 ;
        RECT 55.230 130.525 55.490 130.785 ;
        RECT 54.830 130.465 55.490 130.525 ;
        RECT 54.830 130.385 55.430 130.465 ;
        RECT 54.830 129.765 54.970 130.385 ;
        RECT 54.770 129.445 55.030 129.765 ;
        RECT 57.990 129.105 58.250 129.425 ;
        RECT 58.050 127.045 58.190 129.105 ;
        RECT 57.990 126.725 58.250 127.045 ;
        RECT 58.510 126.025 58.650 134.885 ;
        RECT 58.970 126.365 59.110 136.585 ;
        RECT 59.430 134.185 59.570 138.965 ;
        RECT 60.350 134.185 60.490 142.365 ;
        RECT 60.810 142.345 60.950 148.065 ;
        RECT 61.210 147.805 61.470 148.125 ;
        RECT 61.730 147.785 61.870 163.445 ;
        RECT 62.190 150.925 62.330 164.125 ;
        RECT 62.650 164.105 62.790 167.185 ;
        RECT 63.050 166.165 63.310 166.485 ;
        RECT 62.590 163.785 62.850 164.105 ;
        RECT 63.110 161.725 63.250 166.165 ;
        RECT 63.050 161.405 63.310 161.725 ;
        RECT 63.570 159.345 63.710 183.425 ;
        RECT 67.650 183.165 67.910 183.485 ;
        RECT 68.110 183.165 68.370 183.485 ;
        RECT 63.970 182.825 64.230 183.145 ;
        RECT 66.730 182.825 66.990 183.145 ;
        RECT 64.030 178.045 64.170 182.825 ;
        RECT 64.430 180.445 64.690 180.765 ;
        RECT 63.970 177.725 64.230 178.045 ;
        RECT 64.030 175.325 64.170 177.725 ;
        RECT 64.490 177.705 64.630 180.445 ;
        RECT 66.790 180.085 66.930 182.825 ;
        RECT 67.710 181.105 67.850 183.165 ;
        RECT 68.170 181.445 68.310 183.165 ;
        RECT 68.110 181.125 68.370 181.445 ;
        RECT 67.650 180.785 67.910 181.105 ;
        RECT 67.650 180.105 67.910 180.425 ;
        RECT 66.730 179.995 66.990 180.085 ;
        RECT 66.730 179.855 67.390 179.995 ;
        RECT 66.730 179.765 66.990 179.855 ;
        RECT 64.910 178.890 66.790 179.260 ;
        RECT 66.730 178.405 66.990 178.725 ;
        RECT 66.260 177.870 66.540 178.240 ;
        RECT 66.270 177.725 66.530 177.870 ;
        RECT 64.430 177.385 64.690 177.705 ;
        RECT 65.350 177.275 65.610 177.365 ;
        RECT 65.350 177.135 66.010 177.275 ;
        RECT 65.350 177.045 65.610 177.135 ;
        RECT 64.890 176.705 65.150 177.025 ;
        RECT 63.970 175.005 64.230 175.325 ;
        RECT 64.030 172.605 64.170 175.005 ;
        RECT 64.430 174.665 64.690 174.985 ;
        RECT 64.950 174.840 65.090 176.705 ;
        RECT 65.350 175.685 65.610 176.005 ;
        RECT 64.490 172.605 64.630 174.665 ;
        RECT 64.880 174.470 65.160 174.840 ;
        RECT 65.410 174.305 65.550 175.685 ;
        RECT 65.870 175.405 66.010 177.135 ;
        RECT 66.790 176.005 66.930 178.405 ;
        RECT 67.250 178.240 67.390 179.855 ;
        RECT 67.710 178.725 67.850 180.105 ;
        RECT 68.170 180.085 68.310 181.125 ;
        RECT 68.630 180.765 68.770 183.505 ;
        RECT 69.550 183.145 69.690 190.985 ;
        RECT 70.010 188.585 70.150 193.365 ;
        RECT 70.410 193.025 70.670 193.345 ;
        RECT 69.950 188.265 70.210 188.585 ;
        RECT 69.490 182.825 69.750 183.145 ;
        RECT 68.570 180.445 68.830 180.765 ;
        RECT 68.110 179.765 68.370 180.085 ;
        RECT 67.650 178.405 67.910 178.725 ;
        RECT 68.170 178.385 68.310 179.765 ;
        RECT 68.570 179.425 68.830 179.745 ;
        RECT 67.180 177.870 67.460 178.240 ;
        RECT 68.110 178.065 68.370 178.385 ;
        RECT 68.170 177.705 68.310 178.065 ;
        RECT 68.110 177.385 68.370 177.705 ;
        RECT 68.110 176.705 68.370 177.025 ;
        RECT 66.730 175.685 66.990 176.005 ;
        RECT 66.260 175.405 66.540 175.520 ;
        RECT 65.870 175.265 66.540 175.405 ;
        RECT 66.260 175.150 66.540 175.265 ;
        RECT 66.330 174.985 66.470 175.150 ;
        RECT 66.270 174.665 66.530 174.985 ;
        RECT 67.650 174.665 67.910 174.985 ;
        RECT 65.350 173.985 65.610 174.305 ;
        RECT 64.910 173.450 66.790 173.820 ;
        RECT 63.970 172.285 64.230 172.605 ;
        RECT 64.430 172.285 64.690 172.605 ;
        RECT 64.430 169.565 64.690 169.885 ;
        RECT 64.490 165.125 64.630 169.565 ;
        RECT 67.190 168.885 67.450 169.205 ;
        RECT 64.910 168.010 66.790 168.380 ;
        RECT 67.250 167.505 67.390 168.885 ;
        RECT 67.190 167.185 67.450 167.505 ;
        RECT 67.710 167.165 67.850 174.665 ;
        RECT 67.650 166.845 67.910 167.165 ;
        RECT 67.190 166.505 67.450 166.825 ;
        RECT 64.430 164.805 64.690 165.125 ;
        RECT 67.250 164.105 67.390 166.505 ;
        RECT 64.430 163.785 64.690 164.105 ;
        RECT 67.190 163.785 67.450 164.105 ;
        RECT 64.490 161.240 64.630 163.785 ;
        RECT 64.910 162.570 66.790 162.940 ;
        RECT 67.250 162.405 67.390 163.785 ;
        RECT 67.190 162.085 67.450 162.405 ;
        RECT 67.190 161.405 67.450 161.725 ;
        RECT 67.250 161.240 67.390 161.405 ;
        RECT 64.420 160.870 64.700 161.240 ;
        RECT 67.180 160.870 67.460 161.240 ;
        RECT 63.970 160.385 64.230 160.705 ;
        RECT 67.190 160.385 67.450 160.705 ;
        RECT 64.030 159.685 64.170 160.385 ;
        RECT 63.970 159.365 64.230 159.685 ;
        RECT 66.730 159.365 66.990 159.685 ;
        RECT 63.510 159.085 63.770 159.345 ;
        RECT 63.510 159.025 64.170 159.085 ;
        RECT 63.570 158.945 64.170 159.025 ;
        RECT 63.510 158.005 63.770 158.325 ;
        RECT 63.570 156.480 63.710 158.005 ;
        RECT 63.050 155.965 63.310 156.285 ;
        RECT 63.500 156.110 63.780 156.480 ;
        RECT 64.030 156.285 64.170 158.945 ;
        RECT 66.790 157.985 66.930 159.365 ;
        RECT 67.250 158.665 67.390 160.385 ;
        RECT 67.190 158.345 67.450 158.665 ;
        RECT 66.730 157.665 66.990 157.985 ;
        RECT 64.910 157.130 66.790 157.500 ;
        RECT 67.710 156.625 67.850 166.845 ;
        RECT 67.650 156.535 67.910 156.625 ;
        RECT 67.250 156.395 67.910 156.535 ;
        RECT 63.970 155.965 64.230 156.285 ;
        RECT 63.110 154.245 63.250 155.965 ;
        RECT 66.720 155.430 67.000 155.800 ;
        RECT 66.790 155.265 66.930 155.430 ;
        RECT 66.730 154.945 66.990 155.265 ;
        RECT 63.050 153.925 63.310 154.245 ;
        RECT 67.250 153.565 67.390 156.395 ;
        RECT 67.650 156.305 67.910 156.395 ;
        RECT 68.170 155.855 68.310 176.705 ;
        RECT 68.630 156.285 68.770 179.425 ;
        RECT 69.490 177.560 69.750 177.705 ;
        RECT 69.030 177.045 69.290 177.365 ;
        RECT 69.480 177.190 69.760 177.560 ;
        RECT 69.090 166.825 69.230 177.045 ;
        RECT 69.480 175.150 69.760 175.520 ;
        RECT 69.550 174.985 69.690 175.150 ;
        RECT 69.490 174.665 69.750 174.985 ;
        RECT 69.550 169.545 69.690 174.665 ;
        RECT 69.950 173.985 70.210 174.305 ;
        RECT 69.490 169.225 69.750 169.545 ;
        RECT 69.550 167.165 69.690 169.225 ;
        RECT 69.490 166.845 69.750 167.165 ;
        RECT 69.030 166.505 69.290 166.825 ;
        RECT 69.550 164.445 69.690 166.845 ;
        RECT 69.490 164.125 69.750 164.445 ;
        RECT 69.490 162.085 69.750 162.405 ;
        RECT 69.550 160.705 69.690 162.085 ;
        RECT 69.030 160.385 69.290 160.705 ;
        RECT 69.490 160.385 69.750 160.705 ;
        RECT 68.570 155.965 68.830 156.285 ;
        RECT 67.710 155.715 68.310 155.855 ;
        RECT 67.190 153.245 67.450 153.565 ;
        RECT 64.910 151.690 66.790 152.060 ;
        RECT 62.190 150.785 62.790 150.925 ;
        RECT 63.050 150.865 63.310 151.185 ;
        RECT 62.130 149.845 62.390 150.165 ;
        RECT 61.670 147.465 61.930 147.785 ;
        RECT 61.210 142.705 61.470 143.025 ;
        RECT 60.750 142.255 61.010 142.345 ;
        RECT 61.270 142.255 61.410 142.705 ;
        RECT 61.730 142.345 61.870 147.465 ;
        RECT 60.750 142.115 61.410 142.255 ;
        RECT 60.750 142.025 61.010 142.115 ;
        RECT 61.270 140.305 61.410 142.115 ;
        RECT 61.670 142.025 61.930 142.345 ;
        RECT 61.210 139.985 61.470 140.305 ;
        RECT 60.750 139.645 61.010 139.965 ;
        RECT 59.370 133.865 59.630 134.185 ;
        RECT 60.290 133.865 60.550 134.185 ;
        RECT 59.430 131.805 59.570 133.865 ;
        RECT 59.370 131.485 59.630 131.805 ;
        RECT 60.350 131.125 60.490 133.865 ;
        RECT 60.810 133.505 60.950 139.645 ;
        RECT 60.750 133.185 61.010 133.505 ;
        RECT 60.810 131.805 60.950 133.185 ;
        RECT 60.750 131.485 61.010 131.805 ;
        RECT 60.290 130.805 60.550 131.125 ;
        RECT 60.350 129.085 60.490 130.805 ;
        RECT 60.290 128.765 60.550 129.085 ;
        RECT 60.750 128.765 61.010 129.085 ;
        RECT 58.910 126.045 59.170 126.365 ;
        RECT 58.450 125.705 58.710 126.025 ;
        RECT 58.970 123.645 59.110 126.045 ;
        RECT 60.350 123.645 60.490 128.765 ;
        RECT 60.810 127.045 60.950 128.765 ;
        RECT 60.750 126.725 61.010 127.045 ;
        RECT 58.910 123.325 59.170 123.645 ;
        RECT 60.290 123.325 60.550 123.645 ;
        RECT 54.310 122.305 54.570 122.625 ;
        RECT 54.370 120.245 54.510 122.305 ;
        RECT 57.990 120.605 58.250 120.925 ;
        RECT 54.310 119.925 54.570 120.245 ;
        RECT 58.050 118.885 58.190 120.605 ;
        RECT 57.990 118.565 58.250 118.885 ;
        RECT 58.450 115.165 58.710 115.485 ;
        RECT 52.470 112.445 52.730 112.765 ;
        RECT 48.790 112.105 49.050 112.425 ;
        RECT 56.610 112.105 56.870 112.425 ;
        RECT 46.950 110.405 47.210 110.725 ;
        RECT 48.330 109.045 48.590 109.365 ;
        RECT 48.390 106.825 48.530 109.045 ;
        RECT 48.850 107.325 48.990 112.105 ;
        RECT 53.390 111.425 53.650 111.745 ;
        RECT 49.910 110.890 51.790 111.260 ;
        RECT 53.450 110.045 53.590 111.425 ;
        RECT 53.390 109.725 53.650 110.045 ;
        RECT 53.390 109.045 53.650 109.365 ;
        RECT 53.450 108.005 53.590 109.045 ;
        RECT 53.850 108.705 54.110 109.025 ;
        RECT 53.390 107.685 53.650 108.005 ;
        RECT 53.910 107.325 54.050 108.705 ;
        RECT 48.790 107.005 49.050 107.325 ;
        RECT 53.850 107.005 54.110 107.325 ;
        RECT 48.390 106.685 48.990 106.825 ;
        RECT 12.440 93.885 12.720 95.885 ;
        RECT 17.960 93.885 18.240 95.885 ;
        RECT 23.480 93.885 23.760 95.885 ;
        RECT 29.000 93.885 29.280 95.885 ;
        RECT 34.520 93.885 34.800 95.885 ;
        RECT 40.040 93.885 40.320 95.885 ;
        RECT 45.560 93.885 45.840 95.885 ;
        RECT 48.850 95.845 48.990 106.685 ;
        RECT 49.910 105.450 51.790 105.820 ;
        RECT 50.690 96.385 51.290 96.525 ;
        RECT 50.690 95.845 50.830 96.385 ;
        RECT 51.150 95.885 51.290 96.385 ;
        RECT 56.670 95.885 56.810 112.105 ;
        RECT 58.510 109.365 58.650 115.165 ;
        RECT 58.970 115.145 59.110 123.325 ;
        RECT 60.350 120.925 60.490 123.325 ;
        RECT 60.290 120.605 60.550 120.925 ;
        RECT 58.910 114.825 59.170 115.145 ;
        RECT 59.820 113.270 60.100 113.640 ;
        RECT 58.910 112.785 59.170 113.105 ;
        RECT 58.450 109.045 58.710 109.365 ;
        RECT 58.510 107.325 58.650 109.045 ;
        RECT 58.970 108.005 59.110 112.785 ;
        RECT 59.890 109.705 60.030 113.270 ;
        RECT 60.350 112.425 60.490 120.605 ;
        RECT 62.190 113.445 62.330 149.845 ;
        RECT 62.650 120.585 62.790 150.785 ;
        RECT 63.110 148.805 63.250 150.865 ;
        RECT 65.350 150.185 65.610 150.505 ;
        RECT 65.410 148.805 65.550 150.185 ;
        RECT 63.050 148.485 63.310 148.805 ;
        RECT 65.350 148.485 65.610 148.805 ;
        RECT 66.730 148.145 66.990 148.465 ;
        RECT 64.430 147.465 64.690 147.785 ;
        RECT 66.790 147.640 66.930 148.145 ;
        RECT 64.490 146.085 64.630 147.465 ;
        RECT 66.720 147.270 67.000 147.640 ;
        RECT 66.730 147.125 66.990 147.270 ;
        RECT 64.910 146.250 66.790 146.620 ;
        RECT 64.430 145.765 64.690 146.085 ;
        RECT 65.350 145.425 65.610 145.745 ;
        RECT 65.410 143.365 65.550 145.425 ;
        RECT 65.350 143.045 65.610 143.365 ;
        RECT 63.510 142.025 63.770 142.345 ;
        RECT 63.570 136.905 63.710 142.025 ;
        RECT 64.430 141.685 64.690 142.005 ;
        RECT 64.490 140.645 64.630 141.685 ;
        RECT 64.910 140.810 66.790 141.180 ;
        RECT 64.430 140.325 64.690 140.645 ;
        RECT 64.430 137.265 64.690 137.585 ;
        RECT 63.510 136.585 63.770 136.905 ;
        RECT 63.510 135.905 63.770 136.225 ;
        RECT 63.570 134.865 63.710 135.905 ;
        RECT 63.510 134.545 63.770 134.865 ;
        RECT 64.490 133.505 64.630 137.265 ;
        RECT 64.910 135.370 66.790 135.740 ;
        RECT 66.270 134.205 66.530 134.525 ;
        RECT 64.430 133.185 64.690 133.505 ;
        RECT 66.330 132.145 66.470 134.205 ;
        RECT 66.270 131.825 66.530 132.145 ;
        RECT 67.250 131.805 67.390 153.245 ;
        RECT 67.710 136.905 67.850 155.715 ;
        RECT 68.100 154.750 68.380 155.120 ;
        RECT 68.170 148.125 68.310 154.750 ;
        RECT 68.630 154.245 68.770 155.965 ;
        RECT 68.570 153.925 68.830 154.245 ;
        RECT 68.570 150.185 68.830 150.505 ;
        RECT 68.110 147.805 68.370 148.125 ;
        RECT 68.110 147.125 68.370 147.445 ;
        RECT 68.170 146.085 68.310 147.125 ;
        RECT 68.110 145.765 68.370 146.085 ;
        RECT 68.630 145.405 68.770 150.185 ;
        RECT 69.090 147.785 69.230 160.385 ;
        RECT 69.490 158.685 69.750 159.005 ;
        RECT 69.030 147.465 69.290 147.785 ;
        RECT 68.570 145.085 68.830 145.405 ;
        RECT 68.110 144.745 68.370 145.065 ;
        RECT 68.170 143.365 68.310 144.745 ;
        RECT 68.110 143.045 68.370 143.365 ;
        RECT 69.550 136.905 69.690 158.685 ;
        RECT 70.010 150.505 70.150 173.985 ;
        RECT 70.470 166.485 70.610 193.025 ;
        RECT 71.390 192.325 71.530 196.765 ;
        RECT 71.850 194.025 71.990 196.765 ;
        RECT 72.310 196.405 72.450 196.765 ;
        RECT 72.250 196.085 72.510 196.405 ;
        RECT 72.310 194.365 72.450 196.085 ;
        RECT 72.770 196.065 72.910 198.805 ;
        RECT 72.710 195.745 72.970 196.065 ;
        RECT 73.170 195.745 73.430 196.065 ;
        RECT 72.250 194.045 72.510 194.365 ;
        RECT 71.790 193.705 72.050 194.025 ;
        RECT 71.330 192.005 71.590 192.325 ;
        RECT 71.390 183.825 71.530 192.005 ;
        RECT 71.850 191.305 71.990 193.705 ;
        RECT 72.710 193.025 72.970 193.345 ;
        RECT 72.770 191.305 72.910 193.025 ;
        RECT 73.230 192.325 73.370 195.745 ;
        RECT 76.910 195.045 77.050 199.145 ;
        RECT 76.850 194.725 77.110 195.045 ;
        RECT 78.290 194.705 78.430 199.145 ;
        RECT 79.150 198.805 79.410 199.125 ;
        RECT 80.980 198.950 81.260 199.320 ;
        RECT 79.210 196.405 79.350 198.805 ;
        RECT 79.910 197.930 81.790 198.300 ;
        RECT 81.970 197.085 82.110 201.185 ;
        RECT 94.910 200.650 96.790 201.020 ;
        RECT 86.050 199.485 86.310 199.805 ;
        RECT 82.370 198.465 82.630 198.785 ;
        RECT 82.430 197.425 82.570 198.465 ;
        RECT 82.370 197.105 82.630 197.425 ;
        RECT 81.910 196.765 82.170 197.085 ;
        RECT 79.150 196.085 79.410 196.405 ;
        RECT 75.010 194.385 75.270 194.705 ;
        RECT 78.230 194.385 78.490 194.705 ;
        RECT 73.170 192.005 73.430 192.325 ;
        RECT 75.070 191.985 75.210 194.385 ;
        RECT 76.390 194.045 76.650 194.365 ;
        RECT 76.450 192.325 76.590 194.045 ;
        RECT 81.970 194.025 82.110 196.765 ;
        RECT 86.110 195.045 86.250 199.485 ;
        RECT 109.910 197.930 111.790 198.300 ;
        RECT 99.390 197.105 99.650 197.425 ;
        RECT 97.550 196.085 97.810 196.405 ;
        RECT 94.910 195.210 96.790 195.580 ;
        RECT 97.610 195.045 97.750 196.085 ;
        RECT 86.050 194.725 86.310 195.045 ;
        RECT 97.550 194.725 97.810 195.045 ;
        RECT 86.110 194.365 86.250 194.725 ;
        RECT 82.370 194.045 82.630 194.365 ;
        RECT 86.050 194.045 86.310 194.365 ;
        RECT 81.910 193.705 82.170 194.025 ;
        RECT 79.910 192.490 81.790 192.860 ;
        RECT 76.390 192.005 76.650 192.325 ;
        RECT 75.010 191.665 75.270 191.985 ;
        RECT 71.790 190.985 72.050 191.305 ;
        RECT 72.710 190.985 72.970 191.305 ;
        RECT 77.310 190.305 77.570 190.625 ;
        RECT 77.370 189.605 77.510 190.305 ;
        RECT 82.430 189.605 82.570 194.045 ;
        RECT 86.510 193.705 86.770 194.025 ;
        RECT 88.810 193.705 89.070 194.025 ;
        RECT 98.930 193.705 99.190 194.025 ;
        RECT 84.210 193.025 84.470 193.345 ;
        RECT 84.270 191.645 84.410 193.025 ;
        RECT 84.210 191.325 84.470 191.645 ;
        RECT 86.570 191.305 86.710 193.705 ;
        RECT 88.870 192.325 89.010 193.705 ;
        RECT 93.870 193.025 94.130 193.345 ;
        RECT 88.810 192.005 89.070 192.325 ;
        RECT 93.410 191.325 93.670 191.645 ;
        RECT 86.510 190.985 86.770 191.305 ;
        RECT 83.290 190.645 83.550 190.965 ;
        RECT 83.350 189.605 83.490 190.645 ;
        RECT 77.310 189.285 77.570 189.605 ;
        RECT 82.370 189.285 82.630 189.605 ;
        RECT 83.290 189.285 83.550 189.605 ;
        RECT 75.470 188.945 75.730 189.265 ;
        RECT 75.530 185.185 75.670 188.945 ;
        RECT 75.470 184.865 75.730 185.185 ;
        RECT 71.330 183.505 71.590 183.825 ;
        RECT 73.170 183.165 73.430 183.485 ;
        RECT 71.330 182.825 71.590 183.145 ;
        RECT 70.870 179.765 71.130 180.085 ;
        RECT 70.930 176.005 71.070 179.765 ;
        RECT 71.390 178.045 71.530 182.825 ;
        RECT 72.250 182.485 72.510 182.805 ;
        RECT 72.310 181.445 72.450 182.485 ;
        RECT 72.710 182.145 72.970 182.465 ;
        RECT 72.250 181.125 72.510 181.445 ;
        RECT 72.250 180.105 72.510 180.425 ;
        RECT 72.310 178.045 72.450 180.105 ;
        RECT 72.770 178.385 72.910 182.145 ;
        RECT 73.230 181.445 73.370 183.165 ;
        RECT 75.530 183.145 75.670 184.865 ;
        RECT 75.470 182.825 75.730 183.145 ;
        RECT 73.170 181.125 73.430 181.445 ;
        RECT 72.710 178.065 72.970 178.385 ;
        RECT 71.330 177.725 71.590 178.045 ;
        RECT 72.250 177.725 72.510 178.045 ;
        RECT 74.550 177.725 74.810 178.045 ;
        RECT 73.170 176.880 73.430 177.025 ;
        RECT 73.160 176.510 73.440 176.880 ;
        RECT 74.610 176.005 74.750 177.725 ;
        RECT 70.870 175.685 71.130 176.005 ;
        RECT 73.170 175.685 73.430 176.005 ;
        RECT 74.550 175.685 74.810 176.005 ;
        RECT 70.930 175.325 72.450 175.405 ;
        RECT 72.710 175.345 72.970 175.665 ;
        RECT 70.930 175.265 72.510 175.325 ;
        RECT 70.930 174.985 71.070 175.265 ;
        RECT 72.250 175.005 72.510 175.265 ;
        RECT 70.870 174.665 71.130 174.985 ;
        RECT 71.330 174.840 71.590 174.985 ;
        RECT 71.320 174.470 71.600 174.840 ;
        RECT 71.790 174.725 72.050 174.985 ;
        RECT 72.770 174.725 72.910 175.345 ;
        RECT 73.230 175.325 73.370 175.685 ;
        RECT 73.170 175.005 73.430 175.325 ;
        RECT 75.530 174.985 75.670 182.825 ;
        RECT 75.930 180.105 76.190 180.425 ;
        RECT 75.990 178.045 76.130 180.105 ;
        RECT 75.930 177.725 76.190 178.045 ;
        RECT 76.390 177.725 76.650 178.045 ;
        RECT 76.450 174.985 76.590 177.725 ;
        RECT 77.370 175.665 77.510 189.285 ;
        RECT 78.230 188.605 78.490 188.925 ;
        RECT 85.130 188.605 85.390 188.925 ;
        RECT 77.770 187.585 78.030 187.905 ;
        RECT 77.830 185.525 77.970 187.585 ;
        RECT 77.770 185.205 78.030 185.525 ;
        RECT 78.290 183.485 78.430 188.605 ;
        RECT 78.690 188.265 78.950 188.585 ;
        RECT 78.230 183.165 78.490 183.485 ;
        RECT 78.750 183.145 78.890 188.265 ;
        RECT 79.910 187.050 81.790 187.420 ;
        RECT 85.190 186.545 85.330 188.605 ;
        RECT 85.130 186.285 85.390 186.545 ;
        RECT 84.730 186.225 85.390 186.285 ;
        RECT 84.730 186.145 85.330 186.225 ;
        RECT 86.570 186.205 86.710 190.985 ;
        RECT 92.490 190.305 92.750 190.625 ;
        RECT 92.550 189.605 92.690 190.305 ;
        RECT 92.490 189.285 92.750 189.605 ;
        RECT 89.730 187.585 89.990 187.905 ;
        RECT 81.910 183.165 82.170 183.485 ;
        RECT 82.830 183.165 83.090 183.485 ;
        RECT 77.770 182.825 78.030 183.145 ;
        RECT 78.690 182.825 78.950 183.145 ;
        RECT 79.610 182.885 79.870 183.145 ;
        RECT 79.210 182.825 79.870 182.885 ;
        RECT 77.830 180.085 77.970 182.825 ;
        RECT 78.750 181.445 78.890 182.825 ;
        RECT 79.210 182.745 79.810 182.825 ;
        RECT 78.690 181.125 78.950 181.445 ;
        RECT 77.770 179.765 78.030 180.085 ;
        RECT 79.210 178.045 79.350 182.745 ;
        RECT 79.910 181.610 81.790 181.980 ;
        RECT 79.150 177.725 79.410 178.045 ;
        RECT 78.690 177.385 78.950 177.705 ;
        RECT 77.310 175.345 77.570 175.665 ;
        RECT 78.750 174.985 78.890 177.385 ;
        RECT 79.910 176.170 81.790 176.540 ;
        RECT 81.970 175.325 82.110 183.165 ;
        RECT 82.890 178.725 83.030 183.165 ;
        RECT 84.210 182.145 84.470 182.465 ;
        RECT 84.270 180.765 84.410 182.145 ;
        RECT 84.210 180.445 84.470 180.765 ;
        RECT 84.730 180.165 84.870 186.145 ;
        RECT 86.510 185.885 86.770 186.205 ;
        RECT 87.430 185.885 87.690 186.205 ;
        RECT 86.050 185.545 86.310 185.865 ;
        RECT 86.110 184.165 86.250 185.545 ;
        RECT 86.050 183.845 86.310 184.165 ;
        RECT 86.570 183.145 86.710 185.885 ;
        RECT 86.510 182.825 86.770 183.145 ;
        RECT 85.590 182.145 85.850 182.465 ;
        RECT 84.270 180.025 84.870 180.165 ;
        RECT 82.830 178.405 83.090 178.725 ;
        RECT 84.270 177.705 84.410 180.025 ;
        RECT 85.650 178.725 85.790 182.145 ;
        RECT 86.050 180.675 86.310 180.765 ;
        RECT 86.570 180.675 86.710 182.825 ;
        RECT 86.050 180.535 86.710 180.675 ;
        RECT 86.050 180.445 86.310 180.535 ;
        RECT 85.590 178.405 85.850 178.725 ;
        RECT 84.210 177.385 84.470 177.705 ;
        RECT 81.910 175.005 82.170 175.325 ;
        RECT 84.270 174.985 84.410 177.385 ;
        RECT 71.790 174.665 72.910 174.725 ;
        RECT 75.010 174.665 75.270 174.985 ;
        RECT 75.470 174.665 75.730 174.985 ;
        RECT 76.390 174.665 76.650 174.985 ;
        RECT 78.690 174.665 78.950 174.985 ;
        RECT 84.210 174.665 84.470 174.985 ;
        RECT 71.850 174.585 72.910 174.665 ;
        RECT 71.390 171.585 71.530 174.470 ;
        RECT 73.170 174.160 73.430 174.305 ;
        RECT 73.160 173.790 73.440 174.160 ;
        RECT 73.630 172.625 73.890 172.945 ;
        RECT 71.330 171.265 71.590 171.585 ;
        RECT 73.170 169.565 73.430 169.885 ;
        RECT 71.330 168.885 71.590 169.205 ;
        RECT 71.390 167.505 71.530 168.885 ;
        RECT 71.330 167.185 71.590 167.505 ;
        RECT 70.410 166.165 70.670 166.485 ;
        RECT 71.390 163.765 71.530 167.185 ;
        RECT 73.230 166.825 73.370 169.565 ;
        RECT 73.690 167.845 73.830 172.625 ;
        RECT 74.090 171.605 74.350 171.925 ;
        RECT 73.630 167.525 73.890 167.845 ;
        RECT 74.150 166.825 74.290 171.605 ;
        RECT 75.070 171.585 75.210 174.665 ;
        RECT 75.930 173.985 76.190 174.305 ;
        RECT 75.010 171.265 75.270 171.585 ;
        RECT 73.170 166.505 73.430 166.825 ;
        RECT 74.090 166.505 74.350 166.825 ;
        RECT 73.230 164.445 73.370 166.505 ;
        RECT 73.170 164.125 73.430 164.445 ;
        RECT 71.330 163.445 71.590 163.765 ;
        RECT 70.410 163.105 70.670 163.425 ;
        RECT 70.470 161.725 70.610 163.105 ;
        RECT 71.390 161.725 71.530 163.445 ;
        RECT 72.710 161.745 72.970 162.065 ;
        RECT 70.410 161.405 70.670 161.725 ;
        RECT 70.870 161.405 71.130 161.725 ;
        RECT 71.330 161.405 71.590 161.725 ;
        RECT 70.470 158.665 70.610 161.405 ;
        RECT 70.930 160.560 71.070 161.405 ;
        RECT 70.860 160.190 71.140 160.560 ;
        RECT 70.410 158.520 70.670 158.665 ;
        RECT 70.400 158.150 70.680 158.520 ;
        RECT 70.930 158.235 71.070 160.190 ;
        RECT 72.250 159.025 72.510 159.345 ;
        RECT 71.790 158.685 72.050 159.005 ;
        RECT 71.330 158.235 71.590 158.325 ;
        RECT 70.470 156.965 70.610 158.150 ;
        RECT 70.930 158.095 71.590 158.235 ;
        RECT 71.330 158.005 71.590 158.095 ;
        RECT 70.410 156.645 70.670 156.965 ;
        RECT 71.390 156.625 71.530 158.005 ;
        RECT 71.330 156.305 71.590 156.625 ;
        RECT 71.850 156.285 71.990 158.685 ;
        RECT 70.410 155.965 70.670 156.285 ;
        RECT 71.790 155.965 72.050 156.285 ;
        RECT 70.470 155.120 70.610 155.965 ;
        RECT 70.400 154.750 70.680 155.120 ;
        RECT 71.330 154.945 71.590 155.265 ;
        RECT 70.410 153.925 70.670 154.245 ;
        RECT 69.950 150.185 70.210 150.505 ;
        RECT 69.950 149.505 70.210 149.825 ;
        RECT 67.650 136.585 67.910 136.905 ;
        RECT 69.490 136.585 69.750 136.905 ;
        RECT 67.190 131.485 67.450 131.805 ;
        RECT 64.430 130.465 64.690 130.785 ;
        RECT 64.490 129.085 64.630 130.465 ;
        RECT 64.910 129.930 66.790 130.300 ;
        RECT 64.430 128.765 64.690 129.085 ;
        RECT 64.910 124.490 66.790 124.860 ;
        RECT 65.350 123.665 65.610 123.985 ;
        RECT 63.510 122.985 63.770 123.305 ;
        RECT 62.590 120.265 62.850 120.585 ;
        RECT 62.650 118.545 62.790 120.265 ;
        RECT 63.570 118.885 63.710 122.985 ;
        RECT 65.410 121.605 65.550 123.665 ;
        RECT 65.350 121.285 65.610 121.605 ;
        RECT 64.910 119.050 66.790 119.420 ;
        RECT 63.510 118.565 63.770 118.885 ;
        RECT 62.590 118.225 62.850 118.545 ;
        RECT 67.250 116.165 67.390 131.485 ;
        RECT 67.710 131.465 67.850 136.585 ;
        RECT 67.650 131.145 67.910 131.465 ;
        RECT 68.570 130.465 68.830 130.785 ;
        RECT 68.630 129.085 68.770 130.465 ;
        RECT 68.570 128.765 68.830 129.085 ;
        RECT 68.630 126.705 68.770 128.765 ;
        RECT 69.490 128.425 69.750 128.745 ;
        RECT 68.570 126.385 68.830 126.705 ;
        RECT 69.550 125.345 69.690 128.425 ;
        RECT 68.570 125.025 68.830 125.345 ;
        RECT 69.490 125.025 69.750 125.345 ;
        RECT 68.630 118.205 68.770 125.025 ;
        RECT 69.550 123.645 69.690 125.025 ;
        RECT 69.490 123.325 69.750 123.645 ;
        RECT 69.550 121.605 69.690 123.325 ;
        RECT 69.490 121.285 69.750 121.605 ;
        RECT 69.490 119.925 69.750 120.245 ;
        RECT 69.550 118.885 69.690 119.925 ;
        RECT 69.490 118.565 69.750 118.885 ;
        RECT 68.570 117.885 68.830 118.205 ;
        RECT 67.190 115.845 67.450 116.165 ;
        RECT 70.010 115.145 70.150 149.505 ;
        RECT 70.470 148.125 70.610 153.925 ;
        RECT 71.390 152.545 71.530 154.945 ;
        RECT 71.330 152.225 71.590 152.545 ;
        RECT 71.790 150.755 72.050 150.845 ;
        RECT 72.310 150.755 72.450 159.025 ;
        RECT 72.770 156.285 72.910 161.745 ;
        RECT 73.230 161.385 73.370 164.125 ;
        RECT 73.630 161.405 73.890 161.725 ;
        RECT 73.170 161.065 73.430 161.385 ;
        RECT 73.690 158.665 73.830 161.405 ;
        RECT 74.150 159.685 74.290 166.505 ;
        RECT 75.470 163.785 75.730 164.105 ;
        RECT 74.550 163.105 74.810 163.425 ;
        RECT 74.610 161.385 74.750 163.105 ;
        RECT 74.550 161.065 74.810 161.385 ;
        RECT 74.090 159.365 74.350 159.685 ;
        RECT 73.630 158.345 73.890 158.665 ;
        RECT 74.610 158.325 74.750 161.065 ;
        RECT 75.530 159.685 75.670 163.785 ;
        RECT 75.470 159.365 75.730 159.685 ;
        RECT 74.550 158.005 74.810 158.325 ;
        RECT 72.710 155.965 72.970 156.285 ;
        RECT 74.090 155.965 74.350 156.285 ;
        RECT 74.150 155.800 74.290 155.965 ;
        RECT 74.080 155.430 74.360 155.800 ;
        RECT 74.550 155.515 74.810 155.605 ;
        RECT 74.550 155.375 75.210 155.515 ;
        RECT 74.550 155.285 74.810 155.375 ;
        RECT 73.170 154.945 73.430 155.265 ;
        RECT 71.790 150.615 72.450 150.755 ;
        RECT 71.790 150.525 72.050 150.615 ;
        RECT 72.250 149.505 72.510 149.825 ;
        RECT 71.330 148.485 71.590 148.805 ;
        RECT 70.410 147.805 70.670 148.125 ;
        RECT 70.410 137.605 70.670 137.925 ;
        RECT 70.470 129.765 70.610 137.605 ;
        RECT 70.410 129.445 70.670 129.765 ;
        RECT 71.390 127.045 71.530 148.485 ;
        RECT 71.780 147.950 72.060 148.320 ;
        RECT 71.790 147.805 72.050 147.950 ;
        RECT 71.780 140.470 72.060 140.840 ;
        RECT 71.850 137.245 71.990 140.470 ;
        RECT 71.790 136.925 72.050 137.245 ;
        RECT 71.790 135.905 72.050 136.225 ;
        RECT 71.330 126.725 71.590 127.045 ;
        RECT 69.950 114.825 70.210 115.145 ;
        RECT 69.030 114.145 69.290 114.465 ;
        RECT 70.870 114.145 71.130 114.465 ;
        RECT 64.910 113.610 66.790 113.980 ;
        RECT 62.130 113.125 62.390 113.445 ;
        RECT 61.210 112.785 61.470 113.105 ;
        RECT 60.290 112.105 60.550 112.425 ;
        RECT 60.350 110.045 60.490 112.105 ;
        RECT 61.270 110.725 61.410 112.785 ;
        RECT 69.090 112.765 69.230 114.145 ;
        RECT 70.930 113.445 71.070 114.145 ;
        RECT 70.870 113.125 71.130 113.445 ;
        RECT 69.030 112.445 69.290 112.765 ;
        RECT 67.650 112.105 67.910 112.425 ;
        RECT 65.350 111.425 65.610 111.745 ;
        RECT 61.210 110.405 61.470 110.725 ;
        RECT 65.410 110.045 65.550 111.425 ;
        RECT 60.290 109.725 60.550 110.045 ;
        RECT 65.350 109.725 65.610 110.045 ;
        RECT 59.830 109.385 60.090 109.705 ;
        RECT 62.130 109.045 62.390 109.365 ;
        RECT 58.910 107.685 59.170 108.005 ;
        RECT 58.450 107.005 58.710 107.325 ;
        RECT 62.190 95.885 62.330 109.045 ;
        RECT 64.910 108.170 66.790 108.540 ;
        RECT 67.710 95.885 67.850 112.105 ;
        RECT 71.850 111.745 71.990 135.905 ;
        RECT 72.310 132.485 72.450 149.505 ;
        RECT 72.710 134.885 72.970 135.205 ;
        RECT 72.250 132.165 72.510 132.485 ;
        RECT 72.250 127.745 72.510 128.065 ;
        RECT 72.310 126.705 72.450 127.745 ;
        RECT 72.250 126.385 72.510 126.705 ;
        RECT 72.310 123.305 72.450 126.385 ;
        RECT 72.250 122.985 72.510 123.305 ;
        RECT 72.250 117.545 72.510 117.865 ;
        RECT 72.310 115.145 72.450 117.545 ;
        RECT 72.770 115.825 72.910 134.885 ;
        RECT 73.230 134.525 73.370 154.945 ;
        RECT 74.090 150.525 74.350 150.845 ;
        RECT 74.550 150.525 74.810 150.845 ;
        RECT 74.150 148.465 74.290 150.525 ;
        RECT 74.090 148.145 74.350 148.465 ;
        RECT 74.610 147.785 74.750 150.525 ;
        RECT 75.070 148.465 75.210 155.375 ;
        RECT 75.460 152.710 75.740 153.080 ;
        RECT 75.530 152.545 75.670 152.710 ;
        RECT 75.470 152.225 75.730 152.545 ;
        RECT 75.470 150.525 75.730 150.845 ;
        RECT 75.010 148.145 75.270 148.465 ;
        RECT 73.630 147.465 73.890 147.785 ;
        RECT 74.550 147.465 74.810 147.785 ;
        RECT 73.170 134.205 73.430 134.525 ;
        RECT 72.710 115.505 72.970 115.825 ;
        RECT 72.250 114.825 72.510 115.145 ;
        RECT 73.690 113.015 73.830 147.465 ;
        RECT 74.610 139.965 74.750 147.465 ;
        RECT 75.070 139.965 75.210 148.145 ;
        RECT 75.530 147.785 75.670 150.525 ;
        RECT 75.470 147.465 75.730 147.785 ;
        RECT 75.530 146.085 75.670 147.465 ;
        RECT 75.470 145.765 75.730 146.085 ;
        RECT 75.530 140.305 75.670 145.765 ;
        RECT 75.470 139.985 75.730 140.305 ;
        RECT 74.550 139.645 74.810 139.965 ;
        RECT 75.010 139.645 75.270 139.965 ;
        RECT 74.610 137.585 74.750 139.645 ;
        RECT 75.070 137.925 75.210 139.645 ;
        RECT 75.010 137.605 75.270 137.925 ;
        RECT 74.550 137.265 74.810 137.585 ;
        RECT 75.530 136.905 75.670 139.985 ;
        RECT 75.470 136.585 75.730 136.905 ;
        RECT 75.990 134.185 76.130 173.985 ;
        RECT 78.230 171.605 78.490 171.925 ;
        RECT 77.770 168.885 78.030 169.205 ;
        RECT 77.830 167.845 77.970 168.885 ;
        RECT 78.290 168.865 78.430 171.605 ;
        RECT 78.750 171.585 78.890 174.665 ;
        RECT 86.570 172.605 86.710 180.535 ;
        RECT 87.490 180.425 87.630 185.885 ;
        RECT 89.790 185.525 89.930 187.585 ;
        RECT 89.730 185.205 89.990 185.525 ;
        RECT 88.810 184.865 89.070 185.185 ;
        RECT 88.870 183.825 89.010 184.865 ;
        RECT 88.810 183.505 89.070 183.825 ;
        RECT 92.950 183.165 93.210 183.485 ;
        RECT 92.490 182.825 92.750 183.145 ;
        RECT 87.430 180.105 87.690 180.425 ;
        RECT 87.490 178.385 87.630 180.105 ;
        RECT 92.550 179.745 92.690 182.825 ;
        RECT 93.010 180.425 93.150 183.165 ;
        RECT 93.470 182.805 93.610 191.325 ;
        RECT 93.930 188.585 94.070 193.025 ;
        RECT 98.990 191.645 99.130 193.705 ;
        RECT 98.930 191.325 99.190 191.645 ;
        RECT 97.090 190.305 97.350 190.625 ;
        RECT 94.910 189.770 96.790 190.140 ;
        RECT 97.150 188.925 97.290 190.305 ;
        RECT 97.090 188.605 97.350 188.925 ;
        RECT 93.870 188.265 94.130 188.585 ;
        RECT 98.930 188.265 99.190 188.585 ;
        RECT 93.410 182.485 93.670 182.805 ;
        RECT 93.470 180.765 93.610 182.485 ;
        RECT 93.930 180.765 94.070 188.265 ;
        RECT 97.090 187.585 97.350 187.905 ;
        RECT 94.910 184.330 96.790 184.700 ;
        RECT 97.150 184.165 97.290 187.585 ;
        RECT 97.550 185.205 97.810 185.525 ;
        RECT 97.090 183.845 97.350 184.165 ;
        RECT 97.090 182.485 97.350 182.805 ;
        RECT 93.410 180.445 93.670 180.765 ;
        RECT 93.870 180.445 94.130 180.765 ;
        RECT 92.950 180.105 93.210 180.425 ;
        RECT 94.330 180.165 94.590 180.425 ;
        RECT 93.930 180.105 94.590 180.165 ;
        RECT 93.930 180.025 94.530 180.105 ;
        RECT 90.190 179.425 90.450 179.745 ;
        RECT 92.490 179.425 92.750 179.745 ;
        RECT 92.950 179.425 93.210 179.745 ;
        RECT 87.430 178.065 87.690 178.385 ;
        RECT 90.250 178.045 90.390 179.425 ;
        RECT 90.190 177.725 90.450 178.045 ;
        RECT 87.890 177.385 88.150 177.705 ;
        RECT 91.570 177.385 91.830 177.705 ;
        RECT 87.950 172.945 88.090 177.385 ;
        RECT 88.810 176.705 89.070 177.025 ;
        RECT 88.350 173.985 88.610 174.305 ;
        RECT 88.410 172.945 88.550 173.985 ;
        RECT 87.890 172.625 88.150 172.945 ;
        RECT 88.350 172.625 88.610 172.945 ;
        RECT 86.510 172.285 86.770 172.605 ;
        RECT 84.670 171.945 84.930 172.265 ;
        RECT 78.690 171.265 78.950 171.585 ;
        RECT 79.910 170.730 81.790 171.100 ;
        RECT 84.730 170.565 84.870 171.945 ;
        RECT 84.670 170.245 84.930 170.565 ;
        RECT 86.570 169.885 86.710 172.285 ;
        RECT 88.350 171.945 88.610 172.265 ;
        RECT 88.410 170.565 88.550 171.945 ;
        RECT 88.350 170.245 88.610 170.565 ;
        RECT 78.690 169.565 78.950 169.885 ;
        RECT 86.510 169.565 86.770 169.885 ;
        RECT 78.230 168.545 78.490 168.865 ;
        RECT 77.770 167.525 78.030 167.845 ;
        RECT 78.230 166.845 78.490 167.165 ;
        RECT 78.290 161.725 78.430 166.845 ;
        RECT 78.750 165.125 78.890 169.565 ;
        RECT 79.150 169.225 79.410 169.545 ;
        RECT 79.210 167.845 79.350 169.225 ;
        RECT 86.570 167.845 86.710 169.565 ;
        RECT 79.150 167.525 79.410 167.845 ;
        RECT 86.510 167.525 86.770 167.845 ;
        RECT 79.140 166.990 79.420 167.360 ;
        RECT 79.150 166.845 79.410 166.990 ;
        RECT 78.690 164.805 78.950 165.125 ;
        RECT 79.210 163.960 79.350 166.845 ;
        RECT 79.910 165.290 81.790 165.660 ;
        RECT 79.140 163.590 79.420 163.960 ;
        RECT 84.210 163.105 84.470 163.425 ;
        RECT 84.270 162.065 84.410 163.105 ;
        RECT 84.210 161.745 84.470 162.065 ;
        RECT 86.050 161.745 86.310 162.065 ;
        RECT 78.230 161.635 78.490 161.725 ;
        RECT 77.830 161.495 78.490 161.635 ;
        RECT 77.830 159.005 77.970 161.495 ;
        RECT 78.230 161.405 78.490 161.495 ;
        RECT 78.230 160.385 78.490 160.705 ;
        RECT 78.690 160.385 78.950 160.705 ;
        RECT 82.370 160.385 82.630 160.705 ;
        RECT 77.770 158.685 78.030 159.005 ;
        RECT 78.290 156.625 78.430 160.385 ;
        RECT 78.750 158.325 78.890 160.385 ;
        RECT 79.910 159.850 81.790 160.220 ;
        RECT 82.430 159.005 82.570 160.385 ;
        RECT 86.110 159.685 86.250 161.745 ;
        RECT 86.570 161.385 86.710 167.525 ;
        RECT 86.510 161.065 86.770 161.385 ;
        RECT 86.050 159.365 86.310 159.685 ;
        RECT 86.570 159.005 86.710 161.065 ;
        RECT 82.370 158.685 82.630 159.005 ;
        RECT 86.510 158.685 86.770 159.005 ;
        RECT 86.970 158.345 87.230 158.665 ;
        RECT 78.690 158.005 78.950 158.325 ;
        RECT 78.230 156.305 78.490 156.625 ;
        RECT 79.910 154.410 81.790 154.780 ;
        RECT 76.390 153.245 76.650 153.565 ;
        RECT 76.450 142.685 76.590 153.245 ;
        RECT 78.230 152.905 78.490 153.225 ;
        RECT 76.850 152.225 77.110 152.545 ;
        RECT 77.770 152.225 78.030 152.545 ;
        RECT 76.910 151.185 77.050 152.225 ;
        RECT 76.850 150.865 77.110 151.185 ;
        RECT 77.830 148.125 77.970 152.225 ;
        RECT 78.290 151.525 78.430 152.905 ;
        RECT 79.150 152.565 79.410 152.885 ;
        RECT 78.230 151.205 78.490 151.525 ;
        RECT 77.770 147.805 78.030 148.125 ;
        RECT 77.830 146.085 77.970 147.805 ;
        RECT 79.210 147.785 79.350 152.565 ;
        RECT 84.670 152.225 84.930 152.545 ;
        RECT 86.050 152.225 86.310 152.545 ;
        RECT 84.730 150.845 84.870 152.225 ;
        RECT 86.110 151.525 86.250 152.225 ;
        RECT 86.050 151.205 86.310 151.525 ;
        RECT 84.670 150.525 84.930 150.845 ;
        RECT 86.510 150.185 86.770 150.505 ;
        RECT 79.910 148.970 81.790 149.340 ;
        RECT 79.150 147.465 79.410 147.785 ;
        RECT 81.910 147.465 82.170 147.785 ;
        RECT 77.770 145.765 78.030 146.085 ;
        RECT 77.830 142.685 77.970 145.765 ;
        RECT 76.390 142.365 76.650 142.685 ;
        RECT 77.770 142.365 78.030 142.685 ;
        RECT 76.450 139.365 76.590 142.365 ;
        RECT 77.770 141.345 78.030 141.665 ;
        RECT 77.310 139.645 77.570 139.965 ;
        RECT 76.450 139.225 77.050 139.365 ;
        RECT 76.390 138.625 76.650 138.945 ;
        RECT 76.450 134.865 76.590 138.625 ;
        RECT 76.910 137.925 77.050 139.225 ;
        RECT 76.850 137.605 77.110 137.925 ;
        RECT 76.390 134.545 76.650 134.865 ;
        RECT 76.910 134.185 77.050 137.605 ;
        RECT 77.370 135.205 77.510 139.645 ;
        RECT 77.830 136.225 77.970 141.345 ;
        RECT 79.210 139.965 79.350 147.465 ;
        RECT 80.070 146.785 80.330 147.105 ;
        RECT 80.130 145.745 80.270 146.785 ;
        RECT 80.070 145.425 80.330 145.745 ;
        RECT 79.910 143.530 81.790 143.900 ;
        RECT 81.970 143.365 82.110 147.465 ;
        RECT 84.670 146.785 84.930 147.105 ;
        RECT 84.730 145.405 84.870 146.785 ;
        RECT 84.670 145.085 84.930 145.405 ;
        RECT 86.570 145.065 86.710 150.185 ;
        RECT 87.030 147.785 87.170 158.345 ;
        RECT 87.890 150.865 88.150 151.185 ;
        RECT 87.950 148.805 88.090 150.865 ;
        RECT 88.350 150.185 88.610 150.505 ;
        RECT 88.410 148.805 88.550 150.185 ;
        RECT 87.890 148.485 88.150 148.805 ;
        RECT 88.350 148.485 88.610 148.805 ;
        RECT 86.970 147.465 87.230 147.785 ;
        RECT 87.030 146.085 87.170 147.465 ;
        RECT 86.970 145.765 87.230 146.085 ;
        RECT 86.510 144.745 86.770 145.065 ;
        RECT 81.910 143.045 82.170 143.365 ;
        RECT 84.670 139.985 84.930 140.305 ;
        RECT 79.150 139.645 79.410 139.965 ;
        RECT 78.230 138.625 78.490 138.945 ;
        RECT 78.690 138.625 78.950 138.945 ;
        RECT 78.290 137.245 78.430 138.625 ;
        RECT 78.230 136.925 78.490 137.245 ;
        RECT 78.750 136.565 78.890 138.625 ;
        RECT 78.690 136.245 78.950 136.565 ;
        RECT 77.770 135.905 78.030 136.225 ;
        RECT 77.310 134.885 77.570 135.205 ;
        RECT 79.210 134.605 79.350 139.645 ;
        RECT 79.910 138.090 81.790 138.460 ;
        RECT 84.210 136.585 84.470 136.905 ;
        RECT 79.610 135.905 79.870 136.225 ;
        RECT 79.670 135.205 79.810 135.905 ;
        RECT 79.610 134.885 79.870 135.205 ;
        RECT 79.210 134.525 79.810 134.605 ;
        RECT 79.210 134.465 79.870 134.525 ;
        RECT 79.610 134.205 79.870 134.465 ;
        RECT 75.930 133.865 76.190 134.185 ;
        RECT 76.850 133.865 77.110 134.185 ;
        RECT 77.310 133.185 77.570 133.505 ;
        RECT 74.550 131.485 74.810 131.805 ;
        RECT 74.610 129.765 74.750 131.485 ;
        RECT 77.370 129.765 77.510 133.185 ;
        RECT 79.910 132.650 81.790 133.020 ;
        RECT 84.270 132.485 84.410 136.585 ;
        RECT 84.730 135.205 84.870 139.985 ;
        RECT 86.570 139.625 86.710 144.745 ;
        RECT 88.870 142.685 89.010 176.705 ;
        RECT 91.630 173.285 91.770 177.385 ;
        RECT 92.550 175.325 92.690 179.425 ;
        RECT 92.490 175.005 92.750 175.325 ;
        RECT 92.490 173.985 92.750 174.305 ;
        RECT 92.550 173.285 92.690 173.985 ;
        RECT 91.570 172.965 91.830 173.285 ;
        RECT 92.490 172.965 92.750 173.285 ;
        RECT 91.110 169.905 91.370 170.225 ;
        RECT 90.640 166.990 90.920 167.360 ;
        RECT 90.650 166.845 90.910 166.990 ;
        RECT 89.730 165.825 89.990 166.145 ;
        RECT 89.270 164.125 89.530 164.445 ;
        RECT 89.330 159.685 89.470 164.125 ;
        RECT 89.790 163.765 89.930 165.825 ;
        RECT 89.730 163.445 89.990 163.765 ;
        RECT 89.270 159.365 89.530 159.685 ;
        RECT 91.170 158.665 91.310 169.905 ;
        RECT 92.550 169.885 92.690 172.965 ;
        RECT 92.490 169.565 92.750 169.885 ;
        RECT 92.490 168.885 92.750 169.205 ;
        RECT 92.550 165.125 92.690 168.885 ;
        RECT 92.490 164.805 92.750 165.125 ;
        RECT 91.570 159.365 91.830 159.685 ;
        RECT 91.110 158.345 91.370 158.665 ;
        RECT 90.650 157.665 90.910 157.985 ;
        RECT 90.710 156.195 90.850 157.665 ;
        RECT 91.110 156.195 91.370 156.285 ;
        RECT 90.710 156.055 91.370 156.195 ;
        RECT 91.110 155.965 91.370 156.055 ;
        RECT 89.730 154.945 89.990 155.265 ;
        RECT 89.270 152.225 89.530 152.545 ;
        RECT 89.330 147.785 89.470 152.225 ;
        RECT 89.270 147.465 89.530 147.785 ;
        RECT 88.810 142.365 89.070 142.685 ;
        RECT 89.790 142.345 89.930 154.945 ;
        RECT 91.110 144.745 91.370 145.065 ;
        RECT 90.190 143.045 90.450 143.365 ;
        RECT 89.730 142.025 89.990 142.345 ;
        RECT 86.970 141.345 87.230 141.665 ;
        RECT 86.510 139.305 86.770 139.625 ;
        RECT 86.050 138.625 86.310 138.945 ;
        RECT 86.110 137.245 86.250 138.625 ;
        RECT 86.570 137.245 86.710 139.305 ;
        RECT 86.050 136.925 86.310 137.245 ;
        RECT 86.510 136.925 86.770 137.245 ;
        RECT 84.670 134.885 84.930 135.205 ;
        RECT 86.110 134.865 86.250 136.925 ;
        RECT 86.050 134.545 86.310 134.865 ;
        RECT 85.130 134.205 85.390 134.525 ;
        RECT 85.190 132.485 85.330 134.205 ;
        RECT 85.590 133.185 85.850 133.505 ;
        RECT 84.210 132.165 84.470 132.485 ;
        RECT 85.130 132.165 85.390 132.485 ;
        RECT 74.550 129.445 74.810 129.765 ;
        RECT 77.310 129.445 77.570 129.765 ;
        RECT 74.090 128.425 74.350 128.745 ;
        RECT 74.150 126.365 74.290 128.425 ;
        RECT 74.610 127.045 74.750 129.445 ;
        RECT 84.270 128.745 84.410 132.165 ;
        RECT 84.660 131.630 84.940 132.000 ;
        RECT 84.730 131.465 84.870 131.630 ;
        RECT 84.670 131.145 84.930 131.465 ;
        RECT 85.650 129.085 85.790 133.185 ;
        RECT 85.590 128.765 85.850 129.085 ;
        RECT 79.150 128.425 79.410 128.745 ;
        RECT 84.210 128.425 84.470 128.745 ;
        RECT 76.390 127.745 76.650 128.065 ;
        RECT 76.450 127.045 76.590 127.745 ;
        RECT 74.550 126.725 74.810 127.045 ;
        RECT 76.390 126.725 76.650 127.045 ;
        RECT 74.090 126.045 74.350 126.365 ;
        RECT 74.150 123.985 74.290 126.045 ;
        RECT 78.230 125.365 78.490 125.685 ;
        RECT 78.290 124.325 78.430 125.365 ;
        RECT 78.230 124.005 78.490 124.325 ;
        RECT 74.090 123.665 74.350 123.985 ;
        RECT 78.230 123.325 78.490 123.645 ;
        RECT 76.390 122.305 76.650 122.625 ;
        RECT 76.450 120.585 76.590 122.305 ;
        RECT 76.390 120.265 76.650 120.585 ;
        RECT 78.290 118.545 78.430 123.325 ;
        RECT 79.210 123.305 79.350 128.425 ;
        RECT 79.910 127.210 81.790 127.580 ;
        RECT 84.270 126.705 84.410 128.425 ;
        RECT 84.210 126.385 84.470 126.705 ;
        RECT 79.150 122.985 79.410 123.305 ;
        RECT 79.210 121.605 79.350 122.985 ;
        RECT 79.910 121.770 81.790 122.140 ;
        RECT 79.150 121.285 79.410 121.605 ;
        RECT 81.910 120.605 82.170 120.925 ;
        RECT 84.270 120.835 84.410 126.385 ;
        RECT 86.050 123.665 86.310 123.985 ;
        RECT 84.670 120.835 84.930 120.925 ;
        RECT 84.270 120.695 84.930 120.835 ;
        RECT 84.670 120.605 84.930 120.695 ;
        RECT 81.450 119.925 81.710 120.245 ;
        RECT 81.510 118.885 81.650 119.925 ;
        RECT 81.450 118.565 81.710 118.885 ;
        RECT 78.230 118.225 78.490 118.545 ;
        RECT 79.910 116.330 81.790 116.700 ;
        RECT 78.230 114.485 78.490 114.805 ;
        RECT 75.010 113.015 75.270 113.105 ;
        RECT 73.690 112.875 75.270 113.015 ;
        RECT 75.010 112.785 75.270 112.875 ;
        RECT 74.550 112.105 74.810 112.425 ;
        RECT 71.790 111.425 72.050 111.745 ;
        RECT 74.610 110.045 74.750 112.105 ;
        RECT 77.310 111.425 77.570 111.745 ;
        RECT 74.550 109.725 74.810 110.045 ;
        RECT 74.610 106.985 74.750 109.725 ;
        RECT 77.370 107.665 77.510 111.425 ;
        RECT 78.290 109.025 78.430 114.485 ;
        RECT 81.970 113.105 82.110 120.605 ;
        RECT 86.110 118.885 86.250 123.665 ;
        RECT 86.510 122.305 86.770 122.625 ;
        RECT 86.570 120.925 86.710 122.305 ;
        RECT 86.510 120.605 86.770 120.925 ;
        RECT 86.050 118.565 86.310 118.885 ;
        RECT 87.030 115.145 87.170 141.345 ;
        RECT 87.430 139.645 87.690 139.965 ;
        RECT 87.490 135.205 87.630 139.645 ;
        RECT 88.350 135.905 88.610 136.225 ;
        RECT 87.430 134.885 87.690 135.205 ;
        RECT 88.410 134.525 88.550 135.905 ;
        RECT 88.350 134.205 88.610 134.525 ;
        RECT 90.250 134.185 90.390 143.045 ;
        RECT 91.170 142.345 91.310 144.745 ;
        RECT 91.110 142.025 91.370 142.345 ;
        RECT 91.110 136.585 91.370 136.905 ;
        RECT 90.650 134.425 90.910 134.525 ;
        RECT 91.170 134.425 91.310 136.585 ;
        RECT 90.650 134.285 91.310 134.425 ;
        RECT 90.650 134.205 90.910 134.285 ;
        RECT 90.190 133.865 90.450 134.185 ;
        RECT 87.890 129.105 88.150 129.425 ;
        RECT 87.950 127.045 88.090 129.105 ;
        RECT 87.890 126.725 88.150 127.045 ;
        RECT 91.170 126.025 91.310 134.285 ;
        RECT 91.630 133.505 91.770 159.365 ;
        RECT 92.030 158.345 92.290 158.665 ;
        RECT 92.090 156.965 92.230 158.345 ;
        RECT 92.030 156.645 92.290 156.965 ;
        RECT 92.030 156.195 92.290 156.285 ;
        RECT 92.550 156.195 92.690 164.805 ;
        RECT 93.010 159.005 93.150 179.425 ;
        RECT 93.930 177.365 94.070 180.025 ;
        RECT 94.910 178.890 96.790 179.260 ;
        RECT 97.150 178.045 97.290 182.485 ;
        RECT 97.610 181.445 97.750 185.205 ;
        RECT 98.990 182.805 99.130 188.265 ;
        RECT 98.930 182.485 99.190 182.805 ;
        RECT 97.550 181.125 97.810 181.445 ;
        RECT 98.470 180.105 98.730 180.425 ;
        RECT 98.010 179.765 98.270 180.085 ;
        RECT 98.070 178.385 98.210 179.765 ;
        RECT 98.010 178.065 98.270 178.385 ;
        RECT 98.530 178.045 98.670 180.105 ;
        RECT 99.450 178.045 99.590 197.105 ;
        RECT 99.850 196.765 100.110 197.085 ;
        RECT 99.910 189.605 100.050 196.765 ;
        RECT 109.510 196.425 109.770 196.745 ;
        RECT 100.310 195.745 100.570 196.065 ;
        RECT 100.370 195.045 100.510 195.745 ;
        RECT 100.310 194.725 100.570 195.045 ;
        RECT 100.370 190.965 100.510 194.725 ;
        RECT 100.770 194.045 101.030 194.365 ;
        RECT 100.310 190.645 100.570 190.965 ;
        RECT 99.850 189.285 100.110 189.605 ;
        RECT 100.830 188.925 100.970 194.045 ;
        RECT 101.690 193.705 101.950 194.025 ;
        RECT 101.750 190.625 101.890 193.705 ;
        RECT 107.210 193.025 107.470 193.345 ;
        RECT 108.590 193.025 108.850 193.345 ;
        RECT 107.270 190.965 107.410 193.025 ;
        RECT 108.650 191.645 108.790 193.025 ;
        RECT 108.590 191.325 108.850 191.645 ;
        RECT 109.570 191.215 109.710 196.425 ;
        RECT 109.910 192.490 111.790 192.860 ;
        RECT 109.970 191.215 110.230 191.305 ;
        RECT 109.570 191.075 110.230 191.215 ;
        RECT 107.210 190.645 107.470 190.965 ;
        RECT 101.690 190.305 101.950 190.625 ;
        RECT 100.770 188.605 101.030 188.925 ;
        RECT 101.750 188.585 101.890 190.305 ;
        RECT 101.690 188.265 101.950 188.585 ;
        RECT 107.210 188.265 107.470 188.585 ;
        RECT 100.770 187.585 101.030 187.905 ;
        RECT 101.690 187.585 101.950 187.905 ;
        RECT 103.990 187.585 104.250 187.905 ;
        RECT 100.310 185.205 100.570 185.525 ;
        RECT 100.370 184.165 100.510 185.205 ;
        RECT 100.310 183.845 100.570 184.165 ;
        RECT 100.830 183.825 100.970 187.585 ;
        RECT 101.750 185.525 101.890 187.585 ;
        RECT 103.530 185.885 103.790 186.205 ;
        RECT 101.690 185.205 101.950 185.525 ;
        RECT 100.770 183.505 101.030 183.825 ;
        RECT 99.850 182.145 100.110 182.465 ;
        RECT 99.910 180.425 100.050 182.145 ;
        RECT 99.850 180.105 100.110 180.425 ;
        RECT 103.590 179.745 103.730 185.885 ;
        RECT 104.050 179.745 104.190 187.585 ;
        RECT 104.450 182.145 104.710 182.465 ;
        RECT 104.510 180.765 104.650 182.145 ;
        RECT 104.450 180.445 104.710 180.765 ;
        RECT 107.270 180.425 107.410 188.265 ;
        RECT 109.570 185.185 109.710 191.075 ;
        RECT 109.970 190.985 110.230 191.075 ;
        RECT 109.910 187.050 111.790 187.420 ;
        RECT 111.350 185.205 111.610 185.525 ;
        RECT 109.510 184.865 109.770 185.185 ;
        RECT 111.410 182.725 111.550 185.205 ;
        RECT 111.810 184.865 112.070 185.185 ;
        RECT 111.870 183.485 112.010 184.865 ;
        RECT 111.810 183.165 112.070 183.485 ;
        RECT 113.190 183.165 113.450 183.485 ;
        RECT 111.410 182.585 112.470 182.725 ;
        RECT 109.910 181.610 111.790 181.980 ;
        RECT 112.330 181.445 112.470 182.585 ;
        RECT 112.730 182.145 112.990 182.465 ;
        RECT 112.270 181.125 112.530 181.445 ;
        RECT 112.790 181.105 112.930 182.145 ;
        RECT 112.730 180.785 112.990 181.105 ;
        RECT 107.210 180.105 107.470 180.425 ;
        RECT 108.130 180.105 108.390 180.425 ;
        RECT 112.270 180.105 112.530 180.425 ;
        RECT 103.530 179.425 103.790 179.745 ;
        RECT 103.990 179.425 104.250 179.745 ;
        RECT 105.830 179.425 106.090 179.745 ;
        RECT 94.330 177.725 94.590 178.045 ;
        RECT 95.710 177.725 95.970 178.045 ;
        RECT 97.090 177.725 97.350 178.045 ;
        RECT 97.550 177.725 97.810 178.045 ;
        RECT 98.470 177.725 98.730 178.045 ;
        RECT 99.390 177.725 99.650 178.045 ;
        RECT 100.310 177.725 100.570 178.045 ;
        RECT 93.870 177.045 94.130 177.365 ;
        RECT 94.390 175.325 94.530 177.725 ;
        RECT 95.770 177.365 95.910 177.725 ;
        RECT 95.710 177.045 95.970 177.365 ;
        RECT 97.610 175.325 97.750 177.725 ;
        RECT 98.930 177.045 99.190 177.365 ;
        RECT 98.470 176.705 98.730 177.025 ;
        RECT 94.330 175.005 94.590 175.325 ;
        RECT 97.550 175.005 97.810 175.325 ;
        RECT 93.870 174.665 94.130 174.985 ;
        RECT 93.410 171.945 93.670 172.265 ;
        RECT 93.470 169.885 93.610 171.945 ;
        RECT 93.930 171.585 94.070 174.665 ;
        RECT 93.870 171.265 94.130 171.585 ;
        RECT 93.870 170.475 94.130 170.565 ;
        RECT 94.390 170.475 94.530 175.005 ;
        RECT 97.090 173.985 97.350 174.305 ;
        RECT 94.910 173.450 96.790 173.820 ;
        RECT 97.150 172.605 97.290 173.985 ;
        RECT 97.090 172.285 97.350 172.605 ;
        RECT 97.090 171.265 97.350 171.585 ;
        RECT 93.870 170.335 94.530 170.475 ;
        RECT 93.870 170.245 94.130 170.335 ;
        RECT 93.410 169.565 93.670 169.885 ;
        RECT 93.470 164.105 93.610 169.565 ;
        RECT 94.330 168.885 94.590 169.205 ;
        RECT 93.410 163.785 93.670 164.105 ;
        RECT 93.410 163.105 93.670 163.425 ;
        RECT 93.470 161.725 93.610 163.105 ;
        RECT 94.390 162.065 94.530 168.885 ;
        RECT 94.910 168.010 96.790 168.380 ;
        RECT 94.910 162.570 96.790 162.940 ;
        RECT 94.330 161.745 94.590 162.065 ;
        RECT 93.410 161.405 93.670 161.725 ;
        RECT 92.950 158.685 93.210 159.005 ;
        RECT 93.870 158.345 94.130 158.665 ;
        RECT 92.950 158.005 93.210 158.325 ;
        RECT 93.410 158.005 93.670 158.325 ;
        RECT 93.010 156.625 93.150 158.005 ;
        RECT 92.950 156.305 93.210 156.625 ;
        RECT 92.030 156.055 92.690 156.195 ;
        RECT 92.030 155.965 92.290 156.055 ;
        RECT 93.470 154.245 93.610 158.005 ;
        RECT 93.930 156.285 94.070 158.345 ;
        RECT 94.330 157.665 94.590 157.985 ;
        RECT 93.870 155.965 94.130 156.285 ;
        RECT 93.930 155.265 94.070 155.965 ;
        RECT 93.870 154.945 94.130 155.265 ;
        RECT 93.410 153.925 93.670 154.245 ;
        RECT 93.930 153.225 94.070 154.945 ;
        RECT 92.020 152.710 92.300 153.080 ;
        RECT 93.870 152.905 94.130 153.225 ;
        RECT 92.090 142.345 92.230 152.710 ;
        RECT 93.870 152.225 94.130 152.545 ;
        RECT 93.930 147.785 94.070 152.225 ;
        RECT 93.870 147.465 94.130 147.785 ;
        RECT 93.410 147.125 93.670 147.445 ;
        RECT 92.950 146.785 93.210 147.105 ;
        RECT 92.030 142.025 92.290 142.345 ;
        RECT 92.490 142.025 92.750 142.345 ;
        RECT 92.550 140.645 92.690 142.025 ;
        RECT 92.490 140.325 92.750 140.645 ;
        RECT 92.030 139.985 92.290 140.305 ;
        RECT 92.090 137.925 92.230 139.985 ;
        RECT 92.030 137.605 92.290 137.925 ;
        RECT 92.550 136.565 92.690 140.325 ;
        RECT 92.490 136.245 92.750 136.565 ;
        RECT 92.030 133.865 92.290 134.185 ;
        RECT 91.570 133.185 91.830 133.505 ;
        RECT 92.090 126.025 92.230 133.865 ;
        RECT 92.490 132.165 92.750 132.485 ;
        RECT 91.110 125.705 91.370 126.025 ;
        RECT 92.030 125.935 92.290 126.025 ;
        RECT 91.630 125.795 92.290 125.935 ;
        RECT 90.650 125.025 90.910 125.345 ;
        RECT 90.710 120.585 90.850 125.025 ;
        RECT 91.170 121.265 91.310 125.705 ;
        RECT 91.630 124.325 91.770 125.795 ;
        RECT 92.030 125.705 92.290 125.795 ;
        RECT 92.030 125.025 92.290 125.345 ;
        RECT 91.570 124.005 91.830 124.325 ;
        RECT 92.090 123.305 92.230 125.025 ;
        RECT 92.550 123.645 92.690 132.165 ;
        RECT 92.490 123.325 92.750 123.645 ;
        RECT 91.570 122.985 91.830 123.305 ;
        RECT 92.030 122.985 92.290 123.305 ;
        RECT 91.630 121.605 91.770 122.985 ;
        RECT 92.090 121.605 92.230 122.985 ;
        RECT 91.570 121.285 91.830 121.605 ;
        RECT 92.030 121.285 92.290 121.605 ;
        RECT 91.110 120.945 91.370 121.265 ;
        RECT 90.650 120.265 90.910 120.585 ;
        RECT 93.010 115.485 93.150 146.785 ;
        RECT 93.470 145.065 93.610 147.125 ;
        RECT 94.390 145.405 94.530 157.665 ;
        RECT 94.910 157.130 96.790 157.500 ;
        RECT 95.710 156.195 95.970 156.285 ;
        RECT 96.630 156.195 96.890 156.285 ;
        RECT 97.150 156.195 97.290 171.265 ;
        RECT 98.010 163.105 98.270 163.425 ;
        RECT 98.070 161.725 98.210 163.105 ;
        RECT 98.010 161.635 98.270 161.725 ;
        RECT 97.610 161.495 98.270 161.635 ;
        RECT 97.610 158.665 97.750 161.495 ;
        RECT 98.010 161.405 98.270 161.495 ;
        RECT 98.530 161.125 98.670 176.705 ;
        RECT 98.990 174.985 99.130 177.045 ;
        RECT 100.370 175.325 100.510 177.725 ;
        RECT 103.070 176.705 103.330 177.025 ;
        RECT 100.310 175.005 100.570 175.325 ;
        RECT 98.930 174.665 99.190 174.985 ;
        RECT 99.850 174.665 100.110 174.985 ;
        RECT 98.930 171.265 99.190 171.585 ;
        RECT 98.990 163.765 99.130 171.265 ;
        RECT 99.390 166.505 99.650 166.825 ;
        RECT 99.450 164.445 99.590 166.505 ;
        RECT 99.390 164.125 99.650 164.445 ;
        RECT 98.930 163.445 99.190 163.765 ;
        RECT 98.930 161.405 99.190 161.725 ;
        RECT 98.070 160.985 98.670 161.125 ;
        RECT 97.550 158.345 97.810 158.665 ;
        RECT 95.710 156.055 96.370 156.195 ;
        RECT 95.710 155.965 95.970 156.055 ;
        RECT 95.710 155.285 95.970 155.605 ;
        RECT 95.770 153.225 95.910 155.285 ;
        RECT 96.230 153.565 96.370 156.055 ;
        RECT 96.630 156.055 97.290 156.195 ;
        RECT 96.630 155.965 96.890 156.055 ;
        RECT 98.070 155.125 98.210 160.985 ;
        RECT 98.990 160.615 99.130 161.405 ;
        RECT 99.390 160.725 99.650 161.045 ;
        RECT 98.530 160.475 99.130 160.615 ;
        RECT 98.530 158.665 98.670 160.475 ;
        RECT 99.450 159.005 99.590 160.725 ;
        RECT 99.390 158.685 99.650 159.005 ;
        RECT 99.910 158.665 100.050 174.665 ;
        RECT 102.610 173.985 102.870 174.305 ;
        RECT 101.690 172.285 101.950 172.605 ;
        RECT 101.750 167.505 101.890 172.285 ;
        RECT 102.150 169.905 102.410 170.225 ;
        RECT 101.690 167.185 101.950 167.505 ;
        RECT 100.310 161.405 100.570 161.725 ;
        RECT 98.470 158.345 98.730 158.665 ;
        RECT 99.850 158.345 100.110 158.665 ;
        RECT 98.530 156.965 98.670 158.345 ;
        RECT 100.370 157.985 100.510 161.405 ;
        RECT 100.770 160.385 101.030 160.705 ;
        RECT 99.850 157.665 100.110 157.985 ;
        RECT 100.310 157.665 100.570 157.985 ;
        RECT 98.470 156.645 98.730 156.965 ;
        RECT 98.470 155.965 98.730 156.285 ;
        RECT 98.930 155.965 99.190 156.285 ;
        RECT 97.610 154.985 98.210 155.125 ;
        RECT 97.090 153.925 97.350 154.245 ;
        RECT 96.170 153.245 96.430 153.565 ;
        RECT 97.150 153.225 97.290 153.925 ;
        RECT 95.710 152.905 95.970 153.225 ;
        RECT 97.090 152.905 97.350 153.225 ;
        RECT 94.910 151.690 96.790 152.060 ;
        RECT 97.150 151.435 97.290 152.905 ;
        RECT 96.690 151.295 97.290 151.435 ;
        RECT 94.780 150.670 95.060 151.040 ;
        RECT 94.850 148.125 94.990 150.670 ;
        RECT 94.790 147.805 95.050 148.125 ;
        RECT 96.690 147.785 96.830 151.295 ;
        RECT 97.090 148.485 97.350 148.805 ;
        RECT 96.630 147.465 96.890 147.785 ;
        RECT 94.910 146.250 96.790 146.620 ;
        RECT 94.330 145.085 94.590 145.405 ;
        RECT 93.410 144.745 93.670 145.065 ;
        RECT 93.410 144.065 93.670 144.385 ;
        RECT 93.870 144.065 94.130 144.385 ;
        RECT 92.950 115.165 93.210 115.485 ;
        RECT 93.470 115.145 93.610 144.065 ;
        RECT 93.930 129.765 94.070 144.065 ;
        RECT 94.330 141.345 94.590 141.665 ;
        RECT 94.390 136.905 94.530 141.345 ;
        RECT 94.910 140.810 96.790 141.180 ;
        RECT 95.250 139.305 95.510 139.625 ;
        RECT 95.310 137.925 95.450 139.305 ;
        RECT 97.150 137.925 97.290 148.485 ;
        RECT 97.610 144.725 97.750 154.985 ;
        RECT 98.530 153.905 98.670 155.965 ;
        RECT 98.470 153.585 98.730 153.905 ;
        RECT 98.010 153.080 98.270 153.225 ;
        RECT 98.000 152.710 98.280 153.080 ;
        RECT 98.470 152.905 98.730 153.225 ;
        RECT 98.990 153.080 99.130 155.965 ;
        RECT 99.910 155.945 100.050 157.665 ;
        RECT 100.310 155.965 100.570 156.285 ;
        RECT 99.850 155.625 100.110 155.945 ;
        RECT 99.390 155.285 99.650 155.605 ;
        RECT 99.450 153.225 99.590 155.285 ;
        RECT 99.850 154.945 100.110 155.265 ;
        RECT 98.070 147.105 98.210 152.710 ;
        RECT 98.530 150.505 98.670 152.905 ;
        RECT 98.920 152.710 99.200 153.080 ;
        RECT 99.390 152.905 99.650 153.225 ;
        RECT 98.470 150.185 98.730 150.505 ;
        RECT 98.470 148.485 98.730 148.805 ;
        RECT 98.530 147.785 98.670 148.485 ;
        RECT 98.470 147.465 98.730 147.785 ;
        RECT 98.930 147.695 99.190 147.785 ;
        RECT 99.450 147.695 99.590 152.905 ;
        RECT 99.910 151.185 100.050 154.945 ;
        RECT 100.370 154.245 100.510 155.965 ;
        RECT 100.310 153.925 100.570 154.245 ;
        RECT 99.850 150.865 100.110 151.185 ;
        RECT 99.850 149.505 100.110 149.825 ;
        RECT 98.930 147.555 99.590 147.695 ;
        RECT 98.930 147.465 99.190 147.555 ;
        RECT 98.010 147.015 98.270 147.105 ;
        RECT 98.010 146.875 99.130 147.015 ;
        RECT 98.010 146.785 98.270 146.875 ;
        RECT 98.990 145.745 99.130 146.875 ;
        RECT 98.930 145.425 99.190 145.745 ;
        RECT 99.450 145.405 99.590 147.555 ;
        RECT 98.470 145.315 98.730 145.405 ;
        RECT 98.070 145.175 98.730 145.315 ;
        RECT 97.550 144.405 97.810 144.725 ;
        RECT 98.070 141.665 98.210 145.175 ;
        RECT 98.470 145.085 98.730 145.175 ;
        RECT 99.390 145.085 99.650 145.405 ;
        RECT 99.450 143.025 99.590 145.085 ;
        RECT 99.390 142.705 99.650 143.025 ;
        RECT 98.010 141.345 98.270 141.665 ;
        RECT 97.550 139.305 97.810 139.625 ;
        RECT 95.250 137.605 95.510 137.925 ;
        RECT 97.090 137.605 97.350 137.925 ;
        RECT 94.330 136.585 94.590 136.905 ;
        RECT 97.090 136.585 97.350 136.905 ;
        RECT 94.330 135.905 94.590 136.225 ;
        RECT 94.390 135.205 94.530 135.905 ;
        RECT 94.910 135.370 96.790 135.740 ;
        RECT 94.330 134.885 94.590 135.205 ;
        RECT 94.330 134.205 94.590 134.525 ;
        RECT 94.390 131.465 94.530 134.205 ;
        RECT 94.330 131.145 94.590 131.465 ;
        RECT 93.870 129.445 94.130 129.765 ;
        RECT 94.390 129.425 94.530 131.145 ;
        RECT 94.910 129.930 96.790 130.300 ;
        RECT 94.330 129.105 94.590 129.425 ;
        RECT 97.150 128.405 97.290 136.585 ;
        RECT 97.610 134.865 97.750 139.305 ;
        RECT 98.070 137.585 98.210 141.345 ;
        RECT 99.390 138.625 99.650 138.945 ;
        RECT 98.010 137.265 98.270 137.585 ;
        RECT 97.550 134.545 97.810 134.865 ;
        RECT 97.610 132.485 97.750 134.545 ;
        RECT 98.010 133.865 98.270 134.185 ;
        RECT 97.550 132.165 97.810 132.485 ;
        RECT 97.550 128.425 97.810 128.745 ;
        RECT 97.090 128.085 97.350 128.405 ;
        RECT 97.150 126.365 97.290 128.085 ;
        RECT 97.090 126.045 97.350 126.365 ;
        RECT 94.910 124.490 96.790 124.860 ;
        RECT 97.610 123.645 97.750 128.425 ;
        RECT 98.070 125.345 98.210 133.865 ;
        RECT 98.470 131.485 98.730 131.805 ;
        RECT 98.920 131.630 99.200 132.000 ;
        RECT 98.530 128.745 98.670 131.485 ;
        RECT 98.990 131.465 99.130 131.630 ;
        RECT 98.930 131.145 99.190 131.465 ;
        RECT 98.470 128.425 98.730 128.745 ;
        RECT 98.530 126.705 98.670 128.425 ;
        RECT 99.450 127.805 99.590 138.625 ;
        RECT 99.910 132.485 100.050 149.505 ;
        RECT 100.310 147.465 100.570 147.785 ;
        RECT 100.370 142.005 100.510 147.465 ;
        RECT 100.310 141.685 100.570 142.005 ;
        RECT 100.830 139.965 100.970 160.385 ;
        RECT 101.230 157.665 101.490 157.985 ;
        RECT 101.290 150.845 101.430 157.665 ;
        RECT 102.210 156.285 102.350 169.905 ;
        RECT 102.150 155.965 102.410 156.285 ;
        RECT 102.150 152.565 102.410 152.885 ;
        RECT 102.210 151.525 102.350 152.565 ;
        RECT 102.150 151.205 102.410 151.525 ;
        RECT 101.230 150.525 101.490 150.845 ;
        RECT 101.230 148.145 101.490 148.465 ;
        RECT 101.290 147.785 101.430 148.145 ;
        RECT 101.230 147.465 101.490 147.785 ;
        RECT 102.150 147.015 102.410 147.105 ;
        RECT 101.750 146.875 102.410 147.015 ;
        RECT 101.750 140.305 101.890 146.875 ;
        RECT 102.150 146.785 102.410 146.875 ;
        RECT 102.150 141.345 102.410 141.665 ;
        RECT 101.690 139.985 101.950 140.305 ;
        RECT 100.770 139.645 101.030 139.965 ;
        RECT 100.310 138.625 100.570 138.945 ;
        RECT 100.370 135.205 100.510 138.625 ;
        RECT 102.210 136.905 102.350 141.345 ;
        RECT 102.670 139.965 102.810 173.985 ;
        RECT 103.130 150.505 103.270 176.705 ;
        RECT 103.590 175.665 103.730 179.425 ;
        RECT 105.890 178.045 106.030 179.425 ;
        RECT 108.190 178.385 108.330 180.105 ;
        RECT 109.510 179.425 109.770 179.745 ;
        RECT 108.130 178.065 108.390 178.385 ;
        RECT 105.830 177.725 106.090 178.045 ;
        RECT 109.050 177.725 109.310 178.045 ;
        RECT 103.530 175.345 103.790 175.665 ;
        RECT 103.990 173.985 104.250 174.305 ;
        RECT 104.050 172.265 104.190 173.985 ;
        RECT 103.990 171.945 104.250 172.265 ;
        RECT 104.050 169.545 104.190 171.945 ;
        RECT 105.830 171.605 106.090 171.925 ;
        RECT 104.910 169.565 105.170 169.885 ;
        RECT 103.990 169.225 104.250 169.545 ;
        RECT 104.450 168.885 104.710 169.205 ;
        RECT 103.990 165.825 104.250 166.145 ;
        RECT 104.050 164.445 104.190 165.825 ;
        RECT 104.510 165.125 104.650 168.885 ;
        RECT 104.450 164.805 104.710 165.125 ;
        RECT 103.990 164.125 104.250 164.445 ;
        RECT 104.050 162.065 104.190 164.125 ;
        RECT 104.510 162.065 104.650 164.805 ;
        RECT 103.990 161.745 104.250 162.065 ;
        RECT 104.450 161.745 104.710 162.065 ;
        RECT 104.970 161.385 105.110 169.565 ;
        RECT 105.890 169.205 106.030 171.605 ;
        RECT 109.110 170.565 109.250 177.725 ;
        RECT 109.050 170.245 109.310 170.565 ;
        RECT 105.830 168.885 106.090 169.205 ;
        RECT 108.130 168.885 108.390 169.205 ;
        RECT 105.890 161.725 106.030 168.885 ;
        RECT 107.210 163.445 107.470 163.765 ;
        RECT 105.830 161.405 106.090 161.725 ;
        RECT 104.910 161.065 105.170 161.385 ;
        RECT 103.990 158.005 104.250 158.325 ;
        RECT 103.530 153.245 103.790 153.565 ;
        RECT 103.590 150.505 103.730 153.245 ;
        RECT 103.070 150.185 103.330 150.505 ;
        RECT 103.530 150.185 103.790 150.505 ;
        RECT 103.070 148.485 103.330 148.805 ;
        RECT 103.130 142.345 103.270 148.485 ;
        RECT 103.590 142.685 103.730 150.185 ;
        RECT 103.530 142.365 103.790 142.685 ;
        RECT 103.070 142.025 103.330 142.345 ;
        RECT 102.610 139.645 102.870 139.965 ;
        RECT 103.590 137.245 103.730 142.365 ;
        RECT 103.530 136.925 103.790 137.245 ;
        RECT 102.150 136.585 102.410 136.905 ;
        RECT 100.310 134.885 100.570 135.205 ;
        RECT 100.310 134.205 100.570 134.525 ;
        RECT 99.850 132.165 100.110 132.485 ;
        RECT 100.370 131.465 100.510 134.205 ;
        RECT 104.050 131.465 104.190 158.005 ;
        RECT 104.910 155.625 105.170 155.945 ;
        RECT 104.970 154.245 105.110 155.625 ;
        RECT 104.910 153.925 105.170 154.245 ;
        RECT 105.370 153.585 105.630 153.905 ;
        RECT 105.430 150.845 105.570 153.585 ;
        RECT 105.890 153.225 106.030 161.405 ;
        RECT 107.270 156.965 107.410 163.445 ;
        RECT 108.190 161.725 108.330 168.885 ;
        RECT 109.050 161.745 109.310 162.065 ;
        RECT 108.130 161.405 108.390 161.725 ;
        RECT 107.670 160.385 107.930 160.705 ;
        RECT 107.730 159.005 107.870 160.385 ;
        RECT 108.190 159.685 108.330 161.405 ;
        RECT 108.590 161.065 108.850 161.385 ;
        RECT 108.650 159.685 108.790 161.065 ;
        RECT 108.130 159.365 108.390 159.685 ;
        RECT 108.590 159.365 108.850 159.685 ;
        RECT 107.670 158.685 107.930 159.005 ;
        RECT 107.210 156.645 107.470 156.965 ;
        RECT 109.110 156.285 109.250 161.745 ;
        RECT 109.050 155.965 109.310 156.285 ;
        RECT 108.130 155.285 108.390 155.605 ;
        RECT 107.210 154.945 107.470 155.265 ;
        RECT 107.270 153.225 107.410 154.945 ;
        RECT 105.830 152.905 106.090 153.225 ;
        RECT 107.210 152.905 107.470 153.225 ;
        RECT 107.670 152.225 107.930 152.545 ;
        RECT 107.730 151.525 107.870 152.225 ;
        RECT 107.670 151.205 107.930 151.525 ;
        RECT 105.370 150.525 105.630 150.845 ;
        RECT 106.750 150.185 107.010 150.505 ;
        RECT 106.810 148.805 106.950 150.185 ;
        RECT 106.750 148.485 107.010 148.805 ;
        RECT 107.670 147.125 107.930 147.445 ;
        RECT 107.730 146.085 107.870 147.125 ;
        RECT 107.670 145.765 107.930 146.085 ;
        RECT 106.290 144.065 106.550 144.385 ;
        RECT 104.450 141.345 104.710 141.665 ;
        RECT 104.510 140.645 104.650 141.345 ;
        RECT 104.450 140.325 104.710 140.645 ;
        RECT 106.350 140.305 106.490 144.065 ;
        RECT 106.290 139.985 106.550 140.305 ;
        RECT 104.450 138.625 104.710 138.945 ;
        RECT 104.510 137.245 104.650 138.625 ;
        RECT 104.450 136.925 104.710 137.245 ;
        RECT 108.190 134.425 108.330 155.285 ;
        RECT 108.590 149.505 108.850 149.825 ;
        RECT 107.730 134.285 108.330 134.425 ;
        RECT 99.850 131.145 100.110 131.465 ;
        RECT 100.310 131.145 100.570 131.465 ;
        RECT 103.990 131.145 104.250 131.465 ;
        RECT 99.910 129.845 100.050 131.145 ;
        RECT 100.370 130.525 100.510 131.145 ;
        RECT 100.370 130.385 100.970 130.525 ;
        RECT 103.530 130.465 103.790 130.785 ;
        RECT 99.910 129.705 100.510 129.845 ;
        RECT 100.370 129.085 100.510 129.705 ;
        RECT 100.310 128.765 100.570 129.085 ;
        RECT 98.990 127.665 99.590 127.805 ;
        RECT 98.470 126.385 98.730 126.705 ;
        RECT 98.010 125.025 98.270 125.345 ;
        RECT 98.070 124.325 98.210 125.025 ;
        RECT 98.010 124.005 98.270 124.325 ;
        RECT 94.790 123.325 95.050 123.645 ;
        RECT 97.550 123.325 97.810 123.645 ;
        RECT 94.850 121.605 94.990 123.325 ;
        RECT 98.530 123.305 98.670 126.385 ;
        RECT 98.470 122.985 98.730 123.305 ;
        RECT 95.250 122.305 95.510 122.625 ;
        RECT 94.790 121.285 95.050 121.605 ;
        RECT 95.310 120.245 95.450 122.305 ;
        RECT 95.250 119.925 95.510 120.245 ;
        RECT 94.910 119.050 96.790 119.420 ;
        RECT 98.990 115.145 99.130 127.665 ;
        RECT 100.370 127.045 100.510 128.765 ;
        RECT 100.830 128.745 100.970 130.385 ;
        RECT 100.770 128.425 101.030 128.745 ;
        RECT 103.590 128.405 103.730 130.465 ;
        RECT 104.050 129.085 104.190 131.145 ;
        RECT 103.990 128.765 104.250 129.085 ;
        RECT 103.530 128.085 103.790 128.405 ;
        RECT 101.230 127.745 101.490 128.065 ;
        RECT 100.310 126.725 100.570 127.045 ;
        RECT 101.290 123.645 101.430 127.745 ;
        RECT 102.150 126.045 102.410 126.365 ;
        RECT 102.210 124.325 102.350 126.045 ;
        RECT 102.150 124.005 102.410 124.325 ;
        RECT 101.230 123.325 101.490 123.645 ;
        RECT 99.850 122.305 100.110 122.625 ;
        RECT 99.390 120.265 99.650 120.585 ;
        RECT 99.450 118.885 99.590 120.265 ;
        RECT 99.390 118.565 99.650 118.885 ;
        RECT 99.910 118.205 100.050 122.305 ;
        RECT 104.050 121.605 104.190 128.765 ;
        RECT 104.450 127.745 104.710 128.065 ;
        RECT 104.510 125.685 104.650 127.745 ;
        RECT 104.450 125.365 104.710 125.685 ;
        RECT 106.290 123.665 106.550 123.985 ;
        RECT 106.350 121.605 106.490 123.665 ;
        RECT 103.990 121.285 104.250 121.605 ;
        RECT 106.290 121.285 106.550 121.605 ;
        RECT 104.050 120.585 104.190 121.285 ;
        RECT 103.990 120.265 104.250 120.585 ;
        RECT 105.830 118.565 106.090 118.885 ;
        RECT 99.850 117.885 100.110 118.205 ;
        RECT 105.370 117.205 105.630 117.525 ;
        RECT 101.690 115.505 101.950 115.825 ;
        RECT 86.970 114.825 87.230 115.145 ;
        RECT 93.410 114.825 93.670 115.145 ;
        RECT 98.930 114.825 99.190 115.145 ;
        RECT 89.730 114.145 89.990 114.465 ;
        RECT 92.950 114.145 93.210 114.465 ;
        RECT 100.310 114.145 100.570 114.465 ;
        RECT 89.790 113.105 89.930 114.145 ;
        RECT 81.910 112.785 82.170 113.105 ;
        RECT 86.970 112.785 87.230 113.105 ;
        RECT 89.730 112.785 89.990 113.105 ;
        RECT 81.970 112.425 82.110 112.785 ;
        RECT 83.290 112.445 83.550 112.765 ;
        RECT 81.910 112.105 82.170 112.425 ;
        RECT 79.910 110.890 81.790 111.260 ;
        RECT 78.690 109.725 78.950 110.045 ;
        RECT 78.230 108.705 78.490 109.025 ;
        RECT 77.310 107.345 77.570 107.665 ;
        RECT 78.290 107.325 78.430 108.705 ;
        RECT 78.230 107.005 78.490 107.325 ;
        RECT 73.170 106.665 73.430 106.985 ;
        RECT 74.550 106.665 74.810 106.985 ;
        RECT 73.230 95.885 73.370 106.665 ;
        RECT 78.750 95.885 78.890 109.725 ;
        RECT 80.990 109.045 81.250 109.365 ;
        RECT 81.050 108.005 81.190 109.045 ;
        RECT 80.990 107.685 81.250 108.005 ;
        RECT 83.350 106.825 83.490 112.445 ;
        RECT 86.050 112.105 86.310 112.425 ;
        RECT 84.670 111.425 84.930 111.745 ;
        RECT 84.730 110.045 84.870 111.425 ;
        RECT 86.110 110.045 86.250 112.105 ;
        RECT 87.030 110.725 87.170 112.785 ;
        RECT 86.970 110.405 87.230 110.725 ;
        RECT 93.010 110.045 93.150 114.145 ;
        RECT 94.910 113.610 96.790 113.980 ;
        RECT 100.370 113.105 100.510 114.145 ;
        RECT 97.090 112.785 97.350 113.105 ;
        RECT 100.310 112.785 100.570 113.105 ;
        RECT 94.330 112.105 94.590 112.425 ;
        RECT 84.670 109.725 84.930 110.045 ;
        RECT 86.050 109.725 86.310 110.045 ;
        RECT 92.950 109.725 93.210 110.045 ;
        RECT 89.730 109.045 89.990 109.365 ;
        RECT 83.350 106.685 84.410 106.825 ;
        RECT 79.910 105.450 81.790 105.820 ;
        RECT 84.270 95.885 84.410 106.685 ;
        RECT 89.790 95.885 89.930 109.045 ;
        RECT 94.390 104.685 94.530 112.105 ;
        RECT 94.910 108.170 96.790 108.540 ;
        RECT 97.150 108.005 97.290 112.785 ;
        RECT 101.750 110.045 101.890 115.505 ;
        RECT 105.430 115.485 105.570 117.205 ;
        RECT 103.070 115.165 103.330 115.485 ;
        RECT 105.370 115.165 105.630 115.485 ;
        RECT 103.130 112.765 103.270 115.165 ;
        RECT 104.450 114.145 104.710 114.465 ;
        RECT 104.510 113.105 104.650 114.145 ;
        RECT 104.450 112.785 104.710 113.105 ;
        RECT 103.070 112.445 103.330 112.765 ;
        RECT 103.130 110.385 103.270 112.445 ;
        RECT 103.070 110.065 103.330 110.385 ;
        RECT 101.230 109.725 101.490 110.045 ;
        RECT 101.690 109.725 101.950 110.045 ;
        RECT 100.770 109.045 101.030 109.365 ;
        RECT 100.830 108.005 100.970 109.045 ;
        RECT 97.090 107.685 97.350 108.005 ;
        RECT 100.770 107.685 101.030 108.005 ;
        RECT 101.290 106.825 101.430 109.725 ;
        RECT 103.130 107.325 103.270 110.065 ;
        RECT 105.890 107.665 106.030 118.565 ;
        RECT 107.730 118.545 107.870 134.285 ;
        RECT 108.130 130.465 108.390 130.785 ;
        RECT 108.190 129.425 108.330 130.465 ;
        RECT 108.130 129.105 108.390 129.425 ;
        RECT 107.670 118.225 107.930 118.545 ;
        RECT 108.650 118.205 108.790 149.505 ;
        RECT 109.110 145.405 109.250 155.965 ;
        RECT 109.570 151.040 109.710 179.425 ;
        RECT 112.330 178.725 112.470 180.105 ;
        RECT 112.270 178.405 112.530 178.725 ;
        RECT 112.270 176.705 112.530 177.025 ;
        RECT 109.910 176.170 111.790 176.540 ;
        RECT 112.330 172.945 112.470 176.705 ;
        RECT 113.250 175.325 113.390 183.165 ;
        RECT 113.190 175.005 113.450 175.325 ;
        RECT 112.730 173.985 112.990 174.305 ;
        RECT 112.270 172.625 112.530 172.945 ;
        RECT 109.910 170.730 111.790 171.100 ;
        RECT 112.790 170.565 112.930 173.985 ;
        RECT 113.250 172.605 113.390 175.005 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 113.190 172.285 113.450 172.605 ;
        RECT 112.730 170.245 112.990 170.565 ;
        RECT 112.270 167.185 112.530 167.505 ;
        RECT 109.910 165.290 111.790 165.660 ;
        RECT 112.330 162.405 112.470 167.185 ;
        RECT 113.250 167.075 113.390 172.285 ;
        RECT 114.110 171.265 114.370 171.585 ;
        RECT 114.170 169.545 114.310 171.265 ;
        RECT 116.400 170.390 116.680 170.760 ;
        RECT 114.110 169.225 114.370 169.545 ;
        RECT 116.470 169.205 116.610 170.390 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 116.410 168.885 116.670 169.205 ;
        RECT 113.650 167.075 113.910 167.165 ;
        RECT 113.250 166.935 113.910 167.075 ;
        RECT 113.250 164.105 113.390 166.935 ;
        RECT 113.650 166.845 113.910 166.935 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 113.190 163.785 113.450 164.105 ;
        RECT 112.270 162.085 112.530 162.405 ;
        RECT 109.910 159.850 111.790 160.220 ;
        RECT 112.730 154.945 112.990 155.265 ;
        RECT 109.910 154.410 111.790 154.780 ;
        RECT 112.790 153.565 112.930 154.945 ;
        RECT 112.730 153.245 112.990 153.565 ;
        RECT 113.250 152.885 113.390 163.785 ;
        RECT 113.190 152.565 113.450 152.885 ;
        RECT 109.500 150.670 109.780 151.040 ;
        RECT 112.270 149.505 112.530 149.825 ;
        RECT 109.910 148.970 111.790 149.340 ;
        RECT 112.330 148.125 112.470 149.505 ;
        RECT 112.270 147.805 112.530 148.125 ;
        RECT 114.110 147.465 114.370 147.785 ;
        RECT 109.050 145.085 109.310 145.405 ;
        RECT 109.510 144.065 109.770 144.385 ;
        RECT 109.570 142.005 109.710 144.065 ;
        RECT 109.910 143.530 111.790 143.900 ;
        RECT 114.170 142.685 114.310 147.465 ;
        RECT 114.110 142.365 114.370 142.685 ;
        RECT 112.730 142.025 112.990 142.345 ;
        RECT 109.510 141.685 109.770 142.005 ;
        RECT 112.790 140.645 112.930 142.025 ;
        RECT 112.730 140.325 112.990 140.645 ;
        RECT 112.730 139.645 112.990 139.965 ;
        RECT 109.910 138.090 111.790 138.460 ;
        RECT 112.790 137.925 112.930 139.645 ;
        RECT 114.170 139.625 114.310 142.365 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 114.110 139.305 114.370 139.625 ;
        RECT 112.730 137.605 112.990 137.925 ;
        RECT 109.910 132.650 111.790 133.020 ;
        RECT 112.270 130.465 112.530 130.785 ;
        RECT 112.330 129.085 112.470 130.465 ;
        RECT 114.170 129.085 114.310 139.305 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 112.270 128.765 112.530 129.085 ;
        RECT 114.110 128.765 114.370 129.085 ;
        RECT 109.910 127.210 111.790 127.580 ;
        RECT 114.170 126.365 114.310 128.765 ;
        RECT 109.050 126.045 109.310 126.365 ;
        RECT 114.110 126.045 114.370 126.365 ;
        RECT 109.110 120.245 109.250 126.045 ;
        RECT 110.430 125.025 110.690 125.345 ;
        RECT 110.490 123.645 110.630 125.025 ;
        RECT 114.170 123.645 114.310 126.045 ;
        RECT 110.430 123.325 110.690 123.645 ;
        RECT 114.110 123.325 114.370 123.645 ;
        RECT 109.910 121.770 111.790 122.140 ;
        RECT 109.050 119.925 109.310 120.245 ;
        RECT 108.130 117.885 108.390 118.205 ;
        RECT 108.590 117.885 108.850 118.205 ;
        RECT 106.290 112.105 106.550 112.425 ;
        RECT 105.830 107.345 106.090 107.665 ;
        RECT 103.070 107.005 103.330 107.325 ;
        RECT 100.830 106.685 101.430 106.825 ;
        RECT 94.390 104.545 95.450 104.685 ;
        RECT 95.310 95.885 95.450 104.545 ;
        RECT 100.830 95.885 100.970 106.685 ;
        RECT 106.350 95.885 106.490 112.105 ;
        RECT 108.190 111.655 108.330 117.885 ;
        RECT 108.590 116.865 108.850 117.185 ;
        RECT 108.650 114.805 108.790 116.865 ;
        RECT 109.110 116.165 109.250 119.925 ;
        RECT 114.110 117.885 114.370 118.205 ;
        RECT 109.910 116.330 111.790 116.700 ;
        RECT 109.050 115.845 109.310 116.165 ;
        RECT 108.590 114.485 108.850 114.805 ;
        RECT 108.190 111.515 108.790 111.655 ;
        RECT 108.650 108.005 108.790 111.515 ;
        RECT 109.110 110.725 109.250 115.845 ;
        RECT 112.270 112.785 112.530 113.105 ;
        RECT 109.910 110.890 111.790 111.260 ;
        RECT 112.330 110.725 112.470 112.785 ;
        RECT 114.170 110.920 114.310 117.885 ;
        RECT 117.330 114.485 117.590 114.805 ;
        RECT 109.050 110.405 109.310 110.725 ;
        RECT 112.270 110.405 112.530 110.725 ;
        RECT 114.100 110.550 114.380 110.920 ;
        RECT 112.270 109.385 112.530 109.705 ;
        RECT 112.330 108.005 112.470 109.385 ;
        RECT 113.190 108.705 113.450 109.025 ;
        RECT 108.590 107.685 108.850 108.005 ;
        RECT 112.270 107.685 112.530 108.005 ;
        RECT 113.250 107.665 113.390 108.705 ;
        RECT 113.190 107.345 113.450 107.665 ;
        RECT 112.270 106.665 112.530 106.985 ;
        RECT 109.910 105.450 111.790 105.820 ;
        RECT 112.330 104.685 112.470 106.665 ;
        RECT 111.870 104.545 112.470 104.685 ;
        RECT 111.870 95.885 112.010 104.545 ;
        RECT 117.390 95.885 117.530 114.485 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 48.850 95.705 50.830 95.845 ;
        RECT 51.080 93.885 51.360 95.885 ;
        RECT 56.600 93.885 56.880 95.885 ;
        RECT 62.120 93.885 62.400 95.885 ;
        RECT 67.640 93.885 67.920 95.885 ;
        RECT 73.160 93.885 73.440 95.885 ;
        RECT 78.680 93.885 78.960 95.885 ;
        RECT 84.200 93.885 84.480 95.885 ;
        RECT 89.720 93.885 90.000 95.885 ;
        RECT 95.240 93.885 95.520 95.885 ;
        RECT 100.760 93.885 101.040 95.885 ;
        RECT 106.280 93.885 106.560 95.885 ;
        RECT 111.800 93.885 112.080 95.885 ;
        RECT 117.320 93.885 117.600 95.885 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 34.860 206.110 36.840 206.440 ;
        RECT 64.860 206.110 66.840 206.440 ;
        RECT 94.860 206.110 96.840 206.440 ;
        RECT 19.860 203.390 21.840 203.720 ;
        RECT 49.860 203.390 51.840 203.720 ;
        RECT 79.860 203.390 81.840 203.720 ;
        RECT 109.860 203.390 111.840 203.720 ;
        RECT 34.860 200.670 36.840 201.000 ;
        RECT 64.860 200.670 66.840 201.000 ;
        RECT 94.860 200.670 96.840 201.000 ;
        RECT 76.355 199.285 76.685 199.300 ;
        RECT 80.955 199.285 81.285 199.300 ;
        RECT 76.355 198.985 81.285 199.285 ;
        RECT 76.355 198.970 76.685 198.985 ;
        RECT 80.955 198.970 81.285 198.985 ;
        RECT 19.860 197.950 21.840 198.280 ;
        RECT 49.860 197.950 51.840 198.280 ;
        RECT 79.860 197.950 81.840 198.280 ;
        RECT 109.860 197.950 111.840 198.280 ;
        RECT 34.860 195.230 36.840 195.560 ;
        RECT 64.860 195.230 66.840 195.560 ;
        RECT 94.860 195.230 96.840 195.560 ;
        RECT 19.860 192.510 21.840 192.840 ;
        RECT 49.860 192.510 51.840 192.840 ;
        RECT 79.860 192.510 81.840 192.840 ;
        RECT 109.860 192.510 111.840 192.840 ;
        RECT 34.860 189.790 36.840 190.120 ;
        RECT 64.860 189.790 66.840 190.120 ;
        RECT 94.860 189.790 96.840 190.120 ;
        RECT 19.860 187.070 21.840 187.400 ;
        RECT 49.860 187.070 51.840 187.400 ;
        RECT 79.860 187.070 81.840 187.400 ;
        RECT 109.860 187.070 111.840 187.400 ;
        RECT 35.875 185.685 36.205 185.700 ;
        RECT 39.095 185.685 39.425 185.700 ;
        RECT 35.875 185.385 39.425 185.685 ;
        RECT 35.875 185.370 36.205 185.385 ;
        RECT 39.095 185.370 39.425 185.385 ;
        RECT 34.860 184.350 36.840 184.680 ;
        RECT 64.860 184.350 66.840 184.680 ;
        RECT 94.860 184.350 96.840 184.680 ;
        RECT 19.860 181.630 21.840 181.960 ;
        RECT 49.860 181.630 51.840 181.960 ;
        RECT 79.860 181.630 81.840 181.960 ;
        RECT 109.860 181.630 111.840 181.960 ;
        RECT 34.860 178.910 36.840 179.240 ;
        RECT 64.860 178.910 66.840 179.240 ;
        RECT 94.860 178.910 96.840 179.240 ;
        RECT 66.235 178.205 66.565 178.220 ;
        RECT 67.155 178.205 67.485 178.220 ;
        RECT 66.235 177.905 67.485 178.205 ;
        RECT 66.235 177.890 66.565 177.905 ;
        RECT 67.155 177.890 67.485 177.905 ;
        RECT 62.555 177.525 62.885 177.540 ;
        RECT 69.455 177.525 69.785 177.540 ;
        RECT 62.555 177.225 69.785 177.525 ;
        RECT 62.555 177.210 62.885 177.225 ;
        RECT 69.455 177.210 69.785 177.225 ;
        RECT 71.960 176.845 72.340 176.855 ;
        RECT 73.135 176.845 73.465 176.860 ;
        RECT 71.960 176.545 73.465 176.845 ;
        RECT 71.960 176.535 72.340 176.545 ;
        RECT 73.135 176.530 73.465 176.545 ;
        RECT 19.860 176.190 21.840 176.520 ;
        RECT 49.860 176.190 51.840 176.520 ;
        RECT 79.860 176.190 81.840 176.520 ;
        RECT 109.860 176.190 111.840 176.520 ;
        RECT 66.235 175.485 66.565 175.500 ;
        RECT 69.455 175.485 69.785 175.500 ;
        RECT 66.235 175.185 69.785 175.485 ;
        RECT 66.235 175.170 66.565 175.185 ;
        RECT 69.455 175.170 69.785 175.185 ;
        RECT 49.215 174.805 49.545 174.820 ;
        RECT 64.855 174.805 65.185 174.820 ;
        RECT 71.295 174.805 71.625 174.820 ;
        RECT 49.215 174.505 71.625 174.805 ;
        RECT 49.215 174.490 49.545 174.505 ;
        RECT 64.855 174.490 65.185 174.505 ;
        RECT 71.295 174.490 71.625 174.505 ;
        RECT 73.135 174.135 73.465 174.140 ;
        RECT 72.880 174.125 73.465 174.135 ;
        RECT 72.880 173.825 73.690 174.125 ;
        RECT 72.880 173.815 73.465 173.825 ;
        RECT 73.135 173.810 73.465 173.815 ;
        RECT 34.860 173.470 36.840 173.800 ;
        RECT 64.860 173.470 66.840 173.800 ;
        RECT 94.860 173.470 96.840 173.800 ;
        RECT 32.195 172.765 32.525 172.780 ;
        RECT 39.095 172.765 39.425 172.780 ;
        RECT 63.015 172.765 63.345 172.780 ;
        RECT 32.195 172.465 63.345 172.765 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 32.195 172.450 32.525 172.465 ;
        RECT 39.095 172.450 39.425 172.465 ;
        RECT 63.015 172.450 63.345 172.465 ;
        RECT 19.860 170.750 21.840 171.080 ;
        RECT 49.860 170.750 51.840 171.080 ;
        RECT 79.860 170.750 81.840 171.080 ;
        RECT 109.860 170.750 111.840 171.080 ;
        RECT 116.375 170.725 116.705 170.740 ;
        RECT 119.370 170.725 121.370 170.875 ;
        RECT 116.375 170.425 121.370 170.725 ;
        RECT 116.375 170.410 116.705 170.425 ;
        RECT 119.370 170.275 121.370 170.425 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 44.155 170.045 44.485 170.060 ;
        RECT 51.055 170.045 51.385 170.060 ;
        RECT 44.155 169.745 51.385 170.045 ;
        RECT 44.155 169.730 44.485 169.745 ;
        RECT 51.055 169.730 51.385 169.745 ;
        RECT 34.860 168.030 36.840 168.360 ;
        RECT 64.860 168.030 66.840 168.360 ;
        RECT 94.860 168.030 96.840 168.360 ;
        RECT 79.115 167.325 79.445 167.340 ;
        RECT 86.680 167.325 87.060 167.335 ;
        RECT 90.615 167.325 90.945 167.340 ;
        RECT 79.115 167.025 90.945 167.325 ;
        RECT 79.115 167.010 79.445 167.025 ;
        RECT 86.680 167.015 87.060 167.025 ;
        RECT 90.615 167.010 90.945 167.025 ;
        RECT 40.935 166.645 41.265 166.660 ;
        RECT 41.600 166.645 41.980 166.655 ;
        RECT 40.935 166.345 41.980 166.645 ;
        RECT 40.935 166.330 41.265 166.345 ;
        RECT 41.600 166.335 41.980 166.345 ;
        RECT 19.860 165.310 21.840 165.640 ;
        RECT 49.860 165.310 51.840 165.640 ;
        RECT 79.860 165.310 81.840 165.640 ;
        RECT 109.860 165.310 111.840 165.640 ;
        RECT 36.795 164.605 37.125 164.620 ;
        RECT 39.095 164.605 39.425 164.620 ;
        RECT 42.775 164.605 43.105 164.620 ;
        RECT 36.795 164.305 43.105 164.605 ;
        RECT 36.795 164.290 37.125 164.305 ;
        RECT 39.095 164.290 39.425 164.305 ;
        RECT 42.775 164.290 43.105 164.305 ;
        RECT 54.735 163.925 55.065 163.940 ;
        RECT 79.115 163.925 79.445 163.940 ;
        RECT 54.735 163.625 79.445 163.925 ;
        RECT 54.735 163.610 55.065 163.625 ;
        RECT 79.115 163.610 79.445 163.625 ;
        RECT 34.860 162.590 36.840 162.920 ;
        RECT 64.860 162.590 66.840 162.920 ;
        RECT 94.860 162.590 96.840 162.920 ;
        RECT 64.395 161.205 64.725 161.220 ;
        RECT 67.155 161.215 67.485 161.220 ;
        RECT 67.155 161.205 67.740 161.215 ;
        RECT 64.395 160.905 67.740 161.205 ;
        RECT 64.395 160.890 64.725 160.905 ;
        RECT 67.155 160.895 67.740 160.905 ;
        RECT 67.155 160.890 67.485 160.895 ;
        RECT 59.795 160.525 60.125 160.540 ;
        RECT 70.835 160.525 71.165 160.540 ;
        RECT 59.795 160.225 71.165 160.525 ;
        RECT 59.795 160.210 60.125 160.225 ;
        RECT 70.835 160.210 71.165 160.225 ;
        RECT 19.860 159.870 21.840 160.200 ;
        RECT 49.860 159.870 51.840 160.200 ;
        RECT 79.860 159.870 81.840 160.200 ;
        RECT 109.860 159.870 111.840 160.200 ;
        RECT 41.600 159.165 41.980 159.175 ;
        RECT 54.735 159.165 55.065 159.180 ;
        RECT 41.600 158.865 55.065 159.165 ;
        RECT 41.600 158.855 41.980 158.865 ;
        RECT 54.735 158.850 55.065 158.865 ;
        RECT 50.595 158.485 50.925 158.500 ;
        RECT 70.375 158.485 70.705 158.500 ;
        RECT 50.595 158.185 70.705 158.485 ;
        RECT 50.595 158.170 50.925 158.185 ;
        RECT 70.375 158.170 70.705 158.185 ;
        RECT 34.860 157.150 36.840 157.480 ;
        RECT 64.860 157.150 66.840 157.480 ;
        RECT 94.860 157.150 96.840 157.480 ;
        RECT 63.475 156.445 63.805 156.460 ;
        RECT 104.160 156.445 104.540 156.455 ;
        RECT 63.475 156.145 104.540 156.445 ;
        RECT 63.475 156.130 63.805 156.145 ;
        RECT 104.160 156.135 104.540 156.145 ;
        RECT 66.695 155.765 67.025 155.780 ;
        RECT 74.055 155.765 74.385 155.780 ;
        RECT 66.695 155.465 74.385 155.765 ;
        RECT 66.695 155.450 67.025 155.465 ;
        RECT 74.055 155.450 74.385 155.465 ;
        RECT 67.360 155.085 67.740 155.095 ;
        RECT 68.075 155.085 68.405 155.100 ;
        RECT 70.375 155.085 70.705 155.100 ;
        RECT 67.360 154.785 70.705 155.085 ;
        RECT 67.360 154.775 67.740 154.785 ;
        RECT 68.075 154.770 68.405 154.785 ;
        RECT 70.375 154.770 70.705 154.785 ;
        RECT 19.860 154.430 21.840 154.760 ;
        RECT 49.860 154.430 51.840 154.760 ;
        RECT 79.860 154.430 81.840 154.760 ;
        RECT 109.860 154.430 111.840 154.760 ;
        RECT 29.435 153.045 29.765 153.060 ;
        RECT 36.795 153.045 37.125 153.060 ;
        RECT 29.435 152.745 37.125 153.045 ;
        RECT 29.435 152.730 29.765 152.745 ;
        RECT 36.795 152.730 37.125 152.745 ;
        RECT 59.335 153.045 59.665 153.060 ;
        RECT 75.435 153.045 75.765 153.060 ;
        RECT 91.995 153.045 92.325 153.060 ;
        RECT 97.975 153.045 98.305 153.060 ;
        RECT 98.895 153.045 99.225 153.060 ;
        RECT 59.335 152.745 99.225 153.045 ;
        RECT 59.335 152.730 59.665 152.745 ;
        RECT 75.435 152.730 75.765 152.745 ;
        RECT 91.995 152.730 92.325 152.745 ;
        RECT 97.975 152.730 98.305 152.745 ;
        RECT 98.895 152.730 99.225 152.745 ;
        RECT 41.855 152.365 42.185 152.380 ;
        RECT 60.000 152.365 60.380 152.375 ;
        RECT 41.855 152.065 60.380 152.365 ;
        RECT 41.855 152.050 42.185 152.065 ;
        RECT 60.000 152.055 60.380 152.065 ;
        RECT 34.860 151.710 36.840 152.040 ;
        RECT 64.860 151.710 66.840 152.040 ;
        RECT 94.860 151.710 96.840 152.040 ;
        RECT 33.575 151.005 33.905 151.020 ;
        RECT 36.795 151.005 37.125 151.020 ;
        RECT 57.955 151.005 58.285 151.020 ;
        RECT 33.575 150.705 58.285 151.005 ;
        RECT 33.575 150.690 33.905 150.705 ;
        RECT 36.795 150.690 37.125 150.705 ;
        RECT 57.955 150.690 58.285 150.705 ;
        RECT 94.755 151.005 95.085 151.020 ;
        RECT 109.475 151.005 109.805 151.020 ;
        RECT 94.755 150.705 109.805 151.005 ;
        RECT 94.755 150.690 95.085 150.705 ;
        RECT 109.475 150.690 109.805 150.705 ;
        RECT 19.860 148.990 21.840 149.320 ;
        RECT 49.860 148.990 51.840 149.320 ;
        RECT 79.860 148.990 81.840 149.320 ;
        RECT 109.860 148.990 111.840 149.320 ;
        RECT 46.455 148.285 46.785 148.300 ;
        RECT 50.595 148.285 50.925 148.300 ;
        RECT 46.455 147.985 50.925 148.285 ;
        RECT 46.455 147.970 46.785 147.985 ;
        RECT 50.595 147.970 50.925 147.985 ;
        RECT 71.755 148.285 72.085 148.300 ;
        RECT 72.880 148.285 73.260 148.295 ;
        RECT 71.755 147.985 73.260 148.285 ;
        RECT 71.755 147.970 72.085 147.985 ;
        RECT 72.880 147.975 73.260 147.985 ;
        RECT 48.755 147.605 49.085 147.620 ;
        RECT 51.515 147.605 51.845 147.620 ;
        RECT 66.695 147.605 67.025 147.620 ;
        RECT 48.755 147.305 67.025 147.605 ;
        RECT 48.755 147.290 49.085 147.305 ;
        RECT 51.515 147.290 51.845 147.305 ;
        RECT 66.695 147.290 67.025 147.305 ;
        RECT 34.860 146.270 36.840 146.600 ;
        RECT 64.860 146.270 66.840 146.600 ;
        RECT 94.860 146.270 96.840 146.600 ;
        RECT 19.860 143.550 21.840 143.880 ;
        RECT 49.860 143.550 51.840 143.880 ;
        RECT 79.860 143.550 81.840 143.880 ;
        RECT 109.860 143.550 111.840 143.880 ;
        RECT 34.860 140.830 36.840 141.160 ;
        RECT 64.860 140.830 66.840 141.160 ;
        RECT 94.860 140.830 96.840 141.160 ;
        RECT 71.755 140.815 72.085 140.820 ;
        RECT 71.755 140.805 72.340 140.815 ;
        RECT 104.160 140.805 104.540 140.815 ;
        RECT 119.370 140.805 121.370 140.955 ;
        RECT 71.755 140.505 72.540 140.805 ;
        RECT 104.160 140.505 121.370 140.805 ;
        RECT 71.755 140.495 72.340 140.505 ;
        RECT 104.160 140.495 104.540 140.505 ;
        RECT 71.755 140.490 72.085 140.495 ;
        RECT 119.370 140.355 121.370 140.505 ;
        RECT 19.860 138.110 21.840 138.440 ;
        RECT 49.860 138.110 51.840 138.440 ;
        RECT 79.860 138.110 81.840 138.440 ;
        RECT 109.860 138.110 111.840 138.440 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 34.860 135.390 36.840 135.720 ;
        RECT 64.860 135.390 66.840 135.720 ;
        RECT 94.860 135.390 96.840 135.720 ;
        RECT 19.860 132.670 21.840 133.000 ;
        RECT 49.860 132.670 51.840 133.000 ;
        RECT 79.860 132.670 81.840 133.000 ;
        RECT 109.860 132.670 111.840 133.000 ;
        RECT 84.635 131.965 84.965 131.980 ;
        RECT 86.680 131.965 87.060 131.975 ;
        RECT 98.895 131.965 99.225 131.980 ;
        RECT 84.635 131.665 99.225 131.965 ;
        RECT 84.635 131.650 84.965 131.665 ;
        RECT 86.680 131.655 87.060 131.665 ;
        RECT 98.895 131.650 99.225 131.665 ;
        RECT 34.860 129.950 36.840 130.280 ;
        RECT 64.860 129.950 66.840 130.280 ;
        RECT 94.860 129.950 96.840 130.280 ;
        RECT 41.395 129.935 41.725 129.940 ;
        RECT 41.395 129.925 41.980 129.935 ;
        RECT 41.170 129.625 41.980 129.925 ;
        RECT 41.395 129.615 41.980 129.625 ;
        RECT 41.395 129.610 41.725 129.615 ;
        RECT 19.860 127.230 21.840 127.560 ;
        RECT 49.860 127.230 51.840 127.560 ;
        RECT 79.860 127.230 81.840 127.560 ;
        RECT 109.860 127.230 111.840 127.560 ;
        RECT 34.860 124.510 36.840 124.840 ;
        RECT 64.860 124.510 66.840 124.840 ;
        RECT 94.860 124.510 96.840 124.840 ;
        RECT 19.860 121.790 21.840 122.120 ;
        RECT 49.860 121.790 51.840 122.120 ;
        RECT 79.860 121.790 81.840 122.120 ;
        RECT 109.860 121.790 111.840 122.120 ;
        RECT 34.860 119.070 36.840 119.400 ;
        RECT 64.860 119.070 66.840 119.400 ;
        RECT 94.860 119.070 96.840 119.400 ;
        RECT 19.860 116.350 21.840 116.680 ;
        RECT 49.860 116.350 51.840 116.680 ;
        RECT 79.860 116.350 81.840 116.680 ;
        RECT 109.860 116.350 111.840 116.680 ;
        RECT 34.860 113.630 36.840 113.960 ;
        RECT 64.860 113.630 66.840 113.960 ;
        RECT 94.860 113.630 96.840 113.960 ;
        RECT 59.795 113.615 60.125 113.620 ;
        RECT 59.795 113.605 60.380 113.615 ;
        RECT 59.795 113.305 60.580 113.605 ;
        RECT 59.795 113.295 60.380 113.305 ;
        RECT 59.795 113.290 60.125 113.295 ;
        RECT 19.860 110.910 21.840 111.240 ;
        RECT 49.860 110.910 51.840 111.240 ;
        RECT 79.860 110.910 81.840 111.240 ;
        RECT 109.860 110.910 111.840 111.240 ;
        RECT 114.075 110.885 114.405 110.900 ;
        RECT 119.370 110.885 121.370 111.035 ;
        RECT 114.075 110.585 121.370 110.885 ;
        RECT 114.075 110.570 114.405 110.585 ;
        RECT 119.370 110.435 121.370 110.585 ;
        RECT 34.860 108.190 36.840 108.520 ;
        RECT 64.860 108.190 66.840 108.520 ;
        RECT 94.860 108.190 96.840 108.520 ;
        RECT 19.860 105.470 21.840 105.800 ;
        RECT 49.860 105.470 51.840 105.800 ;
        RECT 79.860 105.470 81.840 105.800 ;
        RECT 109.860 105.470 111.840 105.800 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 19.850 105.395 21.850 206.515 ;
        RECT 34.850 105.395 36.850 206.515 ;
        RECT 41.625 166.330 41.955 166.660 ;
        RECT 41.640 159.180 41.940 166.330 ;
        RECT 41.625 158.850 41.955 159.180 ;
        RECT 41.640 129.940 41.940 158.850 ;
        RECT 41.625 129.610 41.955 129.940 ;
        RECT 49.850 105.395 51.850 206.515 ;
        RECT 60.025 152.050 60.355 152.380 ;
        RECT 60.040 113.620 60.340 152.050 ;
        RECT 60.025 113.290 60.355 113.620 ;
        RECT 64.850 105.395 66.850 206.515 ;
        RECT 71.985 176.530 72.315 176.860 ;
        RECT 67.385 160.890 67.715 161.220 ;
        RECT 67.400 155.100 67.700 160.890 ;
        RECT 67.385 154.770 67.715 155.100 ;
        RECT 72.000 140.820 72.300 176.530 ;
        RECT 72.905 173.810 73.235 174.140 ;
        RECT 72.920 148.300 73.220 173.810 ;
        RECT 72.905 147.970 73.235 148.300 ;
        RECT 71.985 140.490 72.315 140.820 ;
        RECT 79.850 105.395 81.850 206.515 ;
        RECT 86.705 167.010 87.035 167.340 ;
        RECT 86.720 131.980 87.020 167.010 ;
        RECT 86.705 131.650 87.035 131.980 ;
        RECT 94.850 105.395 96.850 206.515 ;
        RECT 104.185 156.130 104.515 156.460 ;
        RECT 104.200 140.820 104.500 156.130 ;
        RECT 104.185 140.490 104.515 140.820 ;
        RECT 109.850 105.395 111.850 206.515 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

