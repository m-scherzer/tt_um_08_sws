MACRO digital_top
  CLASS BLOCK ;
  FOREIGN digital_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 129.675 BY 140.395 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.520 10.640 26.520 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.520 10.640 86.520 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.520 10.640 116.520 128.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.520 10.640 11.520 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.520 10.640 41.520 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 10.640 71.520 128.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.520 10.640 101.520 128.080 ;
    END
  END VPWR
  PIN i_dem_dis
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 2.000 120.320 ;
    END
  END i_dem_dis
  PIN i_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.000 52.320 ;
    END
  END i_reset
  PIN i_sys_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END i_sys_clk
  PIN o_cs_cell_hi[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 3.310 138.395 3.590 140.395 ;
    END
  END o_cs_cell_hi[0]
  PIN o_cs_cell_hi[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 138.395 10.030 140.395 ;
    END
  END o_cs_cell_hi[1]
  PIN o_cs_cell_hi[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 138.395 16.470 140.395 ;
    END
  END o_cs_cell_hi[2]
  PIN o_cs_cell_hi[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 138.395 22.910 140.395 ;
    END
  END o_cs_cell_hi[3]
  PIN o_cs_cell_hi[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 138.395 29.350 140.395 ;
    END
  END o_cs_cell_hi[4]
  PIN o_cs_cell_hi[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 138.395 35.790 140.395 ;
    END
  END o_cs_cell_hi[5]
  PIN o_cs_cell_hi[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 138.395 42.230 140.395 ;
    END
  END o_cs_cell_hi[6]
  PIN o_cs_cell_hi[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 138.395 48.670 140.395 ;
    END
  END o_cs_cell_hi[7]
  PIN o_cs_cell_hi[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 138.395 55.110 140.395 ;
    END
  END o_cs_cell_hi[8]
  PIN o_cs_cell_hi[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 138.395 61.550 140.395 ;
    END
  END o_cs_cell_hi[9]
  PIN o_cs_cell_lo[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 138.395 67.990 140.395 ;
    END
  END o_cs_cell_lo[0]
  PIN o_cs_cell_lo[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 138.395 74.430 140.395 ;
    END
  END o_cs_cell_lo[1]
  PIN o_cs_cell_lo[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 138.395 80.870 140.395 ;
    END
  END o_cs_cell_lo[2]
  PIN o_cs_cell_lo[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 138.395 87.310 140.395 ;
    END
  END o_cs_cell_lo[3]
  PIN o_cs_cell_lo[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 138.395 93.750 140.395 ;
    END
  END o_cs_cell_lo[4]
  PIN o_cs_cell_lo[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 138.395 100.190 140.395 ;
    END
  END o_cs_cell_lo[5]
  PIN o_cs_cell_lo[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 138.395 106.630 140.395 ;
    END
  END o_cs_cell_lo[6]
  PIN o_cs_cell_lo[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 138.395 113.070 140.395 ;
    END
  END o_cs_cell_lo[7]
  PIN o_cs_cell_lo[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 138.395 119.510 140.395 ;
    END
  END o_cs_cell_lo[8]
  PIN o_cs_cell_lo[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 138.395 125.950 140.395 ;
    END
  END o_cs_cell_lo[9]
  OBS
      LAYER nwell ;
        RECT 5.330 126.425 123.930 128.030 ;
      LAYER pwell ;
        RECT 5.525 125.225 6.895 126.035 ;
        RECT 6.905 125.225 12.415 126.035 ;
        RECT 12.425 125.225 17.935 126.035 ;
        RECT 18.415 125.310 18.845 126.095 ;
        RECT 18.865 125.225 24.375 126.035 ;
        RECT 24.385 125.225 29.895 126.035 ;
        RECT 29.905 125.225 31.275 126.035 ;
        RECT 31.295 125.310 31.725 126.095 ;
        RECT 31.745 125.225 37.255 126.035 ;
        RECT 37.265 125.225 42.775 126.035 ;
        RECT 42.785 125.225 44.155 126.035 ;
        RECT 44.175 125.310 44.605 126.095 ;
        RECT 44.625 125.225 50.135 126.035 ;
        RECT 50.145 125.225 55.655 126.035 ;
        RECT 55.665 125.225 57.035 126.035 ;
        RECT 57.055 125.310 57.485 126.095 ;
        RECT 57.505 125.225 63.015 126.035 ;
        RECT 63.025 125.225 68.535 126.035 ;
        RECT 68.545 125.225 69.915 126.035 ;
        RECT 69.935 125.310 70.365 126.095 ;
        RECT 70.385 125.225 75.895 126.035 ;
        RECT 75.905 125.225 81.415 126.035 ;
        RECT 81.425 125.225 82.795 126.035 ;
        RECT 82.815 125.310 83.245 126.095 ;
        RECT 83.265 125.225 88.775 126.035 ;
        RECT 88.785 125.225 94.295 126.035 ;
        RECT 94.305 125.225 95.675 126.035 ;
        RECT 95.695 125.310 96.125 126.095 ;
        RECT 96.145 125.225 101.655 126.035 ;
        RECT 101.665 125.225 107.175 126.035 ;
        RECT 107.185 125.225 108.555 126.035 ;
        RECT 108.575 125.310 109.005 126.095 ;
        RECT 109.025 125.225 111.775 126.035 ;
        RECT 116.755 125.905 117.685 126.125 ;
        RECT 120.515 125.905 121.435 126.135 ;
        RECT 112.245 125.225 121.435 125.905 ;
        RECT 121.455 125.310 121.885 126.095 ;
        RECT 122.365 125.225 123.735 126.035 ;
        RECT 5.665 125.015 5.835 125.225 ;
        RECT 7.045 125.205 7.215 125.225 ;
        RECT 7.045 125.035 7.225 125.205 ;
        RECT 7.055 125.015 7.225 125.035 ;
        RECT 8.425 125.015 8.595 125.205 ;
        RECT 12.100 125.065 12.220 125.175 ;
        RECT 12.565 125.035 12.735 125.225 ;
        RECT 18.080 125.065 18.200 125.175 ;
        RECT 19.005 125.035 19.175 125.225 ;
        RECT 21.305 125.015 21.475 125.205 ;
        RECT 21.765 125.015 21.935 125.205 ;
        RECT 24.525 125.035 24.695 125.225 ;
        RECT 25.440 125.065 25.560 125.175 ;
        RECT 25.905 125.015 26.075 125.205 ;
        RECT 27.285 125.015 27.455 125.205 ;
        RECT 29.120 125.065 29.240 125.175 ;
        RECT 29.585 125.015 29.755 125.205 ;
        RECT 30.045 125.035 30.215 125.225 ;
        RECT 30.960 125.065 31.080 125.175 ;
        RECT 31.885 125.015 32.055 125.225 ;
        RECT 37.405 125.015 37.575 125.225 ;
        RECT 38.785 125.015 38.955 125.205 ;
        RECT 42.925 125.035 43.095 125.225 ;
        RECT 44.765 125.035 44.935 125.225 ;
        RECT 47.985 125.015 48.155 125.205 ;
        RECT 50.285 125.035 50.455 125.225 ;
        RECT 55.805 125.035 55.975 125.225 ;
        RECT 57.645 125.015 57.815 125.225 ;
        RECT 63.165 125.035 63.335 125.225 ;
        RECT 66.840 125.065 66.960 125.175 ;
        RECT 67.305 125.015 67.475 125.205 ;
        RECT 68.685 125.035 68.855 125.225 ;
        RECT 70.525 125.035 70.695 125.225 ;
        RECT 76.045 125.035 76.215 125.225 ;
        RECT 76.505 125.015 76.675 125.205 ;
        RECT 81.565 125.035 81.735 125.225 ;
        RECT 82.035 125.060 82.195 125.170 ;
        RECT 83.405 125.015 83.575 125.225 ;
        RECT 88.925 125.035 89.095 125.225 ;
        RECT 94.445 125.035 94.615 125.225 ;
        RECT 96.285 125.035 96.455 125.225 ;
        RECT 101.345 125.015 101.515 125.205 ;
        RECT 101.805 125.015 101.975 125.225 ;
        RECT 107.325 125.015 107.495 125.225 ;
        RECT 109.165 125.035 109.335 125.225 ;
        RECT 111.920 125.065 112.040 125.175 ;
        RECT 112.385 125.035 112.555 125.225 ;
        RECT 117.905 125.015 118.075 125.205 ;
        RECT 118.365 125.015 118.535 125.205 ;
        RECT 122.040 125.065 122.160 125.175 ;
        RECT 123.425 125.015 123.595 125.225 ;
        RECT 5.525 124.205 6.895 125.015 ;
        RECT 6.905 124.235 8.275 125.015 ;
        RECT 8.285 124.205 11.955 125.015 ;
        RECT 12.425 124.335 21.615 125.015 ;
        RECT 12.425 124.105 13.345 124.335 ;
        RECT 16.175 124.115 17.105 124.335 ;
        RECT 21.625 124.205 25.295 125.015 ;
        RECT 25.775 124.105 27.125 125.015 ;
        RECT 27.145 124.205 28.975 125.015 ;
        RECT 29.455 124.105 30.805 125.015 ;
        RECT 31.295 124.145 31.725 124.930 ;
        RECT 31.745 124.205 37.255 125.015 ;
        RECT 37.265 124.205 38.635 125.015 ;
        RECT 38.645 124.335 47.835 125.015 ;
        RECT 47.845 124.335 57.035 125.015 ;
        RECT 43.155 124.115 44.085 124.335 ;
        RECT 46.915 124.105 47.835 124.335 ;
        RECT 52.355 124.115 53.285 124.335 ;
        RECT 56.115 124.105 57.035 124.335 ;
        RECT 57.055 124.145 57.485 124.930 ;
        RECT 57.505 124.335 66.695 125.015 ;
        RECT 67.165 124.335 76.355 125.015 ;
        RECT 62.015 124.115 62.945 124.335 ;
        RECT 65.775 124.105 66.695 124.335 ;
        RECT 71.675 124.115 72.605 124.335 ;
        RECT 75.435 124.105 76.355 124.335 ;
        RECT 76.365 124.205 81.875 125.015 ;
        RECT 82.815 124.145 83.245 124.930 ;
        RECT 83.265 124.335 92.455 125.015 ;
        RECT 87.775 124.115 88.705 124.335 ;
        RECT 91.535 124.105 92.455 124.335 ;
        RECT 92.465 124.335 101.655 125.015 ;
        RECT 92.465 124.105 93.385 124.335 ;
        RECT 96.215 124.115 97.145 124.335 ;
        RECT 101.665 124.205 107.175 125.015 ;
        RECT 107.185 124.205 108.555 125.015 ;
        RECT 108.575 124.145 109.005 124.930 ;
        RECT 109.025 124.335 118.215 125.015 ;
        RECT 109.025 124.105 109.945 124.335 ;
        RECT 112.775 124.115 113.705 124.335 ;
        RECT 118.225 124.205 121.895 125.015 ;
        RECT 122.365 124.205 123.735 125.015 ;
      LAYER nwell ;
        RECT 5.330 120.985 123.930 123.815 ;
      LAYER pwell ;
        RECT 5.525 119.785 6.895 120.595 ;
        RECT 11.415 120.465 12.345 120.685 ;
        RECT 15.175 120.465 16.095 120.695 ;
        RECT 6.905 119.785 16.095 120.465 ;
        RECT 16.115 119.785 17.465 120.695 ;
        RECT 18.415 119.870 18.845 120.655 ;
        RECT 18.875 119.785 20.225 120.695 ;
        RECT 20.245 119.785 23.915 120.595 ;
        RECT 28.895 120.465 29.825 120.685 ;
        RECT 32.655 120.465 33.575 120.695 ;
        RECT 24.385 119.785 33.575 120.465 ;
        RECT 33.595 119.785 34.945 120.695 ;
        RECT 39.475 120.465 40.405 120.685 ;
        RECT 43.235 120.465 44.155 120.695 ;
        RECT 34.965 119.785 44.155 120.465 ;
        RECT 44.175 119.870 44.605 120.655 ;
        RECT 44.635 119.785 45.985 120.695 ;
        RECT 46.925 119.785 48.295 120.565 ;
        RECT 48.315 119.785 49.665 120.695 ;
        RECT 49.685 119.785 53.355 120.595 ;
        RECT 53.365 119.785 54.735 120.565 ;
        RECT 54.745 119.785 56.115 120.565 ;
        RECT 56.135 119.785 57.485 120.695 ;
        RECT 57.515 119.785 58.865 120.695 ;
        RECT 58.885 119.785 64.395 120.595 ;
        RECT 64.405 119.785 69.915 120.595 ;
        RECT 69.935 119.870 70.365 120.655 ;
        RECT 71.315 119.785 72.665 120.695 ;
        RECT 72.695 119.785 74.045 120.695 ;
        RECT 79.035 120.465 79.965 120.685 ;
        RECT 82.795 120.465 83.715 120.695 ;
        RECT 74.525 119.785 83.715 120.465 ;
        RECT 83.735 119.785 85.085 120.695 ;
        RECT 85.105 119.785 87.855 120.595 ;
        RECT 87.865 119.785 89.235 120.565 ;
        RECT 89.255 119.785 90.605 120.695 ;
        RECT 90.625 119.785 92.455 120.595 ;
        RECT 92.475 119.785 93.825 120.695 ;
        RECT 93.845 119.785 95.675 120.595 ;
        RECT 95.695 119.870 96.125 120.655 ;
        RECT 100.655 120.465 101.585 120.685 ;
        RECT 104.415 120.465 105.335 120.695 ;
        RECT 96.145 119.785 105.335 120.465 ;
        RECT 105.355 119.785 106.705 120.695 ;
        RECT 111.235 120.465 112.165 120.685 ;
        RECT 114.995 120.465 115.915 120.695 ;
        RECT 106.725 119.785 115.915 120.465 ;
        RECT 115.935 119.785 117.285 120.695 ;
        RECT 117.315 119.785 118.665 120.695 ;
        RECT 118.685 119.785 121.435 120.595 ;
        RECT 121.455 119.870 121.885 120.655 ;
        RECT 122.365 119.785 123.735 120.595 ;
        RECT 5.665 119.575 5.835 119.785 ;
        RECT 7.045 119.595 7.215 119.785 ;
        RECT 16.705 119.575 16.875 119.765 ;
        RECT 17.165 119.595 17.335 119.785 ;
        RECT 17.635 119.630 17.795 119.740 ;
        RECT 18.085 119.575 18.255 119.765 ;
        RECT 18.555 119.620 18.715 119.730 ;
        RECT 19.925 119.595 20.095 119.785 ;
        RECT 20.385 119.575 20.555 119.785 ;
        RECT 24.060 119.625 24.180 119.735 ;
        RECT 24.525 119.595 24.695 119.785 ;
        RECT 29.585 119.575 29.755 119.765 ;
        RECT 30.965 119.575 31.135 119.765 ;
        RECT 31.885 119.575 32.055 119.765 ;
        RECT 33.725 119.595 33.895 119.785 ;
        RECT 35.105 119.595 35.275 119.785 ;
        RECT 41.080 119.625 41.200 119.735 ;
        RECT 42.465 119.575 42.635 119.765 ;
        RECT 42.925 119.575 43.095 119.765 ;
        RECT 45.685 119.595 45.855 119.785 ;
        RECT 46.155 119.630 46.315 119.740 ;
        RECT 47.985 119.595 48.155 119.785 ;
        RECT 48.440 119.625 48.560 119.735 ;
        RECT 49.365 119.595 49.535 119.785 ;
        RECT 49.825 119.595 49.995 119.785 ;
        RECT 51.200 119.575 51.370 119.765 ;
        RECT 51.665 119.575 51.835 119.765 ;
        RECT 54.425 119.595 54.595 119.785 ;
        RECT 54.885 119.595 55.055 119.785 ;
        RECT 56.265 119.595 56.435 119.785 ;
        RECT 57.645 119.575 57.815 119.785 ;
        RECT 59.025 119.575 59.195 119.785 ;
        RECT 60.405 119.575 60.575 119.765 ;
        RECT 64.080 119.625 64.200 119.735 ;
        RECT 64.545 119.595 64.715 119.785 ;
        RECT 70.535 119.630 70.695 119.740 ;
        RECT 72.365 119.595 72.535 119.785 ;
        RECT 73.745 119.765 73.915 119.785 ;
        RECT 73.285 119.575 73.455 119.765 ;
        RECT 73.745 119.595 73.920 119.765 ;
        RECT 74.200 119.625 74.320 119.735 ;
        RECT 74.665 119.595 74.835 119.785 ;
        RECT 73.750 119.575 73.920 119.595 ;
        RECT 76.505 119.575 76.675 119.765 ;
        RECT 80.185 119.575 80.355 119.765 ;
        RECT 80.645 119.575 80.815 119.765 ;
        RECT 82.480 119.625 82.600 119.735 ;
        RECT 83.405 119.575 83.575 119.765 ;
        RECT 84.785 119.595 84.955 119.785 ;
        RECT 85.245 119.595 85.415 119.785 ;
        RECT 88.925 119.575 89.095 119.785 ;
        RECT 90.305 119.595 90.475 119.785 ;
        RECT 90.765 119.735 90.935 119.785 ;
        RECT 90.760 119.625 90.935 119.735 ;
        RECT 90.765 119.595 90.935 119.625 ;
        RECT 91.225 119.575 91.395 119.765 ;
        RECT 92.605 119.575 92.775 119.785 ;
        RECT 93.985 119.595 94.155 119.785 ;
        RECT 95.360 119.625 95.480 119.735 ;
        RECT 95.825 119.575 95.995 119.765 ;
        RECT 96.285 119.595 96.455 119.785 ;
        RECT 97.205 119.575 97.375 119.765 ;
        RECT 99.045 119.575 99.215 119.765 ;
        RECT 100.425 119.575 100.595 119.765 ;
        RECT 102.265 119.575 102.435 119.765 ;
        RECT 103.645 119.575 103.815 119.765 ;
        RECT 105.485 119.735 105.655 119.785 ;
        RECT 105.480 119.625 105.655 119.735 ;
        RECT 105.485 119.595 105.655 119.625 ;
        RECT 105.945 119.575 106.115 119.765 ;
        RECT 106.865 119.595 107.035 119.785 ;
        RECT 107.325 119.575 107.495 119.765 ;
        RECT 109.165 119.575 109.335 119.765 ;
        RECT 116.985 119.595 117.155 119.785 ;
        RECT 117.445 119.595 117.615 119.785 ;
        RECT 118.365 119.575 118.535 119.765 ;
        RECT 118.825 119.595 118.995 119.785 ;
        RECT 122.040 119.625 122.160 119.735 ;
        RECT 123.425 119.575 123.595 119.785 ;
        RECT 5.525 118.765 6.895 119.575 ;
        RECT 7.825 118.895 17.015 119.575 ;
        RECT 7.825 118.665 8.745 118.895 ;
        RECT 11.575 118.675 12.505 118.895 ;
        RECT 17.035 118.665 18.385 119.575 ;
        RECT 19.325 118.795 20.695 119.575 ;
        RECT 20.705 118.895 29.895 119.575 ;
        RECT 20.705 118.665 21.625 118.895 ;
        RECT 24.455 118.675 25.385 118.895 ;
        RECT 29.905 118.795 31.275 119.575 ;
        RECT 31.295 118.705 31.725 119.490 ;
        RECT 31.745 118.895 40.935 119.575 ;
        RECT 36.255 118.675 37.185 118.895 ;
        RECT 40.015 118.665 40.935 118.895 ;
        RECT 41.405 118.795 42.775 119.575 ;
        RECT 42.785 118.765 48.295 119.575 ;
        RECT 48.905 118.665 51.515 119.575 ;
        RECT 51.525 118.765 57.035 119.575 ;
        RECT 57.055 118.705 57.485 119.490 ;
        RECT 57.505 118.765 58.875 119.575 ;
        RECT 58.895 118.665 60.245 119.575 ;
        RECT 60.265 118.765 63.935 119.575 ;
        RECT 64.405 118.895 73.595 119.575 ;
        RECT 64.405 118.665 65.325 118.895 ;
        RECT 68.155 118.675 69.085 118.895 ;
        RECT 73.605 118.665 76.215 119.575 ;
        RECT 76.365 118.765 79.115 119.575 ;
        RECT 79.125 118.795 80.495 119.575 ;
        RECT 80.505 118.765 82.335 119.575 ;
        RECT 82.815 118.705 83.245 119.490 ;
        RECT 83.265 118.765 88.775 119.575 ;
        RECT 88.785 118.765 90.615 119.575 ;
        RECT 91.085 118.795 92.455 119.575 ;
        RECT 92.465 118.765 95.215 119.575 ;
        RECT 95.685 118.795 97.055 119.575 ;
        RECT 97.065 118.765 98.895 119.575 ;
        RECT 98.915 118.665 100.265 119.575 ;
        RECT 100.285 118.765 102.115 119.575 ;
        RECT 102.125 118.795 103.495 119.575 ;
        RECT 103.505 118.765 105.335 119.575 ;
        RECT 105.805 118.795 107.175 119.575 ;
        RECT 107.185 118.795 108.555 119.575 ;
        RECT 108.575 118.705 109.005 119.490 ;
        RECT 109.025 118.895 118.215 119.575 ;
        RECT 113.535 118.675 114.465 118.895 ;
        RECT 117.295 118.665 118.215 118.895 ;
        RECT 118.225 118.765 121.895 119.575 ;
        RECT 122.365 118.765 123.735 119.575 ;
      LAYER nwell ;
        RECT 5.330 115.545 123.930 118.375 ;
      LAYER pwell ;
        RECT 5.525 114.345 6.895 115.155 ;
        RECT 6.905 114.345 9.655 115.155 ;
        RECT 10.125 114.345 11.495 115.125 ;
        RECT 11.505 114.345 12.875 115.125 ;
        RECT 12.885 114.345 18.395 115.155 ;
        RECT 18.415 114.430 18.845 115.215 ;
        RECT 18.865 114.345 22.535 115.155 ;
        RECT 22.545 114.345 23.915 115.155 ;
        RECT 23.925 114.345 25.295 115.125 ;
        RECT 25.305 114.345 30.815 115.155 ;
        RECT 30.825 114.345 33.575 115.155 ;
        RECT 33.585 114.345 34.955 115.125 ;
        RECT 34.965 114.345 40.475 115.155 ;
        RECT 40.485 114.345 44.155 115.155 ;
        RECT 44.175 114.430 44.605 115.215 ;
        RECT 44.625 114.345 50.135 115.155 ;
        RECT 50.145 114.345 55.655 115.155 ;
        RECT 55.665 114.345 61.175 115.155 ;
        RECT 61.185 114.345 66.695 115.155 ;
        RECT 66.705 114.345 68.535 115.155 ;
        RECT 68.545 114.345 69.915 115.125 ;
        RECT 69.935 114.430 70.365 115.215 ;
        RECT 71.305 114.345 72.675 115.125 ;
        RECT 72.685 114.345 75.435 115.155 ;
        RECT 77.265 115.025 78.185 115.245 ;
        RECT 84.265 115.145 85.185 115.255 ;
        RECT 82.850 115.025 85.185 115.145 ;
        RECT 75.905 114.345 85.185 115.025 ;
        RECT 85.565 114.345 91.075 115.155 ;
        RECT 91.085 114.345 94.755 115.155 ;
        RECT 95.695 114.430 96.125 115.215 ;
        RECT 96.145 114.345 101.655 115.155 ;
        RECT 101.665 114.345 107.175 115.155 ;
        RECT 107.185 114.345 112.695 115.155 ;
        RECT 113.635 114.345 114.985 115.255 ;
        RECT 115.005 114.345 120.515 115.155 ;
        RECT 121.455 114.430 121.885 115.215 ;
        RECT 122.365 114.345 123.735 115.155 ;
        RECT 5.665 114.135 5.835 114.345 ;
        RECT 7.045 114.135 7.215 114.345 ;
        RECT 9.800 114.185 9.920 114.295 ;
        RECT 10.725 114.135 10.895 114.325 ;
        RECT 11.185 114.155 11.355 114.345 ;
        RECT 12.565 114.155 12.735 114.345 ;
        RECT 13.025 114.155 13.195 114.345 ;
        RECT 19.005 114.155 19.175 114.345 ;
        RECT 20.385 114.135 20.555 114.325 ;
        RECT 22.685 114.155 22.855 114.345 ;
        RECT 24.985 114.155 25.155 114.345 ;
        RECT 25.445 114.155 25.615 114.345 ;
        RECT 25.905 114.135 26.075 114.325 ;
        RECT 30.505 114.135 30.675 114.325 ;
        RECT 30.965 114.295 31.135 114.345 ;
        RECT 30.960 114.185 31.135 114.295 ;
        RECT 30.965 114.155 31.135 114.185 ;
        RECT 32.805 114.135 32.975 114.325 ;
        RECT 33.265 114.135 33.435 114.325 ;
        RECT 34.645 114.155 34.815 114.345 ;
        RECT 35.105 114.155 35.275 114.345 ;
        RECT 38.795 114.180 38.955 114.290 ;
        RECT 39.705 114.135 39.875 114.325 ;
        RECT 40.625 114.155 40.795 114.345 ;
        RECT 44.765 114.155 44.935 114.345 ;
        RECT 49.365 114.135 49.535 114.325 ;
        RECT 50.285 114.155 50.455 114.345 ;
        RECT 54.885 114.135 55.055 114.325 ;
        RECT 55.805 114.155 55.975 114.345 ;
        RECT 56.720 114.185 56.840 114.295 ;
        RECT 61.325 114.155 61.495 114.345 ;
        RECT 66.845 114.135 67.015 114.345 ;
        RECT 67.305 114.135 67.475 114.325 ;
        RECT 69.605 114.155 69.775 114.345 ;
        RECT 70.535 114.190 70.695 114.300 ;
        RECT 72.365 114.155 72.535 114.345 ;
        RECT 72.825 114.135 72.995 114.345 ;
        RECT 75.580 114.185 75.700 114.295 ;
        RECT 76.045 114.155 76.215 114.345 ;
        RECT 76.505 114.135 76.675 114.325 ;
        RECT 78.805 114.135 78.975 114.325 ;
        RECT 79.265 114.135 79.435 114.325 ;
        RECT 80.645 114.135 80.815 114.325 ;
        RECT 82.035 114.180 82.195 114.290 ;
        RECT 83.680 114.135 83.850 114.325 ;
        RECT 85.705 114.155 85.875 114.345 ;
        RECT 88.465 114.135 88.635 114.325 ;
        RECT 89.845 114.135 90.015 114.325 ;
        RECT 90.305 114.135 90.475 114.325 ;
        RECT 91.225 114.155 91.395 114.345 ;
        RECT 92.140 114.185 92.260 114.295 ;
        RECT 92.605 114.135 92.775 114.325 ;
        RECT 93.985 114.135 94.155 114.325 ;
        RECT 94.915 114.190 95.075 114.300 ;
        RECT 95.365 114.135 95.535 114.325 ;
        RECT 96.285 114.155 96.455 114.345 ;
        RECT 101.805 114.155 101.975 114.345 ;
        RECT 105.025 114.135 105.195 114.325 ;
        RECT 106.405 114.135 106.575 114.325 ;
        RECT 107.325 114.155 107.495 114.345 ;
        RECT 108.240 114.185 108.360 114.295 ;
        RECT 109.165 114.135 109.335 114.325 ;
        RECT 112.855 114.190 113.015 114.300 ;
        RECT 113.765 114.155 113.935 114.345 ;
        RECT 114.685 114.135 114.855 114.325 ;
        RECT 115.145 114.155 115.315 114.345 ;
        RECT 120.205 114.135 120.375 114.325 ;
        RECT 120.675 114.190 120.835 114.300 ;
        RECT 122.040 114.185 122.160 114.295 ;
        RECT 123.425 114.135 123.595 114.345 ;
        RECT 5.525 113.325 6.895 114.135 ;
        RECT 6.905 113.325 10.575 114.135 ;
        RECT 10.585 113.455 19.865 114.135 ;
        RECT 11.945 113.235 12.865 113.455 ;
        RECT 17.530 113.335 19.865 113.455 ;
        RECT 18.945 113.225 19.865 113.335 ;
        RECT 20.245 113.325 25.755 114.135 ;
        RECT 25.765 113.325 29.435 114.135 ;
        RECT 29.445 113.355 30.815 114.135 ;
        RECT 31.295 113.265 31.725 114.050 ;
        RECT 31.755 113.225 33.105 114.135 ;
        RECT 33.125 113.325 38.635 114.135 ;
        RECT 39.565 113.455 48.845 114.135 ;
        RECT 40.925 113.235 41.845 113.455 ;
        RECT 46.510 113.335 48.845 113.455 ;
        RECT 47.925 113.225 48.845 113.335 ;
        RECT 49.225 113.325 54.735 114.135 ;
        RECT 54.745 113.325 56.575 114.135 ;
        RECT 57.055 113.265 57.485 114.050 ;
        RECT 57.875 113.455 67.155 114.135 ;
        RECT 57.875 113.335 60.210 113.455 ;
        RECT 57.875 113.225 58.795 113.335 ;
        RECT 64.875 113.235 65.795 113.455 ;
        RECT 67.165 113.325 72.675 114.135 ;
        RECT 72.685 113.325 76.355 114.135 ;
        RECT 76.365 113.325 77.735 114.135 ;
        RECT 77.745 113.355 79.115 114.135 ;
        RECT 79.125 113.325 80.495 114.135 ;
        RECT 80.515 113.225 81.865 114.135 ;
        RECT 82.815 113.265 83.245 114.050 ;
        RECT 83.265 113.455 87.165 114.135 ;
        RECT 83.265 113.225 84.195 113.455 ;
        RECT 87.405 113.355 88.775 114.135 ;
        RECT 88.795 113.225 90.145 114.135 ;
        RECT 90.165 113.325 91.995 114.135 ;
        RECT 92.465 113.355 93.835 114.135 ;
        RECT 93.855 113.225 95.205 114.135 ;
        RECT 95.225 113.455 104.505 114.135 ;
        RECT 96.585 113.235 97.505 113.455 ;
        RECT 102.170 113.335 104.505 113.455 ;
        RECT 104.885 113.355 106.255 114.135 ;
        RECT 103.585 113.225 104.505 113.335 ;
        RECT 106.265 113.325 108.095 114.135 ;
        RECT 108.575 113.265 109.005 114.050 ;
        RECT 109.025 113.325 114.535 114.135 ;
        RECT 114.545 113.325 120.055 114.135 ;
        RECT 120.065 113.325 121.895 114.135 ;
        RECT 122.365 113.325 123.735 114.135 ;
      LAYER nwell ;
        RECT 5.330 110.105 123.930 112.935 ;
      LAYER pwell ;
        RECT 5.525 108.905 6.895 109.715 ;
        RECT 6.905 108.905 12.415 109.715 ;
        RECT 12.425 108.905 14.255 109.715 ;
        RECT 14.265 108.905 15.635 109.685 ;
        RECT 15.655 108.905 17.005 109.815 ;
        RECT 17.025 108.905 18.395 109.715 ;
        RECT 18.415 108.990 18.845 109.775 ;
        RECT 18.865 109.585 19.795 109.815 ;
        RECT 18.865 108.905 22.765 109.585 ;
        RECT 23.005 108.905 24.835 109.715 ;
        RECT 24.855 108.905 26.205 109.815 ;
        RECT 27.585 109.585 28.505 109.805 ;
        RECT 34.585 109.705 35.505 109.815 ;
        RECT 33.170 109.585 35.505 109.705 ;
        RECT 26.225 108.905 35.505 109.585 ;
        RECT 35.885 108.905 41.395 109.715 ;
        RECT 41.405 108.905 42.775 109.685 ;
        RECT 42.785 108.905 44.155 109.715 ;
        RECT 44.175 108.990 44.605 109.775 ;
        RECT 44.635 108.905 45.985 109.815 ;
        RECT 46.005 108.905 47.835 109.715 ;
        RECT 48.305 108.905 49.675 109.685 ;
        RECT 50.155 108.905 51.505 109.815 ;
        RECT 52.445 108.905 53.815 109.685 ;
        RECT 53.825 109.585 54.755 109.815 ;
        RECT 53.825 108.905 57.725 109.585 ;
        RECT 57.965 108.905 59.335 109.685 ;
        RECT 60.705 109.585 61.625 109.805 ;
        RECT 67.705 109.705 68.625 109.815 ;
        RECT 66.290 109.585 68.625 109.705 ;
        RECT 59.345 108.905 68.625 109.585 ;
        RECT 69.935 108.990 70.365 109.775 ;
        RECT 72.205 109.585 73.125 109.805 ;
        RECT 79.205 109.705 80.125 109.815 ;
        RECT 77.790 109.585 80.125 109.705 ;
        RECT 93.825 109.585 94.755 109.815 ;
        RECT 70.845 108.905 80.125 109.585 ;
        RECT 81.510 108.905 90.615 109.585 ;
        RECT 90.855 108.905 94.755 109.585 ;
        RECT 95.695 108.990 96.125 109.775 ;
        RECT 99.345 109.585 100.275 109.815 ;
        RECT 96.375 108.905 100.275 109.585 ;
        RECT 100.285 108.905 101.655 109.685 ;
        RECT 101.675 108.905 103.025 109.815 ;
        RECT 106.705 109.585 107.635 109.815 ;
        RECT 109.005 109.585 109.925 109.805 ;
        RECT 116.005 109.705 116.925 109.815 ;
        RECT 114.590 109.585 116.925 109.705 ;
        RECT 103.735 108.905 107.635 109.585 ;
        RECT 107.645 108.905 116.925 109.585 ;
        RECT 117.315 108.905 118.665 109.815 ;
        RECT 118.685 108.905 121.435 109.715 ;
        RECT 121.455 108.990 121.885 109.775 ;
        RECT 122.365 108.905 123.735 109.715 ;
        RECT 5.665 108.695 5.835 108.905 ;
        RECT 7.045 108.695 7.215 108.905 ;
        RECT 12.565 108.695 12.735 108.905 ;
        RECT 15.325 108.715 15.495 108.905 ;
        RECT 16.705 108.715 16.875 108.905 ;
        RECT 17.165 108.715 17.335 108.905 ;
        RECT 18.095 108.740 18.255 108.850 ;
        RECT 19.005 108.695 19.175 108.885 ;
        RECT 19.280 108.715 19.450 108.905 ;
        RECT 20.385 108.695 20.555 108.885 ;
        RECT 23.145 108.715 23.315 108.905 ;
        RECT 24.985 108.715 25.155 108.905 ;
        RECT 26.365 108.715 26.535 108.905 ;
        RECT 30.045 108.695 30.215 108.885 ;
        RECT 31.895 108.740 32.055 108.850 ;
        RECT 32.805 108.695 32.975 108.885 ;
        RECT 34.185 108.695 34.355 108.885 ;
        RECT 36.025 108.715 36.195 108.905 ;
        RECT 42.465 108.715 42.635 108.905 ;
        RECT 42.925 108.715 43.095 108.905 ;
        RECT 44.765 108.695 44.935 108.885 ;
        RECT 45.220 108.745 45.340 108.855 ;
        RECT 45.685 108.695 45.855 108.905 ;
        RECT 46.145 108.715 46.315 108.905 ;
        RECT 47.980 108.745 48.100 108.855 ;
        RECT 49.365 108.715 49.535 108.905 ;
        RECT 49.820 108.745 49.940 108.855 ;
        RECT 50.285 108.715 50.455 108.905 ;
        RECT 51.675 108.750 51.835 108.860 ;
        RECT 52.585 108.715 52.755 108.905 ;
        RECT 54.240 108.715 54.410 108.905 ;
        RECT 55.345 108.695 55.515 108.885 ;
        RECT 57.655 108.740 57.815 108.850 ;
        RECT 58.105 108.715 58.275 108.905 ;
        RECT 58.565 108.695 58.735 108.885 ;
        RECT 59.485 108.715 59.655 108.905 ;
        RECT 60.220 108.695 60.390 108.885 ;
        RECT 64.080 108.745 64.200 108.855 ;
        RECT 65.465 108.695 65.635 108.885 ;
        RECT 65.925 108.695 66.095 108.885 ;
        RECT 69.155 108.750 69.315 108.860 ;
        RECT 70.520 108.745 70.640 108.855 ;
        RECT 70.985 108.715 71.155 108.905 ;
        RECT 71.445 108.695 71.615 108.885 ;
        RECT 73.745 108.695 73.915 108.885 ;
        RECT 74.210 108.695 74.380 108.885 ;
        RECT 76.975 108.740 77.135 108.850 ;
        RECT 78.160 108.695 78.330 108.885 ;
        RECT 80.655 108.750 80.815 108.860 ;
        RECT 82.035 108.740 82.195 108.850 ;
        RECT 83.410 108.695 83.580 108.885 ;
        RECT 90.305 108.715 90.475 108.905 ;
        RECT 94.170 108.715 94.340 108.905 ;
        RECT 94.915 108.750 95.075 108.860 ;
        RECT 99.690 108.715 99.860 108.905 ;
        RECT 101.345 108.715 101.515 108.905 ;
        RECT 102.725 108.715 102.895 108.905 ;
        RECT 103.180 108.745 103.300 108.855 ;
        RECT 103.645 108.695 103.815 108.885 ;
        RECT 104.105 108.695 104.275 108.885 ;
        RECT 106.865 108.695 107.035 108.885 ;
        RECT 107.050 108.715 107.220 108.905 ;
        RECT 107.785 108.715 107.955 108.905 ;
        RECT 108.240 108.745 108.360 108.855 ;
        RECT 109.165 108.695 109.335 108.885 ;
        RECT 110.545 108.695 110.715 108.885 ;
        RECT 111.925 108.695 112.095 108.885 ;
        RECT 117.445 108.715 117.615 108.905 ;
        RECT 118.825 108.715 118.995 108.905 ;
        RECT 121.595 108.740 121.755 108.850 ;
        RECT 122.040 108.745 122.160 108.855 ;
        RECT 123.425 108.695 123.595 108.905 ;
        RECT 5.525 107.885 6.895 108.695 ;
        RECT 6.905 107.885 12.415 108.695 ;
        RECT 12.425 107.885 17.935 108.695 ;
        RECT 18.865 107.915 20.235 108.695 ;
        RECT 20.245 108.015 29.525 108.695 ;
        RECT 21.605 107.795 22.525 108.015 ;
        RECT 27.190 107.895 29.525 108.015 ;
        RECT 28.605 107.785 29.525 107.895 ;
        RECT 29.905 107.885 31.275 108.695 ;
        RECT 31.295 107.825 31.725 108.610 ;
        RECT 32.665 107.915 34.035 108.695 ;
        RECT 34.045 108.015 43.325 108.695 ;
        RECT 35.405 107.795 36.325 108.015 ;
        RECT 40.990 107.895 43.325 108.015 ;
        RECT 42.405 107.785 43.325 107.895 ;
        RECT 43.715 107.785 45.065 108.695 ;
        RECT 45.545 108.015 54.825 108.695 ;
        RECT 46.905 107.795 47.825 108.015 ;
        RECT 52.490 107.895 54.825 108.015 ;
        RECT 53.905 107.785 54.825 107.895 ;
        RECT 55.205 107.885 57.035 108.695 ;
        RECT 57.055 107.825 57.485 108.610 ;
        RECT 58.435 107.785 59.785 108.695 ;
        RECT 59.805 108.015 63.705 108.695 ;
        RECT 59.805 107.785 60.735 108.015 ;
        RECT 64.415 107.785 65.765 108.695 ;
        RECT 65.785 107.885 71.295 108.695 ;
        RECT 71.305 107.885 72.675 108.695 ;
        RECT 72.685 107.915 74.055 108.695 ;
        RECT 74.065 107.785 76.675 108.695 ;
        RECT 77.745 108.015 81.645 108.695 ;
        RECT 77.745 107.785 78.675 108.015 ;
        RECT 82.815 107.825 83.245 108.610 ;
        RECT 83.265 107.785 94.275 108.695 ;
        RECT 94.675 108.015 103.955 108.695 ;
        RECT 94.675 107.895 97.010 108.015 ;
        RECT 94.675 107.785 95.595 107.895 ;
        RECT 101.675 107.795 102.595 108.015 ;
        RECT 103.965 107.885 106.715 108.695 ;
        RECT 106.725 107.915 108.095 108.695 ;
        RECT 108.575 107.825 109.005 108.610 ;
        RECT 109.025 107.885 110.395 108.695 ;
        RECT 110.405 107.915 111.775 108.695 ;
        RECT 111.785 108.015 121.065 108.695 ;
        RECT 113.145 107.795 114.065 108.015 ;
        RECT 118.730 107.895 121.065 108.015 ;
        RECT 120.145 107.785 121.065 107.895 ;
        RECT 122.365 107.885 123.735 108.695 ;
      LAYER nwell ;
        RECT 5.330 104.665 123.930 107.495 ;
      LAYER pwell ;
        RECT 5.525 103.465 6.895 104.275 ;
        RECT 6.905 103.465 10.575 104.275 ;
        RECT 11.505 103.465 12.875 104.245 ;
        RECT 12.895 103.465 14.245 104.375 ;
        RECT 14.265 104.145 15.195 104.375 ;
        RECT 14.265 103.465 18.165 104.145 ;
        RECT 18.415 103.550 18.845 104.335 ;
        RECT 18.865 103.465 20.695 104.275 ;
        RECT 21.165 104.145 22.095 104.375 ;
        RECT 21.165 103.465 25.065 104.145 ;
        RECT 25.305 103.465 34.410 104.145 ;
        RECT 34.505 103.465 35.875 104.275 ;
        RECT 35.885 104.145 36.815 104.375 ;
        RECT 35.885 103.465 39.785 104.145 ;
        RECT 40.025 103.465 41.395 104.275 ;
        RECT 41.405 103.465 44.145 104.145 ;
        RECT 44.175 103.550 44.605 104.335 ;
        RECT 53.825 104.145 54.755 104.375 ;
        RECT 58.165 104.285 59.115 104.375 ;
        RECT 44.625 103.465 53.730 104.145 ;
        RECT 53.825 103.465 57.725 104.145 ;
        RECT 58.165 103.465 60.095 104.285 ;
        RECT 60.265 103.465 65.775 104.275 ;
        RECT 65.795 103.465 68.535 104.145 ;
        RECT 68.545 103.465 69.915 104.275 ;
        RECT 69.935 103.550 70.365 104.335 ;
        RECT 70.385 103.465 71.755 104.275 ;
        RECT 71.765 103.465 74.505 104.145 ;
        RECT 74.525 103.465 75.895 104.275 ;
        RECT 75.915 103.465 77.265 104.375 ;
        RECT 79.805 104.285 80.755 104.375 ;
        RECT 77.285 103.465 78.655 104.275 ;
        RECT 78.825 103.465 80.755 104.285 ;
        RECT 82.325 104.145 83.245 104.365 ;
        RECT 89.325 104.265 90.245 104.375 ;
        RECT 87.910 104.145 90.245 104.265 ;
        RECT 80.965 103.465 90.245 104.145 ;
        RECT 90.825 104.285 91.775 104.375 ;
        RECT 90.825 103.465 92.755 104.285 ;
        RECT 92.925 103.465 95.675 104.275 ;
        RECT 95.695 103.550 96.125 104.335 ;
        RECT 96.145 103.465 98.895 104.275 ;
        RECT 98.915 103.465 100.265 104.375 ;
        RECT 100.285 103.465 109.390 104.145 ;
        RECT 109.485 103.465 112.235 104.275 ;
        RECT 112.245 104.145 113.175 104.375 ;
        RECT 112.245 103.465 116.145 104.145 ;
        RECT 116.395 103.465 117.745 104.375 ;
        RECT 117.765 103.465 121.435 104.275 ;
        RECT 121.455 103.550 121.885 104.335 ;
        RECT 122.365 103.465 123.735 104.275 ;
        RECT 5.665 103.255 5.835 103.465 ;
        RECT 7.045 103.255 7.215 103.465 ;
        RECT 8.425 103.255 8.595 103.445 ;
        RECT 10.735 103.310 10.895 103.420 ;
        RECT 12.565 103.275 12.735 103.465 ;
        RECT 13.945 103.275 14.115 103.465 ;
        RECT 14.680 103.275 14.850 103.465 ;
        RECT 18.360 103.255 18.530 103.445 ;
        RECT 19.005 103.275 19.175 103.465 ;
        RECT 20.840 103.305 20.960 103.415 ;
        RECT 21.580 103.275 21.750 103.465 ;
        RECT 23.145 103.255 23.315 103.445 ;
        RECT 23.605 103.255 23.775 103.445 ;
        RECT 25.445 103.275 25.615 103.465 ;
        RECT 26.360 103.305 26.480 103.415 ;
        RECT 26.825 103.275 26.995 103.445 ;
        RECT 26.845 103.255 26.995 103.275 ;
        RECT 29.125 103.255 29.295 103.445 ;
        RECT 30.960 103.305 31.080 103.415 ;
        RECT 32.160 103.255 32.330 103.445 ;
        RECT 34.645 103.275 34.815 103.465 ;
        RECT 36.025 103.255 36.195 103.445 ;
        RECT 36.300 103.275 36.470 103.465 ;
        RECT 40.165 103.275 40.335 103.465 ;
        RECT 41.545 103.255 41.715 103.465 ;
        RECT 44.300 103.305 44.420 103.415 ;
        RECT 44.765 103.275 44.935 103.465 ;
        RECT 45.040 103.255 45.210 103.445 ;
        RECT 48.905 103.255 49.075 103.445 ;
        RECT 50.745 103.275 50.915 103.445 ;
        RECT 53.045 103.275 53.215 103.445 ;
        RECT 54.240 103.275 54.410 103.465 ;
        RECT 59.945 103.445 60.095 103.465 ;
        RECT 50.765 103.255 50.915 103.275 ;
        RECT 53.065 103.255 53.215 103.275 ;
        RECT 55.345 103.255 55.515 103.445 ;
        RECT 59.485 103.275 59.655 103.445 ;
        RECT 59.485 103.255 59.635 103.275 ;
        RECT 59.945 103.255 60.115 103.445 ;
        RECT 60.405 103.275 60.575 103.465 ;
        RECT 65.475 103.300 65.635 103.410 ;
        RECT 66.385 103.275 66.555 103.445 ;
        RECT 68.225 103.275 68.395 103.465 ;
        RECT 66.405 103.255 66.555 103.275 ;
        RECT 68.685 103.255 68.855 103.465 ;
        RECT 70.525 103.255 70.695 103.465 ;
        RECT 71.905 103.275 72.075 103.465 ;
        RECT 74.665 103.275 74.835 103.465 ;
        RECT 76.045 103.255 76.215 103.445 ;
        RECT 76.965 103.275 77.135 103.465 ;
        RECT 77.425 103.275 77.595 103.465 ;
        RECT 78.825 103.445 78.975 103.465 ;
        RECT 78.805 103.275 78.975 103.445 ;
        RECT 81.105 103.275 81.275 103.465 ;
        RECT 92.605 103.445 92.755 103.465 ;
        RECT 81.565 103.255 81.735 103.445 ;
        RECT 83.415 103.300 83.575 103.410 ;
        RECT 84.325 103.275 84.495 103.445 ;
        RECT 84.345 103.255 84.495 103.275 ;
        RECT 86.900 103.255 87.070 103.445 ;
        RECT 90.775 103.300 90.935 103.410 ;
        RECT 92.605 103.275 92.775 103.445 ;
        RECT 93.065 103.275 93.235 103.465 ;
        RECT 93.525 103.275 93.695 103.445 ;
        RECT 93.980 103.305 94.100 103.415 ;
        RECT 96.285 103.275 96.455 103.465 ;
        RECT 96.740 103.305 96.860 103.415 ;
        RECT 93.525 103.255 93.675 103.275 ;
        RECT 96.285 103.255 96.435 103.275 ;
        RECT 97.205 103.255 97.375 103.445 ;
        RECT 99.045 103.275 99.215 103.465 ;
        RECT 100.425 103.275 100.595 103.465 ;
        RECT 106.865 103.255 107.035 103.445 ;
        RECT 109.160 103.305 109.280 103.415 ;
        RECT 109.625 103.275 109.795 103.465 ;
        RECT 109.900 103.255 110.070 103.445 ;
        RECT 112.660 103.275 112.830 103.465 ;
        RECT 114.685 103.255 114.855 103.445 ;
        RECT 115.145 103.255 115.315 103.445 ;
        RECT 116.525 103.275 116.695 103.465 ;
        RECT 117.905 103.275 118.075 103.465 ;
        RECT 120.665 103.255 120.835 103.445 ;
        RECT 122.040 103.305 122.160 103.415 ;
        RECT 123.425 103.255 123.595 103.465 ;
        RECT 5.525 102.445 6.895 103.255 ;
        RECT 6.905 102.475 8.275 103.255 ;
        RECT 8.285 102.575 17.565 103.255 ;
        RECT 9.645 102.355 10.565 102.575 ;
        RECT 15.230 102.455 17.565 102.575 ;
        RECT 16.645 102.345 17.565 102.455 ;
        RECT 17.945 102.575 21.845 103.255 ;
        RECT 17.945 102.345 18.875 102.575 ;
        RECT 22.095 102.345 23.445 103.255 ;
        RECT 23.465 102.445 26.215 103.255 ;
        RECT 26.845 102.435 28.775 103.255 ;
        RECT 28.985 102.445 30.815 103.255 ;
        RECT 27.825 102.345 28.775 102.435 ;
        RECT 31.295 102.385 31.725 103.170 ;
        RECT 31.745 102.575 35.645 103.255 ;
        RECT 31.745 102.345 32.675 102.575 ;
        RECT 35.885 102.445 41.395 103.255 ;
        RECT 41.405 102.445 44.155 103.255 ;
        RECT 44.625 102.575 48.525 103.255 ;
        RECT 44.625 102.345 45.555 102.575 ;
        RECT 48.765 102.445 50.595 103.255 ;
        RECT 50.765 102.435 52.695 103.255 ;
        RECT 53.065 102.435 54.995 103.255 ;
        RECT 55.205 102.445 57.035 103.255 ;
        RECT 51.745 102.345 52.695 102.435 ;
        RECT 54.045 102.345 54.995 102.435 ;
        RECT 57.055 102.385 57.485 103.170 ;
        RECT 57.705 102.435 59.635 103.255 ;
        RECT 59.805 102.445 65.315 103.255 ;
        RECT 66.405 102.435 68.335 103.255 ;
        RECT 68.545 102.575 70.375 103.255 ;
        RECT 70.385 102.445 75.895 103.255 ;
        RECT 75.905 102.445 81.415 103.255 ;
        RECT 81.425 102.445 82.795 103.255 ;
        RECT 57.705 102.345 58.655 102.435 ;
        RECT 67.385 102.345 68.335 102.435 ;
        RECT 82.815 102.385 83.245 103.170 ;
        RECT 84.345 102.435 86.275 103.255 ;
        RECT 85.325 102.345 86.275 102.435 ;
        RECT 86.485 102.575 90.385 103.255 ;
        RECT 86.485 102.345 87.415 102.575 ;
        RECT 91.745 102.435 93.675 103.255 ;
        RECT 94.505 102.435 96.435 103.255 ;
        RECT 97.065 102.575 106.345 103.255 ;
        RECT 91.745 102.345 92.695 102.435 ;
        RECT 94.505 102.345 95.455 102.435 ;
        RECT 98.425 102.355 99.345 102.575 ;
        RECT 104.010 102.455 106.345 102.575 ;
        RECT 105.425 102.345 106.345 102.455 ;
        RECT 106.725 102.445 108.555 103.255 ;
        RECT 108.575 102.385 109.005 103.170 ;
        RECT 109.485 102.575 113.385 103.255 ;
        RECT 109.485 102.345 110.415 102.575 ;
        RECT 113.635 102.345 114.985 103.255 ;
        RECT 115.005 102.445 120.515 103.255 ;
        RECT 120.525 102.445 122.355 103.255 ;
        RECT 122.365 102.445 123.735 103.255 ;
      LAYER nwell ;
        RECT 5.330 99.225 123.930 102.055 ;
      LAYER pwell ;
        RECT 5.525 98.025 6.895 98.835 ;
        RECT 9.185 98.705 10.105 98.925 ;
        RECT 16.185 98.825 17.105 98.935 ;
        RECT 14.770 98.705 17.105 98.825 ;
        RECT 7.825 98.025 17.105 98.705 ;
        RECT 18.415 98.110 18.845 98.895 ;
        RECT 23.685 98.845 24.635 98.935 ;
        RECT 18.865 98.025 22.535 98.835 ;
        RECT 22.705 98.025 24.635 98.845 ;
        RECT 25.045 98.845 25.995 98.935 ;
        RECT 28.285 98.845 29.235 98.935 ;
        RECT 25.045 98.025 26.975 98.845 ;
        RECT 5.665 97.815 5.835 98.025 ;
        RECT 7.045 97.815 7.215 98.005 ;
        RECT 7.965 97.835 8.135 98.025 ;
        RECT 12.565 97.815 12.735 98.005 ;
        RECT 17.635 97.870 17.795 97.980 ;
        RECT 18.085 97.815 18.255 98.005 ;
        RECT 19.005 97.835 19.175 98.025 ;
        RECT 22.705 98.005 22.855 98.025 ;
        RECT 26.825 98.005 26.975 98.025 ;
        RECT 27.305 98.025 29.235 98.845 ;
        RECT 34.705 98.845 35.655 98.935 ;
        RECT 29.445 98.025 33.115 98.835 ;
        RECT 33.125 98.025 34.495 98.835 ;
        RECT 34.705 98.025 36.635 98.845 ;
        RECT 36.805 98.025 42.315 98.835 ;
        RECT 42.325 98.025 44.155 98.835 ;
        RECT 44.175 98.110 44.605 98.895 ;
        RECT 44.635 98.025 45.985 98.935 ;
        RECT 46.005 98.025 51.515 98.835 ;
        RECT 51.525 98.025 57.035 98.835 ;
        RECT 57.045 98.025 62.555 98.835 ;
        RECT 62.565 98.025 66.235 98.835 ;
        RECT 66.705 98.025 68.535 98.705 ;
        RECT 68.545 98.025 69.915 98.835 ;
        RECT 69.935 98.110 70.365 98.895 ;
        RECT 70.395 98.025 71.745 98.935 ;
        RECT 71.765 98.025 73.595 98.835 ;
        RECT 73.605 98.025 74.975 98.805 ;
        RECT 74.985 98.025 80.495 98.835 ;
        RECT 80.505 98.025 86.015 98.835 ;
        RECT 86.025 98.025 91.535 98.835 ;
        RECT 91.545 98.025 95.215 98.835 ;
        RECT 95.695 98.110 96.125 98.895 ;
        RECT 96.345 98.845 97.295 98.935 ;
        RECT 96.345 98.025 98.275 98.845 ;
        RECT 98.905 98.025 100.275 98.805 ;
        RECT 100.285 98.705 101.215 98.935 ;
        RECT 100.285 98.025 104.185 98.705 ;
        RECT 104.425 98.025 107.175 98.835 ;
        RECT 109.005 98.705 109.925 98.925 ;
        RECT 116.005 98.825 116.925 98.935 ;
        RECT 114.590 98.705 116.925 98.825 ;
        RECT 107.645 98.025 116.925 98.705 ;
        RECT 117.315 98.025 118.665 98.935 ;
        RECT 118.685 98.025 121.435 98.835 ;
        RECT 121.455 98.110 121.885 98.895 ;
        RECT 122.365 98.025 123.735 98.835 ;
        RECT 27.305 98.005 27.455 98.025 ;
        RECT 22.685 97.835 22.855 98.005 ;
        RECT 22.685 97.815 22.835 97.835 ;
        RECT 24.065 97.815 24.235 98.005 ;
        RECT 24.525 97.815 24.695 98.005 ;
        RECT 26.365 97.815 26.535 98.005 ;
        RECT 26.825 97.835 26.995 98.005 ;
        RECT 27.285 97.835 27.455 98.005 ;
        RECT 27.745 97.815 27.915 98.005 ;
        RECT 29.585 97.835 29.755 98.025 ;
        RECT 31.895 97.860 32.055 97.970 ;
        RECT 32.805 97.815 32.975 98.005 ;
        RECT 33.265 97.835 33.435 98.025 ;
        RECT 36.485 98.005 36.635 98.025 ;
        RECT 34.185 97.815 34.355 98.005 ;
        RECT 36.020 97.865 36.140 97.975 ;
        RECT 36.485 97.835 36.655 98.005 ;
        RECT 36.945 97.835 37.115 98.025 ;
        RECT 37.405 97.815 37.575 98.005 ;
        RECT 37.865 97.815 38.035 98.005 ;
        RECT 39.245 97.815 39.415 98.005 ;
        RECT 40.625 97.815 40.795 98.005 ;
        RECT 42.465 97.835 42.635 98.025 ;
        RECT 44.765 97.835 44.935 98.025 ;
        RECT 46.145 97.835 46.315 98.025 ;
        RECT 50.285 97.815 50.455 98.005 ;
        RECT 51.665 97.835 51.835 98.025 ;
        RECT 53.040 97.865 53.160 97.975 ;
        RECT 5.525 97.005 6.895 97.815 ;
        RECT 6.905 97.005 12.415 97.815 ;
        RECT 12.425 97.005 17.935 97.815 ;
        RECT 17.945 97.005 20.695 97.815 ;
        RECT 20.905 96.995 22.835 97.815 ;
        RECT 23.005 97.035 24.375 97.815 ;
        RECT 24.385 97.005 26.215 97.815 ;
        RECT 20.905 96.905 21.855 96.995 ;
        RECT 26.235 96.905 27.585 97.815 ;
        RECT 27.605 97.005 31.275 97.815 ;
        RECT 31.295 96.945 31.725 97.730 ;
        RECT 32.665 97.035 34.035 97.815 ;
        RECT 34.045 97.005 35.875 97.815 ;
        RECT 36.355 96.905 37.705 97.815 ;
        RECT 37.725 97.005 39.095 97.815 ;
        RECT 39.105 97.035 40.475 97.815 ;
        RECT 40.485 97.135 49.765 97.815 ;
        RECT 41.845 96.915 42.765 97.135 ;
        RECT 47.430 97.015 49.765 97.135 ;
        RECT 48.845 96.905 49.765 97.015 ;
        RECT 50.145 97.005 52.895 97.815 ;
        RECT 53.365 97.785 54.310 97.815 ;
        RECT 55.800 97.785 55.970 98.005 ;
        RECT 56.275 97.860 56.435 97.970 ;
        RECT 57.185 97.835 57.355 98.025 ;
        RECT 57.645 97.815 57.815 98.005 ;
        RECT 60.405 97.815 60.575 98.005 ;
        RECT 62.705 97.835 62.875 98.025 ;
        RECT 66.380 97.865 66.500 97.975 ;
        RECT 66.845 97.835 67.015 98.025 ;
        RECT 68.685 97.835 68.855 98.025 ;
        RECT 70.065 97.815 70.235 98.005 ;
        RECT 71.445 97.835 71.615 98.025 ;
        RECT 71.905 97.835 72.075 98.025 ;
        RECT 74.665 97.835 74.835 98.025 ;
        RECT 75.125 97.835 75.295 98.025 ;
        RECT 79.725 97.815 79.895 98.005 ;
        RECT 80.645 97.835 80.815 98.025 ;
        RECT 82.480 97.865 82.600 97.975 ;
        RECT 83.405 97.815 83.575 98.005 ;
        RECT 86.165 97.835 86.335 98.025 ;
        RECT 88.925 97.815 89.095 98.005 ;
        RECT 91.685 97.835 91.855 98.025 ;
        RECT 98.125 98.005 98.275 98.025 ;
        RECT 94.445 97.815 94.615 98.005 ;
        RECT 95.360 97.865 95.480 97.975 ;
        RECT 98.125 97.815 98.295 98.005 ;
        RECT 98.580 97.865 98.700 97.975 ;
        RECT 99.505 97.835 99.675 98.005 ;
        RECT 99.965 97.835 100.135 98.025 ;
        RECT 100.700 97.835 100.870 98.025 ;
        RECT 99.525 97.815 99.675 97.835 ;
        RECT 101.805 97.815 101.975 98.005 ;
        RECT 104.565 97.835 104.735 98.025 ;
        RECT 107.325 97.975 107.495 98.005 ;
        RECT 107.320 97.865 107.495 97.975 ;
        RECT 107.325 97.815 107.495 97.865 ;
        RECT 107.785 97.835 107.955 98.025 ;
        RECT 110.085 97.815 110.255 98.005 ;
        RECT 110.545 97.815 110.715 98.005 ;
        RECT 111.925 97.815 112.095 98.005 ;
        RECT 117.445 97.835 117.615 98.025 ;
        RECT 118.825 97.835 118.995 98.025 ;
        RECT 121.595 97.860 121.755 97.970 ;
        RECT 122.040 97.865 122.160 97.975 ;
        RECT 123.425 97.815 123.595 98.025 ;
        RECT 53.365 97.105 56.115 97.785 ;
        RECT 53.365 96.905 54.310 97.105 ;
        RECT 57.055 96.945 57.485 97.730 ;
        RECT 57.505 97.005 60.255 97.815 ;
        RECT 60.265 97.135 69.545 97.815 ;
        RECT 69.925 97.135 79.205 97.815 ;
        RECT 61.625 96.915 62.545 97.135 ;
        RECT 67.210 97.015 69.545 97.135 ;
        RECT 68.625 96.905 69.545 97.015 ;
        RECT 71.285 96.915 72.205 97.135 ;
        RECT 76.870 97.015 79.205 97.135 ;
        RECT 78.285 96.905 79.205 97.015 ;
        RECT 79.585 97.005 82.335 97.815 ;
        RECT 82.815 96.945 83.245 97.730 ;
        RECT 83.265 97.005 88.775 97.815 ;
        RECT 88.785 97.005 94.295 97.815 ;
        RECT 94.305 97.005 97.975 97.815 ;
        RECT 97.985 97.005 99.355 97.815 ;
        RECT 99.525 96.995 101.455 97.815 ;
        RECT 101.665 97.005 107.175 97.815 ;
        RECT 107.185 97.005 108.555 97.815 ;
        RECT 100.505 96.905 101.455 96.995 ;
        RECT 108.575 96.945 109.005 97.730 ;
        RECT 109.025 97.035 110.395 97.815 ;
        RECT 110.405 97.035 111.775 97.815 ;
        RECT 111.785 97.135 121.065 97.815 ;
        RECT 113.145 96.915 114.065 97.135 ;
        RECT 118.730 97.015 121.065 97.135 ;
        RECT 120.145 96.905 121.065 97.015 ;
        RECT 122.365 97.005 123.735 97.815 ;
      LAYER nwell ;
        RECT 5.330 93.785 123.930 96.615 ;
      LAYER pwell ;
        RECT 5.525 92.585 6.895 93.395 ;
        RECT 6.905 92.585 12.415 93.395 ;
        RECT 12.425 92.585 17.935 93.395 ;
        RECT 18.415 92.670 18.845 93.455 ;
        RECT 18.865 92.585 21.615 93.395 ;
        RECT 22.985 93.265 23.905 93.485 ;
        RECT 29.985 93.385 30.905 93.495 ;
        RECT 28.570 93.265 30.905 93.385 ;
        RECT 32.645 93.265 33.565 93.485 ;
        RECT 39.645 93.385 40.565 93.495 ;
        RECT 38.230 93.265 40.565 93.385 ;
        RECT 21.625 92.585 30.905 93.265 ;
        RECT 31.285 92.585 40.565 93.265 ;
        RECT 40.945 92.585 43.695 93.395 ;
        RECT 44.175 92.670 44.605 93.455 ;
        RECT 44.625 93.265 45.555 93.495 ;
        RECT 44.625 92.585 48.525 93.265 ;
        RECT 48.765 92.585 50.595 93.395 ;
        RECT 51.260 92.585 54.735 93.495 ;
        RECT 54.745 92.585 56.575 93.395 ;
        RECT 57.945 93.265 58.865 93.485 ;
        RECT 64.945 93.385 65.865 93.495 ;
        RECT 63.530 93.265 65.865 93.385 ;
        RECT 56.585 92.585 65.865 93.265 ;
        RECT 66.245 92.585 67.615 93.365 ;
        RECT 67.625 92.585 68.995 93.365 ;
        RECT 69.935 92.670 70.365 93.455 ;
        RECT 70.385 93.265 71.315 93.495 ;
        RECT 70.385 92.585 74.285 93.265 ;
        RECT 74.535 92.585 75.885 93.495 ;
        RECT 76.825 93.265 77.755 93.495 ;
        RECT 76.825 92.585 80.725 93.265 ;
        RECT 80.965 92.585 82.795 93.395 ;
        RECT 83.000 92.585 86.475 93.495 ;
        RECT 86.680 92.585 90.155 93.495 ;
        RECT 90.165 92.585 91.995 93.395 ;
        RECT 92.465 93.295 93.410 93.495 ;
        RECT 92.465 92.615 95.215 93.295 ;
        RECT 95.695 92.670 96.125 93.455 ;
        RECT 97.950 93.295 98.895 93.495 ;
        RECT 101.885 93.405 102.835 93.495 ;
        RECT 96.145 92.615 98.895 93.295 ;
        RECT 92.465 92.585 93.410 92.615 ;
        RECT 5.665 92.375 5.835 92.585 ;
        RECT 7.045 92.375 7.215 92.585 ;
        RECT 10.735 92.420 10.895 92.530 ;
        RECT 12.565 92.375 12.735 92.585 ;
        RECT 13.025 92.375 13.195 92.565 ;
        RECT 14.680 92.375 14.850 92.565 ;
        RECT 18.080 92.425 18.200 92.535 ;
        RECT 18.545 92.375 18.715 92.565 ;
        RECT 19.005 92.395 19.175 92.585 ;
        RECT 21.765 92.395 21.935 92.585 ;
        RECT 22.225 92.375 22.395 92.565 ;
        RECT 23.880 92.375 24.050 92.565 ;
        RECT 27.745 92.375 27.915 92.565 ;
        RECT 31.425 92.395 31.595 92.585 ;
        RECT 31.895 92.420 32.055 92.530 ;
        RECT 33.080 92.375 33.250 92.565 ;
        RECT 36.945 92.375 37.115 92.565 ;
        RECT 38.780 92.425 38.900 92.535 ;
        RECT 39.245 92.375 39.415 92.565 ;
        RECT 40.625 92.375 40.795 92.565 ;
        RECT 41.085 92.395 41.255 92.585 ;
        RECT 43.840 92.425 43.960 92.535 ;
        RECT 45.040 92.395 45.210 92.585 ;
        RECT 48.905 92.395 49.075 92.585 ;
        RECT 50.740 92.425 50.860 92.535 ;
        RECT 53.500 92.375 53.670 92.565 ;
        RECT 5.525 91.565 6.895 92.375 ;
        RECT 6.905 91.565 10.575 92.375 ;
        RECT 11.505 91.595 12.875 92.375 ;
        RECT 12.885 91.565 14.255 92.375 ;
        RECT 14.265 91.695 18.165 92.375 ;
        RECT 14.265 91.465 15.195 91.695 ;
        RECT 18.405 91.565 22.075 92.375 ;
        RECT 22.085 91.565 23.455 92.375 ;
        RECT 23.465 91.695 27.365 92.375 ;
        RECT 23.465 91.465 24.395 91.695 ;
        RECT 27.605 91.565 31.275 92.375 ;
        RECT 31.295 91.505 31.725 92.290 ;
        RECT 32.665 91.695 36.565 92.375 ;
        RECT 32.665 91.465 33.595 91.695 ;
        RECT 36.805 91.565 38.635 92.375 ;
        RECT 39.105 91.595 40.475 92.375 ;
        RECT 40.485 91.695 49.765 92.375 ;
        RECT 41.845 91.475 42.765 91.695 ;
        RECT 47.430 91.575 49.765 91.695 ;
        RECT 48.845 91.465 49.765 91.575 ;
        RECT 50.340 91.465 53.815 92.375 ;
        RECT 53.970 92.345 54.140 92.565 ;
        RECT 54.420 92.395 54.590 92.585 ;
        RECT 54.885 92.395 55.055 92.585 ;
        RECT 56.725 92.535 56.895 92.585 ;
        RECT 56.720 92.425 56.895 92.535 ;
        RECT 56.725 92.395 56.895 92.425 ;
        RECT 57.645 92.375 57.815 92.565 ;
        RECT 61.325 92.375 61.495 92.565 ;
        RECT 62.700 92.425 62.820 92.535 ;
        RECT 66.570 92.375 66.740 92.565 ;
        RECT 67.305 92.375 67.475 92.585 ;
        RECT 68.685 92.395 68.855 92.585 ;
        RECT 69.155 92.430 69.315 92.540 ;
        RECT 70.800 92.395 70.970 92.585 ;
        RECT 72.825 92.375 72.995 92.565 ;
        RECT 74.665 92.395 74.835 92.585 ;
        RECT 76.055 92.430 76.215 92.540 ;
        RECT 77.240 92.395 77.410 92.585 ;
        RECT 78.345 92.375 78.515 92.565 ;
        RECT 80.180 92.425 80.300 92.535 ;
        RECT 81.105 92.395 81.275 92.585 ;
        RECT 81.565 92.375 81.735 92.565 ;
        RECT 82.035 92.420 82.195 92.530 ;
        RECT 83.680 92.375 83.850 92.565 ;
        RECT 86.160 92.395 86.330 92.585 ;
        RECT 89.840 92.395 90.010 92.585 ;
        RECT 90.305 92.395 90.475 92.585 ;
        RECT 90.760 92.375 90.930 92.565 ;
        RECT 55.630 92.345 56.575 92.375 ;
        RECT 53.825 91.665 56.575 92.345 ;
        RECT 55.630 91.465 56.575 91.665 ;
        RECT 57.055 91.505 57.485 92.290 ;
        RECT 57.505 91.565 61.175 92.375 ;
        RECT 61.195 91.465 62.545 92.375 ;
        RECT 63.255 91.695 67.155 92.375 ;
        RECT 66.225 91.465 67.155 91.695 ;
        RECT 67.165 91.565 72.675 92.375 ;
        RECT 72.685 91.565 78.195 92.375 ;
        RECT 78.205 91.565 80.035 92.375 ;
        RECT 80.505 91.595 81.875 92.375 ;
        RECT 82.815 91.505 83.245 92.290 ;
        RECT 83.265 91.695 87.165 92.375 ;
        RECT 83.265 91.465 84.195 91.695 ;
        RECT 87.600 91.465 91.075 92.375 ;
        RECT 91.230 92.345 91.400 92.565 ;
        RECT 92.140 92.425 92.260 92.535 ;
        RECT 93.985 92.375 94.155 92.565 ;
        RECT 94.900 92.395 95.070 92.615 ;
        RECT 95.360 92.425 95.480 92.535 ;
        RECT 96.290 92.395 96.460 92.615 ;
        RECT 97.950 92.585 98.895 92.615 ;
        RECT 98.905 92.585 100.735 93.395 ;
        RECT 100.905 92.585 102.835 93.405 ;
        RECT 103.245 93.405 104.195 93.495 ;
        RECT 105.545 93.405 106.495 93.495 ;
        RECT 103.245 92.585 105.175 93.405 ;
        RECT 105.545 92.585 107.475 93.405 ;
        RECT 107.645 92.585 111.315 93.395 ;
        RECT 111.325 92.585 112.695 93.395 ;
        RECT 112.705 93.265 113.635 93.495 ;
        RECT 112.705 92.585 116.605 93.265 ;
        RECT 116.845 92.585 120.515 93.395 ;
        RECT 121.455 92.670 121.885 93.455 ;
        RECT 122.365 92.585 123.735 93.395 ;
        RECT 99.045 92.395 99.215 92.585 ;
        RECT 100.905 92.565 101.055 92.585 ;
        RECT 99.505 92.375 99.675 92.565 ;
        RECT 100.885 92.395 101.055 92.565 ;
        RECT 105.025 92.565 105.175 92.585 ;
        RECT 107.325 92.565 107.475 92.585 ;
        RECT 105.025 92.375 105.195 92.565 ;
        RECT 107.325 92.395 107.495 92.565 ;
        RECT 107.785 92.395 107.955 92.585 ;
        RECT 109.165 92.375 109.335 92.565 ;
        RECT 111.465 92.395 111.635 92.585 ;
        RECT 113.120 92.395 113.290 92.585 ;
        RECT 114.685 92.375 114.855 92.565 ;
        RECT 116.985 92.395 117.155 92.585 ;
        RECT 120.205 92.375 120.375 92.565 ;
        RECT 120.675 92.430 120.835 92.540 ;
        RECT 122.040 92.425 122.160 92.535 ;
        RECT 123.425 92.375 123.595 92.585 ;
        RECT 92.890 92.345 93.835 92.375 ;
        RECT 91.085 91.665 93.835 92.345 ;
        RECT 92.890 91.465 93.835 91.665 ;
        RECT 93.845 91.565 99.355 92.375 ;
        RECT 99.365 91.565 104.875 92.375 ;
        RECT 104.885 91.565 108.555 92.375 ;
        RECT 108.575 91.505 109.005 92.290 ;
        RECT 109.025 91.565 114.535 92.375 ;
        RECT 114.545 91.565 120.055 92.375 ;
        RECT 120.065 91.565 121.895 92.375 ;
        RECT 122.365 91.565 123.735 92.375 ;
      LAYER nwell ;
        RECT 5.330 88.345 123.930 91.175 ;
      LAYER pwell ;
        RECT 5.525 87.145 6.895 87.955 ;
        RECT 6.905 87.145 8.735 87.955 ;
        RECT 10.105 87.825 11.025 88.045 ;
        RECT 17.105 87.945 18.025 88.055 ;
        RECT 15.690 87.825 18.025 87.945 ;
        RECT 8.745 87.145 18.025 87.825 ;
        RECT 18.415 87.230 18.845 88.015 ;
        RECT 18.865 87.145 24.375 87.955 ;
        RECT 26.190 87.855 27.135 88.055 ;
        RECT 24.385 87.175 27.135 87.855 ;
        RECT 5.665 86.935 5.835 87.145 ;
        RECT 7.045 86.955 7.215 87.145 ;
        RECT 7.965 86.935 8.135 87.125 ;
        RECT 8.885 86.955 9.055 87.145 ;
        RECT 17.900 86.935 18.070 87.125 ;
        RECT 19.005 86.955 19.175 87.145 ;
        RECT 21.765 86.935 21.935 87.125 ;
        RECT 24.530 86.955 24.700 87.175 ;
        RECT 26.190 87.145 27.135 87.175 ;
        RECT 27.145 87.145 32.655 87.955 ;
        RECT 32.665 87.145 34.035 87.955 ;
        RECT 35.850 87.855 36.795 88.055 ;
        RECT 34.045 87.175 36.795 87.855 ;
        RECT 27.285 86.955 27.455 87.145 ;
        RECT 27.740 86.935 27.910 87.125 ;
        RECT 5.525 86.125 6.895 86.935 ;
        RECT 7.825 86.255 17.105 86.935 ;
        RECT 9.185 86.035 10.105 86.255 ;
        RECT 14.770 86.135 17.105 86.255 ;
        RECT 16.185 86.025 17.105 86.135 ;
        RECT 17.485 86.255 21.385 86.935 ;
        RECT 17.485 86.025 18.415 86.255 ;
        RECT 21.625 86.125 24.375 86.935 ;
        RECT 24.580 86.025 28.055 86.935 ;
        RECT 28.210 86.905 28.380 87.125 ;
        RECT 30.960 86.985 31.080 87.095 ;
        RECT 32.805 86.955 32.975 87.145 ;
        RECT 34.190 86.955 34.360 87.175 ;
        RECT 35.850 87.145 36.795 87.175 ;
        RECT 36.805 87.145 42.315 87.955 ;
        RECT 42.795 87.145 44.145 88.055 ;
        RECT 44.175 87.230 44.605 88.015 ;
        RECT 45.545 87.825 46.475 88.055 ;
        RECT 45.545 87.145 49.445 87.825 ;
        RECT 49.685 87.145 55.195 87.955 ;
        RECT 55.205 87.145 58.875 87.955 ;
        RECT 59.345 87.145 60.715 87.925 ;
        RECT 60.725 87.145 66.235 87.955 ;
        RECT 66.440 87.145 69.915 88.055 ;
        RECT 69.935 87.230 70.365 88.015 ;
        RECT 70.385 87.145 75.895 87.955 ;
        RECT 75.905 87.145 77.735 87.955 ;
        RECT 79.565 87.825 80.485 88.045 ;
        RECT 86.565 87.945 87.485 88.055 ;
        RECT 85.150 87.825 87.485 87.945 ;
        RECT 78.205 87.145 87.485 87.825 ;
        RECT 87.875 87.145 89.225 88.055 ;
        RECT 89.245 87.145 94.755 87.955 ;
        RECT 95.695 87.230 96.125 88.015 ;
        RECT 96.145 87.145 99.815 87.955 ;
        RECT 102.090 87.855 103.035 88.055 ;
        RECT 104.850 87.855 105.795 88.055 ;
        RECT 100.285 87.175 103.035 87.855 ;
        RECT 103.045 87.175 105.795 87.855 ;
        RECT 35.100 86.935 35.270 87.125 ;
        RECT 35.565 86.935 35.735 87.125 ;
        RECT 36.945 86.955 37.115 87.145 ;
        RECT 41.085 86.935 41.255 87.125 ;
        RECT 42.460 86.985 42.580 87.095 ;
        RECT 42.925 86.955 43.095 87.145 ;
        RECT 44.775 86.990 44.935 87.100 ;
        RECT 45.960 86.955 46.130 87.145 ;
        RECT 46.605 86.935 46.775 87.125 ;
        RECT 49.825 86.955 49.995 87.145 ;
        RECT 52.125 86.935 52.295 87.125 ;
        RECT 55.345 86.955 55.515 87.145 ;
        RECT 55.805 86.935 55.975 87.125 ;
        RECT 57.645 86.935 57.815 87.125 ;
        RECT 59.020 86.985 59.140 87.095 ;
        RECT 60.405 86.955 60.575 87.145 ;
        RECT 60.865 86.955 61.035 87.145 ;
        RECT 67.300 86.985 67.420 87.095 ;
        RECT 69.600 86.955 69.770 87.145 ;
        RECT 70.525 86.955 70.695 87.145 ;
        RECT 70.980 86.935 71.150 87.125 ;
        RECT 71.445 86.935 71.615 87.125 ;
        RECT 76.045 86.955 76.215 87.145 ;
        RECT 76.965 86.935 77.135 87.125 ;
        RECT 77.880 86.985 78.000 87.095 ;
        RECT 78.345 86.955 78.515 87.145 ;
        RECT 82.480 86.985 82.600 87.095 ;
        RECT 83.405 86.935 83.575 87.125 ;
        RECT 84.785 86.935 84.955 87.125 ;
        RECT 88.925 86.955 89.095 87.145 ;
        RECT 89.385 86.955 89.555 87.145 ;
        RECT 94.915 86.990 95.075 87.100 ;
        RECT 95.365 86.935 95.535 87.125 ;
        RECT 95.825 86.935 95.995 87.125 ;
        RECT 96.285 86.955 96.455 87.145 ;
        RECT 99.970 87.095 100.140 87.125 ;
        RECT 99.500 86.985 99.620 87.095 ;
        RECT 99.960 86.985 100.140 87.095 ;
        RECT 29.870 86.905 30.815 86.935 ;
        RECT 28.065 86.225 30.815 86.905 ;
        RECT 29.870 86.025 30.815 86.225 ;
        RECT 31.295 86.065 31.725 86.850 ;
        RECT 31.940 86.025 35.415 86.935 ;
        RECT 35.425 86.125 40.935 86.935 ;
        RECT 40.945 86.125 46.455 86.935 ;
        RECT 46.465 86.125 51.975 86.935 ;
        RECT 51.985 86.125 55.655 86.935 ;
        RECT 55.665 86.125 57.035 86.935 ;
        RECT 57.055 86.065 57.485 86.850 ;
        RECT 57.505 86.255 66.785 86.935 ;
        RECT 58.865 86.035 59.785 86.255 ;
        RECT 64.450 86.135 66.785 86.255 ;
        RECT 65.865 86.025 66.785 86.135 ;
        RECT 67.820 86.025 71.295 86.935 ;
        RECT 71.305 86.125 76.815 86.935 ;
        RECT 76.825 86.125 82.335 86.935 ;
        RECT 82.815 86.065 83.245 86.850 ;
        RECT 83.265 86.155 84.635 86.935 ;
        RECT 84.645 86.255 93.925 86.935 ;
        RECT 86.005 86.035 86.925 86.255 ;
        RECT 91.590 86.135 93.925 86.255 ;
        RECT 93.005 86.025 93.925 86.135 ;
        RECT 94.315 86.025 95.665 86.935 ;
        RECT 95.685 86.125 99.355 86.935 ;
        RECT 99.970 86.905 100.140 86.985 ;
        RECT 100.430 86.955 100.600 87.175 ;
        RECT 102.090 87.145 103.035 87.175 ;
        RECT 101.630 86.905 102.575 86.935 ;
        RECT 102.730 86.905 102.900 87.125 ;
        RECT 103.190 86.955 103.360 87.175 ;
        RECT 104.850 87.145 105.795 87.175 ;
        RECT 105.805 87.145 111.315 87.955 ;
        RECT 111.325 87.145 112.695 87.955 ;
        RECT 112.705 87.145 114.075 87.925 ;
        RECT 114.095 87.145 115.445 88.055 ;
        RECT 115.465 87.145 120.975 87.955 ;
        RECT 121.455 87.230 121.885 88.015 ;
        RECT 122.365 87.145 123.735 87.955 ;
        RECT 105.485 86.935 105.655 87.125 ;
        RECT 105.945 86.955 106.115 87.145 ;
        RECT 108.240 86.985 108.360 87.095 ;
        RECT 109.165 86.935 109.335 87.125 ;
        RECT 111.465 86.955 111.635 87.145 ;
        RECT 112.845 86.955 113.015 87.145 ;
        RECT 115.145 86.955 115.315 87.145 ;
        RECT 115.605 86.955 115.775 87.145 ;
        RECT 118.825 86.935 118.995 87.125 ;
        RECT 120.205 86.935 120.375 87.125 ;
        RECT 121.120 86.985 121.240 87.095 ;
        RECT 122.040 86.985 122.160 87.095 ;
        RECT 123.425 86.935 123.595 87.145 ;
        RECT 104.390 86.905 105.335 86.935 ;
        RECT 99.825 86.225 102.575 86.905 ;
        RECT 102.585 86.225 105.335 86.905 ;
        RECT 101.630 86.025 102.575 86.225 ;
        RECT 104.390 86.025 105.335 86.225 ;
        RECT 105.345 86.125 108.095 86.935 ;
        RECT 108.575 86.065 109.005 86.850 ;
        RECT 109.025 86.255 118.305 86.935 ;
        RECT 110.385 86.035 111.305 86.255 ;
        RECT 115.970 86.135 118.305 86.255 ;
        RECT 117.385 86.025 118.305 86.135 ;
        RECT 118.695 86.025 120.045 86.935 ;
        RECT 120.065 86.125 121.895 86.935 ;
        RECT 122.365 86.125 123.735 86.935 ;
      LAYER nwell ;
        RECT 5.330 82.905 123.930 85.735 ;
      LAYER pwell ;
        RECT 5.525 81.705 6.895 82.515 ;
        RECT 6.905 81.705 10.575 82.515 ;
        RECT 10.585 81.705 11.955 82.485 ;
        RECT 12.895 81.705 14.245 82.615 ;
        RECT 14.275 81.705 15.625 82.615 ;
        RECT 15.645 81.705 18.395 82.515 ;
        RECT 18.415 81.790 18.845 82.575 ;
        RECT 18.865 81.705 21.615 82.515 ;
        RECT 22.280 81.705 25.755 82.615 ;
        RECT 25.765 81.705 31.275 82.515 ;
        RECT 31.285 81.705 36.795 82.515 ;
        RECT 36.805 81.705 39.555 82.515 ;
        RECT 40.025 82.385 40.955 82.615 ;
        RECT 40.025 81.705 43.925 82.385 ;
        RECT 44.175 81.790 44.605 82.575 ;
        RECT 44.625 82.385 45.555 82.615 ;
        RECT 44.625 81.705 48.525 82.385 ;
        RECT 48.765 81.705 50.595 82.515 ;
        RECT 51.260 81.705 54.735 82.615 ;
        RECT 54.745 82.415 55.690 82.615 ;
        RECT 54.745 81.735 57.495 82.415 ;
        RECT 54.745 81.705 55.690 81.735 ;
        RECT 5.665 81.495 5.835 81.705 ;
        RECT 7.045 81.495 7.215 81.705 ;
        RECT 11.645 81.515 11.815 81.705 ;
        RECT 12.115 81.550 12.275 81.660 ;
        RECT 12.565 81.495 12.735 81.685 ;
        RECT 13.945 81.515 14.115 81.705 ;
        RECT 15.325 81.515 15.495 81.705 ;
        RECT 15.785 81.515 15.955 81.705 ;
        RECT 18.095 81.540 18.255 81.650 ;
        RECT 19.005 81.515 19.175 81.705 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.685 12.415 81.495 ;
        RECT 12.425 80.685 17.935 81.495 ;
        RECT 18.865 81.465 19.810 81.495 ;
        RECT 21.300 81.465 21.470 81.685 ;
        RECT 21.770 81.655 21.940 81.685 ;
        RECT 21.760 81.545 21.940 81.655 ;
        RECT 21.770 81.495 21.940 81.545 ;
        RECT 25.440 81.515 25.610 81.705 ;
        RECT 25.905 81.515 26.075 81.705 ;
        RECT 28.660 81.495 28.830 81.685 ;
        RECT 29.125 81.495 29.295 81.685 ;
        RECT 30.960 81.545 31.080 81.655 ;
        RECT 31.425 81.515 31.595 81.705 ;
        RECT 31.885 81.495 32.055 81.685 ;
        RECT 35.565 81.495 35.735 81.685 ;
        RECT 36.945 81.515 37.115 81.705 ;
        RECT 37.865 81.495 38.035 81.685 ;
        RECT 38.325 81.495 38.495 81.685 ;
        RECT 39.705 81.655 39.875 81.685 ;
        RECT 39.700 81.545 39.875 81.655 ;
        RECT 39.705 81.495 39.875 81.545 ;
        RECT 40.440 81.515 40.610 81.705 ;
        RECT 45.040 81.515 45.210 81.705 ;
        RECT 48.905 81.515 49.075 81.705 ;
        RECT 54.420 81.685 54.590 81.705 ;
        RECT 49.365 81.495 49.535 81.685 ;
        RECT 50.740 81.545 50.860 81.655 ;
        RECT 53.960 81.495 54.130 81.685 ;
        RECT 54.420 81.515 54.600 81.685 ;
        RECT 57.180 81.515 57.350 81.735 ;
        RECT 57.505 81.705 60.255 82.515 ;
        RECT 60.275 81.705 61.625 82.615 ;
        RECT 62.105 82.385 63.035 82.615 ;
        RECT 62.105 81.705 66.005 82.385 ;
        RECT 66.440 81.705 69.915 82.615 ;
        RECT 69.935 81.790 70.365 82.575 ;
        RECT 70.385 81.705 73.595 82.615 ;
        RECT 73.605 81.705 79.115 82.515 ;
        RECT 79.125 81.705 81.875 82.515 ;
        RECT 82.345 82.385 83.275 82.615 ;
        RECT 82.345 81.705 86.245 82.385 ;
        RECT 86.485 81.705 91.995 82.515 ;
        RECT 92.005 81.705 95.675 82.515 ;
        RECT 95.695 81.790 96.125 82.575 ;
        RECT 96.145 81.705 98.895 82.515 ;
        RECT 99.560 81.705 103.035 82.615 ;
        RECT 103.045 81.705 106.520 82.615 ;
        RECT 110.845 82.385 111.775 82.615 ;
        RECT 113.145 82.385 114.065 82.605 ;
        RECT 120.145 82.505 121.065 82.615 ;
        RECT 118.730 82.385 121.065 82.505 ;
        RECT 107.875 81.705 111.775 82.385 ;
        RECT 111.785 81.705 121.065 82.385 ;
        RECT 121.455 81.790 121.885 82.575 ;
        RECT 122.365 81.705 123.735 82.515 ;
        RECT 18.865 80.785 21.615 81.465 ;
        RECT 18.865 80.585 19.810 80.785 ;
        RECT 21.625 80.585 25.100 81.495 ;
        RECT 25.500 80.585 28.975 81.495 ;
        RECT 28.985 80.685 30.815 81.495 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 31.745 80.685 35.415 81.495 ;
        RECT 35.425 80.685 36.795 81.495 ;
        RECT 36.805 80.715 38.175 81.495 ;
        RECT 38.185 80.715 39.555 81.495 ;
        RECT 39.565 80.815 48.845 81.495 ;
        RECT 40.925 80.595 41.845 80.815 ;
        RECT 46.510 80.695 48.845 80.815 ;
        RECT 47.925 80.585 48.845 80.695 ;
        RECT 49.225 80.685 50.595 81.495 ;
        RECT 50.800 80.585 54.275 81.495 ;
        RECT 54.430 81.465 54.600 81.515 ;
        RECT 57.645 81.495 57.815 81.705 ;
        RECT 60.405 81.515 60.575 81.705 ;
        RECT 61.780 81.545 61.900 81.655 ;
        RECT 62.520 81.515 62.690 81.705 ;
        RECT 63.165 81.495 63.335 81.685 ;
        RECT 65.925 81.495 66.095 81.685 ;
        RECT 69.600 81.515 69.770 81.705 ;
        RECT 73.285 81.515 73.455 81.705 ;
        RECT 73.745 81.515 73.915 81.705 ;
        RECT 75.585 81.495 75.755 81.685 ;
        RECT 76.965 81.495 77.135 81.685 ;
        RECT 79.265 81.495 79.435 81.705 ;
        RECT 79.725 81.495 79.895 81.685 ;
        RECT 82.025 81.655 82.195 81.685 ;
        RECT 82.020 81.545 82.195 81.655 ;
        RECT 82.480 81.545 82.600 81.655 ;
        RECT 82.025 81.495 82.195 81.545 ;
        RECT 82.760 81.515 82.930 81.705 ;
        RECT 83.400 81.545 83.520 81.655 ;
        RECT 86.625 81.515 86.795 81.705 ;
        RECT 87.080 81.495 87.250 81.685 ;
        RECT 56.090 81.465 57.035 81.495 ;
        RECT 54.285 80.785 57.035 81.465 ;
        RECT 56.090 80.585 57.035 80.785 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 57.505 80.685 63.015 81.495 ;
        RECT 63.025 80.685 65.775 81.495 ;
        RECT 65.785 80.815 75.065 81.495 ;
        RECT 67.145 80.595 68.065 80.815 ;
        RECT 72.730 80.695 75.065 80.815 ;
        RECT 74.145 80.585 75.065 80.695 ;
        RECT 75.455 80.585 76.805 81.495 ;
        RECT 76.825 80.685 78.195 81.495 ;
        RECT 78.205 80.715 79.575 81.495 ;
        RECT 79.585 80.685 80.955 81.495 ;
        RECT 80.975 80.585 82.325 81.495 ;
        RECT 82.815 80.625 83.245 81.410 ;
        RECT 83.920 80.585 87.395 81.495 ;
        RECT 87.550 81.465 87.720 81.685 ;
        RECT 90.305 81.495 90.475 81.685 ;
        RECT 92.145 81.515 92.315 81.705 ;
        RECT 95.830 81.495 96.000 81.685 ;
        RECT 96.285 81.515 96.455 81.705 ;
        RECT 99.040 81.545 99.160 81.655 ;
        RECT 102.720 81.495 102.890 81.705 ;
        RECT 103.190 81.685 103.360 81.705 ;
        RECT 103.185 81.515 103.360 81.685 ;
        RECT 106.875 81.550 107.035 81.660 ;
        RECT 103.185 81.495 103.355 81.515 ;
        RECT 109.165 81.495 109.335 81.685 ;
        RECT 110.545 81.495 110.715 81.685 ;
        RECT 111.190 81.515 111.360 81.705 ;
        RECT 111.925 81.515 112.095 81.705 ;
        RECT 112.200 81.495 112.370 81.685 ;
        RECT 116.985 81.495 117.155 81.685 ;
        RECT 117.445 81.495 117.615 81.685 ;
        RECT 121.125 81.495 121.295 81.685 ;
        RECT 122.040 81.545 122.160 81.655 ;
        RECT 123.425 81.495 123.595 81.705 ;
        RECT 89.210 81.465 90.155 81.495 ;
        RECT 87.405 80.785 90.155 81.465 ;
        RECT 89.210 80.585 90.155 80.785 ;
        RECT 90.165 80.685 95.675 81.495 ;
        RECT 95.685 80.585 99.160 81.495 ;
        RECT 99.560 80.585 103.035 81.495 ;
        RECT 103.045 80.685 108.555 81.495 ;
        RECT 108.575 80.625 109.005 81.410 ;
        RECT 109.025 80.715 110.395 81.495 ;
        RECT 110.405 80.685 111.775 81.495 ;
        RECT 111.785 80.815 115.685 81.495 ;
        RECT 111.785 80.585 112.715 80.815 ;
        RECT 115.935 80.585 117.285 81.495 ;
        RECT 117.305 80.685 120.975 81.495 ;
        RECT 120.985 80.685 122.355 81.495 ;
        RECT 122.365 80.685 123.735 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 123.930 80.295 ;
      LAYER pwell ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 6.905 76.265 12.415 77.075 ;
        RECT 13.345 76.945 14.275 77.175 ;
        RECT 13.345 76.265 17.245 76.945 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 19.325 76.975 20.270 77.175 ;
        RECT 19.325 76.295 22.075 76.975 ;
        RECT 19.325 76.265 20.270 76.295 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 7.045 76.055 7.215 76.265 ;
        RECT 9.800 76.105 9.920 76.215 ;
        RECT 11.185 76.055 11.355 76.245 ;
        RECT 12.565 76.055 12.735 76.245 ;
        RECT 13.760 76.075 13.930 76.265 ;
        RECT 13.945 76.055 14.115 76.245 ;
        RECT 14.400 76.105 14.520 76.215 ;
        RECT 15.140 76.055 15.310 76.245 ;
        RECT 17.635 76.110 17.795 76.220 ;
        RECT 19.005 76.215 19.175 76.245 ;
        RECT 19.000 76.105 19.175 76.215 ;
        RECT 19.005 76.055 19.175 76.105 ;
        RECT 21.760 76.075 21.930 76.295 ;
        RECT 22.085 76.265 25.560 77.175 ;
        RECT 25.765 76.265 27.135 77.075 ;
        RECT 27.145 76.975 28.090 77.175 ;
        RECT 27.145 76.295 29.895 76.975 ;
        RECT 27.145 76.265 28.090 76.295 ;
        RECT 22.230 76.075 22.400 76.265 ;
        RECT 22.680 76.105 22.800 76.215 ;
        RECT 23.150 76.055 23.320 76.245 ;
        RECT 25.905 76.075 26.075 76.265 ;
        RECT 26.830 76.055 27.000 76.245 ;
        RECT 29.580 76.075 29.750 76.295 ;
        RECT 29.905 76.265 33.575 77.075 ;
        RECT 33.585 76.265 34.955 77.075 ;
        RECT 39.475 76.945 40.405 77.165 ;
        RECT 43.235 76.945 44.155 77.175 ;
        RECT 34.965 76.265 44.155 76.945 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 44.635 76.265 45.985 77.175 ;
        RECT 46.005 76.265 51.515 77.075 ;
        RECT 51.525 76.265 57.035 77.075 ;
        RECT 57.045 76.265 62.555 77.075 ;
        RECT 62.565 76.265 65.315 77.075 ;
        RECT 65.325 76.945 66.670 77.175 ;
        RECT 65.325 76.265 67.155 76.945 ;
        RECT 67.165 76.265 69.915 77.075 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 70.580 76.265 74.055 77.175 ;
        RECT 74.065 76.265 75.895 77.075 ;
        RECT 77.265 76.945 78.185 77.165 ;
        RECT 84.265 77.065 85.185 77.175 ;
        RECT 82.850 76.945 85.185 77.065 ;
        RECT 75.905 76.265 85.185 76.945 ;
        RECT 85.565 76.945 86.495 77.175 ;
        RECT 85.565 76.265 89.465 76.945 ;
        RECT 89.705 76.265 95.215 77.075 ;
        RECT 95.695 76.350 96.125 77.135 ;
        RECT 96.145 76.265 101.655 77.075 ;
        RECT 101.665 76.265 107.175 77.075 ;
        RECT 107.185 76.265 109.015 77.075 ;
        RECT 109.485 76.265 110.855 77.045 ;
        RECT 112.225 76.945 113.145 77.165 ;
        RECT 119.225 77.065 120.145 77.175 ;
        RECT 117.810 76.945 120.145 77.065 ;
        RECT 110.865 76.265 120.145 76.945 ;
        RECT 121.455 76.350 121.885 77.135 ;
        RECT 122.365 76.265 123.735 77.075 ;
        RECT 30.045 76.075 30.215 76.265 ;
        RECT 30.515 76.100 30.675 76.210 ;
        RECT 31.885 76.055 32.055 76.245 ;
        RECT 33.725 76.075 33.895 76.265 ;
        RECT 35.105 76.075 35.275 76.265 ;
        RECT 37.405 76.055 37.575 76.245 ;
        RECT 39.240 76.105 39.360 76.215 ;
        RECT 39.705 76.055 39.875 76.245 ;
        RECT 41.085 76.055 41.255 76.245 ;
        RECT 44.765 76.075 44.935 76.265 ;
        RECT 46.145 76.075 46.315 76.265 ;
        RECT 46.605 76.055 46.775 76.245 ;
        RECT 51.665 76.075 51.835 76.265 ;
        RECT 52.135 76.100 52.295 76.210 ;
        RECT 56.260 76.055 56.430 76.245 ;
        RECT 56.720 76.105 56.840 76.215 ;
        RECT 57.185 76.075 57.355 76.265 ;
        RECT 59.945 76.055 60.115 76.245 ;
        RECT 60.405 76.055 60.575 76.245 ;
        RECT 62.705 76.075 62.875 76.265 ;
        RECT 63.625 76.055 63.795 76.245 ;
        RECT 64.085 76.055 64.255 76.245 ;
        RECT 66.845 76.075 67.015 76.265 ;
        RECT 67.305 76.075 67.475 76.265 ;
        RECT 73.285 76.055 73.455 76.245 ;
        RECT 73.740 76.075 73.910 76.265 ;
        RECT 74.205 76.075 74.375 76.265 ;
        RECT 76.045 76.075 76.215 76.265 ;
        RECT 78.800 76.105 78.920 76.215 ;
        RECT 82.480 76.055 82.650 76.245 ;
        RECT 85.980 76.075 86.150 76.265 ;
        RECT 89.845 76.245 90.015 76.265 ;
        RECT 86.620 76.055 86.790 76.245 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 6.905 75.245 9.655 76.055 ;
        RECT 10.125 75.275 11.495 76.055 ;
        RECT 11.505 75.275 12.875 76.055 ;
        RECT 12.895 75.145 14.245 76.055 ;
        RECT 14.725 75.375 18.625 76.055 ;
        RECT 14.725 75.145 15.655 75.375 ;
        RECT 18.865 75.245 22.535 76.055 ;
        RECT 23.005 75.145 26.480 76.055 ;
        RECT 26.685 75.145 30.160 76.055 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 31.745 75.245 37.255 76.055 ;
        RECT 37.265 75.245 39.095 76.055 ;
        RECT 39.575 75.145 40.925 76.055 ;
        RECT 40.945 75.245 46.455 76.055 ;
        RECT 46.465 75.245 51.975 76.055 ;
        RECT 53.100 75.145 56.575 76.055 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.515 75.375 60.255 76.055 ;
        RECT 60.265 75.245 62.095 76.055 ;
        RECT 62.105 75.375 63.935 76.055 ;
        RECT 63.945 75.375 73.050 76.055 ;
        RECT 62.105 75.145 63.450 75.375 ;
        RECT 73.145 75.245 78.655 76.055 ;
        RECT 79.320 75.145 82.795 76.055 ;
        RECT 82.815 75.185 83.245 75.970 ;
        RECT 83.460 75.145 86.935 76.055 ;
        RECT 87.090 76.025 87.260 76.245 ;
        RECT 89.845 76.075 90.020 76.245 ;
        RECT 88.750 76.025 89.695 76.055 ;
        RECT 89.850 76.025 90.020 76.075 ;
        RECT 92.605 76.055 92.775 76.245 ;
        RECT 93.990 76.055 94.160 76.245 ;
        RECT 95.360 76.105 95.480 76.215 ;
        RECT 96.285 76.075 96.455 76.265 ;
        RECT 97.670 76.055 97.840 76.245 ;
        RECT 101.805 76.075 101.975 76.265 ;
        RECT 102.265 76.055 102.435 76.245 ;
        RECT 102.725 76.055 102.895 76.245 ;
        RECT 107.325 76.075 107.495 76.265 ;
        RECT 109.165 76.215 109.335 76.245 ;
        RECT 108.240 76.105 108.360 76.215 ;
        RECT 109.160 76.105 109.335 76.215 ;
        RECT 109.165 76.055 109.335 76.105 ;
        RECT 109.625 76.075 109.795 76.265 ;
        RECT 111.005 76.075 111.175 76.265 ;
        RECT 111.920 76.105 112.040 76.215 ;
        RECT 112.660 76.055 112.830 76.245 ;
        RECT 116.525 76.055 116.695 76.245 ;
        RECT 120.675 76.110 120.835 76.220 ;
        RECT 122.040 76.105 122.160 76.215 ;
        RECT 123.425 76.055 123.595 76.265 ;
        RECT 91.510 76.025 92.455 76.055 ;
        RECT 86.945 75.345 89.695 76.025 ;
        RECT 89.705 75.345 92.455 76.025 ;
        RECT 88.750 75.145 89.695 75.345 ;
        RECT 91.510 75.145 92.455 75.345 ;
        RECT 92.465 75.245 93.835 76.055 ;
        RECT 93.845 75.145 97.320 76.055 ;
        RECT 97.525 75.145 101.000 76.055 ;
        RECT 101.205 75.275 102.575 76.055 ;
        RECT 102.585 75.245 108.095 76.055 ;
        RECT 108.575 75.185 109.005 75.970 ;
        RECT 109.025 75.245 111.775 76.055 ;
        RECT 112.245 75.375 116.145 76.055 ;
        RECT 112.245 75.145 113.175 75.375 ;
        RECT 116.385 75.245 121.895 76.055 ;
        RECT 122.365 75.245 123.735 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 123.930 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 8.725 71.505 9.645 71.725 ;
        RECT 15.725 71.625 16.645 71.735 ;
        RECT 14.310 71.505 16.645 71.625 ;
        RECT 7.365 70.825 16.645 71.505 ;
        RECT 17.035 70.825 18.385 71.735 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 18.865 70.825 22.535 71.635 ;
        RECT 22.545 70.825 23.915 71.635 ;
        RECT 23.925 70.825 27.400 71.735 ;
        RECT 27.800 70.825 31.275 71.735 ;
        RECT 31.285 70.825 33.115 71.635 ;
        RECT 33.320 70.825 36.795 71.735 ;
        RECT 36.805 70.825 42.315 71.635 ;
        RECT 42.325 70.825 44.155 71.635 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.625 70.825 48.295 71.635 ;
        RECT 48.775 70.825 50.125 71.735 ;
        RECT 50.340 70.825 53.815 71.735 ;
        RECT 54.020 70.825 57.495 71.735 ;
        RECT 57.505 70.825 60.980 71.735 ;
        RECT 61.185 70.825 63.015 71.635 ;
        RECT 63.025 70.825 65.765 71.505 ;
        RECT 65.785 70.825 67.155 71.635 ;
        RECT 67.650 71.505 68.995 71.735 ;
        RECT 67.165 70.825 68.995 71.505 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 71.305 71.505 72.235 71.735 ;
        RECT 71.305 70.825 75.205 71.505 ;
        RECT 75.445 70.825 80.955 71.635 ;
        RECT 80.965 70.825 86.475 71.635 ;
        RECT 86.485 70.825 88.315 71.635 ;
        RECT 88.980 70.825 92.455 71.735 ;
        RECT 92.465 70.825 95.215 71.635 ;
        RECT 95.695 70.910 96.125 71.695 ;
        RECT 96.145 70.825 98.895 71.635 ;
        RECT 100.725 71.505 101.645 71.725 ;
        RECT 107.725 71.625 108.645 71.735 ;
        RECT 106.310 71.505 108.645 71.625 ;
        RECT 99.365 70.825 108.645 71.505 ;
        RECT 109.035 70.825 110.385 71.735 ;
        RECT 110.405 70.825 112.235 71.635 ;
        RECT 115.905 71.505 116.835 71.735 ;
        RECT 112.935 70.825 116.835 71.505 ;
        RECT 116.845 70.825 118.215 71.605 ;
        RECT 118.225 70.825 120.975 71.635 ;
        RECT 121.455 70.910 121.885 71.695 ;
        RECT 122.365 70.825 123.735 71.635 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.045 70.775 7.215 70.805 ;
        RECT 7.040 70.665 7.215 70.775 ;
        RECT 7.045 70.615 7.215 70.665 ;
        RECT 7.505 70.635 7.675 70.825 ;
        RECT 8.425 70.615 8.595 70.805 ;
        RECT 18.085 70.635 18.255 70.825 ;
        RECT 19.005 70.635 19.175 70.825 ;
        RECT 19.920 70.615 20.090 70.805 ;
        RECT 20.385 70.615 20.555 70.805 ;
        RECT 22.685 70.635 22.855 70.825 ;
        RECT 24.070 70.615 24.240 70.825 ;
        RECT 27.745 70.615 27.915 70.805 ;
        RECT 30.960 70.635 31.130 70.825 ;
        RECT 31.425 70.635 31.595 70.825 ;
        RECT 31.885 70.615 32.055 70.805 ;
        RECT 35.565 70.615 35.735 70.805 ;
        RECT 36.480 70.635 36.650 70.825 ;
        RECT 36.945 70.635 37.115 70.825 ;
        RECT 37.865 70.615 38.035 70.805 ;
        RECT 38.325 70.615 38.495 70.805 ;
        RECT 41.085 70.615 41.255 70.805 ;
        RECT 41.545 70.615 41.715 70.805 ;
        RECT 42.465 70.635 42.635 70.825 ;
        RECT 44.300 70.665 44.420 70.775 ;
        RECT 44.765 70.615 44.935 70.825 ;
        RECT 48.440 70.665 48.560 70.775 ;
        RECT 48.905 70.635 49.075 70.825 ;
        RECT 53.500 70.635 53.670 70.825 ;
        RECT 54.425 70.615 54.595 70.805 ;
        RECT 57.180 70.635 57.350 70.825 ;
        RECT 57.650 70.805 57.820 70.825 ;
        RECT 57.645 70.635 57.820 70.805 ;
        RECT 60.400 70.665 60.520 70.775 ;
        RECT 61.325 70.635 61.495 70.825 ;
        RECT 57.645 70.615 57.815 70.635 ;
        RECT 63.165 70.615 63.335 70.825 ;
        RECT 63.620 70.665 63.740 70.775 ;
        RECT 65.465 70.615 65.635 70.805 ;
        RECT 65.925 70.615 66.095 70.825 ;
        RECT 67.305 70.635 67.475 70.825 ;
        RECT 67.765 70.615 67.935 70.805 ;
        RECT 69.155 70.670 69.315 70.780 ;
        RECT 69.605 70.615 69.775 70.805 ;
        RECT 70.535 70.670 70.695 70.780 ;
        RECT 71.445 70.615 71.615 70.805 ;
        RECT 71.720 70.635 71.890 70.825 ;
        RECT 72.825 70.615 72.995 70.805 ;
        RECT 75.585 70.635 75.755 70.825 ;
        RECT 76.780 70.615 76.950 70.805 ;
        RECT 81.105 70.635 81.275 70.825 ;
        RECT 81.565 70.615 81.735 70.805 ;
        RECT 82.035 70.660 82.195 70.770 ;
        RECT 83.405 70.615 83.575 70.805 ;
        RECT 86.625 70.635 86.795 70.825 ;
        RECT 88.460 70.665 88.580 70.775 ;
        RECT 88.925 70.615 89.095 70.805 ;
        RECT 90.770 70.615 90.940 70.805 ;
        RECT 92.140 70.635 92.310 70.825 ;
        RECT 92.605 70.635 92.775 70.825 ;
        RECT 94.450 70.615 94.620 70.805 ;
        RECT 95.360 70.665 95.480 70.775 ;
        RECT 96.285 70.635 96.455 70.825 ;
        RECT 99.040 70.665 99.160 70.775 ;
        RECT 99.505 70.635 99.675 70.825 ;
        RECT 101.340 70.615 101.510 70.805 ;
        RECT 102.080 70.615 102.250 70.805 ;
        RECT 105.945 70.615 106.115 70.805 ;
        RECT 109.165 70.615 109.335 70.805 ;
        RECT 110.085 70.635 110.255 70.825 ;
        RECT 110.545 70.635 110.715 70.825 ;
        RECT 111.000 70.665 111.120 70.775 ;
        RECT 111.465 70.615 111.635 70.805 ;
        RECT 112.380 70.665 112.500 70.775 ;
        RECT 116.250 70.635 116.420 70.825 ;
        RECT 117.905 70.635 118.075 70.825 ;
        RECT 118.365 70.635 118.535 70.825 ;
        RECT 121.125 70.775 121.295 70.805 ;
        RECT 121.120 70.665 121.295 70.775 ;
        RECT 122.040 70.665 122.160 70.775 ;
        RECT 121.125 70.615 121.295 70.665 ;
        RECT 123.425 70.615 123.595 70.825 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 6.905 69.805 8.275 70.615 ;
        RECT 8.285 69.935 17.475 70.615 ;
        RECT 12.795 69.715 13.725 69.935 ;
        RECT 16.555 69.705 17.475 69.935 ;
        RECT 17.625 69.705 20.235 70.615 ;
        RECT 20.245 69.805 23.915 70.615 ;
        RECT 23.925 69.705 27.400 70.615 ;
        RECT 27.605 69.805 31.275 70.615 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 31.745 69.805 35.415 70.615 ;
        RECT 35.425 69.805 36.795 70.615 ;
        RECT 36.805 69.835 38.175 70.615 ;
        RECT 38.185 69.805 40.015 70.615 ;
        RECT 40.035 69.705 41.385 70.615 ;
        RECT 41.405 69.805 44.155 70.615 ;
        RECT 44.625 69.935 53.905 70.615 ;
        RECT 45.985 69.715 46.905 69.935 ;
        RECT 51.570 69.815 53.905 69.935 ;
        RECT 52.985 69.705 53.905 69.815 ;
        RECT 54.285 69.805 57.035 70.615 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.505 69.805 60.255 70.615 ;
        RECT 60.755 69.705 63.475 70.615 ;
        RECT 63.945 69.935 65.775 70.615 ;
        RECT 65.785 69.935 67.615 70.615 ;
        RECT 67.625 69.935 69.455 70.615 ;
        RECT 69.465 69.935 71.295 70.615 ;
        RECT 63.945 69.705 65.290 69.935 ;
        RECT 66.270 69.705 67.615 69.935 ;
        RECT 68.110 69.705 69.455 69.935 ;
        RECT 69.950 69.705 71.295 69.935 ;
        RECT 71.305 69.835 72.675 70.615 ;
        RECT 72.685 69.805 76.355 70.615 ;
        RECT 76.365 69.935 80.265 70.615 ;
        RECT 76.365 69.705 77.295 69.935 ;
        RECT 80.515 69.705 81.865 70.615 ;
        RECT 82.815 69.745 83.245 70.530 ;
        RECT 83.265 69.805 88.775 70.615 ;
        RECT 88.785 69.805 90.615 70.615 ;
        RECT 90.625 69.705 94.100 70.615 ;
        RECT 94.305 69.705 97.780 70.615 ;
        RECT 98.180 69.705 101.655 70.615 ;
        RECT 101.665 69.935 105.565 70.615 ;
        RECT 101.665 69.705 102.595 69.935 ;
        RECT 105.805 69.805 108.555 70.615 ;
        RECT 108.575 69.745 109.005 70.530 ;
        RECT 109.025 69.805 110.855 70.615 ;
        RECT 111.325 69.935 120.605 70.615 ;
        RECT 112.685 69.715 113.605 69.935 ;
        RECT 118.270 69.815 120.605 69.935 ;
        RECT 119.685 69.705 120.605 69.815 ;
        RECT 120.985 69.805 122.355 70.615 ;
        RECT 122.365 69.805 123.735 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 123.930 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 6.905 65.385 12.415 66.195 ;
        RECT 12.425 65.385 17.935 66.195 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 18.865 65.385 24.375 66.195 ;
        RECT 24.385 65.385 28.055 66.195 ;
        RECT 28.065 65.385 29.435 66.165 ;
        RECT 29.445 66.065 30.375 66.295 ;
        RECT 35.865 66.065 36.785 66.285 ;
        RECT 42.865 66.185 43.785 66.295 ;
        RECT 41.450 66.065 43.785 66.185 ;
        RECT 29.445 65.385 33.345 66.065 ;
        RECT 34.505 65.385 43.785 66.065 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.625 65.385 47.375 66.195 ;
        RECT 47.385 65.385 48.755 66.165 ;
        RECT 48.765 66.065 49.695 66.295 ;
        RECT 48.765 65.385 52.665 66.065 ;
        RECT 52.905 65.385 58.415 66.195 ;
        RECT 58.425 65.385 62.095 66.195 ;
        RECT 62.565 66.065 63.910 66.295 ;
        RECT 64.405 66.065 65.750 66.295 ;
        RECT 62.565 65.385 64.395 66.065 ;
        RECT 64.405 65.385 66.235 66.065 ;
        RECT 66.245 65.385 67.615 66.195 ;
        RECT 67.625 66.065 68.970 66.295 ;
        RECT 67.625 65.385 69.455 66.065 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 70.385 65.385 72.215 66.195 ;
        RECT 72.225 65.385 73.595 66.165 ;
        RECT 74.965 66.065 75.885 66.285 ;
        RECT 81.965 66.185 82.885 66.295 ;
        RECT 80.550 66.065 82.885 66.185 ;
        RECT 73.605 65.385 82.885 66.065 ;
        RECT 83.265 65.385 85.875 66.295 ;
        RECT 86.025 65.385 89.695 66.195 ;
        RECT 90.165 66.065 91.095 66.295 ;
        RECT 90.165 65.385 94.065 66.065 ;
        RECT 94.305 65.385 95.675 66.195 ;
        RECT 95.695 65.470 96.125 66.255 ;
        RECT 96.145 65.385 101.655 66.195 ;
        RECT 101.665 65.385 107.175 66.195 ;
        RECT 107.185 65.385 112.695 66.195 ;
        RECT 115.905 66.065 116.835 66.295 ;
        RECT 112.935 65.385 116.835 66.065 ;
        RECT 116.855 65.385 118.205 66.295 ;
        RECT 118.225 65.385 120.975 66.195 ;
        RECT 121.455 65.470 121.885 66.255 ;
        RECT 122.365 65.385 123.735 66.195 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.045 65.175 7.215 65.385 ;
        RECT 10.725 65.175 10.895 65.365 ;
        RECT 12.565 65.195 12.735 65.385 ;
        RECT 13.025 65.175 13.195 65.365 ;
        RECT 13.490 65.175 13.660 65.365 ;
        RECT 16.255 65.220 16.415 65.330 ;
        RECT 17.440 65.175 17.610 65.365 ;
        RECT 18.080 65.225 18.200 65.335 ;
        RECT 19.005 65.195 19.175 65.385 ;
        RECT 21.580 65.175 21.750 65.365 ;
        RECT 24.525 65.195 24.695 65.385 ;
        RECT 25.440 65.225 25.560 65.335 ;
        RECT 26.180 65.175 26.350 65.365 ;
        RECT 29.125 65.195 29.295 65.385 ;
        RECT 29.860 65.195 30.030 65.385 ;
        RECT 30.045 65.175 30.215 65.365 ;
        RECT 31.885 65.175 32.055 65.365 ;
        RECT 33.265 65.175 33.435 65.365 ;
        RECT 33.735 65.230 33.895 65.340 ;
        RECT 34.645 65.195 34.815 65.385 ;
        RECT 37.220 65.175 37.390 65.365 ;
        RECT 41.085 65.175 41.255 65.365 ;
        RECT 44.765 65.195 44.935 65.385 ;
        RECT 46.605 65.175 46.775 65.365 ;
        RECT 48.445 65.195 48.615 65.385 ;
        RECT 49.180 65.195 49.350 65.385 ;
        RECT 51.205 65.175 51.375 65.365 ;
        RECT 51.940 65.175 52.110 65.365 ;
        RECT 53.045 65.195 53.215 65.385 ;
        RECT 55.805 65.175 55.975 65.365 ;
        RECT 57.645 65.175 57.815 65.365 ;
        RECT 58.565 65.195 58.735 65.385 ;
        RECT 62.240 65.225 62.360 65.335 ;
        RECT 63.165 65.175 63.335 65.365 ;
        RECT 64.085 65.195 64.255 65.385 ;
        RECT 65.925 65.175 66.095 65.385 ;
        RECT 66.385 65.195 66.555 65.385 ;
        RECT 67.765 65.175 67.935 65.365 ;
        RECT 69.145 65.195 69.315 65.385 ;
        RECT 69.600 65.330 69.720 65.335 ;
        RECT 69.600 65.225 69.775 65.330 ;
        RECT 69.615 65.220 69.775 65.225 ;
        RECT 70.525 65.175 70.695 65.385 ;
        RECT 72.365 65.195 72.535 65.385 ;
        RECT 73.745 65.195 73.915 65.385 ;
        RECT 83.410 65.365 83.580 65.385 ;
        RECT 80.645 65.175 80.815 65.365 ;
        RECT 81.105 65.175 81.275 65.365 ;
        RECT 83.405 65.195 83.580 65.365 ;
        RECT 86.165 65.195 86.335 65.385 ;
        RECT 83.405 65.175 83.575 65.195 ;
        RECT 88.005 65.175 88.175 65.365 ;
        RECT 88.465 65.175 88.635 65.365 ;
        RECT 89.840 65.225 89.960 65.335 ;
        RECT 90.580 65.195 90.750 65.385 ;
        RECT 91.235 65.220 91.395 65.330 ;
        RECT 94.445 65.195 94.615 65.385 ;
        RECT 95.550 65.175 95.720 65.365 ;
        RECT 96.285 65.175 96.455 65.385 ;
        RECT 97.665 65.175 97.835 65.365 ;
        RECT 100.700 65.175 100.870 65.365 ;
        RECT 101.805 65.195 101.975 65.385 ;
        RECT 104.565 65.175 104.735 65.365 ;
        RECT 107.325 65.195 107.495 65.385 ;
        RECT 108.240 65.225 108.360 65.335 ;
        RECT 109.165 65.175 109.335 65.365 ;
        RECT 111.925 65.175 112.095 65.365 ;
        RECT 116.250 65.195 116.420 65.385 ;
        RECT 117.905 65.195 118.075 65.385 ;
        RECT 118.365 65.195 118.535 65.385 ;
        RECT 121.125 65.335 121.295 65.365 ;
        RECT 121.120 65.225 121.295 65.335 ;
        RECT 122.040 65.225 122.160 65.335 ;
        RECT 121.125 65.175 121.295 65.225 ;
        RECT 123.425 65.175 123.595 65.385 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.365 10.575 65.175 ;
        RECT 10.585 64.365 11.955 65.175 ;
        RECT 11.965 64.395 13.335 65.175 ;
        RECT 13.345 64.265 15.955 65.175 ;
        RECT 17.025 64.495 20.925 65.175 ;
        RECT 21.165 64.495 25.065 65.175 ;
        RECT 25.765 64.495 29.665 65.175 ;
        RECT 17.025 64.265 17.955 64.495 ;
        RECT 21.165 64.265 22.095 64.495 ;
        RECT 25.765 64.265 26.695 64.495 ;
        RECT 29.905 64.365 31.275 65.175 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 31.755 64.265 33.105 65.175 ;
        RECT 33.125 64.365 36.795 65.175 ;
        RECT 36.805 64.495 40.705 65.175 ;
        RECT 36.805 64.265 37.735 64.495 ;
        RECT 40.945 64.365 46.455 65.175 ;
        RECT 46.465 64.365 50.135 65.175 ;
        RECT 50.145 64.395 51.515 65.175 ;
        RECT 51.525 64.495 55.425 65.175 ;
        RECT 51.525 64.265 52.455 64.495 ;
        RECT 55.665 64.365 57.035 65.175 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.505 64.365 63.015 65.175 ;
        RECT 63.025 64.365 65.775 65.175 ;
        RECT 65.785 64.495 67.615 65.175 ;
        RECT 67.625 64.495 69.455 65.175 ;
        RECT 70.385 64.495 79.575 65.175 ;
        RECT 66.270 64.265 67.615 64.495 ;
        RECT 68.110 64.265 69.455 64.495 ;
        RECT 74.895 64.275 75.825 64.495 ;
        RECT 78.655 64.265 79.575 64.495 ;
        RECT 79.595 64.265 80.945 65.175 ;
        RECT 80.965 64.365 82.795 65.175 ;
        RECT 82.815 64.305 83.245 65.090 ;
        RECT 83.265 64.365 86.935 65.175 ;
        RECT 86.945 64.395 88.315 65.175 ;
        RECT 88.325 64.495 91.065 65.175 ;
        RECT 92.235 64.495 96.135 65.175 ;
        RECT 95.205 64.265 96.135 64.495 ;
        RECT 96.145 64.395 97.515 65.175 ;
        RECT 97.525 64.365 100.275 65.175 ;
        RECT 100.285 64.495 104.185 65.175 ;
        RECT 100.285 64.265 101.215 64.495 ;
        RECT 104.425 64.365 108.095 65.175 ;
        RECT 108.575 64.305 109.005 65.090 ;
        RECT 109.025 64.365 111.775 65.175 ;
        RECT 111.785 64.495 120.975 65.175 ;
        RECT 116.295 64.275 117.225 64.495 ;
        RECT 120.055 64.265 120.975 64.495 ;
        RECT 120.985 64.365 122.355 65.175 ;
        RECT 122.365 64.365 123.735 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 123.930 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 12.335 60.625 13.265 60.845 ;
        RECT 16.095 60.625 17.015 60.855 ;
        RECT 7.825 59.945 17.015 60.625 ;
        RECT 17.025 59.945 18.395 60.725 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 19.785 60.625 20.715 60.855 ;
        RECT 19.785 59.945 23.685 60.625 ;
        RECT 23.925 59.945 26.675 60.755 ;
        RECT 28.505 60.625 29.425 60.845 ;
        RECT 35.505 60.745 36.425 60.855 ;
        RECT 34.090 60.625 36.425 60.745 ;
        RECT 27.145 59.945 36.425 60.625 ;
        RECT 36.805 59.945 42.315 60.755 ;
        RECT 42.325 59.945 44.155 60.755 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 44.625 59.945 45.995 60.755 ;
        RECT 46.015 59.945 47.365 60.855 ;
        RECT 47.395 59.945 48.745 60.855 ;
        RECT 50.125 60.625 51.045 60.845 ;
        RECT 57.125 60.745 58.045 60.855 ;
        RECT 55.710 60.625 58.045 60.745 ;
        RECT 48.765 59.945 58.045 60.625 ;
        RECT 59.355 59.945 62.095 60.625 ;
        RECT 62.595 59.945 65.315 60.855 ;
        RECT 65.810 60.625 67.155 60.855 ;
        RECT 65.325 59.945 67.155 60.625 ;
        RECT 67.165 59.945 69.915 60.755 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 72.995 60.855 ;
        RECT 73.145 59.945 78.655 60.755 ;
        RECT 78.665 59.945 84.175 60.755 ;
        RECT 89.615 60.625 90.545 60.845 ;
        RECT 93.375 60.625 94.295 60.855 ;
        RECT 85.105 59.945 94.295 60.625 ;
        RECT 94.305 59.945 95.675 60.755 ;
        RECT 95.695 60.030 96.125 60.815 ;
        RECT 100.655 60.625 101.585 60.845 ;
        RECT 104.415 60.625 105.335 60.855 ;
        RECT 109.855 60.625 110.785 60.845 ;
        RECT 113.615 60.625 114.535 60.855 ;
        RECT 96.145 59.945 105.335 60.625 ;
        RECT 105.345 59.945 114.535 60.625 ;
        RECT 114.545 60.625 115.475 60.855 ;
        RECT 114.545 59.945 118.445 60.625 ;
        RECT 118.685 59.945 120.055 60.725 ;
        RECT 120.065 59.945 121.435 60.755 ;
        RECT 121.455 60.030 121.885 60.815 ;
        RECT 122.365 59.945 123.735 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 7.045 59.735 7.215 59.925 ;
        RECT 7.965 59.755 8.135 59.945 ;
        RECT 9.800 59.785 9.920 59.895 ;
        RECT 11.185 59.735 11.355 59.925 ;
        RECT 12.565 59.735 12.735 59.925 ;
        RECT 13.025 59.735 13.195 59.925 ;
        RECT 18.085 59.755 18.255 59.945 ;
        RECT 19.015 59.790 19.175 59.900 ;
        RECT 20.200 59.755 20.370 59.945 ;
        RECT 22.225 59.735 22.395 59.925 ;
        RECT 24.065 59.755 24.235 59.945 ;
        RECT 26.820 59.785 26.940 59.895 ;
        RECT 27.285 59.755 27.455 59.945 ;
        RECT 31.885 59.735 32.055 59.925 ;
        RECT 35.575 59.780 35.735 59.890 ;
        RECT 36.945 59.755 37.115 59.945 ;
        RECT 37.405 59.735 37.575 59.925 ;
        RECT 38.140 59.735 38.310 59.925 ;
        RECT 42.015 59.780 42.175 59.890 ;
        RECT 42.465 59.755 42.635 59.945 ;
        RECT 42.925 59.735 43.095 59.925 ;
        RECT 44.765 59.755 44.935 59.945 ;
        RECT 46.145 59.755 46.315 59.945 ;
        RECT 47.525 59.755 47.695 59.945 ;
        RECT 48.905 59.755 49.075 59.945 ;
        RECT 52.860 59.735 53.030 59.925 ;
        RECT 56.720 59.785 56.840 59.895 ;
        RECT 57.645 59.735 57.815 59.925 ;
        RECT 58.575 59.790 58.735 59.900 ;
        RECT 61.785 59.755 61.955 59.945 ;
        RECT 62.240 59.785 62.360 59.895 ;
        RECT 63.165 59.735 63.335 59.925 ;
        RECT 65.005 59.755 65.175 59.945 ;
        RECT 65.465 59.755 65.635 59.945 ;
        RECT 67.305 59.755 67.475 59.945 ;
        RECT 68.685 59.735 68.855 59.925 ;
        RECT 70.530 59.755 70.700 59.945 ;
        RECT 73.285 59.755 73.455 59.945 ;
        RECT 74.205 59.735 74.375 59.925 ;
        RECT 75.590 59.735 75.760 59.925 ;
        RECT 78.345 59.735 78.515 59.925 ;
        RECT 78.805 59.755 78.975 59.945 ;
        RECT 82.035 59.780 82.195 59.890 ;
        RECT 83.410 59.735 83.580 59.925 ;
        RECT 84.335 59.790 84.495 59.900 ;
        RECT 85.245 59.755 85.415 59.945 ;
        RECT 86.165 59.735 86.335 59.925 ;
        RECT 89.845 59.735 90.015 59.925 ;
        RECT 91.225 59.735 91.395 59.925 ;
        RECT 94.445 59.755 94.615 59.945 ;
        RECT 96.285 59.755 96.455 59.945 ;
        RECT 96.745 59.735 96.915 59.925 ;
        RECT 99.505 59.735 99.675 59.925 ;
        RECT 100.885 59.735 101.055 59.925 ;
        RECT 102.265 59.735 102.435 59.925 ;
        RECT 105.485 59.755 105.655 59.945 ;
        RECT 105.945 59.735 106.115 59.925 ;
        RECT 107.325 59.735 107.495 59.925 ;
        RECT 109.165 59.735 109.335 59.925 ;
        RECT 114.960 59.755 115.130 59.945 ;
        RECT 118.365 59.735 118.535 59.925 ;
        RECT 119.745 59.735 119.915 59.945 ;
        RECT 120.205 59.755 120.375 59.945 ;
        RECT 122.040 59.785 122.160 59.895 ;
        RECT 123.425 59.735 123.595 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 58.925 9.655 59.735 ;
        RECT 10.125 58.955 11.495 59.735 ;
        RECT 11.515 58.825 12.865 59.735 ;
        RECT 12.885 59.055 22.075 59.735 ;
        RECT 22.085 59.055 31.275 59.735 ;
        RECT 17.395 58.835 18.325 59.055 ;
        RECT 21.155 58.825 22.075 59.055 ;
        RECT 26.595 58.835 27.525 59.055 ;
        RECT 30.355 58.825 31.275 59.055 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 58.925 35.415 59.735 ;
        RECT 36.345 58.955 37.715 59.735 ;
        RECT 37.725 59.055 41.625 59.735 ;
        RECT 42.785 59.055 52.065 59.735 ;
        RECT 37.725 58.825 38.655 59.055 ;
        RECT 44.145 58.835 45.065 59.055 ;
        RECT 49.730 58.935 52.065 59.055 ;
        RECT 51.145 58.825 52.065 58.935 ;
        RECT 52.445 59.055 56.345 59.735 ;
        RECT 52.445 58.825 53.375 59.055 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 57.505 58.925 63.015 59.735 ;
        RECT 63.025 58.925 68.535 59.735 ;
        RECT 68.545 58.925 74.055 59.735 ;
        RECT 74.065 58.925 75.435 59.735 ;
        RECT 75.445 58.825 78.055 59.735 ;
        RECT 78.205 58.925 81.875 59.735 ;
        RECT 82.815 58.865 83.245 59.650 ;
        RECT 83.265 58.825 85.875 59.735 ;
        RECT 86.025 58.925 89.695 59.735 ;
        RECT 89.715 58.825 91.065 59.735 ;
        RECT 91.085 58.925 96.595 59.735 ;
        RECT 96.605 58.925 99.355 59.735 ;
        RECT 99.365 58.955 100.735 59.735 ;
        RECT 100.755 58.825 102.105 59.735 ;
        RECT 102.125 58.925 105.795 59.735 ;
        RECT 105.815 58.825 107.165 59.735 ;
        RECT 107.185 58.955 108.555 59.735 ;
        RECT 108.575 58.865 109.005 59.650 ;
        RECT 109.025 59.055 118.215 59.735 ;
        RECT 113.535 58.835 114.465 59.055 ;
        RECT 117.295 58.825 118.215 59.055 ;
        RECT 118.235 58.825 119.585 59.735 ;
        RECT 119.605 58.925 122.355 59.735 ;
        RECT 122.365 58.925 123.735 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 123.930 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 54.505 8.735 55.315 ;
        RECT 13.715 55.185 14.645 55.405 ;
        RECT 17.475 55.185 18.395 55.415 ;
        RECT 9.205 54.505 18.395 55.185 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 18.875 54.505 20.225 55.415 ;
        RECT 20.705 54.505 22.075 55.285 ;
        RECT 38.095 55.185 39.025 55.405 ;
        RECT 41.855 55.185 42.775 55.415 ;
        RECT 22.500 54.505 23.455 55.185 ;
        RECT 23.550 54.505 32.655 55.185 ;
        RECT 33.585 54.505 42.775 55.185 ;
        RECT 42.795 54.505 44.145 55.415 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 44.625 54.505 46.455 55.315 ;
        RECT 46.465 54.505 47.835 55.285 ;
        RECT 47.845 54.505 53.355 55.315 ;
        RECT 53.365 54.505 58.875 55.315 ;
        RECT 58.885 54.505 62.555 55.315 ;
        RECT 63.240 54.735 65.995 55.415 ;
        RECT 63.725 54.505 65.995 54.735 ;
        RECT 66.245 55.185 67.590 55.415 ;
        RECT 66.245 54.505 68.075 55.185 ;
        RECT 68.095 54.505 69.445 55.415 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 70.870 55.185 72.215 55.415 ;
        RECT 70.385 54.505 72.215 55.185 ;
        RECT 72.225 54.505 77.735 55.315 ;
        RECT 77.745 54.505 79.115 55.285 ;
        RECT 79.135 54.505 80.485 55.415 ;
        RECT 80.505 54.505 91.515 55.415 ;
        RECT 91.740 54.505 95.215 55.415 ;
        RECT 95.695 54.590 96.125 55.375 ;
        RECT 96.145 54.505 98.895 55.315 ;
        RECT 99.780 54.505 100.735 55.185 ;
        RECT 100.745 54.505 109.850 55.185 ;
        RECT 109.945 54.505 112.695 55.315 ;
        RECT 113.175 54.505 114.525 55.415 ;
        RECT 114.545 54.505 120.055 55.315 ;
        RECT 120.065 54.505 121.435 55.315 ;
        RECT 121.455 54.590 121.885 55.375 ;
        RECT 122.365 54.505 123.735 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.045 54.295 7.215 54.505 ;
        RECT 8.880 54.345 9.000 54.455 ;
        RECT 9.345 54.315 9.515 54.505 ;
        RECT 9.800 54.345 9.920 54.455 ;
        RECT 10.265 54.295 10.435 54.485 ;
        RECT 12.105 54.295 12.275 54.485 ;
        RECT 13.940 54.345 14.060 54.455 ;
        RECT 15.325 54.295 15.495 54.485 ;
        RECT 15.785 54.295 15.955 54.485 ;
        RECT 19.925 54.315 20.095 54.505 ;
        RECT 20.380 54.345 20.500 54.455 ;
        RECT 20.845 54.315 21.015 54.505 ;
        RECT 21.305 54.295 21.475 54.485 ;
        RECT 22.225 54.315 22.395 54.485 ;
        RECT 26.825 54.295 26.995 54.485 ;
        RECT 30.505 54.295 30.675 54.485 ;
        RECT 30.960 54.345 31.080 54.455 ;
        RECT 31.885 54.295 32.055 54.485 ;
        RECT 32.345 54.315 32.515 54.505 ;
        RECT 32.815 54.350 32.975 54.460 ;
        RECT 33.725 54.315 33.895 54.505 ;
        RECT 37.400 54.345 37.520 54.455 ;
        RECT 37.865 54.315 38.035 54.485 ;
        RECT 43.845 54.315 44.015 54.505 ;
        RECT 44.765 54.315 44.935 54.505 ;
        RECT 47.525 54.315 47.695 54.505 ;
        RECT 47.985 54.295 48.155 54.505 ;
        RECT 48.440 54.345 48.560 54.455 ;
        RECT 52.120 54.295 52.290 54.485 ;
        RECT 52.585 54.295 52.755 54.485 ;
        RECT 53.505 54.315 53.675 54.505 ;
        RECT 56.275 54.340 56.435 54.450 ;
        RECT 57.645 54.295 57.815 54.485 ;
        RECT 59.025 54.315 59.195 54.505 ;
        RECT 65.925 54.485 65.995 54.505 ;
        RECT 61.325 54.295 61.495 54.485 ;
        RECT 62.700 54.345 62.820 54.455 ;
        RECT 65.925 54.295 66.095 54.485 ;
        RECT 67.765 54.315 67.935 54.505 ;
        RECT 68.225 54.315 68.395 54.505 ;
        RECT 69.600 54.345 69.720 54.455 ;
        RECT 70.525 54.295 70.695 54.505 ;
        RECT 72.365 54.295 72.535 54.505 ;
        RECT 73.745 54.295 73.915 54.485 ;
        RECT 78.805 54.315 78.975 54.505 ;
        RECT 80.185 54.315 80.355 54.505 ;
        RECT 80.650 54.315 80.820 54.505 ;
        RECT 92.145 54.295 92.315 54.485 ;
        RECT 92.605 54.295 92.775 54.485 ;
        RECT 94.900 54.315 95.070 54.505 ;
        RECT 95.360 54.345 95.480 54.455 ;
        RECT 96.285 54.315 96.455 54.505 ;
        RECT 99.050 54.455 99.220 54.485 ;
        RECT 98.135 54.340 98.295 54.450 ;
        RECT 99.040 54.345 99.220 54.455 ;
        RECT 99.050 54.295 99.220 54.345 ;
        RECT 99.505 54.315 99.675 54.485 ;
        RECT 100.885 54.315 101.055 54.505 ;
        RECT 102.725 54.295 102.895 54.485 ;
        RECT 108.240 54.345 108.360 54.455 ;
        RECT 109.165 54.295 109.335 54.485 ;
        RECT 110.085 54.315 110.255 54.505 ;
        RECT 112.840 54.345 112.960 54.455 ;
        RECT 113.305 54.315 113.475 54.505 ;
        RECT 114.685 54.295 114.855 54.505 ;
        RECT 120.205 54.295 120.375 54.505 ;
        RECT 122.040 54.345 122.160 54.455 ;
        RECT 123.425 54.295 123.595 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 6.905 53.485 9.655 54.295 ;
        RECT 10.125 53.615 11.955 54.295 ;
        RECT 11.965 53.485 13.795 54.295 ;
        RECT 14.275 53.385 15.625 54.295 ;
        RECT 15.645 53.485 21.155 54.295 ;
        RECT 21.165 53.485 26.675 54.295 ;
        RECT 26.685 53.485 29.435 54.295 ;
        RECT 29.455 53.385 30.805 54.295 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.745 53.485 37.255 54.295 ;
        RECT 38.140 53.615 39.095 54.295 ;
        RECT 39.190 53.615 48.295 54.295 ;
        RECT 48.960 53.385 52.435 54.295 ;
        RECT 52.445 53.485 56.115 54.295 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 57.505 53.485 61.175 54.295 ;
        RECT 61.185 54.065 62.755 54.295 ;
        RECT 64.845 54.255 65.765 54.295 ;
        RECT 64.845 54.065 65.775 54.255 ;
        RECT 61.185 53.705 65.775 54.065 ;
        RECT 61.185 53.615 65.765 53.705 ;
        RECT 62.765 53.385 65.765 53.615 ;
        RECT 65.785 53.385 70.335 54.295 ;
        RECT 70.385 53.615 72.215 54.295 ;
        RECT 70.870 53.385 72.215 53.615 ;
        RECT 72.225 53.485 73.595 54.295 ;
        RECT 73.605 53.615 82.795 54.295 ;
        RECT 78.115 53.395 79.045 53.615 ;
        RECT 81.875 53.385 82.795 53.615 ;
        RECT 82.815 53.425 83.245 54.210 ;
        RECT 83.350 53.615 92.455 54.295 ;
        RECT 92.465 53.485 97.975 54.295 ;
        RECT 98.905 53.385 102.380 54.295 ;
        RECT 102.585 53.485 108.095 54.295 ;
        RECT 108.575 53.425 109.005 54.210 ;
        RECT 109.025 53.485 114.535 54.295 ;
        RECT 114.545 53.485 120.055 54.295 ;
        RECT 120.065 53.485 121.895 54.295 ;
        RECT 122.365 53.485 123.735 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 123.930 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 6.905 49.065 12.415 49.875 ;
        RECT 12.425 49.065 17.935 49.875 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 18.865 49.065 22.535 49.875 ;
        RECT 23.005 49.065 26.480 49.975 ;
        RECT 26.685 49.065 30.160 49.975 ;
        RECT 30.365 49.065 35.875 49.875 ;
        RECT 35.885 49.065 41.395 49.875 ;
        RECT 41.405 49.065 44.155 49.875 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 45.225 49.065 47.835 49.975 ;
        RECT 47.845 49.065 49.675 49.875 ;
        RECT 49.880 49.065 53.355 49.975 ;
        RECT 53.560 49.065 57.035 49.975 ;
        RECT 57.045 49.065 62.555 49.875 ;
        RECT 62.565 49.065 64.395 49.875 ;
        RECT 65.080 49.295 67.835 49.975 ;
        RECT 65.565 49.065 67.835 49.295 ;
        RECT 68.085 49.745 69.430 49.975 ;
        RECT 68.085 49.065 69.915 49.745 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 70.625 49.295 73.380 49.975 ;
        RECT 74.090 49.745 75.435 49.975 ;
        RECT 70.625 49.065 72.895 49.295 ;
        RECT 73.605 49.065 75.435 49.745 ;
        RECT 75.445 49.065 76.815 49.875 ;
        RECT 79.585 49.745 80.515 49.975 ;
        RECT 76.825 49.065 79.565 49.745 ;
        RECT 79.585 49.065 83.485 49.745 ;
        RECT 83.920 49.065 87.395 49.975 ;
        RECT 87.405 49.065 90.880 49.975 ;
        RECT 91.085 49.065 94.560 49.975 ;
        RECT 95.695 49.150 96.125 49.935 ;
        RECT 96.340 49.065 99.815 49.975 ;
        RECT 99.825 49.065 103.300 49.975 ;
        RECT 103.505 49.065 106.980 49.975 ;
        RECT 107.185 49.065 112.695 49.875 ;
        RECT 112.705 49.065 118.215 49.875 ;
        RECT 118.225 49.065 120.975 49.875 ;
        RECT 121.455 49.150 121.885 49.935 ;
        RECT 122.365 49.065 123.735 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.045 48.855 7.215 49.065 ;
        RECT 10.725 48.855 10.895 49.045 ;
        RECT 12.565 48.875 12.735 49.065 ;
        RECT 13.025 48.855 13.195 49.045 ;
        RECT 14.405 48.855 14.575 49.045 ;
        RECT 15.785 48.855 15.955 49.045 ;
        RECT 16.240 48.905 16.360 49.015 ;
        RECT 16.980 48.855 17.150 49.045 ;
        RECT 18.080 48.905 18.200 49.015 ;
        RECT 19.005 48.875 19.175 49.065 ;
        RECT 20.845 48.855 21.015 49.045 ;
        RECT 22.680 48.905 22.800 49.015 ;
        RECT 23.150 48.855 23.320 49.065 ;
        RECT 26.830 48.875 27.000 49.065 ;
        RECT 30.040 48.855 30.210 49.045 ;
        RECT 30.505 48.875 30.675 49.065 ;
        RECT 35.100 48.855 35.270 49.045 ;
        RECT 35.565 48.855 35.735 49.045 ;
        RECT 36.025 48.875 36.195 49.065 ;
        RECT 37.865 48.855 38.035 49.045 ;
        RECT 38.325 48.855 38.495 49.045 ;
        RECT 41.545 48.875 41.715 49.065 ;
        RECT 43.845 48.855 44.015 49.045 ;
        RECT 44.760 48.905 44.880 49.015 ;
        RECT 47.520 48.875 47.690 49.065 ;
        RECT 47.985 48.875 48.155 49.065 ;
        RECT 53.040 49.045 53.210 49.065 ;
        RECT 48.905 48.855 49.075 49.045 ;
        RECT 52.580 48.855 52.750 49.045 ;
        RECT 53.040 48.875 53.215 49.045 ;
        RECT 56.720 48.875 56.890 49.065 ;
        RECT 57.185 48.875 57.355 49.065 ;
        RECT 53.045 48.855 53.215 48.875 ;
        RECT 57.645 48.855 57.815 49.045 ;
        RECT 59.025 48.855 59.195 49.045 ;
        RECT 62.705 48.875 62.875 49.065 ;
        RECT 67.765 49.045 67.835 49.065 ;
        RECT 64.540 49.010 64.660 49.015 ;
        RECT 64.540 48.905 64.715 49.010 ;
        RECT 64.555 48.900 64.715 48.905 ;
        RECT 67.765 48.875 67.935 49.045 ;
        RECT 68.225 48.875 68.395 49.045 ;
        RECT 68.225 48.855 68.295 48.875 ;
        RECT 68.685 48.855 68.855 49.045 ;
        RECT 69.605 48.875 69.775 49.065 ;
        RECT 70.625 49.045 70.695 49.065 ;
        RECT 70.525 48.875 70.695 49.045 ;
        RECT 73.745 48.875 73.915 49.065 ;
        RECT 74.205 48.855 74.375 49.045 ;
        RECT 75.585 48.875 75.755 49.065 ;
        RECT 76.965 48.875 77.135 49.065 ;
        RECT 79.725 48.855 79.895 49.045 ;
        RECT 80.000 48.875 80.170 49.065 ;
        RECT 82.480 48.905 82.600 49.015 ;
        RECT 83.680 48.855 83.850 49.045 ;
        RECT 87.080 48.875 87.250 49.065 ;
        RECT 87.550 48.875 87.720 49.065 ;
        RECT 90.760 48.855 90.930 49.045 ;
        RECT 91.230 48.875 91.400 49.065 ;
        RECT 94.440 48.855 94.610 49.045 ;
        RECT 94.905 48.855 95.075 49.045 ;
        RECT 98.595 48.900 98.755 49.010 ;
        RECT 99.500 48.875 99.670 49.065 ;
        RECT 99.970 48.875 100.140 49.065 ;
        RECT 102.910 48.855 103.080 49.045 ;
        RECT 103.650 48.875 103.820 49.065 ;
        RECT 104.565 48.855 104.735 49.045 ;
        RECT 105.035 48.900 105.195 49.010 ;
        RECT 105.945 48.855 106.115 49.045 ;
        RECT 107.325 48.855 107.495 49.065 ;
        RECT 110.085 48.855 110.255 49.045 ;
        RECT 110.545 48.855 110.715 49.045 ;
        RECT 112.845 48.875 113.015 49.065 ;
        RECT 116.065 48.855 116.235 49.045 ;
        RECT 118.365 48.875 118.535 49.065 ;
        RECT 121.120 48.905 121.240 49.015 ;
        RECT 121.595 48.900 121.755 49.010 ;
        RECT 122.040 48.905 122.160 49.015 ;
        RECT 123.425 48.855 123.595 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.045 10.575 48.855 ;
        RECT 10.585 48.045 11.955 48.855 ;
        RECT 11.965 48.075 13.335 48.855 ;
        RECT 13.345 48.075 14.715 48.855 ;
        RECT 14.735 47.945 16.085 48.855 ;
        RECT 16.565 48.175 20.465 48.855 ;
        RECT 16.565 47.945 17.495 48.175 ;
        RECT 20.705 48.045 22.535 48.855 ;
        RECT 23.005 47.945 26.480 48.855 ;
        RECT 26.880 47.945 30.355 48.855 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 31.940 47.945 35.415 48.855 ;
        RECT 35.425 48.045 36.795 48.855 ;
        RECT 36.805 48.075 38.175 48.855 ;
        RECT 38.185 48.045 43.695 48.855 ;
        RECT 43.705 48.045 46.455 48.855 ;
        RECT 46.475 48.175 49.215 48.855 ;
        RECT 49.420 47.945 52.895 48.855 ;
        RECT 52.905 48.045 56.575 48.855 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.515 47.945 58.865 48.855 ;
        RECT 58.885 48.045 64.395 48.855 ;
        RECT 66.025 48.625 68.295 48.855 ;
        RECT 65.540 47.945 68.295 48.625 ;
        RECT 68.545 48.045 74.055 48.855 ;
        RECT 74.065 48.045 79.575 48.855 ;
        RECT 79.585 48.045 82.335 48.855 ;
        RECT 82.815 47.985 83.245 48.770 ;
        RECT 83.265 48.175 87.165 48.855 ;
        RECT 83.265 47.945 84.195 48.175 ;
        RECT 87.600 47.945 91.075 48.855 ;
        RECT 91.280 47.945 94.755 48.855 ;
        RECT 94.765 48.045 98.435 48.855 ;
        RECT 99.595 48.175 103.495 48.855 ;
        RECT 102.565 47.945 103.495 48.175 ;
        RECT 103.505 48.075 104.875 48.855 ;
        RECT 105.805 48.075 107.175 48.855 ;
        RECT 107.185 48.045 108.555 48.855 ;
        RECT 108.575 47.985 109.005 48.770 ;
        RECT 109.035 47.945 110.385 48.855 ;
        RECT 110.405 48.045 115.915 48.855 ;
        RECT 115.925 48.045 121.435 48.855 ;
        RECT 122.365 48.045 123.735 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 123.930 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 8.735 44.435 ;
        RECT 13.715 44.305 14.645 44.525 ;
        RECT 17.475 44.305 18.395 44.535 ;
        RECT 9.205 43.625 18.395 44.305 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 18.865 44.305 19.795 44.535 ;
        RECT 18.865 43.625 22.765 44.305 ;
        RECT 23.005 43.625 25.755 44.435 ;
        RECT 25.960 43.625 29.435 44.535 ;
        RECT 29.445 43.625 34.955 44.435 ;
        RECT 39.475 44.305 40.405 44.525 ;
        RECT 43.235 44.305 44.155 44.535 ;
        RECT 34.965 43.625 44.155 44.305 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 44.635 43.625 45.985 44.535 ;
        RECT 46.005 43.625 47.375 44.435 ;
        RECT 47.525 43.625 50.135 44.535 ;
        RECT 50.145 43.625 52.895 44.435 ;
        RECT 57.415 44.305 58.345 44.525 ;
        RECT 61.175 44.305 62.095 44.535 ;
        RECT 63.685 44.305 66.685 44.535 ;
        RECT 67.190 44.305 68.535 44.535 ;
        RECT 52.905 43.625 62.095 44.305 ;
        RECT 62.105 44.215 66.685 44.305 ;
        RECT 62.105 43.855 66.695 44.215 ;
        RECT 62.105 43.625 63.675 43.855 ;
        RECT 65.765 43.665 66.695 43.855 ;
        RECT 65.765 43.625 66.685 43.665 ;
        RECT 66.705 43.625 68.535 44.305 ;
        RECT 68.545 43.625 69.915 44.435 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 70.385 43.625 75.895 44.435 ;
        RECT 75.905 43.625 78.655 44.435 ;
        RECT 78.665 43.625 80.035 44.405 ;
        RECT 80.515 43.625 81.865 44.535 ;
        RECT 81.885 43.625 87.395 44.435 ;
        RECT 87.405 43.625 89.235 44.435 ;
        RECT 89.245 43.625 90.615 44.405 ;
        RECT 90.625 44.305 91.555 44.535 ;
        RECT 90.625 43.625 94.525 44.305 ;
        RECT 95.695 43.710 96.125 44.495 ;
        RECT 96.145 43.625 101.655 44.435 ;
        RECT 106.635 44.305 107.565 44.525 ;
        RECT 110.395 44.305 111.315 44.535 ;
        RECT 102.125 43.625 111.315 44.305 ;
        RECT 111.325 43.625 116.835 44.435 ;
        RECT 116.845 43.625 120.515 44.435 ;
        RECT 121.455 43.710 121.885 44.495 ;
        RECT 122.365 43.625 123.735 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.625 ;
        RECT 8.885 43.575 9.055 43.605 ;
        RECT 8.880 43.465 9.055 43.575 ;
        RECT 8.885 43.415 9.055 43.465 ;
        RECT 9.345 43.435 9.515 43.625 ;
        RECT 19.005 43.415 19.175 43.605 ;
        RECT 19.280 43.435 19.450 43.625 ;
        RECT 19.465 43.415 19.635 43.605 ;
        RECT 23.145 43.435 23.315 43.625 ;
        RECT 24.985 43.415 25.155 43.605 ;
        RECT 26.640 43.415 26.810 43.605 ;
        RECT 29.120 43.435 29.290 43.625 ;
        RECT 29.585 43.435 29.755 43.625 ;
        RECT 30.515 43.460 30.675 43.570 ;
        RECT 31.885 43.415 32.055 43.605 ;
        RECT 35.105 43.435 35.275 43.625 ;
        RECT 35.575 43.460 35.735 43.570 ;
        RECT 36.760 43.415 36.930 43.605 ;
        RECT 40.635 43.460 40.795 43.570 ;
        RECT 41.820 43.415 41.990 43.605 ;
        RECT 45.685 43.415 45.855 43.625 ;
        RECT 46.145 43.435 46.315 43.625 ;
        RECT 49.820 43.435 49.990 43.625 ;
        RECT 50.285 43.435 50.455 43.625 ;
        RECT 51.205 43.415 51.375 43.605 ;
        RECT 53.045 43.435 53.215 43.625 ;
        RECT 56.720 43.465 56.840 43.575 ;
        RECT 57.655 43.460 57.815 43.570 ;
        RECT 59.485 43.415 59.655 43.605 ;
        RECT 59.945 43.415 60.115 43.605 ;
        RECT 61.325 43.415 61.495 43.605 ;
        RECT 62.245 43.435 62.415 43.625 ;
        RECT 65.005 43.415 65.175 43.605 ;
        RECT 66.845 43.415 67.015 43.625 ;
        RECT 68.685 43.435 68.855 43.625 ;
        RECT 70.525 43.435 70.695 43.625 ;
        RECT 72.365 43.415 72.535 43.605 ;
        RECT 73.745 43.415 73.915 43.605 ;
        RECT 76.045 43.435 76.215 43.625 ;
        RECT 79.725 43.435 79.895 43.625 ;
        RECT 80.180 43.465 80.300 43.575 ;
        RECT 81.565 43.435 81.735 43.625 ;
        RECT 82.025 43.435 82.195 43.625 ;
        RECT 83.415 43.460 83.575 43.570 ;
        RECT 84.600 43.415 84.770 43.605 ;
        RECT 87.545 43.435 87.715 43.625 ;
        RECT 88.465 43.415 88.635 43.605 ;
        RECT 89.385 43.435 89.555 43.625 ;
        RECT 90.300 43.465 90.420 43.575 ;
        RECT 90.765 43.415 90.935 43.605 ;
        RECT 91.040 43.435 91.210 43.625 ;
        RECT 94.915 43.470 95.075 43.580 ;
        RECT 96.285 43.435 96.455 43.625 ;
        RECT 99.965 43.415 100.135 43.605 ;
        RECT 101.800 43.465 101.920 43.575 ;
        RECT 102.265 43.435 102.435 43.625 ;
        RECT 103.655 43.460 103.815 43.570 ;
        RECT 107.970 43.415 108.140 43.605 ;
        RECT 109.165 43.415 109.335 43.605 ;
        RECT 111.465 43.435 111.635 43.625 ;
        RECT 116.985 43.435 117.155 43.625 ;
        RECT 118.365 43.415 118.535 43.605 ;
        RECT 120.675 43.470 120.835 43.580 ;
        RECT 122.040 43.465 122.160 43.575 ;
        RECT 123.425 43.415 123.595 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 8.735 43.415 ;
        RECT 8.745 42.735 17.935 43.415 ;
        RECT 13.255 42.515 14.185 42.735 ;
        RECT 17.015 42.505 17.935 42.735 ;
        RECT 17.955 42.505 19.305 43.415 ;
        RECT 19.325 42.605 24.835 43.415 ;
        RECT 24.845 42.635 26.215 43.415 ;
        RECT 26.225 42.735 30.125 43.415 ;
        RECT 26.225 42.505 27.155 42.735 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.745 42.605 35.415 43.415 ;
        RECT 36.345 42.735 40.245 43.415 ;
        RECT 41.405 42.735 45.305 43.415 ;
        RECT 36.345 42.505 37.275 42.735 ;
        RECT 41.405 42.505 42.335 42.735 ;
        RECT 45.545 42.605 51.055 43.415 ;
        RECT 51.065 42.605 56.575 43.415 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 58.435 42.505 59.785 43.415 ;
        RECT 59.805 42.605 61.175 43.415 ;
        RECT 61.185 42.735 64.855 43.415 ;
        RECT 64.865 42.735 66.695 43.415 ;
        RECT 63.925 42.505 64.855 42.735 ;
        RECT 66.705 42.605 72.215 43.415 ;
        RECT 72.225 42.605 73.595 43.415 ;
        RECT 73.605 42.735 82.795 43.415 ;
        RECT 78.115 42.515 79.045 42.735 ;
        RECT 81.875 42.505 82.795 42.735 ;
        RECT 82.815 42.545 83.245 43.330 ;
        RECT 84.185 42.735 88.085 43.415 ;
        RECT 84.185 42.505 85.115 42.735 ;
        RECT 88.325 42.605 90.155 43.415 ;
        RECT 90.625 42.735 99.815 43.415 ;
        RECT 95.135 42.515 96.065 42.735 ;
        RECT 98.895 42.505 99.815 42.735 ;
        RECT 99.825 42.605 103.495 43.415 ;
        RECT 104.655 42.735 108.555 43.415 ;
        RECT 107.625 42.505 108.555 42.735 ;
        RECT 108.575 42.545 109.005 43.330 ;
        RECT 109.025 42.735 118.215 43.415 ;
        RECT 113.535 42.515 114.465 42.735 ;
        RECT 117.295 42.505 118.215 42.735 ;
        RECT 118.225 42.605 121.895 43.415 ;
        RECT 122.365 42.605 123.735 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 123.930 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 6.905 38.185 12.415 38.995 ;
        RECT 12.425 38.185 17.935 38.995 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.185 24.375 38.995 ;
        RECT 29.815 38.865 30.745 39.085 ;
        RECT 33.575 38.865 34.495 39.095 ;
        RECT 25.305 38.185 34.495 38.865 ;
        RECT 34.515 38.185 35.865 39.095 ;
        RECT 35.885 38.185 39.555 38.995 ;
        RECT 39.565 38.185 40.935 38.965 ;
        RECT 40.945 38.185 43.695 38.995 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 44.625 38.185 50.135 38.995 ;
        RECT 50.145 38.185 51.515 38.995 ;
        RECT 56.035 38.865 56.965 39.085 ;
        RECT 59.795 38.865 60.715 39.095 ;
        RECT 51.525 38.185 60.715 38.865 ;
        RECT 60.725 38.185 66.235 38.995 ;
        RECT 66.245 38.185 69.915 38.995 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 70.385 38.185 75.895 38.995 ;
        RECT 75.905 38.185 79.575 38.995 ;
        RECT 79.585 38.185 80.955 38.995 ;
        RECT 85.475 38.865 86.405 39.085 ;
        RECT 89.235 38.865 90.155 39.095 ;
        RECT 80.965 38.185 90.155 38.865 ;
        RECT 90.165 38.185 95.675 38.995 ;
        RECT 95.695 38.270 96.125 39.055 ;
        RECT 96.155 38.185 97.505 39.095 ;
        RECT 97.525 38.185 101.195 38.995 ;
        RECT 106.635 38.865 107.565 39.085 ;
        RECT 110.395 38.865 111.315 39.095 ;
        RECT 102.125 38.185 111.315 38.865 ;
        RECT 111.335 38.185 112.685 39.095 ;
        RECT 112.705 38.185 118.215 38.995 ;
        RECT 118.225 38.185 120.975 38.995 ;
        RECT 121.455 38.270 121.885 39.055 ;
        RECT 122.365 38.185 123.735 38.995 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.975 7.215 38.185 ;
        RECT 12.565 37.975 12.735 38.185 ;
        RECT 18.085 38.135 18.255 38.165 ;
        RECT 18.080 38.025 18.255 38.135 ;
        RECT 18.085 37.975 18.255 38.025 ;
        RECT 19.005 37.995 19.175 38.185 ;
        RECT 23.605 37.975 23.775 38.165 ;
        RECT 24.535 38.030 24.695 38.140 ;
        RECT 25.445 37.995 25.615 38.185 ;
        RECT 29.125 37.975 29.295 38.165 ;
        RECT 30.960 38.025 31.080 38.135 ;
        RECT 31.885 37.975 32.055 38.165 ;
        RECT 35.565 37.995 35.735 38.185 ;
        RECT 36.025 37.995 36.195 38.185 ;
        RECT 37.400 38.025 37.520 38.135 ;
        RECT 37.865 37.975 38.035 38.165 ;
        RECT 40.625 37.995 40.795 38.185 ;
        RECT 41.085 37.995 41.255 38.185 ;
        RECT 43.840 38.025 43.960 38.135 ;
        RECT 44.765 37.995 44.935 38.185 ;
        RECT 47.340 37.975 47.510 38.165 ;
        RECT 50.285 37.995 50.455 38.185 ;
        RECT 51.205 37.975 51.375 38.165 ;
        RECT 51.665 37.995 51.835 38.185 ;
        RECT 54.895 38.020 55.055 38.130 ;
        RECT 55.805 37.975 55.975 38.165 ;
        RECT 58.565 37.975 58.735 38.165 ;
        RECT 59.025 37.975 59.195 38.165 ;
        RECT 60.865 37.995 61.035 38.185 ;
        RECT 64.545 37.995 64.715 38.165 ;
        RECT 64.545 37.975 64.710 37.995 ;
        RECT 65.005 37.975 65.175 38.165 ;
        RECT 66.385 37.995 66.555 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.165 12.415 37.975 ;
        RECT 12.425 37.165 17.935 37.975 ;
        RECT 17.945 37.165 23.455 37.975 ;
        RECT 23.465 37.165 28.975 37.975 ;
        RECT 28.985 37.165 30.815 37.975 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.745 37.165 37.255 37.975 ;
        RECT 37.725 37.295 46.915 37.975 ;
        RECT 42.235 37.075 43.165 37.295 ;
        RECT 45.995 37.065 46.915 37.295 ;
        RECT 46.925 37.295 50.825 37.975 ;
        RECT 46.925 37.065 47.855 37.295 ;
        RECT 51.065 37.165 54.735 37.975 ;
        RECT 55.675 37.065 57.025 37.975 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 57.505 37.195 58.875 37.975 ;
        RECT 58.885 37.165 62.555 37.975 ;
        RECT 62.875 37.295 64.710 37.975 ;
        RECT 62.875 37.065 63.805 37.295 ;
        RECT 64.865 37.165 66.695 37.975 ;
        RECT 66.705 37.945 67.650 37.975 ;
        RECT 69.605 37.945 69.775 38.165 ;
        RECT 70.070 37.975 70.240 38.165 ;
        RECT 70.525 37.995 70.695 38.185 ;
        RECT 73.285 37.975 73.455 38.165 ;
        RECT 76.045 37.995 76.215 38.185 ;
        RECT 78.805 37.975 78.975 38.165 ;
        RECT 79.725 37.995 79.895 38.185 ;
        RECT 81.105 37.995 81.275 38.185 ;
        RECT 82.480 38.025 82.600 38.135 ;
        RECT 84.325 37.975 84.495 38.165 ;
        RECT 84.785 37.975 84.955 38.165 ;
        RECT 86.165 37.975 86.335 38.165 ;
        RECT 90.305 37.995 90.475 38.185 ;
        RECT 91.685 37.975 91.855 38.165 ;
        RECT 97.205 38.135 97.375 38.185 ;
        RECT 97.200 38.025 97.375 38.135 ;
        RECT 97.205 37.995 97.375 38.025 ;
        RECT 97.665 37.975 97.835 38.185 ;
        RECT 99.045 37.975 99.215 38.165 ;
        RECT 101.355 38.030 101.515 38.140 ;
        RECT 101.800 38.025 101.920 38.135 ;
        RECT 102.265 37.975 102.435 38.185 ;
        RECT 103.920 37.975 104.090 38.165 ;
        RECT 107.795 38.020 107.955 38.130 ;
        RECT 110.085 37.975 110.255 38.165 ;
        RECT 110.545 37.975 110.715 38.165 ;
        RECT 111.465 37.995 111.635 38.185 ;
        RECT 112.845 37.995 113.015 38.185 ;
        RECT 116.065 37.975 116.235 38.165 ;
        RECT 118.365 37.995 118.535 38.185 ;
        RECT 121.120 38.025 121.240 38.135 ;
        RECT 121.595 38.020 121.755 38.130 ;
        RECT 122.040 38.025 122.160 38.135 ;
        RECT 123.425 37.975 123.595 38.185 ;
        RECT 66.705 37.745 69.775 37.945 ;
        RECT 66.705 37.265 69.915 37.745 ;
        RECT 66.705 37.065 67.650 37.265 ;
        RECT 68.985 37.065 69.915 37.265 ;
        RECT 69.925 37.065 72.845 37.975 ;
        RECT 73.145 37.165 78.655 37.975 ;
        RECT 78.665 37.165 82.335 37.975 ;
        RECT 82.815 37.105 83.245 37.890 ;
        RECT 83.265 37.195 84.635 37.975 ;
        RECT 84.655 37.065 86.005 37.975 ;
        RECT 86.025 37.165 91.535 37.975 ;
        RECT 91.545 37.165 97.055 37.975 ;
        RECT 97.535 37.065 98.885 37.975 ;
        RECT 98.905 37.165 101.655 37.975 ;
        RECT 102.125 37.195 103.495 37.975 ;
        RECT 103.505 37.295 107.405 37.975 ;
        RECT 103.505 37.065 104.435 37.295 ;
        RECT 108.575 37.105 109.005 37.890 ;
        RECT 109.035 37.065 110.385 37.975 ;
        RECT 110.405 37.165 115.915 37.975 ;
        RECT 115.925 37.165 121.435 37.975 ;
        RECT 122.365 37.165 123.735 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 123.930 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 12.415 33.555 ;
        RECT 12.425 32.745 15.175 33.555 ;
        RECT 15.185 32.745 16.555 33.525 ;
        RECT 16.565 32.745 18.395 33.555 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 18.865 33.425 19.795 33.655 ;
        RECT 23.005 33.425 23.935 33.655 ;
        RECT 18.865 32.745 22.765 33.425 ;
        RECT 23.005 32.745 26.905 33.425 ;
        RECT 27.145 32.745 32.655 33.555 ;
        RECT 32.665 32.745 38.175 33.555 ;
        RECT 38.185 32.745 40.935 33.555 ;
        RECT 40.945 32.745 42.315 33.525 ;
        RECT 42.335 32.745 43.685 33.655 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 44.635 32.745 45.985 33.655 ;
        RECT 46.005 32.745 51.515 33.555 ;
        RECT 51.525 32.745 57.035 33.555 ;
        RECT 57.045 32.745 58.875 33.555 ;
        RECT 59.365 32.745 60.715 33.655 ;
        RECT 60.725 33.425 61.645 33.655 ;
        RECT 60.725 32.745 63.015 33.425 ;
        RECT 63.025 32.745 65.315 33.655 ;
        RECT 65.325 33.455 66.255 33.655 ;
        RECT 67.590 33.455 68.535 33.655 ;
        RECT 65.325 32.975 68.535 33.455 ;
        RECT 65.465 32.775 68.535 32.975 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.535 7.215 32.745 ;
        RECT 8.880 32.585 9.000 32.695 ;
        RECT 9.345 32.535 9.515 32.725 ;
        RECT 12.565 32.555 12.735 32.745 ;
        RECT 16.245 32.555 16.415 32.745 ;
        RECT 16.705 32.555 16.875 32.745 ;
        RECT 18.545 32.535 18.715 32.725 ;
        RECT 19.280 32.555 19.450 32.745 ;
        RECT 23.420 32.555 23.590 32.745 ;
        RECT 27.285 32.555 27.455 32.745 ;
        RECT 27.740 32.585 27.860 32.695 ;
        RECT 29.125 32.535 29.295 32.725 ;
        RECT 29.585 32.535 29.755 32.725 ;
        RECT 32.160 32.535 32.330 32.725 ;
        RECT 32.805 32.555 32.975 32.745 ;
        RECT 36.025 32.535 36.195 32.725 ;
        RECT 38.325 32.555 38.495 32.745 ;
        RECT 38.785 32.535 38.955 32.725 ;
        RECT 42.005 32.555 42.175 32.745 ;
        RECT 42.465 32.555 42.635 32.745 ;
        RECT 43.840 32.585 43.960 32.695 ;
        RECT 45.685 32.555 45.855 32.745 ;
        RECT 46.145 32.555 46.315 32.745 ;
        RECT 48.445 32.535 48.615 32.725 ;
        RECT 51.665 32.555 51.835 32.745 ;
        RECT 53.965 32.535 54.135 32.725 ;
        RECT 56.720 32.585 56.840 32.695 ;
        RECT 57.185 32.555 57.355 32.745 ;
        RECT 59.020 32.585 59.140 32.695 ;
        RECT 59.480 32.555 59.650 32.745 ;
        RECT 60.405 32.535 60.575 32.725 ;
        RECT 62.245 32.535 62.415 32.725 ;
        RECT 62.705 32.535 62.875 32.745 ;
        RECT 63.170 32.555 63.340 32.745 ;
        RECT 65.465 32.695 65.635 32.775 ;
        RECT 67.590 32.745 68.535 32.775 ;
        RECT 68.545 32.745 69.915 33.555 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 70.385 33.425 71.305 33.655 ;
        RECT 70.385 32.745 72.675 33.425 ;
        RECT 72.685 32.745 78.195 33.555 ;
        RECT 78.205 32.745 83.715 33.555 ;
        RECT 83.725 32.745 89.235 33.555 ;
        RECT 90.165 33.425 91.095 33.655 ;
        RECT 90.165 32.745 94.065 33.425 ;
        RECT 94.305 32.745 95.675 33.525 ;
        RECT 95.695 32.830 96.125 33.615 ;
        RECT 97.505 33.425 98.425 33.645 ;
        RECT 104.505 33.545 105.425 33.655 ;
        RECT 103.090 33.425 105.425 33.545 ;
        RECT 96.145 32.745 105.425 33.425 ;
        RECT 105.805 32.745 111.315 33.555 ;
        RECT 111.325 32.745 116.835 33.555 ;
        RECT 116.845 32.745 120.515 33.555 ;
        RECT 121.455 32.830 121.885 33.615 ;
        RECT 122.365 32.745 123.735 33.555 ;
        RECT 65.460 32.585 65.635 32.695 ;
        RECT 65.465 32.555 65.635 32.585 ;
        RECT 65.925 32.535 66.095 32.725 ;
        RECT 67.305 32.535 67.475 32.725 ;
        RECT 68.685 32.555 68.855 32.745 ;
        RECT 72.365 32.555 72.535 32.745 ;
        RECT 72.825 32.555 72.995 32.745 ;
        RECT 77.885 32.535 78.055 32.725 ;
        RECT 78.345 32.555 78.515 32.745 ;
        RECT 80.645 32.535 80.815 32.725 ;
        RECT 81.100 32.585 81.220 32.695 ;
        RECT 81.565 32.535 81.735 32.725 ;
        RECT 83.680 32.535 83.850 32.725 ;
        RECT 83.865 32.555 84.035 32.745 ;
        RECT 87.545 32.535 87.715 32.725 ;
        RECT 88.925 32.535 89.095 32.725 ;
        RECT 89.395 32.590 89.555 32.700 ;
        RECT 90.305 32.535 90.475 32.725 ;
        RECT 90.580 32.555 90.750 32.745 ;
        RECT 93.995 32.580 94.155 32.690 ;
        RECT 94.445 32.555 94.615 32.745 ;
        RECT 95.180 32.535 95.350 32.725 ;
        RECT 96.285 32.555 96.455 32.745 ;
        RECT 99.045 32.535 99.215 32.725 ;
        RECT 104.565 32.535 104.735 32.725 ;
        RECT 105.945 32.555 106.115 32.745 ;
        RECT 108.240 32.585 108.360 32.695 ;
        RECT 109.165 32.535 109.335 32.725 ;
        RECT 111.465 32.555 111.635 32.745 ;
        RECT 114.685 32.535 114.855 32.725 ;
        RECT 116.985 32.555 117.155 32.745 ;
        RECT 120.205 32.535 120.375 32.725 ;
        RECT 120.675 32.590 120.835 32.700 ;
        RECT 122.040 32.585 122.160 32.695 ;
        RECT 123.425 32.535 123.595 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.725 8.735 32.535 ;
        RECT 9.205 31.855 18.395 32.535 ;
        RECT 18.405 31.855 27.595 32.535 ;
        RECT 13.715 31.635 14.645 31.855 ;
        RECT 17.475 31.625 18.395 31.855 ;
        RECT 22.915 31.635 23.845 31.855 ;
        RECT 26.675 31.625 27.595 31.855 ;
        RECT 28.065 31.755 29.435 32.535 ;
        RECT 29.445 31.725 31.275 32.535 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.745 31.855 35.645 32.535 ;
        RECT 31.745 31.625 32.675 31.855 ;
        RECT 35.885 31.725 38.635 32.535 ;
        RECT 38.645 31.855 47.925 32.535 ;
        RECT 40.005 31.635 40.925 31.855 ;
        RECT 45.590 31.735 47.925 31.855 ;
        RECT 47.005 31.625 47.925 31.735 ;
        RECT 48.305 31.725 53.815 32.535 ;
        RECT 53.825 31.725 56.575 32.535 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 57.505 31.625 60.615 32.535 ;
        RECT 60.725 31.855 62.555 32.535 ;
        RECT 60.725 31.625 62.070 31.855 ;
        RECT 62.565 31.725 65.315 32.535 ;
        RECT 65.785 31.755 67.155 32.535 ;
        RECT 67.165 31.855 77.535 32.535 ;
        RECT 71.675 31.635 72.605 31.855 ;
        RECT 75.325 31.625 77.535 31.855 ;
        RECT 77.745 31.725 79.575 32.535 ;
        RECT 79.585 31.755 80.955 32.535 ;
        RECT 81.435 31.625 82.785 32.535 ;
        RECT 82.815 31.665 83.245 32.450 ;
        RECT 83.265 31.855 87.165 32.535 ;
        RECT 83.265 31.625 84.195 31.855 ;
        RECT 87.415 31.625 88.765 32.535 ;
        RECT 88.785 31.755 90.155 32.535 ;
        RECT 90.165 31.725 93.835 32.535 ;
        RECT 94.765 31.855 98.665 32.535 ;
        RECT 94.765 31.625 95.695 31.855 ;
        RECT 98.905 31.725 104.415 32.535 ;
        RECT 104.425 31.725 108.095 32.535 ;
        RECT 108.575 31.665 109.005 32.450 ;
        RECT 109.025 31.725 114.535 32.535 ;
        RECT 114.545 31.725 120.055 32.535 ;
        RECT 120.065 31.725 121.895 32.535 ;
        RECT 122.365 31.725 123.735 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 123.930 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 12.415 28.115 ;
        RECT 12.425 27.305 16.095 28.115 ;
        RECT 16.575 27.305 17.925 28.215 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.865 27.305 20.695 28.115 ;
        RECT 21.165 27.305 22.535 28.085 ;
        RECT 23.475 27.305 24.825 28.215 ;
        RECT 29.815 27.985 30.745 28.205 ;
        RECT 33.575 27.985 34.495 28.215 ;
        RECT 25.305 27.305 34.495 27.985 ;
        RECT 34.515 27.305 35.865 28.215 ;
        RECT 35.885 27.305 39.555 28.115 ;
        RECT 40.485 27.305 41.855 28.085 ;
        RECT 42.795 27.305 44.145 28.215 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.625 27.985 45.555 28.215 ;
        RECT 44.625 27.305 48.525 27.985 ;
        RECT 48.765 27.305 51.515 28.115 ;
        RECT 56.035 27.985 56.965 28.205 ;
        RECT 59.795 27.985 60.715 28.215 ;
        RECT 51.525 27.305 60.715 27.985 ;
        RECT 60.725 27.305 66.235 28.115 ;
        RECT 66.245 27.305 69.915 28.115 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 70.855 27.305 72.205 28.215 ;
        RECT 72.225 27.305 75.895 28.115 ;
        RECT 81.335 27.985 82.265 28.205 ;
        RECT 85.095 27.985 86.015 28.215 ;
        RECT 76.825 27.305 86.015 27.985 ;
        RECT 86.025 27.985 86.945 28.215 ;
        RECT 89.775 27.985 90.705 28.205 ;
        RECT 86.025 27.305 95.215 27.985 ;
        RECT 95.695 27.390 96.125 28.175 ;
        RECT 96.145 27.305 101.655 28.115 ;
        RECT 101.665 27.305 107.175 28.115 ;
        RECT 107.185 27.305 112.695 28.115 ;
        RECT 112.705 27.305 118.215 28.115 ;
        RECT 118.225 27.305 120.975 28.115 ;
        RECT 121.455 27.390 121.885 28.175 ;
        RECT 122.365 27.305 123.735 28.115 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.095 7.215 27.305 ;
        RECT 12.565 27.095 12.735 27.305 ;
        RECT 16.240 27.145 16.360 27.255 ;
        RECT 17.625 27.115 17.795 27.305 ;
        RECT 18.085 27.255 18.255 27.285 ;
        RECT 18.080 27.145 18.255 27.255 ;
        RECT 18.085 27.095 18.255 27.145 ;
        RECT 19.005 27.115 19.175 27.305 ;
        RECT 20.840 27.145 20.960 27.255 ;
        RECT 22.225 27.115 22.395 27.305 ;
        RECT 22.695 27.150 22.855 27.260 ;
        RECT 23.605 27.095 23.775 27.305 ;
        RECT 24.980 27.145 25.100 27.255 ;
        RECT 25.445 27.115 25.615 27.305 ;
        RECT 29.125 27.095 29.295 27.285 ;
        RECT 30.960 27.145 31.080 27.255 ;
        RECT 31.885 27.095 32.055 27.285 ;
        RECT 35.565 27.115 35.735 27.305 ;
        RECT 36.025 27.115 36.195 27.305 ;
        RECT 37.415 27.140 37.575 27.250 ;
        RECT 38.325 27.095 38.495 27.285 ;
        RECT 39.715 27.150 39.875 27.260 ;
        RECT 41.545 27.115 41.715 27.305 ;
        RECT 42.015 27.150 42.175 27.260 ;
        RECT 42.925 27.115 43.095 27.305 ;
        RECT 45.040 27.115 45.210 27.305 ;
        RECT 47.985 27.095 48.155 27.285 ;
        RECT 48.905 27.115 49.075 27.305 ;
        RECT 51.665 27.115 51.835 27.305 ;
        RECT 53.505 27.095 53.675 27.285 ;
        RECT 55.340 27.145 55.460 27.255 ;
        RECT 55.805 27.095 55.975 27.285 ;
        RECT 57.645 27.095 57.815 27.285 ;
        RECT 60.865 27.115 61.035 27.305 ;
        RECT 63.165 27.095 63.335 27.285 ;
        RECT 66.385 27.115 66.555 27.305 ;
        RECT 70.520 27.145 70.640 27.255 ;
        RECT 70.985 27.115 71.155 27.305 ;
        RECT 72.365 27.115 72.535 27.305 ;
        RECT 75.585 27.095 75.755 27.285 ;
        RECT 76.045 27.095 76.215 27.285 ;
        RECT 76.965 27.115 77.135 27.305 ;
        RECT 81.565 27.095 81.735 27.285 ;
        RECT 83.405 27.095 83.575 27.285 ;
        RECT 88.925 27.095 89.095 27.285 ;
        RECT 94.445 27.095 94.615 27.285 ;
        RECT 94.905 27.115 95.075 27.305 ;
        RECT 95.360 27.145 95.480 27.255 ;
        RECT 96.285 27.115 96.455 27.305 ;
        RECT 99.965 27.095 100.135 27.285 ;
        RECT 101.805 27.115 101.975 27.305 ;
        RECT 105.485 27.095 105.655 27.285 ;
        RECT 107.325 27.115 107.495 27.305 ;
        RECT 108.240 27.145 108.360 27.255 ;
        RECT 109.165 27.095 109.335 27.285 ;
        RECT 112.845 27.115 113.015 27.305 ;
        RECT 114.685 27.095 114.855 27.285 ;
        RECT 118.365 27.115 118.535 27.305 ;
        RECT 120.205 27.095 120.375 27.285 ;
        RECT 121.120 27.145 121.240 27.255 ;
        RECT 122.040 27.145 122.160 27.255 ;
        RECT 123.425 27.095 123.595 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 6.905 26.285 12.415 27.095 ;
        RECT 12.425 26.285 17.935 27.095 ;
        RECT 17.945 26.285 23.455 27.095 ;
        RECT 23.465 26.285 28.975 27.095 ;
        RECT 28.985 26.285 30.815 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.745 26.285 37.255 27.095 ;
        RECT 38.185 26.415 47.465 27.095 ;
        RECT 39.545 26.195 40.465 26.415 ;
        RECT 45.130 26.295 47.465 26.415 ;
        RECT 46.545 26.185 47.465 26.295 ;
        RECT 47.845 26.285 53.355 27.095 ;
        RECT 53.365 26.285 55.195 27.095 ;
        RECT 55.675 26.185 57.025 27.095 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 57.505 26.285 63.015 27.095 ;
        RECT 63.125 26.185 66.235 27.095 ;
        RECT 66.285 26.415 75.895 27.095 ;
        RECT 66.285 26.185 67.625 26.415 ;
        RECT 70.455 26.195 71.385 26.415 ;
        RECT 75.905 26.285 81.415 27.095 ;
        RECT 81.425 26.285 82.795 27.095 ;
        RECT 82.815 26.225 83.245 27.010 ;
        RECT 83.265 26.285 88.775 27.095 ;
        RECT 88.785 26.285 94.295 27.095 ;
        RECT 94.305 26.285 99.815 27.095 ;
        RECT 99.825 26.285 105.335 27.095 ;
        RECT 105.345 26.285 108.095 27.095 ;
        RECT 108.575 26.225 109.005 27.010 ;
        RECT 109.025 26.285 114.535 27.095 ;
        RECT 114.545 26.285 120.055 27.095 ;
        RECT 120.065 26.285 121.895 27.095 ;
        RECT 122.365 26.285 123.735 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 123.930 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 21.865 12.415 22.675 ;
        RECT 12.425 21.865 17.935 22.675 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 18.865 21.865 24.375 22.675 ;
        RECT 24.385 21.865 29.895 22.675 ;
        RECT 29.905 21.865 35.415 22.675 ;
        RECT 35.425 21.865 40.935 22.675 ;
        RECT 40.945 21.865 43.695 22.675 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 50.135 22.675 ;
        RECT 50.145 21.865 55.655 22.675 ;
        RECT 55.665 21.865 61.175 22.675 ;
        RECT 61.185 21.865 66.695 22.675 ;
        RECT 66.705 21.865 69.455 22.675 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.395 21.865 71.745 22.775 ;
        RECT 71.765 21.865 77.275 22.675 ;
        RECT 77.285 21.865 82.795 22.675 ;
        RECT 82.805 21.865 88.315 22.675 ;
        RECT 88.325 21.865 93.835 22.675 ;
        RECT 93.845 21.865 95.675 22.675 ;
        RECT 95.695 21.950 96.125 22.735 ;
        RECT 96.145 21.865 101.655 22.675 ;
        RECT 101.665 21.865 107.175 22.675 ;
        RECT 107.185 21.865 112.695 22.675 ;
        RECT 112.705 21.865 118.215 22.675 ;
        RECT 118.225 21.865 120.975 22.675 ;
        RECT 121.455 21.950 121.885 22.735 ;
        RECT 122.365 21.865 123.735 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.655 7.215 21.865 ;
        RECT 12.565 21.655 12.735 21.865 ;
        RECT 18.085 21.815 18.255 21.845 ;
        RECT 18.080 21.705 18.255 21.815 ;
        RECT 18.085 21.655 18.255 21.705 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 23.605 21.655 23.775 21.845 ;
        RECT 24.525 21.675 24.695 21.865 ;
        RECT 29.125 21.655 29.295 21.845 ;
        RECT 30.045 21.675 30.215 21.865 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 35.565 21.675 35.735 21.865 ;
        RECT 37.405 21.655 37.575 21.845 ;
        RECT 41.085 21.675 41.255 21.865 ;
        RECT 42.925 21.655 43.095 21.845 ;
        RECT 43.840 21.705 43.960 21.815 ;
        RECT 44.765 21.675 44.935 21.865 ;
        RECT 48.445 21.655 48.615 21.845 ;
        RECT 50.285 21.675 50.455 21.865 ;
        RECT 53.965 21.655 54.135 21.845 ;
        RECT 55.805 21.675 55.975 21.865 ;
        RECT 56.720 21.705 56.840 21.815 ;
        RECT 57.645 21.655 57.815 21.845 ;
        RECT 61.325 21.675 61.495 21.865 ;
        RECT 63.165 21.655 63.335 21.845 ;
        RECT 66.845 21.675 67.015 21.865 ;
        RECT 68.685 21.655 68.855 21.845 ;
        RECT 69.600 21.705 69.720 21.815 ;
        RECT 70.525 21.675 70.695 21.865 ;
        RECT 71.905 21.675 72.075 21.865 ;
        RECT 74.205 21.655 74.375 21.845 ;
        RECT 77.425 21.675 77.595 21.865 ;
        RECT 79.725 21.655 79.895 21.845 ;
        RECT 82.480 21.705 82.600 21.815 ;
        RECT 82.945 21.675 83.115 21.865 ;
        RECT 83.405 21.655 83.575 21.845 ;
        RECT 88.465 21.675 88.635 21.865 ;
        RECT 88.925 21.655 89.095 21.845 ;
        RECT 93.985 21.675 94.155 21.865 ;
        RECT 94.445 21.655 94.615 21.845 ;
        RECT 96.285 21.675 96.455 21.865 ;
        RECT 99.965 21.655 100.135 21.845 ;
        RECT 101.805 21.675 101.975 21.865 ;
        RECT 105.485 21.655 105.655 21.845 ;
        RECT 107.325 21.675 107.495 21.865 ;
        RECT 108.240 21.705 108.360 21.815 ;
        RECT 109.165 21.655 109.335 21.845 ;
        RECT 112.845 21.675 113.015 21.865 ;
        RECT 114.685 21.655 114.855 21.845 ;
        RECT 118.365 21.675 118.535 21.865 ;
        RECT 120.205 21.655 120.375 21.845 ;
        RECT 121.120 21.705 121.240 21.815 ;
        RECT 122.040 21.705 122.160 21.815 ;
        RECT 123.425 21.655 123.595 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.845 12.415 21.655 ;
        RECT 12.425 20.845 17.935 21.655 ;
        RECT 17.945 20.845 23.455 21.655 ;
        RECT 23.465 20.845 28.975 21.655 ;
        RECT 28.985 20.845 30.815 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.265 20.845 42.775 21.655 ;
        RECT 42.785 20.845 48.295 21.655 ;
        RECT 48.305 20.845 53.815 21.655 ;
        RECT 53.825 20.845 56.575 21.655 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.505 20.845 63.015 21.655 ;
        RECT 63.025 20.845 68.535 21.655 ;
        RECT 68.545 20.845 74.055 21.655 ;
        RECT 74.065 20.845 79.575 21.655 ;
        RECT 79.585 20.845 82.335 21.655 ;
        RECT 82.815 20.785 83.245 21.570 ;
        RECT 83.265 20.845 88.775 21.655 ;
        RECT 88.785 20.845 94.295 21.655 ;
        RECT 94.305 20.845 99.815 21.655 ;
        RECT 99.825 20.845 105.335 21.655 ;
        RECT 105.345 20.845 108.095 21.655 ;
        RECT 108.575 20.785 109.005 21.570 ;
        RECT 109.025 20.845 114.535 21.655 ;
        RECT 114.545 20.845 120.055 21.655 ;
        RECT 120.065 20.845 121.895 21.655 ;
        RECT 122.365 20.845 123.735 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 123.930 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 12.415 17.235 ;
        RECT 12.425 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 24.375 17.235 ;
        RECT 24.385 16.425 29.895 17.235 ;
        RECT 29.905 16.425 35.415 17.235 ;
        RECT 35.425 16.425 40.935 17.235 ;
        RECT 40.945 16.425 43.695 17.235 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 44.625 16.425 50.135 17.235 ;
        RECT 50.145 16.425 55.655 17.235 ;
        RECT 55.665 16.425 61.175 17.235 ;
        RECT 61.185 16.425 66.695 17.235 ;
        RECT 66.705 16.425 69.455 17.235 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 70.385 16.425 75.895 17.235 ;
        RECT 75.905 16.425 81.415 17.235 ;
        RECT 81.425 16.425 86.935 17.235 ;
        RECT 86.945 16.425 92.455 17.235 ;
        RECT 92.465 16.425 95.215 17.235 ;
        RECT 95.695 16.510 96.125 17.295 ;
        RECT 96.145 16.425 101.655 17.235 ;
        RECT 101.665 16.425 107.175 17.235 ;
        RECT 107.185 16.425 112.695 17.235 ;
        RECT 112.705 16.425 118.215 17.235 ;
        RECT 118.225 16.425 120.975 17.235 ;
        RECT 121.455 16.510 121.885 17.295 ;
        RECT 122.365 16.425 123.735 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 12.565 16.215 12.735 16.425 ;
        RECT 18.085 16.375 18.255 16.405 ;
        RECT 18.080 16.265 18.255 16.375 ;
        RECT 18.085 16.215 18.255 16.265 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.605 16.215 23.775 16.405 ;
        RECT 24.525 16.235 24.695 16.425 ;
        RECT 29.125 16.215 29.295 16.405 ;
        RECT 30.045 16.235 30.215 16.425 ;
        RECT 30.960 16.265 31.080 16.375 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 35.565 16.235 35.735 16.425 ;
        RECT 37.405 16.215 37.575 16.405 ;
        RECT 41.085 16.235 41.255 16.425 ;
        RECT 42.925 16.215 43.095 16.405 ;
        RECT 43.840 16.265 43.960 16.375 ;
        RECT 44.765 16.235 44.935 16.425 ;
        RECT 48.445 16.215 48.615 16.405 ;
        RECT 50.285 16.235 50.455 16.425 ;
        RECT 53.965 16.215 54.135 16.405 ;
        RECT 55.805 16.235 55.975 16.425 ;
        RECT 56.720 16.265 56.840 16.375 ;
        RECT 57.645 16.215 57.815 16.405 ;
        RECT 61.325 16.235 61.495 16.425 ;
        RECT 63.165 16.215 63.335 16.405 ;
        RECT 66.845 16.235 67.015 16.425 ;
        RECT 68.685 16.215 68.855 16.405 ;
        RECT 69.600 16.265 69.720 16.375 ;
        RECT 70.525 16.235 70.695 16.425 ;
        RECT 74.205 16.215 74.375 16.405 ;
        RECT 76.045 16.235 76.215 16.425 ;
        RECT 79.725 16.215 79.895 16.405 ;
        RECT 81.565 16.235 81.735 16.425 ;
        RECT 82.480 16.265 82.600 16.375 ;
        RECT 83.405 16.215 83.575 16.405 ;
        RECT 87.085 16.235 87.255 16.425 ;
        RECT 88.925 16.215 89.095 16.405 ;
        RECT 92.605 16.235 92.775 16.425 ;
        RECT 94.445 16.215 94.615 16.405 ;
        RECT 95.360 16.265 95.480 16.375 ;
        RECT 96.285 16.235 96.455 16.425 ;
        RECT 99.965 16.215 100.135 16.405 ;
        RECT 101.805 16.235 101.975 16.425 ;
        RECT 105.485 16.215 105.655 16.405 ;
        RECT 107.325 16.235 107.495 16.425 ;
        RECT 108.240 16.265 108.360 16.375 ;
        RECT 109.165 16.215 109.335 16.405 ;
        RECT 112.845 16.235 113.015 16.425 ;
        RECT 114.685 16.215 114.855 16.405 ;
        RECT 118.365 16.235 118.535 16.425 ;
        RECT 120.205 16.215 120.375 16.405 ;
        RECT 121.120 16.265 121.240 16.375 ;
        RECT 122.040 16.265 122.160 16.375 ;
        RECT 123.425 16.215 123.595 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 23.455 16.215 ;
        RECT 23.465 15.405 28.975 16.215 ;
        RECT 28.985 15.405 30.815 16.215 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.745 15.405 37.255 16.215 ;
        RECT 37.265 15.405 42.775 16.215 ;
        RECT 42.785 15.405 48.295 16.215 ;
        RECT 48.305 15.405 53.815 16.215 ;
        RECT 53.825 15.405 56.575 16.215 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.405 63.015 16.215 ;
        RECT 63.025 15.405 68.535 16.215 ;
        RECT 68.545 15.405 74.055 16.215 ;
        RECT 74.065 15.405 79.575 16.215 ;
        RECT 79.585 15.405 82.335 16.215 ;
        RECT 82.815 15.345 83.245 16.130 ;
        RECT 83.265 15.405 88.775 16.215 ;
        RECT 88.785 15.405 94.295 16.215 ;
        RECT 94.305 15.405 99.815 16.215 ;
        RECT 99.825 15.405 105.335 16.215 ;
        RECT 105.345 15.405 108.095 16.215 ;
        RECT 108.575 15.345 109.005 16.130 ;
        RECT 109.025 15.405 114.535 16.215 ;
        RECT 114.545 15.405 120.055 16.215 ;
        RECT 120.065 15.405 121.895 16.215 ;
        RECT 122.365 15.405 123.735 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 123.930 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 12.425 10.985 17.935 11.795 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 18.865 10.985 24.375 11.795 ;
        RECT 24.385 10.985 29.895 11.795 ;
        RECT 29.905 10.985 31.275 11.795 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 31.745 10.985 37.255 11.795 ;
        RECT 37.265 10.985 42.775 11.795 ;
        RECT 42.785 10.985 44.155 11.795 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 44.625 10.985 50.135 11.795 ;
        RECT 50.145 10.985 55.655 11.795 ;
        RECT 55.665 10.985 57.035 11.795 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 57.505 10.985 63.015 11.795 ;
        RECT 63.025 10.985 68.535 11.795 ;
        RECT 68.545 10.985 69.915 11.795 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 70.385 10.985 75.895 11.795 ;
        RECT 75.905 10.985 81.415 11.795 ;
        RECT 81.425 10.985 82.795 11.795 ;
        RECT 82.815 11.070 83.245 11.855 ;
        RECT 83.265 10.985 88.775 11.795 ;
        RECT 88.785 10.985 94.295 11.795 ;
        RECT 94.305 10.985 95.675 11.795 ;
        RECT 95.695 11.070 96.125 11.855 ;
        RECT 96.145 10.985 101.655 11.795 ;
        RECT 101.665 10.985 107.175 11.795 ;
        RECT 107.185 10.985 108.555 11.795 ;
        RECT 108.575 11.070 109.005 11.855 ;
        RECT 109.025 10.985 114.535 11.795 ;
        RECT 114.545 10.985 120.055 11.795 ;
        RECT 120.065 10.985 121.435 11.795 ;
        RECT 121.455 11.070 121.885 11.855 ;
        RECT 122.365 10.985 123.735 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.565 10.795 12.735 10.985 ;
        RECT 18.080 10.825 18.200 10.935 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 31.885 10.795 32.055 10.985 ;
        RECT 37.405 10.795 37.575 10.985 ;
        RECT 42.925 10.795 43.095 10.985 ;
        RECT 44.765 10.795 44.935 10.985 ;
        RECT 50.285 10.795 50.455 10.985 ;
        RECT 55.805 10.795 55.975 10.985 ;
        RECT 57.645 10.795 57.815 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 68.685 10.795 68.855 10.985 ;
        RECT 70.525 10.795 70.695 10.985 ;
        RECT 76.045 10.795 76.215 10.985 ;
        RECT 81.565 10.795 81.735 10.985 ;
        RECT 83.405 10.795 83.575 10.985 ;
        RECT 88.925 10.795 89.095 10.985 ;
        RECT 94.445 10.795 94.615 10.985 ;
        RECT 96.285 10.795 96.455 10.985 ;
        RECT 101.805 10.795 101.975 10.985 ;
        RECT 107.325 10.795 107.495 10.985 ;
        RECT 109.165 10.795 109.335 10.985 ;
        RECT 114.685 10.795 114.855 10.985 ;
        RECT 120.205 10.795 120.375 10.985 ;
        RECT 122.040 10.825 122.160 10.935 ;
        RECT 123.425 10.795 123.595 10.985 ;
      LAYER li1 ;
        RECT 5.520 127.755 123.740 127.925 ;
        RECT 5.605 126.665 6.815 127.755 ;
        RECT 6.985 127.320 12.330 127.755 ;
        RECT 12.505 127.320 17.850 127.755 ;
        RECT 5.605 125.955 6.125 126.495 ;
        RECT 6.295 126.125 6.815 126.665 ;
        RECT 5.605 125.205 6.815 125.955 ;
        RECT 8.570 125.750 8.910 126.580 ;
        RECT 10.390 126.070 10.740 127.320 ;
        RECT 14.090 125.750 14.430 126.580 ;
        RECT 15.910 126.070 16.260 127.320 ;
        RECT 18.485 126.590 18.775 127.755 ;
        RECT 18.945 127.320 24.290 127.755 ;
        RECT 24.465 127.320 29.810 127.755 ;
        RECT 6.985 125.205 12.330 125.750 ;
        RECT 12.505 125.205 17.850 125.750 ;
        RECT 18.485 125.205 18.775 125.930 ;
        RECT 20.530 125.750 20.870 126.580 ;
        RECT 22.350 126.070 22.700 127.320 ;
        RECT 26.050 125.750 26.390 126.580 ;
        RECT 27.870 126.070 28.220 127.320 ;
        RECT 29.985 126.665 31.195 127.755 ;
        RECT 29.985 125.955 30.505 126.495 ;
        RECT 30.675 126.125 31.195 126.665 ;
        RECT 31.365 126.590 31.655 127.755 ;
        RECT 31.825 127.320 37.170 127.755 ;
        RECT 37.345 127.320 42.690 127.755 ;
        RECT 18.945 125.205 24.290 125.750 ;
        RECT 24.465 125.205 29.810 125.750 ;
        RECT 29.985 125.205 31.195 125.955 ;
        RECT 31.365 125.205 31.655 125.930 ;
        RECT 33.410 125.750 33.750 126.580 ;
        RECT 35.230 126.070 35.580 127.320 ;
        RECT 38.930 125.750 39.270 126.580 ;
        RECT 40.750 126.070 41.100 127.320 ;
        RECT 42.865 126.665 44.075 127.755 ;
        RECT 42.865 125.955 43.385 126.495 ;
        RECT 43.555 126.125 44.075 126.665 ;
        RECT 44.245 126.590 44.535 127.755 ;
        RECT 44.705 127.320 50.050 127.755 ;
        RECT 50.225 127.320 55.570 127.755 ;
        RECT 31.825 125.205 37.170 125.750 ;
        RECT 37.345 125.205 42.690 125.750 ;
        RECT 42.865 125.205 44.075 125.955 ;
        RECT 44.245 125.205 44.535 125.930 ;
        RECT 46.290 125.750 46.630 126.580 ;
        RECT 48.110 126.070 48.460 127.320 ;
        RECT 51.810 125.750 52.150 126.580 ;
        RECT 53.630 126.070 53.980 127.320 ;
        RECT 55.745 126.665 56.955 127.755 ;
        RECT 55.745 125.955 56.265 126.495 ;
        RECT 56.435 126.125 56.955 126.665 ;
        RECT 57.125 126.590 57.415 127.755 ;
        RECT 57.585 127.320 62.930 127.755 ;
        RECT 63.105 127.320 68.450 127.755 ;
        RECT 44.705 125.205 50.050 125.750 ;
        RECT 50.225 125.205 55.570 125.750 ;
        RECT 55.745 125.205 56.955 125.955 ;
        RECT 57.125 125.205 57.415 125.930 ;
        RECT 59.170 125.750 59.510 126.580 ;
        RECT 60.990 126.070 61.340 127.320 ;
        RECT 64.690 125.750 65.030 126.580 ;
        RECT 66.510 126.070 66.860 127.320 ;
        RECT 68.625 126.665 69.835 127.755 ;
        RECT 68.625 125.955 69.145 126.495 ;
        RECT 69.315 126.125 69.835 126.665 ;
        RECT 70.005 126.590 70.295 127.755 ;
        RECT 70.465 127.320 75.810 127.755 ;
        RECT 75.985 127.320 81.330 127.755 ;
        RECT 57.585 125.205 62.930 125.750 ;
        RECT 63.105 125.205 68.450 125.750 ;
        RECT 68.625 125.205 69.835 125.955 ;
        RECT 70.005 125.205 70.295 125.930 ;
        RECT 72.050 125.750 72.390 126.580 ;
        RECT 73.870 126.070 74.220 127.320 ;
        RECT 77.570 125.750 77.910 126.580 ;
        RECT 79.390 126.070 79.740 127.320 ;
        RECT 81.505 126.665 82.715 127.755 ;
        RECT 81.505 125.955 82.025 126.495 ;
        RECT 82.195 126.125 82.715 126.665 ;
        RECT 82.885 126.590 83.175 127.755 ;
        RECT 83.345 127.320 88.690 127.755 ;
        RECT 88.865 127.320 94.210 127.755 ;
        RECT 70.465 125.205 75.810 125.750 ;
        RECT 75.985 125.205 81.330 125.750 ;
        RECT 81.505 125.205 82.715 125.955 ;
        RECT 82.885 125.205 83.175 125.930 ;
        RECT 84.930 125.750 85.270 126.580 ;
        RECT 86.750 126.070 87.100 127.320 ;
        RECT 90.450 125.750 90.790 126.580 ;
        RECT 92.270 126.070 92.620 127.320 ;
        RECT 94.385 126.665 95.595 127.755 ;
        RECT 94.385 125.955 94.905 126.495 ;
        RECT 95.075 126.125 95.595 126.665 ;
        RECT 95.765 126.590 96.055 127.755 ;
        RECT 96.225 127.320 101.570 127.755 ;
        RECT 101.745 127.320 107.090 127.755 ;
        RECT 83.345 125.205 88.690 125.750 ;
        RECT 88.865 125.205 94.210 125.750 ;
        RECT 94.385 125.205 95.595 125.955 ;
        RECT 95.765 125.205 96.055 125.930 ;
        RECT 97.810 125.750 98.150 126.580 ;
        RECT 99.630 126.070 99.980 127.320 ;
        RECT 103.330 125.750 103.670 126.580 ;
        RECT 105.150 126.070 105.500 127.320 ;
        RECT 107.265 126.665 108.475 127.755 ;
        RECT 107.265 125.955 107.785 126.495 ;
        RECT 107.955 126.125 108.475 126.665 ;
        RECT 108.645 126.590 108.935 127.755 ;
        RECT 109.105 126.665 111.695 127.755 ;
        RECT 112.330 127.085 112.585 127.585 ;
        RECT 112.755 127.255 113.085 127.755 ;
        RECT 112.330 126.915 113.080 127.085 ;
        RECT 109.105 125.975 110.315 126.495 ;
        RECT 110.485 126.145 111.695 126.665 ;
        RECT 112.330 126.095 112.680 126.745 ;
        RECT 96.225 125.205 101.570 125.750 ;
        RECT 101.745 125.205 107.090 125.750 ;
        RECT 107.265 125.205 108.475 125.955 ;
        RECT 108.645 125.205 108.935 125.930 ;
        RECT 109.105 125.205 111.695 125.975 ;
        RECT 112.850 125.925 113.080 126.915 ;
        RECT 112.330 125.755 113.080 125.925 ;
        RECT 112.330 125.465 112.585 125.755 ;
        RECT 112.755 125.205 113.085 125.585 ;
        RECT 113.255 125.465 113.425 127.585 ;
        RECT 113.595 126.785 113.920 127.570 ;
        RECT 114.090 127.295 114.340 127.755 ;
        RECT 114.510 127.255 114.760 127.585 ;
        RECT 114.975 127.255 115.655 127.585 ;
        RECT 114.510 127.125 114.680 127.255 ;
        RECT 114.285 126.955 114.680 127.125 ;
        RECT 113.655 125.735 114.115 126.785 ;
        RECT 114.285 125.595 114.455 126.955 ;
        RECT 114.850 126.695 115.315 127.085 ;
        RECT 114.625 125.885 114.975 126.505 ;
        RECT 115.145 126.105 115.315 126.695 ;
        RECT 115.485 126.475 115.655 127.255 ;
        RECT 115.825 127.155 115.995 127.495 ;
        RECT 116.230 127.325 116.560 127.755 ;
        RECT 116.730 127.155 116.900 127.495 ;
        RECT 117.195 127.295 117.565 127.755 ;
        RECT 115.825 126.985 116.900 127.155 ;
        RECT 117.735 127.125 117.905 127.585 ;
        RECT 118.140 127.245 119.010 127.585 ;
        RECT 119.180 127.295 119.430 127.755 ;
        RECT 117.345 126.955 117.905 127.125 ;
        RECT 117.345 126.815 117.515 126.955 ;
        RECT 116.015 126.645 117.515 126.815 ;
        RECT 118.210 126.785 118.670 127.075 ;
        RECT 115.485 126.305 117.175 126.475 ;
        RECT 115.145 125.885 115.500 126.105 ;
        RECT 115.670 125.595 115.840 126.305 ;
        RECT 116.045 125.885 116.835 126.135 ;
        RECT 117.005 126.125 117.175 126.305 ;
        RECT 117.345 125.955 117.515 126.645 ;
        RECT 113.785 125.205 114.115 125.565 ;
        RECT 114.285 125.425 114.780 125.595 ;
        RECT 114.985 125.425 115.840 125.595 ;
        RECT 116.715 125.205 117.045 125.665 ;
        RECT 117.255 125.565 117.515 125.955 ;
        RECT 117.705 126.775 118.670 126.785 ;
        RECT 118.840 126.865 119.010 127.245 ;
        RECT 119.600 127.205 119.770 127.495 ;
        RECT 119.950 127.375 120.280 127.755 ;
        RECT 119.600 127.035 120.400 127.205 ;
        RECT 117.705 126.615 118.380 126.775 ;
        RECT 118.840 126.695 120.060 126.865 ;
        RECT 117.705 125.825 117.915 126.615 ;
        RECT 118.840 126.605 119.010 126.695 ;
        RECT 118.085 125.825 118.435 126.445 ;
        RECT 118.605 126.435 119.010 126.605 ;
        RECT 118.605 125.655 118.775 126.435 ;
        RECT 118.945 125.985 119.165 126.265 ;
        RECT 119.345 126.155 119.885 126.525 ;
        RECT 120.230 126.445 120.400 127.035 ;
        RECT 120.620 126.615 120.925 127.755 ;
        RECT 121.095 126.565 121.350 127.445 ;
        RECT 121.525 126.590 121.815 127.755 ;
        RECT 122.445 126.665 123.655 127.755 ;
        RECT 120.230 126.415 120.970 126.445 ;
        RECT 118.945 125.815 119.475 125.985 ;
        RECT 117.255 125.395 117.605 125.565 ;
        RECT 117.825 125.375 118.775 125.655 ;
        RECT 118.945 125.205 119.135 125.645 ;
        RECT 119.305 125.585 119.475 125.815 ;
        RECT 119.645 125.755 119.885 126.155 ;
        RECT 120.055 126.115 120.970 126.415 ;
        RECT 120.055 125.940 120.380 126.115 ;
        RECT 120.055 125.585 120.375 125.940 ;
        RECT 121.140 125.915 121.350 126.565 ;
        RECT 122.445 126.125 122.965 126.665 ;
        RECT 123.135 125.955 123.655 126.495 ;
        RECT 119.305 125.415 120.375 125.585 ;
        RECT 120.620 125.205 120.925 125.665 ;
        RECT 121.095 125.385 121.350 125.915 ;
        RECT 121.525 125.205 121.815 125.930 ;
        RECT 122.445 125.205 123.655 125.955 ;
        RECT 5.520 125.035 123.740 125.205 ;
        RECT 5.605 124.285 6.815 125.035 ;
        RECT 7.075 124.485 7.245 124.865 ;
        RECT 7.425 124.655 7.755 125.035 ;
        RECT 7.075 124.315 7.740 124.485 ;
        RECT 7.935 124.360 8.195 124.865 ;
        RECT 5.605 123.745 6.125 124.285 ;
        RECT 6.295 123.575 6.815 124.115 ;
        RECT 7.005 123.765 7.345 124.135 ;
        RECT 7.570 124.060 7.740 124.315 ;
        RECT 7.570 123.730 7.845 124.060 ;
        RECT 7.570 123.585 7.740 123.730 ;
        RECT 5.605 122.485 6.815 123.575 ;
        RECT 7.065 123.415 7.740 123.585 ;
        RECT 8.015 123.560 8.195 124.360 ;
        RECT 8.365 124.265 11.875 125.035 ;
        RECT 12.510 124.325 12.765 124.855 ;
        RECT 12.935 124.575 13.240 125.035 ;
        RECT 13.485 124.655 14.555 124.825 ;
        RECT 8.365 123.745 10.015 124.265 ;
        RECT 10.185 123.575 11.875 124.095 ;
        RECT 7.065 122.655 7.245 123.415 ;
        RECT 7.425 122.485 7.755 123.245 ;
        RECT 7.925 122.655 8.195 123.560 ;
        RECT 8.365 122.485 11.875 123.575 ;
        RECT 12.510 123.675 12.720 124.325 ;
        RECT 13.485 124.300 13.805 124.655 ;
        RECT 13.480 124.125 13.805 124.300 ;
        RECT 12.890 123.825 13.805 124.125 ;
        RECT 13.975 124.085 14.215 124.485 ;
        RECT 14.385 124.425 14.555 124.655 ;
        RECT 14.725 124.595 14.915 125.035 ;
        RECT 15.085 124.585 16.035 124.865 ;
        RECT 16.255 124.675 16.605 124.845 ;
        RECT 14.385 124.255 14.915 124.425 ;
        RECT 12.890 123.795 13.630 123.825 ;
        RECT 12.510 122.795 12.765 123.675 ;
        RECT 12.935 122.485 13.240 123.625 ;
        RECT 13.460 123.205 13.630 123.795 ;
        RECT 13.975 123.715 14.515 124.085 ;
        RECT 14.695 123.975 14.915 124.255 ;
        RECT 15.085 123.805 15.255 124.585 ;
        RECT 14.850 123.635 15.255 123.805 ;
        RECT 15.425 123.795 15.775 124.415 ;
        RECT 14.850 123.545 15.020 123.635 ;
        RECT 15.945 123.625 16.155 124.415 ;
        RECT 13.800 123.375 15.020 123.545 ;
        RECT 15.480 123.465 16.155 123.625 ;
        RECT 13.460 123.035 14.260 123.205 ;
        RECT 13.580 122.485 13.910 122.865 ;
        RECT 14.090 122.745 14.260 123.035 ;
        RECT 14.850 122.995 15.020 123.375 ;
        RECT 15.190 123.455 16.155 123.465 ;
        RECT 16.345 124.285 16.605 124.675 ;
        RECT 16.815 124.575 17.145 125.035 ;
        RECT 18.020 124.645 18.875 124.815 ;
        RECT 19.080 124.645 19.575 124.815 ;
        RECT 19.745 124.675 20.075 125.035 ;
        RECT 16.345 123.595 16.515 124.285 ;
        RECT 16.685 123.935 16.855 124.115 ;
        RECT 17.025 124.105 17.815 124.355 ;
        RECT 18.020 123.935 18.190 124.645 ;
        RECT 18.360 124.135 18.715 124.355 ;
        RECT 16.685 123.765 18.375 123.935 ;
        RECT 15.190 123.165 15.650 123.455 ;
        RECT 16.345 123.425 17.845 123.595 ;
        RECT 16.345 123.285 16.515 123.425 ;
        RECT 15.955 123.115 16.515 123.285 ;
        RECT 14.430 122.485 14.680 122.945 ;
        RECT 14.850 122.655 15.720 122.995 ;
        RECT 15.955 122.655 16.125 123.115 ;
        RECT 16.960 123.085 18.035 123.255 ;
        RECT 16.295 122.485 16.665 122.945 ;
        RECT 16.960 122.745 17.130 123.085 ;
        RECT 17.300 122.485 17.630 122.915 ;
        RECT 17.865 122.745 18.035 123.085 ;
        RECT 18.205 122.985 18.375 123.765 ;
        RECT 18.545 123.545 18.715 124.135 ;
        RECT 18.885 123.735 19.235 124.355 ;
        RECT 18.545 123.155 19.010 123.545 ;
        RECT 19.405 123.285 19.575 124.645 ;
        RECT 19.745 123.455 20.205 124.505 ;
        RECT 19.180 123.115 19.575 123.285 ;
        RECT 19.180 122.985 19.350 123.115 ;
        RECT 18.205 122.655 18.885 122.985 ;
        RECT 19.100 122.655 19.350 122.985 ;
        RECT 19.520 122.485 19.770 122.945 ;
        RECT 19.940 122.670 20.265 123.455 ;
        RECT 20.435 122.655 20.605 124.775 ;
        RECT 20.775 124.655 21.105 125.035 ;
        RECT 21.275 124.485 21.530 124.775 ;
        RECT 20.780 124.315 21.530 124.485 ;
        RECT 20.780 123.325 21.010 124.315 ;
        RECT 21.705 124.265 25.215 125.035 ;
        RECT 21.180 123.495 21.530 124.145 ;
        RECT 21.705 123.745 23.355 124.265 ;
        RECT 25.885 124.215 26.115 125.035 ;
        RECT 26.285 124.235 26.615 124.865 ;
        RECT 23.525 123.575 25.215 124.095 ;
        RECT 25.865 123.795 26.195 124.045 ;
        RECT 26.365 123.635 26.615 124.235 ;
        RECT 26.785 124.215 26.995 125.035 ;
        RECT 27.225 124.265 28.895 125.035 ;
        RECT 27.225 123.745 27.975 124.265 ;
        RECT 29.565 124.215 29.795 125.035 ;
        RECT 29.965 124.235 30.295 124.865 ;
        RECT 20.780 123.155 21.530 123.325 ;
        RECT 20.775 122.485 21.105 122.985 ;
        RECT 21.275 122.655 21.530 123.155 ;
        RECT 21.705 122.485 25.215 123.575 ;
        RECT 25.885 122.485 26.115 123.625 ;
        RECT 26.285 122.655 26.615 123.635 ;
        RECT 26.785 122.485 26.995 123.625 ;
        RECT 28.145 123.575 28.895 124.095 ;
        RECT 29.545 123.795 29.875 124.045 ;
        RECT 30.045 123.635 30.295 124.235 ;
        RECT 30.465 124.215 30.675 125.035 ;
        RECT 31.365 124.310 31.655 125.035 ;
        RECT 31.825 124.490 37.170 125.035 ;
        RECT 33.410 123.660 33.750 124.490 ;
        RECT 37.345 124.285 38.555 125.035 ;
        RECT 38.730 124.485 38.985 124.775 ;
        RECT 39.155 124.655 39.485 125.035 ;
        RECT 38.730 124.315 39.480 124.485 ;
        RECT 27.225 122.485 28.895 123.575 ;
        RECT 29.565 122.485 29.795 123.625 ;
        RECT 29.965 122.655 30.295 123.635 ;
        RECT 30.465 122.485 30.675 123.625 ;
        RECT 31.365 122.485 31.655 123.650 ;
        RECT 35.230 122.920 35.580 124.170 ;
        RECT 37.345 123.745 37.865 124.285 ;
        RECT 38.035 123.575 38.555 124.115 ;
        RECT 31.825 122.485 37.170 122.920 ;
        RECT 37.345 122.485 38.555 123.575 ;
        RECT 38.730 123.495 39.080 124.145 ;
        RECT 39.250 123.325 39.480 124.315 ;
        RECT 38.730 123.155 39.480 123.325 ;
        RECT 38.730 122.655 38.985 123.155 ;
        RECT 39.155 122.485 39.485 122.985 ;
        RECT 39.655 122.655 39.825 124.775 ;
        RECT 40.185 124.675 40.515 125.035 ;
        RECT 40.685 124.645 41.180 124.815 ;
        RECT 41.385 124.645 42.240 124.815 ;
        RECT 40.055 123.455 40.515 124.505 ;
        RECT 39.995 122.670 40.320 123.455 ;
        RECT 40.685 123.285 40.855 124.645 ;
        RECT 41.025 123.735 41.375 124.355 ;
        RECT 41.545 124.135 41.900 124.355 ;
        RECT 41.545 123.545 41.715 124.135 ;
        RECT 42.070 123.935 42.240 124.645 ;
        RECT 43.115 124.575 43.445 125.035 ;
        RECT 43.655 124.675 44.005 124.845 ;
        RECT 42.445 124.105 43.235 124.355 ;
        RECT 43.655 124.285 43.915 124.675 ;
        RECT 44.225 124.585 45.175 124.865 ;
        RECT 45.345 124.595 45.535 125.035 ;
        RECT 45.705 124.655 46.775 124.825 ;
        RECT 43.405 123.935 43.575 124.115 ;
        RECT 40.685 123.115 41.080 123.285 ;
        RECT 41.250 123.155 41.715 123.545 ;
        RECT 41.885 123.765 43.575 123.935 ;
        RECT 40.910 122.985 41.080 123.115 ;
        RECT 41.885 122.985 42.055 123.765 ;
        RECT 43.745 123.595 43.915 124.285 ;
        RECT 42.415 123.425 43.915 123.595 ;
        RECT 44.105 123.625 44.315 124.415 ;
        RECT 44.485 123.795 44.835 124.415 ;
        RECT 45.005 123.805 45.175 124.585 ;
        RECT 45.705 124.425 45.875 124.655 ;
        RECT 45.345 124.255 45.875 124.425 ;
        RECT 45.345 123.975 45.565 124.255 ;
        RECT 46.045 124.085 46.285 124.485 ;
        RECT 45.005 123.635 45.410 123.805 ;
        RECT 45.745 123.715 46.285 124.085 ;
        RECT 46.455 124.300 46.775 124.655 ;
        RECT 47.020 124.575 47.325 125.035 ;
        RECT 47.495 124.325 47.750 124.855 ;
        RECT 46.455 124.125 46.780 124.300 ;
        RECT 46.455 123.825 47.370 124.125 ;
        RECT 46.630 123.795 47.370 123.825 ;
        RECT 44.105 123.465 44.780 123.625 ;
        RECT 45.240 123.545 45.410 123.635 ;
        RECT 44.105 123.455 45.070 123.465 ;
        RECT 43.745 123.285 43.915 123.425 ;
        RECT 40.490 122.485 40.740 122.945 ;
        RECT 40.910 122.655 41.160 122.985 ;
        RECT 41.375 122.655 42.055 122.985 ;
        RECT 42.225 123.085 43.300 123.255 ;
        RECT 43.745 123.115 44.305 123.285 ;
        RECT 44.610 123.165 45.070 123.455 ;
        RECT 45.240 123.375 46.460 123.545 ;
        RECT 42.225 122.745 42.395 123.085 ;
        RECT 42.630 122.485 42.960 122.915 ;
        RECT 43.130 122.745 43.300 123.085 ;
        RECT 43.595 122.485 43.965 122.945 ;
        RECT 44.135 122.655 44.305 123.115 ;
        RECT 45.240 122.995 45.410 123.375 ;
        RECT 46.630 123.205 46.800 123.795 ;
        RECT 47.540 123.675 47.750 124.325 ;
        RECT 47.930 124.485 48.185 124.775 ;
        RECT 48.355 124.655 48.685 125.035 ;
        RECT 47.930 124.315 48.680 124.485 ;
        RECT 44.540 122.655 45.410 122.995 ;
        RECT 46.000 123.035 46.800 123.205 ;
        RECT 45.580 122.485 45.830 122.945 ;
        RECT 46.000 122.745 46.170 123.035 ;
        RECT 46.350 122.485 46.680 122.865 ;
        RECT 47.020 122.485 47.325 123.625 ;
        RECT 47.495 122.795 47.750 123.675 ;
        RECT 47.930 123.495 48.280 124.145 ;
        RECT 48.450 123.325 48.680 124.315 ;
        RECT 47.930 123.155 48.680 123.325 ;
        RECT 47.930 122.655 48.185 123.155 ;
        RECT 48.355 122.485 48.685 122.985 ;
        RECT 48.855 122.655 49.025 124.775 ;
        RECT 49.385 124.675 49.715 125.035 ;
        RECT 49.885 124.645 50.380 124.815 ;
        RECT 50.585 124.645 51.440 124.815 ;
        RECT 49.255 123.455 49.715 124.505 ;
        RECT 49.195 122.670 49.520 123.455 ;
        RECT 49.885 123.285 50.055 124.645 ;
        RECT 50.225 123.735 50.575 124.355 ;
        RECT 50.745 124.135 51.100 124.355 ;
        RECT 50.745 123.545 50.915 124.135 ;
        RECT 51.270 123.935 51.440 124.645 ;
        RECT 52.315 124.575 52.645 125.035 ;
        RECT 52.855 124.675 53.205 124.845 ;
        RECT 51.645 124.105 52.435 124.355 ;
        RECT 52.855 124.285 53.115 124.675 ;
        RECT 53.425 124.585 54.375 124.865 ;
        RECT 54.545 124.595 54.735 125.035 ;
        RECT 54.905 124.655 55.975 124.825 ;
        RECT 52.605 123.935 52.775 124.115 ;
        RECT 49.885 123.115 50.280 123.285 ;
        RECT 50.450 123.155 50.915 123.545 ;
        RECT 51.085 123.765 52.775 123.935 ;
        RECT 50.110 122.985 50.280 123.115 ;
        RECT 51.085 122.985 51.255 123.765 ;
        RECT 52.945 123.595 53.115 124.285 ;
        RECT 51.615 123.425 53.115 123.595 ;
        RECT 53.305 123.625 53.515 124.415 ;
        RECT 53.685 123.795 54.035 124.415 ;
        RECT 54.205 123.805 54.375 124.585 ;
        RECT 54.905 124.425 55.075 124.655 ;
        RECT 54.545 124.255 55.075 124.425 ;
        RECT 54.545 123.975 54.765 124.255 ;
        RECT 55.245 124.085 55.485 124.485 ;
        RECT 54.205 123.635 54.610 123.805 ;
        RECT 54.945 123.715 55.485 124.085 ;
        RECT 55.655 124.300 55.975 124.655 ;
        RECT 56.220 124.575 56.525 125.035 ;
        RECT 56.695 124.325 56.950 124.855 ;
        RECT 55.655 124.125 55.980 124.300 ;
        RECT 55.655 123.825 56.570 124.125 ;
        RECT 55.830 123.795 56.570 123.825 ;
        RECT 53.305 123.465 53.980 123.625 ;
        RECT 54.440 123.545 54.610 123.635 ;
        RECT 53.305 123.455 54.270 123.465 ;
        RECT 52.945 123.285 53.115 123.425 ;
        RECT 49.690 122.485 49.940 122.945 ;
        RECT 50.110 122.655 50.360 122.985 ;
        RECT 50.575 122.655 51.255 122.985 ;
        RECT 51.425 123.085 52.500 123.255 ;
        RECT 52.945 123.115 53.505 123.285 ;
        RECT 53.810 123.165 54.270 123.455 ;
        RECT 54.440 123.375 55.660 123.545 ;
        RECT 51.425 122.745 51.595 123.085 ;
        RECT 51.830 122.485 52.160 122.915 ;
        RECT 52.330 122.745 52.500 123.085 ;
        RECT 52.795 122.485 53.165 122.945 ;
        RECT 53.335 122.655 53.505 123.115 ;
        RECT 54.440 122.995 54.610 123.375 ;
        RECT 55.830 123.205 56.000 123.795 ;
        RECT 56.740 123.675 56.950 124.325 ;
        RECT 57.125 124.310 57.415 125.035 ;
        RECT 57.590 124.485 57.845 124.775 ;
        RECT 58.015 124.655 58.345 125.035 ;
        RECT 57.590 124.315 58.340 124.485 ;
        RECT 53.740 122.655 54.610 122.995 ;
        RECT 55.200 123.035 56.000 123.205 ;
        RECT 54.780 122.485 55.030 122.945 ;
        RECT 55.200 122.745 55.370 123.035 ;
        RECT 55.550 122.485 55.880 122.865 ;
        RECT 56.220 122.485 56.525 123.625 ;
        RECT 56.695 122.795 56.950 123.675 ;
        RECT 57.125 122.485 57.415 123.650 ;
        RECT 57.590 123.495 57.940 124.145 ;
        RECT 58.110 123.325 58.340 124.315 ;
        RECT 57.590 123.155 58.340 123.325 ;
        RECT 57.590 122.655 57.845 123.155 ;
        RECT 58.015 122.485 58.345 122.985 ;
        RECT 58.515 122.655 58.685 124.775 ;
        RECT 59.045 124.675 59.375 125.035 ;
        RECT 59.545 124.645 60.040 124.815 ;
        RECT 60.245 124.645 61.100 124.815 ;
        RECT 58.915 123.455 59.375 124.505 ;
        RECT 58.855 122.670 59.180 123.455 ;
        RECT 59.545 123.285 59.715 124.645 ;
        RECT 59.885 123.735 60.235 124.355 ;
        RECT 60.405 124.135 60.760 124.355 ;
        RECT 60.405 123.545 60.575 124.135 ;
        RECT 60.930 123.935 61.100 124.645 ;
        RECT 61.975 124.575 62.305 125.035 ;
        RECT 62.515 124.675 62.865 124.845 ;
        RECT 61.305 124.105 62.095 124.355 ;
        RECT 62.515 124.285 62.775 124.675 ;
        RECT 63.085 124.585 64.035 124.865 ;
        RECT 64.205 124.595 64.395 125.035 ;
        RECT 64.565 124.655 65.635 124.825 ;
        RECT 62.265 123.935 62.435 124.115 ;
        RECT 59.545 123.115 59.940 123.285 ;
        RECT 60.110 123.155 60.575 123.545 ;
        RECT 60.745 123.765 62.435 123.935 ;
        RECT 59.770 122.985 59.940 123.115 ;
        RECT 60.745 122.985 60.915 123.765 ;
        RECT 62.605 123.595 62.775 124.285 ;
        RECT 61.275 123.425 62.775 123.595 ;
        RECT 62.965 123.625 63.175 124.415 ;
        RECT 63.345 123.795 63.695 124.415 ;
        RECT 63.865 123.805 64.035 124.585 ;
        RECT 64.565 124.425 64.735 124.655 ;
        RECT 64.205 124.255 64.735 124.425 ;
        RECT 64.205 123.975 64.425 124.255 ;
        RECT 64.905 124.085 65.145 124.485 ;
        RECT 63.865 123.635 64.270 123.805 ;
        RECT 64.605 123.715 65.145 124.085 ;
        RECT 65.315 124.300 65.635 124.655 ;
        RECT 65.880 124.575 66.185 125.035 ;
        RECT 66.355 124.325 66.610 124.855 ;
        RECT 65.315 124.125 65.640 124.300 ;
        RECT 65.315 123.825 66.230 124.125 ;
        RECT 65.490 123.795 66.230 123.825 ;
        RECT 62.965 123.465 63.640 123.625 ;
        RECT 64.100 123.545 64.270 123.635 ;
        RECT 62.965 123.455 63.930 123.465 ;
        RECT 62.605 123.285 62.775 123.425 ;
        RECT 59.350 122.485 59.600 122.945 ;
        RECT 59.770 122.655 60.020 122.985 ;
        RECT 60.235 122.655 60.915 122.985 ;
        RECT 61.085 123.085 62.160 123.255 ;
        RECT 62.605 123.115 63.165 123.285 ;
        RECT 63.470 123.165 63.930 123.455 ;
        RECT 64.100 123.375 65.320 123.545 ;
        RECT 61.085 122.745 61.255 123.085 ;
        RECT 61.490 122.485 61.820 122.915 ;
        RECT 61.990 122.745 62.160 123.085 ;
        RECT 62.455 122.485 62.825 122.945 ;
        RECT 62.995 122.655 63.165 123.115 ;
        RECT 64.100 122.995 64.270 123.375 ;
        RECT 65.490 123.205 65.660 123.795 ;
        RECT 66.400 123.675 66.610 124.325 ;
        RECT 67.250 124.485 67.505 124.775 ;
        RECT 67.675 124.655 68.005 125.035 ;
        RECT 67.250 124.315 68.000 124.485 ;
        RECT 63.400 122.655 64.270 122.995 ;
        RECT 64.860 123.035 65.660 123.205 ;
        RECT 64.440 122.485 64.690 122.945 ;
        RECT 64.860 122.745 65.030 123.035 ;
        RECT 65.210 122.485 65.540 122.865 ;
        RECT 65.880 122.485 66.185 123.625 ;
        RECT 66.355 122.795 66.610 123.675 ;
        RECT 67.250 123.495 67.600 124.145 ;
        RECT 67.770 123.325 68.000 124.315 ;
        RECT 67.250 123.155 68.000 123.325 ;
        RECT 67.250 122.655 67.505 123.155 ;
        RECT 67.675 122.485 68.005 122.985 ;
        RECT 68.175 122.655 68.345 124.775 ;
        RECT 68.705 124.675 69.035 125.035 ;
        RECT 69.205 124.645 69.700 124.815 ;
        RECT 69.905 124.645 70.760 124.815 ;
        RECT 68.575 123.455 69.035 124.505 ;
        RECT 68.515 122.670 68.840 123.455 ;
        RECT 69.205 123.285 69.375 124.645 ;
        RECT 69.545 123.735 69.895 124.355 ;
        RECT 70.065 124.135 70.420 124.355 ;
        RECT 70.065 123.545 70.235 124.135 ;
        RECT 70.590 123.935 70.760 124.645 ;
        RECT 71.635 124.575 71.965 125.035 ;
        RECT 72.175 124.675 72.525 124.845 ;
        RECT 70.965 124.105 71.755 124.355 ;
        RECT 72.175 124.285 72.435 124.675 ;
        RECT 72.745 124.585 73.695 124.865 ;
        RECT 73.865 124.595 74.055 125.035 ;
        RECT 74.225 124.655 75.295 124.825 ;
        RECT 71.925 123.935 72.095 124.115 ;
        RECT 69.205 123.115 69.600 123.285 ;
        RECT 69.770 123.155 70.235 123.545 ;
        RECT 70.405 123.765 72.095 123.935 ;
        RECT 69.430 122.985 69.600 123.115 ;
        RECT 70.405 122.985 70.575 123.765 ;
        RECT 72.265 123.595 72.435 124.285 ;
        RECT 70.935 123.425 72.435 123.595 ;
        RECT 72.625 123.625 72.835 124.415 ;
        RECT 73.005 123.795 73.355 124.415 ;
        RECT 73.525 123.805 73.695 124.585 ;
        RECT 74.225 124.425 74.395 124.655 ;
        RECT 73.865 124.255 74.395 124.425 ;
        RECT 73.865 123.975 74.085 124.255 ;
        RECT 74.565 124.085 74.805 124.485 ;
        RECT 73.525 123.635 73.930 123.805 ;
        RECT 74.265 123.715 74.805 124.085 ;
        RECT 74.975 124.300 75.295 124.655 ;
        RECT 75.540 124.575 75.845 125.035 ;
        RECT 76.015 124.325 76.270 124.855 ;
        RECT 76.445 124.490 81.790 125.035 ;
        RECT 74.975 124.125 75.300 124.300 ;
        RECT 74.975 123.825 75.890 124.125 ;
        RECT 75.150 123.795 75.890 123.825 ;
        RECT 72.625 123.465 73.300 123.625 ;
        RECT 73.760 123.545 73.930 123.635 ;
        RECT 72.625 123.455 73.590 123.465 ;
        RECT 72.265 123.285 72.435 123.425 ;
        RECT 69.010 122.485 69.260 122.945 ;
        RECT 69.430 122.655 69.680 122.985 ;
        RECT 69.895 122.655 70.575 122.985 ;
        RECT 70.745 123.085 71.820 123.255 ;
        RECT 72.265 123.115 72.825 123.285 ;
        RECT 73.130 123.165 73.590 123.455 ;
        RECT 73.760 123.375 74.980 123.545 ;
        RECT 70.745 122.745 70.915 123.085 ;
        RECT 71.150 122.485 71.480 122.915 ;
        RECT 71.650 122.745 71.820 123.085 ;
        RECT 72.115 122.485 72.485 122.945 ;
        RECT 72.655 122.655 72.825 123.115 ;
        RECT 73.760 122.995 73.930 123.375 ;
        RECT 75.150 123.205 75.320 123.795 ;
        RECT 76.060 123.675 76.270 124.325 ;
        RECT 73.060 122.655 73.930 122.995 ;
        RECT 74.520 123.035 75.320 123.205 ;
        RECT 74.100 122.485 74.350 122.945 ;
        RECT 74.520 122.745 74.690 123.035 ;
        RECT 74.870 122.485 75.200 122.865 ;
        RECT 75.540 122.485 75.845 123.625 ;
        RECT 76.015 122.795 76.270 123.675 ;
        RECT 78.030 123.660 78.370 124.490 ;
        RECT 82.885 124.310 83.175 125.035 ;
        RECT 83.350 124.485 83.605 124.775 ;
        RECT 83.775 124.655 84.105 125.035 ;
        RECT 83.350 124.315 84.100 124.485 ;
        RECT 79.850 122.920 80.200 124.170 ;
        RECT 76.445 122.485 81.790 122.920 ;
        RECT 82.885 122.485 83.175 123.650 ;
        RECT 83.350 123.495 83.700 124.145 ;
        RECT 83.870 123.325 84.100 124.315 ;
        RECT 83.350 123.155 84.100 123.325 ;
        RECT 83.350 122.655 83.605 123.155 ;
        RECT 83.775 122.485 84.105 122.985 ;
        RECT 84.275 122.655 84.445 124.775 ;
        RECT 84.805 124.675 85.135 125.035 ;
        RECT 85.305 124.645 85.800 124.815 ;
        RECT 86.005 124.645 86.860 124.815 ;
        RECT 84.675 123.455 85.135 124.505 ;
        RECT 84.615 122.670 84.940 123.455 ;
        RECT 85.305 123.285 85.475 124.645 ;
        RECT 85.645 123.735 85.995 124.355 ;
        RECT 86.165 124.135 86.520 124.355 ;
        RECT 86.165 123.545 86.335 124.135 ;
        RECT 86.690 123.935 86.860 124.645 ;
        RECT 87.735 124.575 88.065 125.035 ;
        RECT 88.275 124.675 88.625 124.845 ;
        RECT 87.065 124.105 87.855 124.355 ;
        RECT 88.275 124.285 88.535 124.675 ;
        RECT 88.845 124.585 89.795 124.865 ;
        RECT 89.965 124.595 90.155 125.035 ;
        RECT 90.325 124.655 91.395 124.825 ;
        RECT 88.025 123.935 88.195 124.115 ;
        RECT 85.305 123.115 85.700 123.285 ;
        RECT 85.870 123.155 86.335 123.545 ;
        RECT 86.505 123.765 88.195 123.935 ;
        RECT 85.530 122.985 85.700 123.115 ;
        RECT 86.505 122.985 86.675 123.765 ;
        RECT 88.365 123.595 88.535 124.285 ;
        RECT 87.035 123.425 88.535 123.595 ;
        RECT 88.725 123.625 88.935 124.415 ;
        RECT 89.105 123.795 89.455 124.415 ;
        RECT 89.625 123.805 89.795 124.585 ;
        RECT 90.325 124.425 90.495 124.655 ;
        RECT 89.965 124.255 90.495 124.425 ;
        RECT 89.965 123.975 90.185 124.255 ;
        RECT 90.665 124.085 90.905 124.485 ;
        RECT 89.625 123.635 90.030 123.805 ;
        RECT 90.365 123.715 90.905 124.085 ;
        RECT 91.075 124.300 91.395 124.655 ;
        RECT 91.640 124.575 91.945 125.035 ;
        RECT 92.115 124.325 92.370 124.855 ;
        RECT 91.075 124.125 91.400 124.300 ;
        RECT 91.075 123.825 91.990 124.125 ;
        RECT 91.250 123.795 91.990 123.825 ;
        RECT 88.725 123.465 89.400 123.625 ;
        RECT 89.860 123.545 90.030 123.635 ;
        RECT 88.725 123.455 89.690 123.465 ;
        RECT 88.365 123.285 88.535 123.425 ;
        RECT 85.110 122.485 85.360 122.945 ;
        RECT 85.530 122.655 85.780 122.985 ;
        RECT 85.995 122.655 86.675 122.985 ;
        RECT 86.845 123.085 87.920 123.255 ;
        RECT 88.365 123.115 88.925 123.285 ;
        RECT 89.230 123.165 89.690 123.455 ;
        RECT 89.860 123.375 91.080 123.545 ;
        RECT 86.845 122.745 87.015 123.085 ;
        RECT 87.250 122.485 87.580 122.915 ;
        RECT 87.750 122.745 87.920 123.085 ;
        RECT 88.215 122.485 88.585 122.945 ;
        RECT 88.755 122.655 88.925 123.115 ;
        RECT 89.860 122.995 90.030 123.375 ;
        RECT 91.250 123.205 91.420 123.795 ;
        RECT 92.160 123.675 92.370 124.325 ;
        RECT 89.160 122.655 90.030 122.995 ;
        RECT 90.620 123.035 91.420 123.205 ;
        RECT 90.200 122.485 90.450 122.945 ;
        RECT 90.620 122.745 90.790 123.035 ;
        RECT 90.970 122.485 91.300 122.865 ;
        RECT 91.640 122.485 91.945 123.625 ;
        RECT 92.115 122.795 92.370 123.675 ;
        RECT 92.550 124.325 92.805 124.855 ;
        RECT 92.975 124.575 93.280 125.035 ;
        RECT 93.525 124.655 94.595 124.825 ;
        RECT 92.550 123.675 92.760 124.325 ;
        RECT 93.525 124.300 93.845 124.655 ;
        RECT 93.520 124.125 93.845 124.300 ;
        RECT 92.930 123.825 93.845 124.125 ;
        RECT 94.015 124.085 94.255 124.485 ;
        RECT 94.425 124.425 94.595 124.655 ;
        RECT 94.765 124.595 94.955 125.035 ;
        RECT 95.125 124.585 96.075 124.865 ;
        RECT 96.295 124.675 96.645 124.845 ;
        RECT 94.425 124.255 94.955 124.425 ;
        RECT 92.930 123.795 93.670 123.825 ;
        RECT 92.550 122.795 92.805 123.675 ;
        RECT 92.975 122.485 93.280 123.625 ;
        RECT 93.500 123.205 93.670 123.795 ;
        RECT 94.015 123.715 94.555 124.085 ;
        RECT 94.735 123.975 94.955 124.255 ;
        RECT 95.125 123.805 95.295 124.585 ;
        RECT 94.890 123.635 95.295 123.805 ;
        RECT 95.465 123.795 95.815 124.415 ;
        RECT 94.890 123.545 95.060 123.635 ;
        RECT 95.985 123.625 96.195 124.415 ;
        RECT 93.840 123.375 95.060 123.545 ;
        RECT 95.520 123.465 96.195 123.625 ;
        RECT 93.500 123.035 94.300 123.205 ;
        RECT 93.620 122.485 93.950 122.865 ;
        RECT 94.130 122.745 94.300 123.035 ;
        RECT 94.890 122.995 95.060 123.375 ;
        RECT 95.230 123.455 96.195 123.465 ;
        RECT 96.385 124.285 96.645 124.675 ;
        RECT 96.855 124.575 97.185 125.035 ;
        RECT 98.060 124.645 98.915 124.815 ;
        RECT 99.120 124.645 99.615 124.815 ;
        RECT 99.785 124.675 100.115 125.035 ;
        RECT 96.385 123.595 96.555 124.285 ;
        RECT 96.725 123.935 96.895 124.115 ;
        RECT 97.065 124.105 97.855 124.355 ;
        RECT 98.060 123.935 98.230 124.645 ;
        RECT 98.400 124.135 98.755 124.355 ;
        RECT 96.725 123.765 98.415 123.935 ;
        RECT 95.230 123.165 95.690 123.455 ;
        RECT 96.385 123.425 97.885 123.595 ;
        RECT 96.385 123.285 96.555 123.425 ;
        RECT 95.995 123.115 96.555 123.285 ;
        RECT 94.470 122.485 94.720 122.945 ;
        RECT 94.890 122.655 95.760 122.995 ;
        RECT 95.995 122.655 96.165 123.115 ;
        RECT 97.000 123.085 98.075 123.255 ;
        RECT 96.335 122.485 96.705 122.945 ;
        RECT 97.000 122.745 97.170 123.085 ;
        RECT 97.340 122.485 97.670 122.915 ;
        RECT 97.905 122.745 98.075 123.085 ;
        RECT 98.245 122.985 98.415 123.765 ;
        RECT 98.585 123.545 98.755 124.135 ;
        RECT 98.925 123.735 99.275 124.355 ;
        RECT 98.585 123.155 99.050 123.545 ;
        RECT 99.445 123.285 99.615 124.645 ;
        RECT 99.785 123.455 100.245 124.505 ;
        RECT 99.220 123.115 99.615 123.285 ;
        RECT 99.220 122.985 99.390 123.115 ;
        RECT 98.245 122.655 98.925 122.985 ;
        RECT 99.140 122.655 99.390 122.985 ;
        RECT 99.560 122.485 99.810 122.945 ;
        RECT 99.980 122.670 100.305 123.455 ;
        RECT 100.475 122.655 100.645 124.775 ;
        RECT 100.815 124.655 101.145 125.035 ;
        RECT 101.315 124.485 101.570 124.775 ;
        RECT 101.745 124.490 107.090 125.035 ;
        RECT 100.820 124.315 101.570 124.485 ;
        RECT 100.820 123.325 101.050 124.315 ;
        RECT 101.220 123.495 101.570 124.145 ;
        RECT 103.330 123.660 103.670 124.490 ;
        RECT 107.265 124.285 108.475 125.035 ;
        RECT 108.645 124.310 108.935 125.035 ;
        RECT 109.110 124.325 109.365 124.855 ;
        RECT 109.535 124.575 109.840 125.035 ;
        RECT 110.085 124.655 111.155 124.825 ;
        RECT 100.820 123.155 101.570 123.325 ;
        RECT 100.815 122.485 101.145 122.985 ;
        RECT 101.315 122.655 101.570 123.155 ;
        RECT 105.150 122.920 105.500 124.170 ;
        RECT 107.265 123.745 107.785 124.285 ;
        RECT 107.955 123.575 108.475 124.115 ;
        RECT 109.110 123.675 109.320 124.325 ;
        RECT 110.085 124.300 110.405 124.655 ;
        RECT 110.080 124.125 110.405 124.300 ;
        RECT 109.490 123.825 110.405 124.125 ;
        RECT 110.575 124.085 110.815 124.485 ;
        RECT 110.985 124.425 111.155 124.655 ;
        RECT 111.325 124.595 111.515 125.035 ;
        RECT 111.685 124.585 112.635 124.865 ;
        RECT 112.855 124.675 113.205 124.845 ;
        RECT 110.985 124.255 111.515 124.425 ;
        RECT 109.490 123.795 110.230 123.825 ;
        RECT 101.745 122.485 107.090 122.920 ;
        RECT 107.265 122.485 108.475 123.575 ;
        RECT 108.645 122.485 108.935 123.650 ;
        RECT 109.110 122.795 109.365 123.675 ;
        RECT 109.535 122.485 109.840 123.625 ;
        RECT 110.060 123.205 110.230 123.795 ;
        RECT 110.575 123.715 111.115 124.085 ;
        RECT 111.295 123.975 111.515 124.255 ;
        RECT 111.685 123.805 111.855 124.585 ;
        RECT 111.450 123.635 111.855 123.805 ;
        RECT 112.025 123.795 112.375 124.415 ;
        RECT 111.450 123.545 111.620 123.635 ;
        RECT 112.545 123.625 112.755 124.415 ;
        RECT 110.400 123.375 111.620 123.545 ;
        RECT 112.080 123.465 112.755 123.625 ;
        RECT 110.060 123.035 110.860 123.205 ;
        RECT 110.180 122.485 110.510 122.865 ;
        RECT 110.690 122.745 110.860 123.035 ;
        RECT 111.450 122.995 111.620 123.375 ;
        RECT 111.790 123.455 112.755 123.465 ;
        RECT 112.945 124.285 113.205 124.675 ;
        RECT 113.415 124.575 113.745 125.035 ;
        RECT 114.620 124.645 115.475 124.815 ;
        RECT 115.680 124.645 116.175 124.815 ;
        RECT 116.345 124.675 116.675 125.035 ;
        RECT 112.945 123.595 113.115 124.285 ;
        RECT 113.285 123.935 113.455 124.115 ;
        RECT 113.625 124.105 114.415 124.355 ;
        RECT 114.620 123.935 114.790 124.645 ;
        RECT 114.960 124.135 115.315 124.355 ;
        RECT 113.285 123.765 114.975 123.935 ;
        RECT 111.790 123.165 112.250 123.455 ;
        RECT 112.945 123.425 114.445 123.595 ;
        RECT 112.945 123.285 113.115 123.425 ;
        RECT 112.555 123.115 113.115 123.285 ;
        RECT 111.030 122.485 111.280 122.945 ;
        RECT 111.450 122.655 112.320 122.995 ;
        RECT 112.555 122.655 112.725 123.115 ;
        RECT 113.560 123.085 114.635 123.255 ;
        RECT 112.895 122.485 113.265 122.945 ;
        RECT 113.560 122.745 113.730 123.085 ;
        RECT 113.900 122.485 114.230 122.915 ;
        RECT 114.465 122.745 114.635 123.085 ;
        RECT 114.805 122.985 114.975 123.765 ;
        RECT 115.145 123.545 115.315 124.135 ;
        RECT 115.485 123.735 115.835 124.355 ;
        RECT 115.145 123.155 115.610 123.545 ;
        RECT 116.005 123.285 116.175 124.645 ;
        RECT 116.345 123.455 116.805 124.505 ;
        RECT 115.780 123.115 116.175 123.285 ;
        RECT 115.780 122.985 115.950 123.115 ;
        RECT 114.805 122.655 115.485 122.985 ;
        RECT 115.700 122.655 115.950 122.985 ;
        RECT 116.120 122.485 116.370 122.945 ;
        RECT 116.540 122.670 116.865 123.455 ;
        RECT 117.035 122.655 117.205 124.775 ;
        RECT 117.375 124.655 117.705 125.035 ;
        RECT 117.875 124.485 118.130 124.775 ;
        RECT 117.380 124.315 118.130 124.485 ;
        RECT 117.380 123.325 117.610 124.315 ;
        RECT 118.305 124.265 121.815 125.035 ;
        RECT 122.445 124.285 123.655 125.035 ;
        RECT 117.780 123.495 118.130 124.145 ;
        RECT 118.305 123.745 119.955 124.265 ;
        RECT 120.125 123.575 121.815 124.095 ;
        RECT 117.380 123.155 118.130 123.325 ;
        RECT 117.375 122.485 117.705 122.985 ;
        RECT 117.875 122.655 118.130 123.155 ;
        RECT 118.305 122.485 121.815 123.575 ;
        RECT 122.445 123.575 122.965 124.115 ;
        RECT 123.135 123.745 123.655 124.285 ;
        RECT 122.445 122.485 123.655 123.575 ;
        RECT 5.520 122.315 123.740 122.485 ;
        RECT 5.605 121.225 6.815 122.315 ;
        RECT 6.990 121.645 7.245 122.145 ;
        RECT 7.415 121.815 7.745 122.315 ;
        RECT 6.990 121.475 7.740 121.645 ;
        RECT 5.605 120.515 6.125 121.055 ;
        RECT 6.295 120.685 6.815 121.225 ;
        RECT 6.990 120.655 7.340 121.305 ;
        RECT 5.605 119.765 6.815 120.515 ;
        RECT 7.510 120.485 7.740 121.475 ;
        RECT 6.990 120.315 7.740 120.485 ;
        RECT 6.990 120.025 7.245 120.315 ;
        RECT 7.415 119.765 7.745 120.145 ;
        RECT 7.915 120.025 8.085 122.145 ;
        RECT 8.255 121.345 8.580 122.130 ;
        RECT 8.750 121.855 9.000 122.315 ;
        RECT 9.170 121.815 9.420 122.145 ;
        RECT 9.635 121.815 10.315 122.145 ;
        RECT 9.170 121.685 9.340 121.815 ;
        RECT 8.945 121.515 9.340 121.685 ;
        RECT 8.315 120.295 8.775 121.345 ;
        RECT 8.945 120.155 9.115 121.515 ;
        RECT 9.510 121.255 9.975 121.645 ;
        RECT 9.285 120.445 9.635 121.065 ;
        RECT 9.805 120.665 9.975 121.255 ;
        RECT 10.145 121.035 10.315 121.815 ;
        RECT 10.485 121.715 10.655 122.055 ;
        RECT 10.890 121.885 11.220 122.315 ;
        RECT 11.390 121.715 11.560 122.055 ;
        RECT 11.855 121.855 12.225 122.315 ;
        RECT 10.485 121.545 11.560 121.715 ;
        RECT 12.395 121.685 12.565 122.145 ;
        RECT 12.800 121.805 13.670 122.145 ;
        RECT 13.840 121.855 14.090 122.315 ;
        RECT 12.005 121.515 12.565 121.685 ;
        RECT 12.005 121.375 12.175 121.515 ;
        RECT 10.675 121.205 12.175 121.375 ;
        RECT 12.870 121.345 13.330 121.635 ;
        RECT 10.145 120.865 11.835 121.035 ;
        RECT 9.805 120.445 10.160 120.665 ;
        RECT 10.330 120.155 10.500 120.865 ;
        RECT 10.705 120.445 11.495 120.695 ;
        RECT 11.665 120.685 11.835 120.865 ;
        RECT 12.005 120.515 12.175 121.205 ;
        RECT 8.445 119.765 8.775 120.125 ;
        RECT 8.945 119.985 9.440 120.155 ;
        RECT 9.645 119.985 10.500 120.155 ;
        RECT 11.375 119.765 11.705 120.225 ;
        RECT 11.915 120.125 12.175 120.515 ;
        RECT 12.365 121.335 13.330 121.345 ;
        RECT 13.500 121.425 13.670 121.805 ;
        RECT 14.260 121.765 14.430 122.055 ;
        RECT 14.610 121.935 14.940 122.315 ;
        RECT 14.260 121.595 15.060 121.765 ;
        RECT 12.365 121.175 13.040 121.335 ;
        RECT 13.500 121.255 14.720 121.425 ;
        RECT 12.365 120.385 12.575 121.175 ;
        RECT 13.500 121.165 13.670 121.255 ;
        RECT 12.745 120.385 13.095 121.005 ;
        RECT 13.265 120.995 13.670 121.165 ;
        RECT 13.265 120.215 13.435 120.995 ;
        RECT 13.605 120.545 13.825 120.825 ;
        RECT 14.005 120.715 14.545 121.085 ;
        RECT 14.890 121.005 15.060 121.595 ;
        RECT 15.280 121.175 15.585 122.315 ;
        RECT 15.755 121.125 16.010 122.005 ;
        RECT 16.245 121.175 16.455 122.315 ;
        RECT 14.890 120.975 15.630 121.005 ;
        RECT 13.605 120.375 14.135 120.545 ;
        RECT 11.915 119.955 12.265 120.125 ;
        RECT 12.485 119.935 13.435 120.215 ;
        RECT 13.605 119.765 13.795 120.205 ;
        RECT 13.965 120.145 14.135 120.375 ;
        RECT 14.305 120.315 14.545 120.715 ;
        RECT 14.715 120.675 15.630 120.975 ;
        RECT 14.715 120.500 15.040 120.675 ;
        RECT 14.715 120.145 15.035 120.500 ;
        RECT 15.800 120.475 16.010 121.125 ;
        RECT 16.625 121.165 16.955 122.145 ;
        RECT 17.125 121.175 17.355 122.315 ;
        RECT 13.965 119.975 15.035 120.145 ;
        RECT 15.280 119.765 15.585 120.225 ;
        RECT 15.755 119.945 16.010 120.475 ;
        RECT 16.245 119.765 16.455 120.585 ;
        RECT 16.625 120.565 16.875 121.165 ;
        RECT 18.485 121.150 18.775 122.315 ;
        RECT 19.005 121.175 19.215 122.315 ;
        RECT 19.385 121.165 19.715 122.145 ;
        RECT 19.885 121.175 20.115 122.315 ;
        RECT 20.325 121.225 23.835 122.315 ;
        RECT 24.470 121.645 24.725 122.145 ;
        RECT 24.895 121.815 25.225 122.315 ;
        RECT 24.470 121.475 25.220 121.645 ;
        RECT 17.045 120.755 17.375 121.005 ;
        RECT 16.625 119.935 16.955 120.565 ;
        RECT 17.125 119.765 17.355 120.585 ;
        RECT 18.485 119.765 18.775 120.490 ;
        RECT 19.005 119.765 19.215 120.585 ;
        RECT 19.385 120.565 19.635 121.165 ;
        RECT 19.805 120.755 20.135 121.005 ;
        RECT 19.385 119.935 19.715 120.565 ;
        RECT 19.885 119.765 20.115 120.585 ;
        RECT 20.325 120.535 21.975 121.055 ;
        RECT 22.145 120.705 23.835 121.225 ;
        RECT 24.470 120.655 24.820 121.305 ;
        RECT 20.325 119.765 23.835 120.535 ;
        RECT 24.990 120.485 25.220 121.475 ;
        RECT 24.470 120.315 25.220 120.485 ;
        RECT 24.470 120.025 24.725 120.315 ;
        RECT 24.895 119.765 25.225 120.145 ;
        RECT 25.395 120.025 25.565 122.145 ;
        RECT 25.735 121.345 26.060 122.130 ;
        RECT 26.230 121.855 26.480 122.315 ;
        RECT 26.650 121.815 26.900 122.145 ;
        RECT 27.115 121.815 27.795 122.145 ;
        RECT 26.650 121.685 26.820 121.815 ;
        RECT 26.425 121.515 26.820 121.685 ;
        RECT 25.795 120.295 26.255 121.345 ;
        RECT 26.425 120.155 26.595 121.515 ;
        RECT 26.990 121.255 27.455 121.645 ;
        RECT 26.765 120.445 27.115 121.065 ;
        RECT 27.285 120.665 27.455 121.255 ;
        RECT 27.625 121.035 27.795 121.815 ;
        RECT 27.965 121.715 28.135 122.055 ;
        RECT 28.370 121.885 28.700 122.315 ;
        RECT 28.870 121.715 29.040 122.055 ;
        RECT 29.335 121.855 29.705 122.315 ;
        RECT 27.965 121.545 29.040 121.715 ;
        RECT 29.875 121.685 30.045 122.145 ;
        RECT 30.280 121.805 31.150 122.145 ;
        RECT 31.320 121.855 31.570 122.315 ;
        RECT 29.485 121.515 30.045 121.685 ;
        RECT 29.485 121.375 29.655 121.515 ;
        RECT 28.155 121.205 29.655 121.375 ;
        RECT 30.350 121.345 30.810 121.635 ;
        RECT 27.625 120.865 29.315 121.035 ;
        RECT 27.285 120.445 27.640 120.665 ;
        RECT 27.810 120.155 27.980 120.865 ;
        RECT 28.185 120.445 28.975 120.695 ;
        RECT 29.145 120.685 29.315 120.865 ;
        RECT 29.485 120.515 29.655 121.205 ;
        RECT 25.925 119.765 26.255 120.125 ;
        RECT 26.425 119.985 26.920 120.155 ;
        RECT 27.125 119.985 27.980 120.155 ;
        RECT 28.855 119.765 29.185 120.225 ;
        RECT 29.395 120.125 29.655 120.515 ;
        RECT 29.845 121.335 30.810 121.345 ;
        RECT 30.980 121.425 31.150 121.805 ;
        RECT 31.740 121.765 31.910 122.055 ;
        RECT 32.090 121.935 32.420 122.315 ;
        RECT 31.740 121.595 32.540 121.765 ;
        RECT 29.845 121.175 30.520 121.335 ;
        RECT 30.980 121.255 32.200 121.425 ;
        RECT 29.845 120.385 30.055 121.175 ;
        RECT 30.980 121.165 31.150 121.255 ;
        RECT 30.225 120.385 30.575 121.005 ;
        RECT 30.745 120.995 31.150 121.165 ;
        RECT 30.745 120.215 30.915 120.995 ;
        RECT 31.085 120.545 31.305 120.825 ;
        RECT 31.485 120.715 32.025 121.085 ;
        RECT 32.370 121.005 32.540 121.595 ;
        RECT 32.760 121.175 33.065 122.315 ;
        RECT 33.235 121.125 33.490 122.005 ;
        RECT 33.705 121.175 33.935 122.315 ;
        RECT 34.105 121.165 34.435 122.145 ;
        RECT 34.605 121.175 34.815 122.315 ;
        RECT 35.050 121.645 35.305 122.145 ;
        RECT 35.475 121.815 35.805 122.315 ;
        RECT 35.050 121.475 35.800 121.645 ;
        RECT 32.370 120.975 33.110 121.005 ;
        RECT 31.085 120.375 31.615 120.545 ;
        RECT 29.395 119.955 29.745 120.125 ;
        RECT 29.965 119.935 30.915 120.215 ;
        RECT 31.085 119.765 31.275 120.205 ;
        RECT 31.445 120.145 31.615 120.375 ;
        RECT 31.785 120.315 32.025 120.715 ;
        RECT 32.195 120.675 33.110 120.975 ;
        RECT 32.195 120.500 32.520 120.675 ;
        RECT 32.195 120.145 32.515 120.500 ;
        RECT 33.280 120.475 33.490 121.125 ;
        RECT 33.685 120.755 34.015 121.005 ;
        RECT 31.445 119.975 32.515 120.145 ;
        RECT 32.760 119.765 33.065 120.225 ;
        RECT 33.235 119.945 33.490 120.475 ;
        RECT 33.705 119.765 33.935 120.585 ;
        RECT 34.185 120.565 34.435 121.165 ;
        RECT 35.050 120.655 35.400 121.305 ;
        RECT 34.105 119.935 34.435 120.565 ;
        RECT 34.605 119.765 34.815 120.585 ;
        RECT 35.570 120.485 35.800 121.475 ;
        RECT 35.050 120.315 35.800 120.485 ;
        RECT 35.050 120.025 35.305 120.315 ;
        RECT 35.475 119.765 35.805 120.145 ;
        RECT 35.975 120.025 36.145 122.145 ;
        RECT 36.315 121.345 36.640 122.130 ;
        RECT 36.810 121.855 37.060 122.315 ;
        RECT 37.230 121.815 37.480 122.145 ;
        RECT 37.695 121.815 38.375 122.145 ;
        RECT 37.230 121.685 37.400 121.815 ;
        RECT 37.005 121.515 37.400 121.685 ;
        RECT 36.375 120.295 36.835 121.345 ;
        RECT 37.005 120.155 37.175 121.515 ;
        RECT 37.570 121.255 38.035 121.645 ;
        RECT 37.345 120.445 37.695 121.065 ;
        RECT 37.865 120.665 38.035 121.255 ;
        RECT 38.205 121.035 38.375 121.815 ;
        RECT 38.545 121.715 38.715 122.055 ;
        RECT 38.950 121.885 39.280 122.315 ;
        RECT 39.450 121.715 39.620 122.055 ;
        RECT 39.915 121.855 40.285 122.315 ;
        RECT 38.545 121.545 39.620 121.715 ;
        RECT 40.455 121.685 40.625 122.145 ;
        RECT 40.860 121.805 41.730 122.145 ;
        RECT 41.900 121.855 42.150 122.315 ;
        RECT 40.065 121.515 40.625 121.685 ;
        RECT 40.065 121.375 40.235 121.515 ;
        RECT 38.735 121.205 40.235 121.375 ;
        RECT 40.930 121.345 41.390 121.635 ;
        RECT 38.205 120.865 39.895 121.035 ;
        RECT 37.865 120.445 38.220 120.665 ;
        RECT 38.390 120.155 38.560 120.865 ;
        RECT 38.765 120.445 39.555 120.695 ;
        RECT 39.725 120.685 39.895 120.865 ;
        RECT 40.065 120.515 40.235 121.205 ;
        RECT 36.505 119.765 36.835 120.125 ;
        RECT 37.005 119.985 37.500 120.155 ;
        RECT 37.705 119.985 38.560 120.155 ;
        RECT 39.435 119.765 39.765 120.225 ;
        RECT 39.975 120.125 40.235 120.515 ;
        RECT 40.425 121.335 41.390 121.345 ;
        RECT 41.560 121.425 41.730 121.805 ;
        RECT 42.320 121.765 42.490 122.055 ;
        RECT 42.670 121.935 43.000 122.315 ;
        RECT 42.320 121.595 43.120 121.765 ;
        RECT 40.425 121.175 41.100 121.335 ;
        RECT 41.560 121.255 42.780 121.425 ;
        RECT 40.425 120.385 40.635 121.175 ;
        RECT 41.560 121.165 41.730 121.255 ;
        RECT 40.805 120.385 41.155 121.005 ;
        RECT 41.325 120.995 41.730 121.165 ;
        RECT 41.325 120.215 41.495 120.995 ;
        RECT 41.665 120.545 41.885 120.825 ;
        RECT 42.065 120.715 42.605 121.085 ;
        RECT 42.950 121.005 43.120 121.595 ;
        RECT 43.340 121.175 43.645 122.315 ;
        RECT 43.815 121.125 44.070 122.005 ;
        RECT 44.245 121.150 44.535 122.315 ;
        RECT 44.765 121.175 44.975 122.315 ;
        RECT 45.145 121.165 45.475 122.145 ;
        RECT 45.645 121.175 45.875 122.315 ;
        RECT 47.005 121.240 47.275 122.145 ;
        RECT 47.445 121.555 47.775 122.315 ;
        RECT 47.955 121.385 48.125 122.145 ;
        RECT 42.950 120.975 43.690 121.005 ;
        RECT 41.665 120.375 42.195 120.545 ;
        RECT 39.975 119.955 40.325 120.125 ;
        RECT 40.545 119.935 41.495 120.215 ;
        RECT 41.665 119.765 41.855 120.205 ;
        RECT 42.025 120.145 42.195 120.375 ;
        RECT 42.365 120.315 42.605 120.715 ;
        RECT 42.775 120.675 43.690 120.975 ;
        RECT 42.775 120.500 43.100 120.675 ;
        RECT 42.775 120.145 43.095 120.500 ;
        RECT 43.860 120.475 44.070 121.125 ;
        RECT 42.025 119.975 43.095 120.145 ;
        RECT 43.340 119.765 43.645 120.225 ;
        RECT 43.815 119.945 44.070 120.475 ;
        RECT 44.245 119.765 44.535 120.490 ;
        RECT 44.765 119.765 44.975 120.585 ;
        RECT 45.145 120.565 45.395 121.165 ;
        RECT 45.565 120.755 45.895 121.005 ;
        RECT 45.145 119.935 45.475 120.565 ;
        RECT 45.645 119.765 45.875 120.585 ;
        RECT 47.005 120.440 47.175 121.240 ;
        RECT 47.460 121.215 48.125 121.385 ;
        RECT 47.460 121.070 47.630 121.215 ;
        RECT 48.445 121.175 48.655 122.315 ;
        RECT 47.345 120.740 47.630 121.070 ;
        RECT 48.825 121.165 49.155 122.145 ;
        RECT 49.325 121.175 49.555 122.315 ;
        RECT 49.765 121.225 53.275 122.315 ;
        RECT 47.460 120.485 47.630 120.740 ;
        RECT 47.865 120.665 48.195 121.035 ;
        RECT 47.005 119.935 47.265 120.440 ;
        RECT 47.460 120.315 48.125 120.485 ;
        RECT 47.445 119.765 47.775 120.145 ;
        RECT 47.955 119.935 48.125 120.315 ;
        RECT 48.445 119.765 48.655 120.585 ;
        RECT 48.825 120.565 49.075 121.165 ;
        RECT 49.245 120.755 49.575 121.005 ;
        RECT 48.825 119.935 49.155 120.565 ;
        RECT 49.325 119.765 49.555 120.585 ;
        RECT 49.765 120.535 51.415 121.055 ;
        RECT 51.585 120.705 53.275 121.225 ;
        RECT 53.445 121.240 53.715 122.145 ;
        RECT 53.885 121.555 54.215 122.315 ;
        RECT 54.395 121.385 54.565 122.145 ;
        RECT 49.765 119.765 53.275 120.535 ;
        RECT 53.445 120.440 53.615 121.240 ;
        RECT 53.900 121.215 54.565 121.385 ;
        RECT 54.915 121.385 55.085 122.145 ;
        RECT 55.265 121.555 55.595 122.315 ;
        RECT 54.915 121.215 55.580 121.385 ;
        RECT 55.765 121.240 56.035 122.145 ;
        RECT 53.900 121.070 54.070 121.215 ;
        RECT 53.785 120.740 54.070 121.070 ;
        RECT 55.410 121.070 55.580 121.215 ;
        RECT 53.900 120.485 54.070 120.740 ;
        RECT 54.305 120.665 54.635 121.035 ;
        RECT 54.845 120.665 55.175 121.035 ;
        RECT 55.410 120.740 55.695 121.070 ;
        RECT 55.410 120.485 55.580 120.740 ;
        RECT 53.445 119.935 53.705 120.440 ;
        RECT 53.900 120.315 54.565 120.485 ;
        RECT 53.885 119.765 54.215 120.145 ;
        RECT 54.395 119.935 54.565 120.315 ;
        RECT 54.915 120.315 55.580 120.485 ;
        RECT 55.865 120.440 56.035 121.240 ;
        RECT 56.245 121.175 56.475 122.315 ;
        RECT 56.645 121.165 56.975 122.145 ;
        RECT 57.145 121.175 57.355 122.315 ;
        RECT 57.625 121.175 57.855 122.315 ;
        RECT 58.025 121.165 58.355 122.145 ;
        RECT 58.525 121.175 58.735 122.315 ;
        RECT 58.965 121.880 64.310 122.315 ;
        RECT 64.485 121.880 69.830 122.315 ;
        RECT 56.225 120.755 56.555 121.005 ;
        RECT 54.915 119.935 55.085 120.315 ;
        RECT 55.265 119.765 55.595 120.145 ;
        RECT 55.775 119.935 56.035 120.440 ;
        RECT 56.245 119.765 56.475 120.585 ;
        RECT 56.725 120.565 56.975 121.165 ;
        RECT 57.605 120.755 57.935 121.005 ;
        RECT 56.645 119.935 56.975 120.565 ;
        RECT 57.145 119.765 57.355 120.585 ;
        RECT 57.625 119.765 57.855 120.585 ;
        RECT 58.105 120.565 58.355 121.165 ;
        RECT 58.025 119.935 58.355 120.565 ;
        RECT 58.525 119.765 58.735 120.585 ;
        RECT 60.550 120.310 60.890 121.140 ;
        RECT 62.370 120.630 62.720 121.880 ;
        RECT 66.070 120.310 66.410 121.140 ;
        RECT 67.890 120.630 68.240 121.880 ;
        RECT 70.005 121.150 70.295 122.315 ;
        RECT 71.445 121.175 71.655 122.315 ;
        RECT 71.825 121.165 72.155 122.145 ;
        RECT 72.325 121.175 72.555 122.315 ;
        RECT 72.825 121.175 73.035 122.315 ;
        RECT 73.205 121.165 73.535 122.145 ;
        RECT 73.705 121.175 73.935 122.315 ;
        RECT 74.610 121.645 74.865 122.145 ;
        RECT 75.035 121.815 75.365 122.315 ;
        RECT 74.610 121.475 75.360 121.645 ;
        RECT 58.965 119.765 64.310 120.310 ;
        RECT 64.485 119.765 69.830 120.310 ;
        RECT 70.005 119.765 70.295 120.490 ;
        RECT 71.445 119.765 71.655 120.585 ;
        RECT 71.825 120.565 72.075 121.165 ;
        RECT 72.245 120.755 72.575 121.005 ;
        RECT 71.825 119.935 72.155 120.565 ;
        RECT 72.325 119.765 72.555 120.585 ;
        RECT 72.825 119.765 73.035 120.585 ;
        RECT 73.205 120.565 73.455 121.165 ;
        RECT 73.625 120.755 73.955 121.005 ;
        RECT 74.610 120.655 74.960 121.305 ;
        RECT 73.205 119.935 73.535 120.565 ;
        RECT 73.705 119.765 73.935 120.585 ;
        RECT 75.130 120.485 75.360 121.475 ;
        RECT 74.610 120.315 75.360 120.485 ;
        RECT 74.610 120.025 74.865 120.315 ;
        RECT 75.035 119.765 75.365 120.145 ;
        RECT 75.535 120.025 75.705 122.145 ;
        RECT 75.875 121.345 76.200 122.130 ;
        RECT 76.370 121.855 76.620 122.315 ;
        RECT 76.790 121.815 77.040 122.145 ;
        RECT 77.255 121.815 77.935 122.145 ;
        RECT 76.790 121.685 76.960 121.815 ;
        RECT 76.565 121.515 76.960 121.685 ;
        RECT 75.935 120.295 76.395 121.345 ;
        RECT 76.565 120.155 76.735 121.515 ;
        RECT 77.130 121.255 77.595 121.645 ;
        RECT 76.905 120.445 77.255 121.065 ;
        RECT 77.425 120.665 77.595 121.255 ;
        RECT 77.765 121.035 77.935 121.815 ;
        RECT 78.105 121.715 78.275 122.055 ;
        RECT 78.510 121.885 78.840 122.315 ;
        RECT 79.010 121.715 79.180 122.055 ;
        RECT 79.475 121.855 79.845 122.315 ;
        RECT 78.105 121.545 79.180 121.715 ;
        RECT 80.015 121.685 80.185 122.145 ;
        RECT 80.420 121.805 81.290 122.145 ;
        RECT 81.460 121.855 81.710 122.315 ;
        RECT 79.625 121.515 80.185 121.685 ;
        RECT 79.625 121.375 79.795 121.515 ;
        RECT 78.295 121.205 79.795 121.375 ;
        RECT 80.490 121.345 80.950 121.635 ;
        RECT 77.765 120.865 79.455 121.035 ;
        RECT 77.425 120.445 77.780 120.665 ;
        RECT 77.950 120.155 78.120 120.865 ;
        RECT 78.325 120.445 79.115 120.695 ;
        RECT 79.285 120.685 79.455 120.865 ;
        RECT 79.625 120.515 79.795 121.205 ;
        RECT 76.065 119.765 76.395 120.125 ;
        RECT 76.565 119.985 77.060 120.155 ;
        RECT 77.265 119.985 78.120 120.155 ;
        RECT 78.995 119.765 79.325 120.225 ;
        RECT 79.535 120.125 79.795 120.515 ;
        RECT 79.985 121.335 80.950 121.345 ;
        RECT 81.120 121.425 81.290 121.805 ;
        RECT 81.880 121.765 82.050 122.055 ;
        RECT 82.230 121.935 82.560 122.315 ;
        RECT 81.880 121.595 82.680 121.765 ;
        RECT 79.985 121.175 80.660 121.335 ;
        RECT 81.120 121.255 82.340 121.425 ;
        RECT 79.985 120.385 80.195 121.175 ;
        RECT 81.120 121.165 81.290 121.255 ;
        RECT 80.365 120.385 80.715 121.005 ;
        RECT 80.885 120.995 81.290 121.165 ;
        RECT 80.885 120.215 81.055 120.995 ;
        RECT 81.225 120.545 81.445 120.825 ;
        RECT 81.625 120.715 82.165 121.085 ;
        RECT 82.510 121.005 82.680 121.595 ;
        RECT 82.900 121.175 83.205 122.315 ;
        RECT 83.375 121.125 83.630 122.005 ;
        RECT 83.865 121.175 84.075 122.315 ;
        RECT 82.510 120.975 83.250 121.005 ;
        RECT 81.225 120.375 81.755 120.545 ;
        RECT 79.535 119.955 79.885 120.125 ;
        RECT 80.105 119.935 81.055 120.215 ;
        RECT 81.225 119.765 81.415 120.205 ;
        RECT 81.585 120.145 81.755 120.375 ;
        RECT 81.925 120.315 82.165 120.715 ;
        RECT 82.335 120.675 83.250 120.975 ;
        RECT 82.335 120.500 82.660 120.675 ;
        RECT 82.335 120.145 82.655 120.500 ;
        RECT 83.420 120.475 83.630 121.125 ;
        RECT 84.245 121.165 84.575 122.145 ;
        RECT 84.745 121.175 84.975 122.315 ;
        RECT 85.185 121.225 87.775 122.315 ;
        RECT 81.585 119.975 82.655 120.145 ;
        RECT 82.900 119.765 83.205 120.225 ;
        RECT 83.375 119.945 83.630 120.475 ;
        RECT 83.865 119.765 84.075 120.585 ;
        RECT 84.245 120.565 84.495 121.165 ;
        RECT 84.665 120.755 84.995 121.005 ;
        RECT 84.245 119.935 84.575 120.565 ;
        RECT 84.745 119.765 84.975 120.585 ;
        RECT 85.185 120.535 86.395 121.055 ;
        RECT 86.565 120.705 87.775 121.225 ;
        RECT 87.945 121.240 88.215 122.145 ;
        RECT 88.385 121.555 88.715 122.315 ;
        RECT 88.895 121.385 89.065 122.145 ;
        RECT 85.185 119.765 87.775 120.535 ;
        RECT 87.945 120.440 88.115 121.240 ;
        RECT 88.400 121.215 89.065 121.385 ;
        RECT 88.400 121.070 88.570 121.215 ;
        RECT 89.385 121.175 89.595 122.315 ;
        RECT 88.285 120.740 88.570 121.070 ;
        RECT 89.765 121.165 90.095 122.145 ;
        RECT 90.265 121.175 90.495 122.315 ;
        RECT 90.705 121.225 92.375 122.315 ;
        RECT 88.400 120.485 88.570 120.740 ;
        RECT 88.805 120.665 89.135 121.035 ;
        RECT 87.945 119.935 88.205 120.440 ;
        RECT 88.400 120.315 89.065 120.485 ;
        RECT 88.385 119.765 88.715 120.145 ;
        RECT 88.895 119.935 89.065 120.315 ;
        RECT 89.385 119.765 89.595 120.585 ;
        RECT 89.765 120.565 90.015 121.165 ;
        RECT 90.185 120.755 90.515 121.005 ;
        RECT 89.765 119.935 90.095 120.565 ;
        RECT 90.265 119.765 90.495 120.585 ;
        RECT 90.705 120.535 91.455 121.055 ;
        RECT 91.625 120.705 92.375 121.225 ;
        RECT 92.585 121.175 92.815 122.315 ;
        RECT 92.985 121.165 93.315 122.145 ;
        RECT 93.485 121.175 93.695 122.315 ;
        RECT 93.925 121.225 95.595 122.315 ;
        RECT 92.565 120.755 92.895 121.005 ;
        RECT 90.705 119.765 92.375 120.535 ;
        RECT 92.585 119.765 92.815 120.585 ;
        RECT 93.065 120.565 93.315 121.165 ;
        RECT 92.985 119.935 93.315 120.565 ;
        RECT 93.485 119.765 93.695 120.585 ;
        RECT 93.925 120.535 94.675 121.055 ;
        RECT 94.845 120.705 95.595 121.225 ;
        RECT 95.765 121.150 96.055 122.315 ;
        RECT 96.230 121.645 96.485 122.145 ;
        RECT 96.655 121.815 96.985 122.315 ;
        RECT 96.230 121.475 96.980 121.645 ;
        RECT 96.230 120.655 96.580 121.305 ;
        RECT 93.925 119.765 95.595 120.535 ;
        RECT 95.765 119.765 96.055 120.490 ;
        RECT 96.750 120.485 96.980 121.475 ;
        RECT 96.230 120.315 96.980 120.485 ;
        RECT 96.230 120.025 96.485 120.315 ;
        RECT 96.655 119.765 96.985 120.145 ;
        RECT 97.155 120.025 97.325 122.145 ;
        RECT 97.495 121.345 97.820 122.130 ;
        RECT 97.990 121.855 98.240 122.315 ;
        RECT 98.410 121.815 98.660 122.145 ;
        RECT 98.875 121.815 99.555 122.145 ;
        RECT 98.410 121.685 98.580 121.815 ;
        RECT 98.185 121.515 98.580 121.685 ;
        RECT 97.555 120.295 98.015 121.345 ;
        RECT 98.185 120.155 98.355 121.515 ;
        RECT 98.750 121.255 99.215 121.645 ;
        RECT 98.525 120.445 98.875 121.065 ;
        RECT 99.045 120.665 99.215 121.255 ;
        RECT 99.385 121.035 99.555 121.815 ;
        RECT 99.725 121.715 99.895 122.055 ;
        RECT 100.130 121.885 100.460 122.315 ;
        RECT 100.630 121.715 100.800 122.055 ;
        RECT 101.095 121.855 101.465 122.315 ;
        RECT 99.725 121.545 100.800 121.715 ;
        RECT 101.635 121.685 101.805 122.145 ;
        RECT 102.040 121.805 102.910 122.145 ;
        RECT 103.080 121.855 103.330 122.315 ;
        RECT 101.245 121.515 101.805 121.685 ;
        RECT 101.245 121.375 101.415 121.515 ;
        RECT 99.915 121.205 101.415 121.375 ;
        RECT 102.110 121.345 102.570 121.635 ;
        RECT 99.385 120.865 101.075 121.035 ;
        RECT 99.045 120.445 99.400 120.665 ;
        RECT 99.570 120.155 99.740 120.865 ;
        RECT 99.945 120.445 100.735 120.695 ;
        RECT 100.905 120.685 101.075 120.865 ;
        RECT 101.245 120.515 101.415 121.205 ;
        RECT 97.685 119.765 98.015 120.125 ;
        RECT 98.185 119.985 98.680 120.155 ;
        RECT 98.885 119.985 99.740 120.155 ;
        RECT 100.615 119.765 100.945 120.225 ;
        RECT 101.155 120.125 101.415 120.515 ;
        RECT 101.605 121.335 102.570 121.345 ;
        RECT 102.740 121.425 102.910 121.805 ;
        RECT 103.500 121.765 103.670 122.055 ;
        RECT 103.850 121.935 104.180 122.315 ;
        RECT 103.500 121.595 104.300 121.765 ;
        RECT 101.605 121.175 102.280 121.335 ;
        RECT 102.740 121.255 103.960 121.425 ;
        RECT 101.605 120.385 101.815 121.175 ;
        RECT 102.740 121.165 102.910 121.255 ;
        RECT 101.985 120.385 102.335 121.005 ;
        RECT 102.505 120.995 102.910 121.165 ;
        RECT 102.505 120.215 102.675 120.995 ;
        RECT 102.845 120.545 103.065 120.825 ;
        RECT 103.245 120.715 103.785 121.085 ;
        RECT 104.130 121.005 104.300 121.595 ;
        RECT 104.520 121.175 104.825 122.315 ;
        RECT 104.995 121.125 105.250 122.005 ;
        RECT 105.465 121.175 105.695 122.315 ;
        RECT 105.865 121.165 106.195 122.145 ;
        RECT 106.365 121.175 106.575 122.315 ;
        RECT 106.810 121.645 107.065 122.145 ;
        RECT 107.235 121.815 107.565 122.315 ;
        RECT 106.810 121.475 107.560 121.645 ;
        RECT 104.130 120.975 104.870 121.005 ;
        RECT 102.845 120.375 103.375 120.545 ;
        RECT 101.155 119.955 101.505 120.125 ;
        RECT 101.725 119.935 102.675 120.215 ;
        RECT 102.845 119.765 103.035 120.205 ;
        RECT 103.205 120.145 103.375 120.375 ;
        RECT 103.545 120.315 103.785 120.715 ;
        RECT 103.955 120.675 104.870 120.975 ;
        RECT 103.955 120.500 104.280 120.675 ;
        RECT 103.955 120.145 104.275 120.500 ;
        RECT 105.040 120.475 105.250 121.125 ;
        RECT 105.445 120.755 105.775 121.005 ;
        RECT 103.205 119.975 104.275 120.145 ;
        RECT 104.520 119.765 104.825 120.225 ;
        RECT 104.995 119.945 105.250 120.475 ;
        RECT 105.465 119.765 105.695 120.585 ;
        RECT 105.945 120.565 106.195 121.165 ;
        RECT 106.810 120.655 107.160 121.305 ;
        RECT 105.865 119.935 106.195 120.565 ;
        RECT 106.365 119.765 106.575 120.585 ;
        RECT 107.330 120.485 107.560 121.475 ;
        RECT 106.810 120.315 107.560 120.485 ;
        RECT 106.810 120.025 107.065 120.315 ;
        RECT 107.235 119.765 107.565 120.145 ;
        RECT 107.735 120.025 107.905 122.145 ;
        RECT 108.075 121.345 108.400 122.130 ;
        RECT 108.570 121.855 108.820 122.315 ;
        RECT 108.990 121.815 109.240 122.145 ;
        RECT 109.455 121.815 110.135 122.145 ;
        RECT 108.990 121.685 109.160 121.815 ;
        RECT 108.765 121.515 109.160 121.685 ;
        RECT 108.135 120.295 108.595 121.345 ;
        RECT 108.765 120.155 108.935 121.515 ;
        RECT 109.330 121.255 109.795 121.645 ;
        RECT 109.105 120.445 109.455 121.065 ;
        RECT 109.625 120.665 109.795 121.255 ;
        RECT 109.965 121.035 110.135 121.815 ;
        RECT 110.305 121.715 110.475 122.055 ;
        RECT 110.710 121.885 111.040 122.315 ;
        RECT 111.210 121.715 111.380 122.055 ;
        RECT 111.675 121.855 112.045 122.315 ;
        RECT 110.305 121.545 111.380 121.715 ;
        RECT 112.215 121.685 112.385 122.145 ;
        RECT 112.620 121.805 113.490 122.145 ;
        RECT 113.660 121.855 113.910 122.315 ;
        RECT 111.825 121.515 112.385 121.685 ;
        RECT 111.825 121.375 111.995 121.515 ;
        RECT 110.495 121.205 111.995 121.375 ;
        RECT 112.690 121.345 113.150 121.635 ;
        RECT 109.965 120.865 111.655 121.035 ;
        RECT 109.625 120.445 109.980 120.665 ;
        RECT 110.150 120.155 110.320 120.865 ;
        RECT 110.525 120.445 111.315 120.695 ;
        RECT 111.485 120.685 111.655 120.865 ;
        RECT 111.825 120.515 111.995 121.205 ;
        RECT 108.265 119.765 108.595 120.125 ;
        RECT 108.765 119.985 109.260 120.155 ;
        RECT 109.465 119.985 110.320 120.155 ;
        RECT 111.195 119.765 111.525 120.225 ;
        RECT 111.735 120.125 111.995 120.515 ;
        RECT 112.185 121.335 113.150 121.345 ;
        RECT 113.320 121.425 113.490 121.805 ;
        RECT 114.080 121.765 114.250 122.055 ;
        RECT 114.430 121.935 114.760 122.315 ;
        RECT 114.080 121.595 114.880 121.765 ;
        RECT 112.185 121.175 112.860 121.335 ;
        RECT 113.320 121.255 114.540 121.425 ;
        RECT 112.185 120.385 112.395 121.175 ;
        RECT 113.320 121.165 113.490 121.255 ;
        RECT 112.565 120.385 112.915 121.005 ;
        RECT 113.085 120.995 113.490 121.165 ;
        RECT 113.085 120.215 113.255 120.995 ;
        RECT 113.425 120.545 113.645 120.825 ;
        RECT 113.825 120.715 114.365 121.085 ;
        RECT 114.710 121.005 114.880 121.595 ;
        RECT 115.100 121.175 115.405 122.315 ;
        RECT 115.575 121.125 115.830 122.005 ;
        RECT 116.065 121.175 116.275 122.315 ;
        RECT 114.710 120.975 115.450 121.005 ;
        RECT 113.425 120.375 113.955 120.545 ;
        RECT 111.735 119.955 112.085 120.125 ;
        RECT 112.305 119.935 113.255 120.215 ;
        RECT 113.425 119.765 113.615 120.205 ;
        RECT 113.785 120.145 113.955 120.375 ;
        RECT 114.125 120.315 114.365 120.715 ;
        RECT 114.535 120.675 115.450 120.975 ;
        RECT 114.535 120.500 114.860 120.675 ;
        RECT 114.535 120.145 114.855 120.500 ;
        RECT 115.620 120.475 115.830 121.125 ;
        RECT 116.445 121.165 116.775 122.145 ;
        RECT 116.945 121.175 117.175 122.315 ;
        RECT 117.425 121.175 117.655 122.315 ;
        RECT 117.825 121.165 118.155 122.145 ;
        RECT 118.325 121.175 118.535 122.315 ;
        RECT 118.765 121.225 121.355 122.315 ;
        RECT 113.785 119.975 114.855 120.145 ;
        RECT 115.100 119.765 115.405 120.225 ;
        RECT 115.575 119.945 115.830 120.475 ;
        RECT 116.065 119.765 116.275 120.585 ;
        RECT 116.445 120.565 116.695 121.165 ;
        RECT 116.865 120.755 117.195 121.005 ;
        RECT 117.405 120.755 117.735 121.005 ;
        RECT 116.445 119.935 116.775 120.565 ;
        RECT 116.945 119.765 117.175 120.585 ;
        RECT 117.425 119.765 117.655 120.585 ;
        RECT 117.905 120.565 118.155 121.165 ;
        RECT 117.825 119.935 118.155 120.565 ;
        RECT 118.325 119.765 118.535 120.585 ;
        RECT 118.765 120.535 119.975 121.055 ;
        RECT 120.145 120.705 121.355 121.225 ;
        RECT 121.525 121.150 121.815 122.315 ;
        RECT 122.445 121.225 123.655 122.315 ;
        RECT 122.445 120.685 122.965 121.225 ;
        RECT 118.765 119.765 121.355 120.535 ;
        RECT 123.135 120.515 123.655 121.055 ;
        RECT 121.525 119.765 121.815 120.490 ;
        RECT 122.445 119.765 123.655 120.515 ;
        RECT 5.520 119.595 123.740 119.765 ;
        RECT 5.605 118.845 6.815 119.595 ;
        RECT 7.910 118.885 8.165 119.415 ;
        RECT 8.335 119.135 8.640 119.595 ;
        RECT 8.885 119.215 9.955 119.385 ;
        RECT 5.605 118.305 6.125 118.845 ;
        RECT 6.295 118.135 6.815 118.675 ;
        RECT 5.605 117.045 6.815 118.135 ;
        RECT 7.910 118.235 8.120 118.885 ;
        RECT 8.885 118.860 9.205 119.215 ;
        RECT 8.880 118.685 9.205 118.860 ;
        RECT 8.290 118.385 9.205 118.685 ;
        RECT 9.375 118.645 9.615 119.045 ;
        RECT 9.785 118.985 9.955 119.215 ;
        RECT 10.125 119.155 10.315 119.595 ;
        RECT 10.485 119.145 11.435 119.425 ;
        RECT 11.655 119.235 12.005 119.405 ;
        RECT 9.785 118.815 10.315 118.985 ;
        RECT 8.290 118.355 9.030 118.385 ;
        RECT 7.910 117.355 8.165 118.235 ;
        RECT 8.335 117.045 8.640 118.185 ;
        RECT 8.860 117.765 9.030 118.355 ;
        RECT 9.375 118.275 9.915 118.645 ;
        RECT 10.095 118.535 10.315 118.815 ;
        RECT 10.485 118.365 10.655 119.145 ;
        RECT 10.250 118.195 10.655 118.365 ;
        RECT 10.825 118.355 11.175 118.975 ;
        RECT 10.250 118.105 10.420 118.195 ;
        RECT 11.345 118.185 11.555 118.975 ;
        RECT 9.200 117.935 10.420 118.105 ;
        RECT 10.880 118.025 11.555 118.185 ;
        RECT 8.860 117.595 9.660 117.765 ;
        RECT 8.980 117.045 9.310 117.425 ;
        RECT 9.490 117.305 9.660 117.595 ;
        RECT 10.250 117.555 10.420 117.935 ;
        RECT 10.590 118.015 11.555 118.025 ;
        RECT 11.745 118.845 12.005 119.235 ;
        RECT 12.215 119.135 12.545 119.595 ;
        RECT 13.420 119.205 14.275 119.375 ;
        RECT 14.480 119.205 14.975 119.375 ;
        RECT 15.145 119.235 15.475 119.595 ;
        RECT 11.745 118.155 11.915 118.845 ;
        RECT 12.085 118.495 12.255 118.675 ;
        RECT 12.425 118.665 13.215 118.915 ;
        RECT 13.420 118.495 13.590 119.205 ;
        RECT 13.760 118.695 14.115 118.915 ;
        RECT 12.085 118.325 13.775 118.495 ;
        RECT 10.590 117.725 11.050 118.015 ;
        RECT 11.745 117.985 13.245 118.155 ;
        RECT 11.745 117.845 11.915 117.985 ;
        RECT 11.355 117.675 11.915 117.845 ;
        RECT 9.830 117.045 10.080 117.505 ;
        RECT 10.250 117.215 11.120 117.555 ;
        RECT 11.355 117.215 11.525 117.675 ;
        RECT 12.360 117.645 13.435 117.815 ;
        RECT 11.695 117.045 12.065 117.505 ;
        RECT 12.360 117.305 12.530 117.645 ;
        RECT 12.700 117.045 13.030 117.475 ;
        RECT 13.265 117.305 13.435 117.645 ;
        RECT 13.605 117.545 13.775 118.325 ;
        RECT 13.945 118.105 14.115 118.695 ;
        RECT 14.285 118.295 14.635 118.915 ;
        RECT 13.945 117.715 14.410 118.105 ;
        RECT 14.805 117.845 14.975 119.205 ;
        RECT 15.145 118.015 15.605 119.065 ;
        RECT 14.580 117.675 14.975 117.845 ;
        RECT 14.580 117.545 14.750 117.675 ;
        RECT 13.605 117.215 14.285 117.545 ;
        RECT 14.500 117.215 14.750 117.545 ;
        RECT 14.920 117.045 15.170 117.505 ;
        RECT 15.340 117.230 15.665 118.015 ;
        RECT 15.835 117.215 16.005 119.335 ;
        RECT 16.175 119.215 16.505 119.595 ;
        RECT 16.675 119.045 16.930 119.335 ;
        RECT 16.180 118.875 16.930 119.045 ;
        RECT 16.180 117.885 16.410 118.875 ;
        RECT 17.165 118.775 17.375 119.595 ;
        RECT 17.545 118.795 17.875 119.425 ;
        RECT 16.580 118.055 16.930 118.705 ;
        RECT 17.545 118.195 17.795 118.795 ;
        RECT 18.045 118.775 18.275 119.595 ;
        RECT 19.405 118.920 19.665 119.425 ;
        RECT 19.845 119.215 20.175 119.595 ;
        RECT 20.355 119.045 20.525 119.425 ;
        RECT 17.965 118.355 18.295 118.605 ;
        RECT 16.180 117.715 16.930 117.885 ;
        RECT 16.175 117.045 16.505 117.545 ;
        RECT 16.675 117.215 16.930 117.715 ;
        RECT 17.165 117.045 17.375 118.185 ;
        RECT 17.545 117.215 17.875 118.195 ;
        RECT 18.045 117.045 18.275 118.185 ;
        RECT 19.405 118.120 19.575 118.920 ;
        RECT 19.860 118.875 20.525 119.045 ;
        RECT 20.790 118.885 21.045 119.415 ;
        RECT 21.215 119.135 21.520 119.595 ;
        RECT 21.765 119.215 22.835 119.385 ;
        RECT 19.860 118.620 20.030 118.875 ;
        RECT 19.745 118.290 20.030 118.620 ;
        RECT 20.265 118.325 20.595 118.695 ;
        RECT 19.860 118.145 20.030 118.290 ;
        RECT 20.790 118.235 21.000 118.885 ;
        RECT 21.765 118.860 22.085 119.215 ;
        RECT 21.760 118.685 22.085 118.860 ;
        RECT 21.170 118.385 22.085 118.685 ;
        RECT 22.255 118.645 22.495 119.045 ;
        RECT 22.665 118.985 22.835 119.215 ;
        RECT 23.005 119.155 23.195 119.595 ;
        RECT 23.365 119.145 24.315 119.425 ;
        RECT 24.535 119.235 24.885 119.405 ;
        RECT 22.665 118.815 23.195 118.985 ;
        RECT 21.170 118.355 21.910 118.385 ;
        RECT 19.405 117.215 19.675 118.120 ;
        RECT 19.860 117.975 20.525 118.145 ;
        RECT 19.845 117.045 20.175 117.805 ;
        RECT 20.355 117.215 20.525 117.975 ;
        RECT 20.790 117.355 21.045 118.235 ;
        RECT 21.215 117.045 21.520 118.185 ;
        RECT 21.740 117.765 21.910 118.355 ;
        RECT 22.255 118.275 22.795 118.645 ;
        RECT 22.975 118.535 23.195 118.815 ;
        RECT 23.365 118.365 23.535 119.145 ;
        RECT 23.130 118.195 23.535 118.365 ;
        RECT 23.705 118.355 24.055 118.975 ;
        RECT 23.130 118.105 23.300 118.195 ;
        RECT 24.225 118.185 24.435 118.975 ;
        RECT 22.080 117.935 23.300 118.105 ;
        RECT 23.760 118.025 24.435 118.185 ;
        RECT 21.740 117.595 22.540 117.765 ;
        RECT 21.860 117.045 22.190 117.425 ;
        RECT 22.370 117.305 22.540 117.595 ;
        RECT 23.130 117.555 23.300 117.935 ;
        RECT 23.470 118.015 24.435 118.025 ;
        RECT 24.625 118.845 24.885 119.235 ;
        RECT 25.095 119.135 25.425 119.595 ;
        RECT 26.300 119.205 27.155 119.375 ;
        RECT 27.360 119.205 27.855 119.375 ;
        RECT 28.025 119.235 28.355 119.595 ;
        RECT 24.625 118.155 24.795 118.845 ;
        RECT 24.965 118.495 25.135 118.675 ;
        RECT 25.305 118.665 26.095 118.915 ;
        RECT 26.300 118.495 26.470 119.205 ;
        RECT 26.640 118.695 26.995 118.915 ;
        RECT 24.965 118.325 26.655 118.495 ;
        RECT 23.470 117.725 23.930 118.015 ;
        RECT 24.625 117.985 26.125 118.155 ;
        RECT 24.625 117.845 24.795 117.985 ;
        RECT 24.235 117.675 24.795 117.845 ;
        RECT 22.710 117.045 22.960 117.505 ;
        RECT 23.130 117.215 24.000 117.555 ;
        RECT 24.235 117.215 24.405 117.675 ;
        RECT 25.240 117.645 26.315 117.815 ;
        RECT 24.575 117.045 24.945 117.505 ;
        RECT 25.240 117.305 25.410 117.645 ;
        RECT 25.580 117.045 25.910 117.475 ;
        RECT 26.145 117.305 26.315 117.645 ;
        RECT 26.485 117.545 26.655 118.325 ;
        RECT 26.825 118.105 26.995 118.695 ;
        RECT 27.165 118.295 27.515 118.915 ;
        RECT 26.825 117.715 27.290 118.105 ;
        RECT 27.685 117.845 27.855 119.205 ;
        RECT 28.025 118.015 28.485 119.065 ;
        RECT 27.460 117.675 27.855 117.845 ;
        RECT 27.460 117.545 27.630 117.675 ;
        RECT 26.485 117.215 27.165 117.545 ;
        RECT 27.380 117.215 27.630 117.545 ;
        RECT 27.800 117.045 28.050 117.505 ;
        RECT 28.220 117.230 28.545 118.015 ;
        RECT 28.715 117.215 28.885 119.335 ;
        RECT 29.055 119.215 29.385 119.595 ;
        RECT 29.555 119.045 29.810 119.335 ;
        RECT 29.060 118.875 29.810 119.045 ;
        RECT 29.985 118.920 30.245 119.425 ;
        RECT 30.425 119.215 30.755 119.595 ;
        RECT 30.935 119.045 31.105 119.425 ;
        RECT 29.060 117.885 29.290 118.875 ;
        RECT 29.460 118.055 29.810 118.705 ;
        RECT 29.985 118.120 30.155 118.920 ;
        RECT 30.440 118.875 31.105 119.045 ;
        RECT 30.440 118.620 30.610 118.875 ;
        RECT 31.365 118.870 31.655 119.595 ;
        RECT 31.830 119.045 32.085 119.335 ;
        RECT 32.255 119.215 32.585 119.595 ;
        RECT 31.830 118.875 32.580 119.045 ;
        RECT 30.325 118.290 30.610 118.620 ;
        RECT 30.845 118.325 31.175 118.695 ;
        RECT 30.440 118.145 30.610 118.290 ;
        RECT 29.060 117.715 29.810 117.885 ;
        RECT 29.055 117.045 29.385 117.545 ;
        RECT 29.555 117.215 29.810 117.715 ;
        RECT 29.985 117.215 30.255 118.120 ;
        RECT 30.440 117.975 31.105 118.145 ;
        RECT 30.425 117.045 30.755 117.805 ;
        RECT 30.935 117.215 31.105 117.975 ;
        RECT 31.365 117.045 31.655 118.210 ;
        RECT 31.830 118.055 32.180 118.705 ;
        RECT 32.350 117.885 32.580 118.875 ;
        RECT 31.830 117.715 32.580 117.885 ;
        RECT 31.830 117.215 32.085 117.715 ;
        RECT 32.255 117.045 32.585 117.545 ;
        RECT 32.755 117.215 32.925 119.335 ;
        RECT 33.285 119.235 33.615 119.595 ;
        RECT 33.785 119.205 34.280 119.375 ;
        RECT 34.485 119.205 35.340 119.375 ;
        RECT 33.155 118.015 33.615 119.065 ;
        RECT 33.095 117.230 33.420 118.015 ;
        RECT 33.785 117.845 33.955 119.205 ;
        RECT 34.125 118.295 34.475 118.915 ;
        RECT 34.645 118.695 35.000 118.915 ;
        RECT 34.645 118.105 34.815 118.695 ;
        RECT 35.170 118.495 35.340 119.205 ;
        RECT 36.215 119.135 36.545 119.595 ;
        RECT 36.755 119.235 37.105 119.405 ;
        RECT 35.545 118.665 36.335 118.915 ;
        RECT 36.755 118.845 37.015 119.235 ;
        RECT 37.325 119.145 38.275 119.425 ;
        RECT 38.445 119.155 38.635 119.595 ;
        RECT 38.805 119.215 39.875 119.385 ;
        RECT 36.505 118.495 36.675 118.675 ;
        RECT 33.785 117.675 34.180 117.845 ;
        RECT 34.350 117.715 34.815 118.105 ;
        RECT 34.985 118.325 36.675 118.495 ;
        RECT 34.010 117.545 34.180 117.675 ;
        RECT 34.985 117.545 35.155 118.325 ;
        RECT 36.845 118.155 37.015 118.845 ;
        RECT 35.515 117.985 37.015 118.155 ;
        RECT 37.205 118.185 37.415 118.975 ;
        RECT 37.585 118.355 37.935 118.975 ;
        RECT 38.105 118.365 38.275 119.145 ;
        RECT 38.805 118.985 38.975 119.215 ;
        RECT 38.445 118.815 38.975 118.985 ;
        RECT 38.445 118.535 38.665 118.815 ;
        RECT 39.145 118.645 39.385 119.045 ;
        RECT 38.105 118.195 38.510 118.365 ;
        RECT 38.845 118.275 39.385 118.645 ;
        RECT 39.555 118.860 39.875 119.215 ;
        RECT 40.120 119.135 40.425 119.595 ;
        RECT 40.595 118.885 40.850 119.415 ;
        RECT 39.555 118.685 39.880 118.860 ;
        RECT 39.555 118.385 40.470 118.685 ;
        RECT 39.730 118.355 40.470 118.385 ;
        RECT 37.205 118.025 37.880 118.185 ;
        RECT 38.340 118.105 38.510 118.195 ;
        RECT 37.205 118.015 38.170 118.025 ;
        RECT 36.845 117.845 37.015 117.985 ;
        RECT 33.590 117.045 33.840 117.505 ;
        RECT 34.010 117.215 34.260 117.545 ;
        RECT 34.475 117.215 35.155 117.545 ;
        RECT 35.325 117.645 36.400 117.815 ;
        RECT 36.845 117.675 37.405 117.845 ;
        RECT 37.710 117.725 38.170 118.015 ;
        RECT 38.340 117.935 39.560 118.105 ;
        RECT 35.325 117.305 35.495 117.645 ;
        RECT 35.730 117.045 36.060 117.475 ;
        RECT 36.230 117.305 36.400 117.645 ;
        RECT 36.695 117.045 37.065 117.505 ;
        RECT 37.235 117.215 37.405 117.675 ;
        RECT 38.340 117.555 38.510 117.935 ;
        RECT 39.730 117.765 39.900 118.355 ;
        RECT 40.640 118.235 40.850 118.885 ;
        RECT 37.640 117.215 38.510 117.555 ;
        RECT 39.100 117.595 39.900 117.765 ;
        RECT 38.680 117.045 38.930 117.505 ;
        RECT 39.100 117.305 39.270 117.595 ;
        RECT 39.450 117.045 39.780 117.425 ;
        RECT 40.120 117.045 40.425 118.185 ;
        RECT 40.595 117.355 40.850 118.235 ;
        RECT 41.485 118.920 41.745 119.425 ;
        RECT 41.925 119.215 42.255 119.595 ;
        RECT 42.435 119.045 42.605 119.425 ;
        RECT 42.865 119.050 48.210 119.595 ;
        RECT 41.485 118.120 41.655 118.920 ;
        RECT 41.940 118.875 42.605 119.045 ;
        RECT 41.940 118.620 42.110 118.875 ;
        RECT 41.825 118.290 42.110 118.620 ;
        RECT 42.345 118.325 42.675 118.695 ;
        RECT 41.940 118.145 42.110 118.290 ;
        RECT 44.450 118.220 44.790 119.050 ;
        RECT 48.995 118.795 49.325 119.595 ;
        RECT 49.495 118.945 49.665 119.425 ;
        RECT 49.835 119.115 50.165 119.595 ;
        RECT 50.335 118.945 50.505 119.425 ;
        RECT 50.755 119.115 50.995 119.595 ;
        RECT 51.175 118.945 51.345 119.425 ;
        RECT 51.605 119.050 56.950 119.595 ;
        RECT 49.495 118.775 50.505 118.945 ;
        RECT 50.710 118.775 51.345 118.945 ;
        RECT 49.495 118.745 49.995 118.775 ;
        RECT 41.485 117.215 41.755 118.120 ;
        RECT 41.940 117.975 42.605 118.145 ;
        RECT 41.925 117.045 42.255 117.805 ;
        RECT 42.435 117.215 42.605 117.975 ;
        RECT 46.270 117.480 46.620 118.730 ;
        RECT 49.495 118.235 49.990 118.745 ;
        RECT 50.710 118.605 50.880 118.775 ;
        RECT 50.380 118.435 50.880 118.605 ;
        RECT 42.865 117.045 48.210 117.480 ;
        RECT 48.995 117.045 49.325 118.195 ;
        RECT 49.495 118.065 50.505 118.235 ;
        RECT 49.495 117.215 49.665 118.065 ;
        RECT 49.835 117.045 50.165 117.845 ;
        RECT 50.335 117.215 50.505 118.065 ;
        RECT 50.710 118.195 50.880 118.435 ;
        RECT 51.050 118.365 51.430 118.605 ;
        RECT 53.190 118.220 53.530 119.050 ;
        RECT 57.125 118.870 57.415 119.595 ;
        RECT 57.585 118.845 58.795 119.595 ;
        RECT 50.710 118.025 51.425 118.195 ;
        RECT 50.685 117.045 50.925 117.845 ;
        RECT 51.095 117.215 51.425 118.025 ;
        RECT 55.010 117.480 55.360 118.730 ;
        RECT 57.585 118.305 58.105 118.845 ;
        RECT 59.005 118.775 59.235 119.595 ;
        RECT 59.405 118.795 59.735 119.425 ;
        RECT 51.605 117.045 56.950 117.480 ;
        RECT 57.125 117.045 57.415 118.210 ;
        RECT 58.275 118.135 58.795 118.675 ;
        RECT 58.985 118.355 59.315 118.605 ;
        RECT 59.485 118.195 59.735 118.795 ;
        RECT 59.905 118.775 60.115 119.595 ;
        RECT 60.345 118.825 63.855 119.595 ;
        RECT 64.490 118.885 64.745 119.415 ;
        RECT 64.915 119.135 65.220 119.595 ;
        RECT 65.465 119.215 66.535 119.385 ;
        RECT 60.345 118.305 61.995 118.825 ;
        RECT 57.585 117.045 58.795 118.135 ;
        RECT 59.005 117.045 59.235 118.185 ;
        RECT 59.405 117.215 59.735 118.195 ;
        RECT 59.905 117.045 60.115 118.185 ;
        RECT 62.165 118.135 63.855 118.655 ;
        RECT 60.345 117.045 63.855 118.135 ;
        RECT 64.490 118.235 64.700 118.885 ;
        RECT 65.465 118.860 65.785 119.215 ;
        RECT 65.460 118.685 65.785 118.860 ;
        RECT 64.870 118.385 65.785 118.685 ;
        RECT 65.955 118.645 66.195 119.045 ;
        RECT 66.365 118.985 66.535 119.215 ;
        RECT 66.705 119.155 66.895 119.595 ;
        RECT 67.065 119.145 68.015 119.425 ;
        RECT 68.235 119.235 68.585 119.405 ;
        RECT 66.365 118.815 66.895 118.985 ;
        RECT 64.870 118.355 65.610 118.385 ;
        RECT 64.490 117.355 64.745 118.235 ;
        RECT 64.915 117.045 65.220 118.185 ;
        RECT 65.440 117.765 65.610 118.355 ;
        RECT 65.955 118.275 66.495 118.645 ;
        RECT 66.675 118.535 66.895 118.815 ;
        RECT 67.065 118.365 67.235 119.145 ;
        RECT 66.830 118.195 67.235 118.365 ;
        RECT 67.405 118.355 67.755 118.975 ;
        RECT 66.830 118.105 67.000 118.195 ;
        RECT 67.925 118.185 68.135 118.975 ;
        RECT 65.780 117.935 67.000 118.105 ;
        RECT 67.460 118.025 68.135 118.185 ;
        RECT 65.440 117.595 66.240 117.765 ;
        RECT 65.560 117.045 65.890 117.425 ;
        RECT 66.070 117.305 66.240 117.595 ;
        RECT 66.830 117.555 67.000 117.935 ;
        RECT 67.170 118.015 68.135 118.025 ;
        RECT 68.325 118.845 68.585 119.235 ;
        RECT 68.795 119.135 69.125 119.595 ;
        RECT 70.000 119.205 70.855 119.375 ;
        RECT 71.060 119.205 71.555 119.375 ;
        RECT 71.725 119.235 72.055 119.595 ;
        RECT 68.325 118.155 68.495 118.845 ;
        RECT 68.665 118.495 68.835 118.675 ;
        RECT 69.005 118.665 69.795 118.915 ;
        RECT 70.000 118.495 70.170 119.205 ;
        RECT 70.340 118.695 70.695 118.915 ;
        RECT 68.665 118.325 70.355 118.495 ;
        RECT 67.170 117.725 67.630 118.015 ;
        RECT 68.325 117.985 69.825 118.155 ;
        RECT 68.325 117.845 68.495 117.985 ;
        RECT 67.935 117.675 68.495 117.845 ;
        RECT 66.410 117.045 66.660 117.505 ;
        RECT 66.830 117.215 67.700 117.555 ;
        RECT 67.935 117.215 68.105 117.675 ;
        RECT 68.940 117.645 70.015 117.815 ;
        RECT 68.275 117.045 68.645 117.505 ;
        RECT 68.940 117.305 69.110 117.645 ;
        RECT 69.280 117.045 69.610 117.475 ;
        RECT 69.845 117.305 70.015 117.645 ;
        RECT 70.185 117.545 70.355 118.325 ;
        RECT 70.525 118.105 70.695 118.695 ;
        RECT 70.865 118.295 71.215 118.915 ;
        RECT 70.525 117.715 70.990 118.105 ;
        RECT 71.385 117.845 71.555 119.205 ;
        RECT 71.725 118.015 72.185 119.065 ;
        RECT 71.160 117.675 71.555 117.845 ;
        RECT 71.160 117.545 71.330 117.675 ;
        RECT 70.185 117.215 70.865 117.545 ;
        RECT 71.080 117.215 71.330 117.545 ;
        RECT 71.500 117.045 71.750 117.505 ;
        RECT 71.920 117.230 72.245 118.015 ;
        RECT 72.415 117.215 72.585 119.335 ;
        RECT 72.755 119.215 73.085 119.595 ;
        RECT 73.255 119.045 73.510 119.335 ;
        RECT 72.760 118.875 73.510 119.045 ;
        RECT 73.775 118.945 73.945 119.425 ;
        RECT 74.125 119.115 74.365 119.595 ;
        RECT 74.615 118.945 74.785 119.425 ;
        RECT 74.955 119.115 75.285 119.595 ;
        RECT 75.455 118.945 75.625 119.425 ;
        RECT 72.760 117.885 72.990 118.875 ;
        RECT 73.775 118.775 74.410 118.945 ;
        RECT 74.615 118.775 75.625 118.945 ;
        RECT 75.795 118.795 76.125 119.595 ;
        RECT 76.445 118.825 79.035 119.595 ;
        RECT 79.205 118.920 79.465 119.425 ;
        RECT 79.645 119.215 79.975 119.595 ;
        RECT 80.155 119.045 80.325 119.425 ;
        RECT 73.160 118.055 73.510 118.705 ;
        RECT 74.240 118.605 74.410 118.775 ;
        RECT 75.125 118.745 75.625 118.775 ;
        RECT 73.690 118.365 74.070 118.605 ;
        RECT 74.240 118.435 74.740 118.605 ;
        RECT 74.240 118.195 74.410 118.435 ;
        RECT 75.130 118.235 75.625 118.745 ;
        RECT 76.445 118.305 77.655 118.825 ;
        RECT 73.695 118.025 74.410 118.195 ;
        RECT 74.615 118.065 75.625 118.235 ;
        RECT 72.760 117.715 73.510 117.885 ;
        RECT 72.755 117.045 73.085 117.545 ;
        RECT 73.255 117.215 73.510 117.715 ;
        RECT 73.695 117.215 74.025 118.025 ;
        RECT 74.195 117.045 74.435 117.845 ;
        RECT 74.615 117.215 74.785 118.065 ;
        RECT 74.955 117.045 75.285 117.845 ;
        RECT 75.455 117.215 75.625 118.065 ;
        RECT 75.795 117.045 76.125 118.195 ;
        RECT 77.825 118.135 79.035 118.655 ;
        RECT 76.445 117.045 79.035 118.135 ;
        RECT 79.205 118.120 79.375 118.920 ;
        RECT 79.660 118.875 80.325 119.045 ;
        RECT 79.660 118.620 79.830 118.875 ;
        RECT 80.585 118.825 82.255 119.595 ;
        RECT 82.885 118.870 83.175 119.595 ;
        RECT 83.345 119.050 88.690 119.595 ;
        RECT 79.545 118.290 79.830 118.620 ;
        RECT 80.065 118.325 80.395 118.695 ;
        RECT 80.585 118.305 81.335 118.825 ;
        RECT 79.660 118.145 79.830 118.290 ;
        RECT 79.205 117.215 79.475 118.120 ;
        RECT 79.660 117.975 80.325 118.145 ;
        RECT 81.505 118.135 82.255 118.655 ;
        RECT 84.930 118.220 85.270 119.050 ;
        RECT 88.865 118.825 90.535 119.595 ;
        RECT 91.255 119.045 91.425 119.425 ;
        RECT 91.605 119.215 91.935 119.595 ;
        RECT 91.255 118.875 91.920 119.045 ;
        RECT 92.115 118.920 92.375 119.425 ;
        RECT 79.645 117.045 79.975 117.805 ;
        RECT 80.155 117.215 80.325 117.975 ;
        RECT 80.585 117.045 82.255 118.135 ;
        RECT 82.885 117.045 83.175 118.210 ;
        RECT 86.750 117.480 87.100 118.730 ;
        RECT 88.865 118.305 89.615 118.825 ;
        RECT 89.785 118.135 90.535 118.655 ;
        RECT 91.185 118.325 91.515 118.695 ;
        RECT 91.750 118.620 91.920 118.875 ;
        RECT 91.750 118.290 92.035 118.620 ;
        RECT 91.750 118.145 91.920 118.290 ;
        RECT 83.345 117.045 88.690 117.480 ;
        RECT 88.865 117.045 90.535 118.135 ;
        RECT 91.255 117.975 91.920 118.145 ;
        RECT 92.205 118.120 92.375 118.920 ;
        RECT 92.545 118.825 95.135 119.595 ;
        RECT 95.855 119.045 96.025 119.425 ;
        RECT 96.205 119.215 96.535 119.595 ;
        RECT 95.855 118.875 96.520 119.045 ;
        RECT 96.715 118.920 96.975 119.425 ;
        RECT 92.545 118.305 93.755 118.825 ;
        RECT 93.925 118.135 95.135 118.655 ;
        RECT 95.785 118.325 96.115 118.695 ;
        RECT 96.350 118.620 96.520 118.875 ;
        RECT 96.350 118.290 96.635 118.620 ;
        RECT 96.350 118.145 96.520 118.290 ;
        RECT 91.255 117.215 91.425 117.975 ;
        RECT 91.605 117.045 91.935 117.805 ;
        RECT 92.105 117.215 92.375 118.120 ;
        RECT 92.545 117.045 95.135 118.135 ;
        RECT 95.855 117.975 96.520 118.145 ;
        RECT 96.805 118.120 96.975 118.920 ;
        RECT 97.145 118.825 98.815 119.595 ;
        RECT 97.145 118.305 97.895 118.825 ;
        RECT 99.025 118.775 99.255 119.595 ;
        RECT 99.425 118.795 99.755 119.425 ;
        RECT 98.065 118.135 98.815 118.655 ;
        RECT 99.005 118.355 99.335 118.605 ;
        RECT 99.505 118.195 99.755 118.795 ;
        RECT 99.925 118.775 100.135 119.595 ;
        RECT 100.365 118.825 102.035 119.595 ;
        RECT 102.295 119.045 102.465 119.425 ;
        RECT 102.645 119.215 102.975 119.595 ;
        RECT 102.295 118.875 102.960 119.045 ;
        RECT 103.155 118.920 103.415 119.425 ;
        RECT 100.365 118.305 101.115 118.825 ;
        RECT 95.855 117.215 96.025 117.975 ;
        RECT 96.205 117.045 96.535 117.805 ;
        RECT 96.705 117.215 96.975 118.120 ;
        RECT 97.145 117.045 98.815 118.135 ;
        RECT 99.025 117.045 99.255 118.185 ;
        RECT 99.425 117.215 99.755 118.195 ;
        RECT 99.925 117.045 100.135 118.185 ;
        RECT 101.285 118.135 102.035 118.655 ;
        RECT 102.225 118.325 102.555 118.695 ;
        RECT 102.790 118.620 102.960 118.875 ;
        RECT 102.790 118.290 103.075 118.620 ;
        RECT 102.790 118.145 102.960 118.290 ;
        RECT 100.365 117.045 102.035 118.135 ;
        RECT 102.295 117.975 102.960 118.145 ;
        RECT 103.245 118.120 103.415 118.920 ;
        RECT 103.585 118.825 105.255 119.595 ;
        RECT 105.975 119.045 106.145 119.425 ;
        RECT 106.325 119.215 106.655 119.595 ;
        RECT 105.975 118.875 106.640 119.045 ;
        RECT 106.835 118.920 107.095 119.425 ;
        RECT 103.585 118.305 104.335 118.825 ;
        RECT 104.505 118.135 105.255 118.655 ;
        RECT 105.905 118.325 106.235 118.695 ;
        RECT 106.470 118.620 106.640 118.875 ;
        RECT 106.470 118.290 106.755 118.620 ;
        RECT 106.470 118.145 106.640 118.290 ;
        RECT 102.295 117.215 102.465 117.975 ;
        RECT 102.645 117.045 102.975 117.805 ;
        RECT 103.145 117.215 103.415 118.120 ;
        RECT 103.585 117.045 105.255 118.135 ;
        RECT 105.975 117.975 106.640 118.145 ;
        RECT 106.925 118.120 107.095 118.920 ;
        RECT 107.355 119.045 107.525 119.425 ;
        RECT 107.705 119.215 108.035 119.595 ;
        RECT 107.355 118.875 108.020 119.045 ;
        RECT 108.215 118.920 108.475 119.425 ;
        RECT 107.285 118.325 107.615 118.695 ;
        RECT 107.850 118.620 108.020 118.875 ;
        RECT 107.850 118.290 108.135 118.620 ;
        RECT 107.850 118.145 108.020 118.290 ;
        RECT 105.975 117.215 106.145 117.975 ;
        RECT 106.325 117.045 106.655 117.805 ;
        RECT 106.825 117.215 107.095 118.120 ;
        RECT 107.355 117.975 108.020 118.145 ;
        RECT 108.305 118.120 108.475 118.920 ;
        RECT 108.645 118.870 108.935 119.595 ;
        RECT 109.110 119.045 109.365 119.335 ;
        RECT 109.535 119.215 109.865 119.595 ;
        RECT 109.110 118.875 109.860 119.045 ;
        RECT 107.355 117.215 107.525 117.975 ;
        RECT 107.705 117.045 108.035 117.805 ;
        RECT 108.205 117.215 108.475 118.120 ;
        RECT 108.645 117.045 108.935 118.210 ;
        RECT 109.110 118.055 109.460 118.705 ;
        RECT 109.630 117.885 109.860 118.875 ;
        RECT 109.110 117.715 109.860 117.885 ;
        RECT 109.110 117.215 109.365 117.715 ;
        RECT 109.535 117.045 109.865 117.545 ;
        RECT 110.035 117.215 110.205 119.335 ;
        RECT 110.565 119.235 110.895 119.595 ;
        RECT 111.065 119.205 111.560 119.375 ;
        RECT 111.765 119.205 112.620 119.375 ;
        RECT 110.435 118.015 110.895 119.065 ;
        RECT 110.375 117.230 110.700 118.015 ;
        RECT 111.065 117.845 111.235 119.205 ;
        RECT 111.405 118.295 111.755 118.915 ;
        RECT 111.925 118.695 112.280 118.915 ;
        RECT 111.925 118.105 112.095 118.695 ;
        RECT 112.450 118.495 112.620 119.205 ;
        RECT 113.495 119.135 113.825 119.595 ;
        RECT 114.035 119.235 114.385 119.405 ;
        RECT 112.825 118.665 113.615 118.915 ;
        RECT 114.035 118.845 114.295 119.235 ;
        RECT 114.605 119.145 115.555 119.425 ;
        RECT 115.725 119.155 115.915 119.595 ;
        RECT 116.085 119.215 117.155 119.385 ;
        RECT 113.785 118.495 113.955 118.675 ;
        RECT 111.065 117.675 111.460 117.845 ;
        RECT 111.630 117.715 112.095 118.105 ;
        RECT 112.265 118.325 113.955 118.495 ;
        RECT 111.290 117.545 111.460 117.675 ;
        RECT 112.265 117.545 112.435 118.325 ;
        RECT 114.125 118.155 114.295 118.845 ;
        RECT 112.795 117.985 114.295 118.155 ;
        RECT 114.485 118.185 114.695 118.975 ;
        RECT 114.865 118.355 115.215 118.975 ;
        RECT 115.385 118.365 115.555 119.145 ;
        RECT 116.085 118.985 116.255 119.215 ;
        RECT 115.725 118.815 116.255 118.985 ;
        RECT 115.725 118.535 115.945 118.815 ;
        RECT 116.425 118.645 116.665 119.045 ;
        RECT 115.385 118.195 115.790 118.365 ;
        RECT 116.125 118.275 116.665 118.645 ;
        RECT 116.835 118.860 117.155 119.215 ;
        RECT 117.400 119.135 117.705 119.595 ;
        RECT 117.875 118.885 118.130 119.415 ;
        RECT 116.835 118.685 117.160 118.860 ;
        RECT 116.835 118.385 117.750 118.685 ;
        RECT 117.010 118.355 117.750 118.385 ;
        RECT 114.485 118.025 115.160 118.185 ;
        RECT 115.620 118.105 115.790 118.195 ;
        RECT 114.485 118.015 115.450 118.025 ;
        RECT 114.125 117.845 114.295 117.985 ;
        RECT 110.870 117.045 111.120 117.505 ;
        RECT 111.290 117.215 111.540 117.545 ;
        RECT 111.755 117.215 112.435 117.545 ;
        RECT 112.605 117.645 113.680 117.815 ;
        RECT 114.125 117.675 114.685 117.845 ;
        RECT 114.990 117.725 115.450 118.015 ;
        RECT 115.620 117.935 116.840 118.105 ;
        RECT 112.605 117.305 112.775 117.645 ;
        RECT 113.010 117.045 113.340 117.475 ;
        RECT 113.510 117.305 113.680 117.645 ;
        RECT 113.975 117.045 114.345 117.505 ;
        RECT 114.515 117.215 114.685 117.675 ;
        RECT 115.620 117.555 115.790 117.935 ;
        RECT 117.010 117.765 117.180 118.355 ;
        RECT 117.920 118.235 118.130 118.885 ;
        RECT 118.305 118.825 121.815 119.595 ;
        RECT 122.445 118.845 123.655 119.595 ;
        RECT 118.305 118.305 119.955 118.825 ;
        RECT 114.920 117.215 115.790 117.555 ;
        RECT 116.380 117.595 117.180 117.765 ;
        RECT 115.960 117.045 116.210 117.505 ;
        RECT 116.380 117.305 116.550 117.595 ;
        RECT 116.730 117.045 117.060 117.425 ;
        RECT 117.400 117.045 117.705 118.185 ;
        RECT 117.875 117.355 118.130 118.235 ;
        RECT 120.125 118.135 121.815 118.655 ;
        RECT 118.305 117.045 121.815 118.135 ;
        RECT 122.445 118.135 122.965 118.675 ;
        RECT 123.135 118.305 123.655 118.845 ;
        RECT 122.445 117.045 123.655 118.135 ;
        RECT 5.520 116.875 123.740 117.045 ;
        RECT 5.605 115.785 6.815 116.875 ;
        RECT 6.985 115.785 9.575 116.875 ;
        RECT 5.605 115.075 6.125 115.615 ;
        RECT 6.295 115.245 6.815 115.785 ;
        RECT 6.985 115.095 8.195 115.615 ;
        RECT 8.365 115.265 9.575 115.785 ;
        RECT 10.205 115.800 10.475 116.705 ;
        RECT 10.645 116.115 10.975 116.875 ;
        RECT 11.155 115.945 11.325 116.705 ;
        RECT 5.605 114.325 6.815 115.075 ;
        RECT 6.985 114.325 9.575 115.095 ;
        RECT 10.205 115.000 10.375 115.800 ;
        RECT 10.660 115.775 11.325 115.945 ;
        RECT 11.585 115.800 11.855 116.705 ;
        RECT 12.025 116.115 12.355 116.875 ;
        RECT 12.535 115.945 12.705 116.705 ;
        RECT 12.965 116.440 18.310 116.875 ;
        RECT 10.660 115.630 10.830 115.775 ;
        RECT 10.545 115.300 10.830 115.630 ;
        RECT 10.660 115.045 10.830 115.300 ;
        RECT 11.065 115.225 11.395 115.595 ;
        RECT 10.205 114.495 10.465 115.000 ;
        RECT 10.660 114.875 11.325 115.045 ;
        RECT 10.645 114.325 10.975 114.705 ;
        RECT 11.155 114.495 11.325 114.875 ;
        RECT 11.585 115.000 11.755 115.800 ;
        RECT 12.040 115.775 12.705 115.945 ;
        RECT 12.040 115.630 12.210 115.775 ;
        RECT 11.925 115.300 12.210 115.630 ;
        RECT 12.040 115.045 12.210 115.300 ;
        RECT 12.445 115.225 12.775 115.595 ;
        RECT 11.585 114.495 11.845 115.000 ;
        RECT 12.040 114.875 12.705 115.045 ;
        RECT 12.025 114.325 12.355 114.705 ;
        RECT 12.535 114.495 12.705 114.875 ;
        RECT 14.550 114.870 14.890 115.700 ;
        RECT 16.370 115.190 16.720 116.440 ;
        RECT 18.485 115.710 18.775 116.875 ;
        RECT 18.945 115.785 22.455 116.875 ;
        RECT 22.625 115.785 23.835 116.875 ;
        RECT 18.945 115.095 20.595 115.615 ;
        RECT 20.765 115.265 22.455 115.785 ;
        RECT 12.965 114.325 18.310 114.870 ;
        RECT 18.485 114.325 18.775 115.050 ;
        RECT 18.945 114.325 22.455 115.095 ;
        RECT 22.625 115.075 23.145 115.615 ;
        RECT 23.315 115.245 23.835 115.785 ;
        RECT 24.005 115.800 24.275 116.705 ;
        RECT 24.445 116.115 24.775 116.875 ;
        RECT 24.955 115.945 25.125 116.705 ;
        RECT 25.385 116.440 30.730 116.875 ;
        RECT 22.625 114.325 23.835 115.075 ;
        RECT 24.005 115.000 24.175 115.800 ;
        RECT 24.460 115.775 25.125 115.945 ;
        RECT 24.460 115.630 24.630 115.775 ;
        RECT 24.345 115.300 24.630 115.630 ;
        RECT 24.460 115.045 24.630 115.300 ;
        RECT 24.865 115.225 25.195 115.595 ;
        RECT 24.005 114.495 24.265 115.000 ;
        RECT 24.460 114.875 25.125 115.045 ;
        RECT 24.445 114.325 24.775 114.705 ;
        RECT 24.955 114.495 25.125 114.875 ;
        RECT 26.970 114.870 27.310 115.700 ;
        RECT 28.790 115.190 29.140 116.440 ;
        RECT 30.905 115.785 33.495 116.875 ;
        RECT 30.905 115.095 32.115 115.615 ;
        RECT 32.285 115.265 33.495 115.785 ;
        RECT 33.665 115.800 33.935 116.705 ;
        RECT 34.105 116.115 34.435 116.875 ;
        RECT 34.615 115.945 34.785 116.705 ;
        RECT 35.045 116.440 40.390 116.875 ;
        RECT 25.385 114.325 30.730 114.870 ;
        RECT 30.905 114.325 33.495 115.095 ;
        RECT 33.665 115.000 33.835 115.800 ;
        RECT 34.120 115.775 34.785 115.945 ;
        RECT 34.120 115.630 34.290 115.775 ;
        RECT 34.005 115.300 34.290 115.630 ;
        RECT 34.120 115.045 34.290 115.300 ;
        RECT 34.525 115.225 34.855 115.595 ;
        RECT 33.665 114.495 33.925 115.000 ;
        RECT 34.120 114.875 34.785 115.045 ;
        RECT 34.105 114.325 34.435 114.705 ;
        RECT 34.615 114.495 34.785 114.875 ;
        RECT 36.630 114.870 36.970 115.700 ;
        RECT 38.450 115.190 38.800 116.440 ;
        RECT 40.565 115.785 44.075 116.875 ;
        RECT 40.565 115.095 42.215 115.615 ;
        RECT 42.385 115.265 44.075 115.785 ;
        RECT 44.245 115.710 44.535 116.875 ;
        RECT 44.705 116.440 50.050 116.875 ;
        RECT 50.225 116.440 55.570 116.875 ;
        RECT 55.745 116.440 61.090 116.875 ;
        RECT 61.265 116.440 66.610 116.875 ;
        RECT 35.045 114.325 40.390 114.870 ;
        RECT 40.565 114.325 44.075 115.095 ;
        RECT 44.245 114.325 44.535 115.050 ;
        RECT 46.290 114.870 46.630 115.700 ;
        RECT 48.110 115.190 48.460 116.440 ;
        RECT 51.810 114.870 52.150 115.700 ;
        RECT 53.630 115.190 53.980 116.440 ;
        RECT 57.330 114.870 57.670 115.700 ;
        RECT 59.150 115.190 59.500 116.440 ;
        RECT 62.850 114.870 63.190 115.700 ;
        RECT 64.670 115.190 65.020 116.440 ;
        RECT 66.785 115.785 68.455 116.875 ;
        RECT 66.785 115.095 67.535 115.615 ;
        RECT 67.705 115.265 68.455 115.785 ;
        RECT 68.625 115.800 68.895 116.705 ;
        RECT 69.065 116.115 69.395 116.875 ;
        RECT 69.575 115.945 69.745 116.705 ;
        RECT 44.705 114.325 50.050 114.870 ;
        RECT 50.225 114.325 55.570 114.870 ;
        RECT 55.745 114.325 61.090 114.870 ;
        RECT 61.265 114.325 66.610 114.870 ;
        RECT 66.785 114.325 68.455 115.095 ;
        RECT 68.625 115.000 68.795 115.800 ;
        RECT 69.080 115.775 69.745 115.945 ;
        RECT 69.080 115.630 69.250 115.775 ;
        RECT 70.005 115.710 70.295 116.875 ;
        RECT 71.385 115.800 71.655 116.705 ;
        RECT 71.825 116.115 72.155 116.875 ;
        RECT 72.335 115.945 72.505 116.705 ;
        RECT 68.965 115.300 69.250 115.630 ;
        RECT 69.080 115.045 69.250 115.300 ;
        RECT 69.485 115.225 69.815 115.595 ;
        RECT 68.625 114.495 68.885 115.000 ;
        RECT 69.080 114.875 69.745 115.045 ;
        RECT 69.065 114.325 69.395 114.705 ;
        RECT 69.575 114.495 69.745 114.875 ;
        RECT 70.005 114.325 70.295 115.050 ;
        RECT 71.385 115.000 71.555 115.800 ;
        RECT 71.840 115.775 72.505 115.945 ;
        RECT 72.765 115.785 75.355 116.875 ;
        RECT 76.075 116.205 76.245 116.705 ;
        RECT 76.415 116.375 76.745 116.875 ;
        RECT 76.075 116.035 76.740 116.205 ;
        RECT 71.840 115.630 72.010 115.775 ;
        RECT 71.725 115.300 72.010 115.630 ;
        RECT 71.840 115.045 72.010 115.300 ;
        RECT 72.245 115.225 72.575 115.595 ;
        RECT 72.765 115.095 73.975 115.615 ;
        RECT 74.145 115.265 75.355 115.785 ;
        RECT 75.990 115.215 76.340 115.865 ;
        RECT 71.385 114.495 71.645 115.000 ;
        RECT 71.840 114.875 72.505 115.045 ;
        RECT 71.825 114.325 72.155 114.705 ;
        RECT 72.335 114.495 72.505 114.875 ;
        RECT 72.765 114.325 75.355 115.095 ;
        RECT 76.510 115.045 76.740 116.035 ;
        RECT 76.075 114.875 76.740 115.045 ;
        RECT 76.075 114.585 76.245 114.875 ;
        RECT 76.415 114.325 76.745 114.705 ;
        RECT 76.915 114.585 77.140 116.705 ;
        RECT 77.355 116.375 77.685 116.875 ;
        RECT 77.855 116.205 78.025 116.705 ;
        RECT 78.260 116.490 79.090 116.660 ;
        RECT 79.330 116.495 79.710 116.875 ;
        RECT 77.330 116.035 78.025 116.205 ;
        RECT 77.330 115.065 77.500 116.035 ;
        RECT 77.670 115.245 78.080 115.865 ;
        RECT 78.250 115.815 78.750 116.195 ;
        RECT 77.330 114.875 78.025 115.065 ;
        RECT 78.250 114.945 78.470 115.815 ;
        RECT 78.920 115.645 79.090 116.490 ;
        RECT 79.890 116.325 80.060 116.615 ;
        RECT 80.230 116.495 80.560 116.875 ;
        RECT 81.030 116.405 81.660 116.655 ;
        RECT 81.840 116.495 82.260 116.875 ;
        RECT 81.490 116.325 81.660 116.405 ;
        RECT 82.460 116.325 82.700 116.615 ;
        RECT 79.260 116.075 80.630 116.325 ;
        RECT 79.260 115.815 79.510 116.075 ;
        RECT 80.020 115.645 80.270 115.805 ;
        RECT 78.920 115.475 80.270 115.645 ;
        RECT 78.920 115.435 79.340 115.475 ;
        RECT 78.650 114.885 79.000 115.255 ;
        RECT 77.355 114.325 77.685 114.705 ;
        RECT 77.855 114.545 78.025 114.875 ;
        RECT 79.170 114.705 79.340 115.435 ;
        RECT 80.440 115.305 80.630 116.075 ;
        RECT 79.510 114.975 79.920 115.305 ;
        RECT 80.210 114.965 80.630 115.305 ;
        RECT 80.800 115.895 81.320 116.205 ;
        RECT 81.490 116.155 82.700 116.325 ;
        RECT 82.930 116.185 83.260 116.875 ;
        RECT 80.800 115.135 80.970 115.895 ;
        RECT 81.140 115.305 81.320 115.715 ;
        RECT 81.490 115.645 81.660 116.155 ;
        RECT 83.430 116.005 83.600 116.615 ;
        RECT 83.870 116.155 84.200 116.665 ;
        RECT 83.430 115.985 83.750 116.005 ;
        RECT 81.830 115.815 83.750 115.985 ;
        RECT 81.490 115.475 83.390 115.645 ;
        RECT 81.720 115.135 82.050 115.255 ;
        RECT 80.800 114.965 82.050 115.135 ;
        RECT 78.325 114.505 79.340 114.705 ;
        RECT 79.510 114.325 79.920 114.765 ;
        RECT 80.210 114.535 80.460 114.965 ;
        RECT 80.660 114.325 80.980 114.785 ;
        RECT 82.220 114.715 82.390 115.475 ;
        RECT 83.060 115.415 83.390 115.475 ;
        RECT 82.580 115.245 82.910 115.305 ;
        RECT 82.580 114.975 83.240 115.245 ;
        RECT 83.560 114.920 83.750 115.815 ;
        RECT 81.540 114.545 82.390 114.715 ;
        RECT 82.590 114.325 83.250 114.805 ;
        RECT 83.430 114.590 83.750 114.920 ;
        RECT 83.950 115.565 84.200 116.155 ;
        RECT 84.380 116.075 84.665 116.875 ;
        RECT 84.845 115.895 85.100 116.565 ;
        RECT 85.645 116.440 90.990 116.875 ;
        RECT 83.950 115.235 84.750 115.565 ;
        RECT 83.950 114.585 84.200 115.235 ;
        RECT 84.920 115.035 85.100 115.895 ;
        RECT 84.845 114.835 85.100 115.035 ;
        RECT 87.230 114.870 87.570 115.700 ;
        RECT 89.050 115.190 89.400 116.440 ;
        RECT 91.165 115.785 94.675 116.875 ;
        RECT 91.165 115.095 92.815 115.615 ;
        RECT 92.985 115.265 94.675 115.785 ;
        RECT 95.765 115.710 96.055 116.875 ;
        RECT 96.225 116.440 101.570 116.875 ;
        RECT 101.745 116.440 107.090 116.875 ;
        RECT 107.265 116.440 112.610 116.875 ;
        RECT 84.380 114.325 84.665 114.785 ;
        RECT 84.845 114.665 85.185 114.835 ;
        RECT 84.845 114.505 85.100 114.665 ;
        RECT 85.645 114.325 90.990 114.870 ;
        RECT 91.165 114.325 94.675 115.095 ;
        RECT 95.765 114.325 96.055 115.050 ;
        RECT 97.810 114.870 98.150 115.700 ;
        RECT 99.630 115.190 99.980 116.440 ;
        RECT 103.330 114.870 103.670 115.700 ;
        RECT 105.150 115.190 105.500 116.440 ;
        RECT 108.850 114.870 109.190 115.700 ;
        RECT 110.670 115.190 111.020 116.440 ;
        RECT 113.745 115.735 113.975 116.875 ;
        RECT 114.145 115.725 114.475 116.705 ;
        RECT 114.645 115.735 114.855 116.875 ;
        RECT 115.085 116.440 120.430 116.875 ;
        RECT 113.725 115.315 114.055 115.565 ;
        RECT 96.225 114.325 101.570 114.870 ;
        RECT 101.745 114.325 107.090 114.870 ;
        RECT 107.265 114.325 112.610 114.870 ;
        RECT 113.745 114.325 113.975 115.145 ;
        RECT 114.225 115.125 114.475 115.725 ;
        RECT 114.145 114.495 114.475 115.125 ;
        RECT 114.645 114.325 114.855 115.145 ;
        RECT 116.670 114.870 117.010 115.700 ;
        RECT 118.490 115.190 118.840 116.440 ;
        RECT 121.525 115.710 121.815 116.875 ;
        RECT 122.445 115.785 123.655 116.875 ;
        RECT 122.445 115.245 122.965 115.785 ;
        RECT 123.135 115.075 123.655 115.615 ;
        RECT 115.085 114.325 120.430 114.870 ;
        RECT 121.525 114.325 121.815 115.050 ;
        RECT 122.445 114.325 123.655 115.075 ;
        RECT 5.520 114.155 123.740 114.325 ;
        RECT 5.605 113.405 6.815 114.155 ;
        RECT 5.605 112.865 6.125 113.405 ;
        RECT 6.985 113.385 10.495 114.155 ;
        RECT 10.755 113.605 10.925 113.895 ;
        RECT 11.095 113.775 11.425 114.155 ;
        RECT 10.755 113.435 11.420 113.605 ;
        RECT 6.295 112.695 6.815 113.235 ;
        RECT 6.985 112.865 8.635 113.385 ;
        RECT 8.805 112.695 10.495 113.215 ;
        RECT 5.605 111.605 6.815 112.695 ;
        RECT 6.985 111.605 10.495 112.695 ;
        RECT 10.670 112.615 11.020 113.265 ;
        RECT 11.190 112.445 11.420 113.435 ;
        RECT 10.755 112.275 11.420 112.445 ;
        RECT 10.755 111.775 10.925 112.275 ;
        RECT 11.095 111.605 11.425 112.105 ;
        RECT 11.595 111.775 11.820 113.895 ;
        RECT 12.035 113.775 12.365 114.155 ;
        RECT 12.535 113.605 12.705 113.935 ;
        RECT 13.005 113.775 14.020 113.975 ;
        RECT 12.010 113.415 12.705 113.605 ;
        RECT 12.010 112.445 12.180 113.415 ;
        RECT 12.350 112.615 12.760 113.235 ;
        RECT 12.930 112.665 13.150 113.535 ;
        RECT 13.330 113.225 13.680 113.595 ;
        RECT 13.850 113.045 14.020 113.775 ;
        RECT 14.190 113.715 14.600 114.155 ;
        RECT 14.890 113.515 15.140 113.945 ;
        RECT 15.340 113.695 15.660 114.155 ;
        RECT 16.220 113.765 17.070 113.935 ;
        RECT 14.190 113.175 14.600 113.505 ;
        RECT 14.890 113.175 15.310 113.515 ;
        RECT 13.600 113.005 14.020 113.045 ;
        RECT 13.600 112.835 14.950 113.005 ;
        RECT 12.010 112.275 12.705 112.445 ;
        RECT 12.930 112.285 13.430 112.665 ;
        RECT 12.035 111.605 12.365 112.105 ;
        RECT 12.535 111.775 12.705 112.275 ;
        RECT 13.600 111.990 13.770 112.835 ;
        RECT 14.700 112.675 14.950 112.835 ;
        RECT 13.940 112.405 14.190 112.665 ;
        RECT 15.120 112.405 15.310 113.175 ;
        RECT 13.940 112.155 15.310 112.405 ;
        RECT 15.480 113.345 16.730 113.515 ;
        RECT 15.480 112.585 15.650 113.345 ;
        RECT 16.400 113.225 16.730 113.345 ;
        RECT 15.820 112.765 16.000 113.175 ;
        RECT 16.900 113.005 17.070 113.765 ;
        RECT 17.270 113.675 17.930 114.155 ;
        RECT 18.110 113.560 18.430 113.890 ;
        RECT 17.260 113.235 17.920 113.505 ;
        RECT 17.260 113.175 17.590 113.235 ;
        RECT 17.740 113.005 18.070 113.065 ;
        RECT 16.170 112.835 18.070 113.005 ;
        RECT 15.480 112.275 16.000 112.585 ;
        RECT 16.170 112.325 16.340 112.835 ;
        RECT 18.240 112.665 18.430 113.560 ;
        RECT 16.510 112.495 18.430 112.665 ;
        RECT 18.110 112.475 18.430 112.495 ;
        RECT 18.630 113.245 18.880 113.895 ;
        RECT 19.060 113.695 19.345 114.155 ;
        RECT 19.525 113.445 19.780 113.975 ;
        RECT 20.325 113.610 25.670 114.155 ;
        RECT 18.630 112.915 19.430 113.245 ;
        RECT 16.170 112.155 17.380 112.325 ;
        RECT 12.940 111.820 13.770 111.990 ;
        RECT 14.010 111.605 14.390 111.985 ;
        RECT 14.570 111.865 14.740 112.155 ;
        RECT 16.170 112.075 16.340 112.155 ;
        RECT 14.910 111.605 15.240 111.985 ;
        RECT 15.710 111.825 16.340 112.075 ;
        RECT 16.520 111.605 16.940 111.985 ;
        RECT 17.140 111.865 17.380 112.155 ;
        RECT 17.610 111.605 17.940 112.295 ;
        RECT 18.110 111.865 18.280 112.475 ;
        RECT 18.630 112.325 18.880 112.915 ;
        RECT 19.600 112.585 19.780 113.445 ;
        RECT 21.910 112.780 22.250 113.610 ;
        RECT 25.845 113.385 29.355 114.155 ;
        RECT 29.525 113.480 29.785 113.985 ;
        RECT 29.965 113.775 30.295 114.155 ;
        RECT 30.475 113.605 30.645 113.985 ;
        RECT 18.550 111.815 18.880 112.325 ;
        RECT 19.060 111.605 19.345 112.405 ;
        RECT 19.525 112.115 19.780 112.585 ;
        RECT 19.525 111.945 19.865 112.115 ;
        RECT 23.730 112.040 24.080 113.290 ;
        RECT 25.845 112.865 27.495 113.385 ;
        RECT 27.665 112.695 29.355 113.215 ;
        RECT 19.525 111.915 19.780 111.945 ;
        RECT 20.325 111.605 25.670 112.040 ;
        RECT 25.845 111.605 29.355 112.695 ;
        RECT 29.525 112.680 29.695 113.480 ;
        RECT 29.980 113.435 30.645 113.605 ;
        RECT 29.980 113.180 30.150 113.435 ;
        RECT 31.365 113.430 31.655 114.155 ;
        RECT 31.885 113.335 32.095 114.155 ;
        RECT 32.265 113.355 32.595 113.985 ;
        RECT 29.865 112.850 30.150 113.180 ;
        RECT 30.385 112.885 30.715 113.255 ;
        RECT 29.980 112.705 30.150 112.850 ;
        RECT 29.525 111.775 29.795 112.680 ;
        RECT 29.980 112.535 30.645 112.705 ;
        RECT 29.965 111.605 30.295 112.365 ;
        RECT 30.475 111.775 30.645 112.535 ;
        RECT 31.365 111.605 31.655 112.770 ;
        RECT 32.265 112.755 32.515 113.355 ;
        RECT 32.765 113.335 32.995 114.155 ;
        RECT 33.205 113.610 38.550 114.155 ;
        RECT 32.685 112.915 33.015 113.165 ;
        RECT 34.790 112.780 35.130 113.610 ;
        RECT 39.735 113.605 39.905 113.895 ;
        RECT 40.075 113.775 40.405 114.155 ;
        RECT 39.735 113.435 40.400 113.605 ;
        RECT 31.885 111.605 32.095 112.745 ;
        RECT 32.265 111.775 32.595 112.755 ;
        RECT 32.765 111.605 32.995 112.745 ;
        RECT 36.610 112.040 36.960 113.290 ;
        RECT 39.650 112.615 40.000 113.265 ;
        RECT 40.170 112.445 40.400 113.435 ;
        RECT 39.735 112.275 40.400 112.445 ;
        RECT 33.205 111.605 38.550 112.040 ;
        RECT 39.735 111.775 39.905 112.275 ;
        RECT 40.075 111.605 40.405 112.105 ;
        RECT 40.575 111.775 40.800 113.895 ;
        RECT 41.015 113.775 41.345 114.155 ;
        RECT 41.515 113.605 41.685 113.935 ;
        RECT 41.985 113.775 43.000 113.975 ;
        RECT 40.990 113.415 41.685 113.605 ;
        RECT 40.990 112.445 41.160 113.415 ;
        RECT 41.330 112.615 41.740 113.235 ;
        RECT 41.910 112.665 42.130 113.535 ;
        RECT 42.310 113.225 42.660 113.595 ;
        RECT 42.830 113.045 43.000 113.775 ;
        RECT 43.170 113.715 43.580 114.155 ;
        RECT 43.870 113.515 44.120 113.945 ;
        RECT 44.320 113.695 44.640 114.155 ;
        RECT 45.200 113.765 46.050 113.935 ;
        RECT 43.170 113.175 43.580 113.505 ;
        RECT 43.870 113.175 44.290 113.515 ;
        RECT 42.580 113.005 43.000 113.045 ;
        RECT 42.580 112.835 43.930 113.005 ;
        RECT 40.990 112.275 41.685 112.445 ;
        RECT 41.910 112.285 42.410 112.665 ;
        RECT 41.015 111.605 41.345 112.105 ;
        RECT 41.515 111.775 41.685 112.275 ;
        RECT 42.580 111.990 42.750 112.835 ;
        RECT 43.680 112.675 43.930 112.835 ;
        RECT 42.920 112.405 43.170 112.665 ;
        RECT 44.100 112.405 44.290 113.175 ;
        RECT 42.920 112.155 44.290 112.405 ;
        RECT 44.460 113.345 45.710 113.515 ;
        RECT 44.460 112.585 44.630 113.345 ;
        RECT 45.380 113.225 45.710 113.345 ;
        RECT 44.800 112.765 44.980 113.175 ;
        RECT 45.880 113.005 46.050 113.765 ;
        RECT 46.250 113.675 46.910 114.155 ;
        RECT 47.090 113.560 47.410 113.890 ;
        RECT 46.240 113.235 46.900 113.505 ;
        RECT 46.240 113.175 46.570 113.235 ;
        RECT 46.720 113.005 47.050 113.065 ;
        RECT 45.150 112.835 47.050 113.005 ;
        RECT 44.460 112.275 44.980 112.585 ;
        RECT 45.150 112.325 45.320 112.835 ;
        RECT 47.220 112.665 47.410 113.560 ;
        RECT 45.490 112.495 47.410 112.665 ;
        RECT 47.090 112.475 47.410 112.495 ;
        RECT 47.610 113.245 47.860 113.895 ;
        RECT 48.040 113.695 48.325 114.155 ;
        RECT 48.505 113.445 48.760 113.975 ;
        RECT 49.305 113.610 54.650 114.155 ;
        RECT 47.610 112.915 48.410 113.245 ;
        RECT 45.150 112.155 46.360 112.325 ;
        RECT 41.920 111.820 42.750 111.990 ;
        RECT 42.990 111.605 43.370 111.985 ;
        RECT 43.550 111.865 43.720 112.155 ;
        RECT 45.150 112.075 45.320 112.155 ;
        RECT 43.890 111.605 44.220 111.985 ;
        RECT 44.690 111.825 45.320 112.075 ;
        RECT 45.500 111.605 45.920 111.985 ;
        RECT 46.120 111.865 46.360 112.155 ;
        RECT 46.590 111.605 46.920 112.295 ;
        RECT 47.090 111.865 47.260 112.475 ;
        RECT 47.610 112.325 47.860 112.915 ;
        RECT 48.580 112.585 48.760 113.445 ;
        RECT 50.890 112.780 51.230 113.610 ;
        RECT 54.825 113.385 56.495 114.155 ;
        RECT 57.125 113.430 57.415 114.155 ;
        RECT 57.960 113.445 58.215 113.975 ;
        RECT 58.395 113.695 58.680 114.155 ;
        RECT 47.530 111.815 47.860 112.325 ;
        RECT 48.040 111.605 48.325 112.405 ;
        RECT 48.505 112.115 48.760 112.585 ;
        RECT 48.505 111.945 48.845 112.115 ;
        RECT 52.710 112.040 53.060 113.290 ;
        RECT 54.825 112.865 55.575 113.385 ;
        RECT 55.745 112.695 56.495 113.215 ;
        RECT 48.505 111.915 48.760 111.945 ;
        RECT 49.305 111.605 54.650 112.040 ;
        RECT 54.825 111.605 56.495 112.695 ;
        RECT 57.125 111.605 57.415 112.770 ;
        RECT 57.960 112.585 58.140 113.445 ;
        RECT 58.860 113.245 59.110 113.895 ;
        RECT 58.310 112.915 59.110 113.245 ;
        RECT 57.960 112.115 58.215 112.585 ;
        RECT 57.875 111.945 58.215 112.115 ;
        RECT 57.960 111.915 58.215 111.945 ;
        RECT 58.395 111.605 58.680 112.405 ;
        RECT 58.860 112.325 59.110 112.915 ;
        RECT 59.310 113.560 59.630 113.890 ;
        RECT 59.810 113.675 60.470 114.155 ;
        RECT 60.670 113.765 61.520 113.935 ;
        RECT 59.310 112.665 59.500 113.560 ;
        RECT 59.820 113.235 60.480 113.505 ;
        RECT 60.150 113.175 60.480 113.235 ;
        RECT 59.670 113.005 60.000 113.065 ;
        RECT 60.670 113.005 60.840 113.765 ;
        RECT 62.080 113.695 62.400 114.155 ;
        RECT 62.600 113.515 62.850 113.945 ;
        RECT 63.140 113.715 63.550 114.155 ;
        RECT 63.720 113.775 64.735 113.975 ;
        RECT 61.010 113.345 62.260 113.515 ;
        RECT 61.010 113.225 61.340 113.345 ;
        RECT 59.670 112.835 61.570 113.005 ;
        RECT 59.310 112.495 61.230 112.665 ;
        RECT 59.310 112.475 59.630 112.495 ;
        RECT 58.860 111.815 59.190 112.325 ;
        RECT 59.460 111.865 59.630 112.475 ;
        RECT 61.400 112.325 61.570 112.835 ;
        RECT 61.740 112.765 61.920 113.175 ;
        RECT 62.090 112.585 62.260 113.345 ;
        RECT 59.800 111.605 60.130 112.295 ;
        RECT 60.360 112.155 61.570 112.325 ;
        RECT 61.740 112.275 62.260 112.585 ;
        RECT 62.430 113.175 62.850 113.515 ;
        RECT 63.140 113.175 63.550 113.505 ;
        RECT 62.430 112.405 62.620 113.175 ;
        RECT 63.720 113.045 63.890 113.775 ;
        RECT 65.035 113.605 65.205 113.935 ;
        RECT 65.375 113.775 65.705 114.155 ;
        RECT 64.060 113.225 64.410 113.595 ;
        RECT 63.720 113.005 64.140 113.045 ;
        RECT 62.790 112.835 64.140 113.005 ;
        RECT 62.790 112.675 63.040 112.835 ;
        RECT 63.550 112.405 63.800 112.665 ;
        RECT 62.430 112.155 63.800 112.405 ;
        RECT 60.360 111.865 60.600 112.155 ;
        RECT 61.400 112.075 61.570 112.155 ;
        RECT 60.800 111.605 61.220 111.985 ;
        RECT 61.400 111.825 62.030 112.075 ;
        RECT 62.500 111.605 62.830 111.985 ;
        RECT 63.000 111.865 63.170 112.155 ;
        RECT 63.970 111.990 64.140 112.835 ;
        RECT 64.590 112.665 64.810 113.535 ;
        RECT 65.035 113.415 65.730 113.605 ;
        RECT 64.310 112.285 64.810 112.665 ;
        RECT 64.980 112.615 65.390 113.235 ;
        RECT 65.560 112.445 65.730 113.415 ;
        RECT 65.035 112.275 65.730 112.445 ;
        RECT 63.350 111.605 63.730 111.985 ;
        RECT 63.970 111.820 64.800 111.990 ;
        RECT 65.035 111.775 65.205 112.275 ;
        RECT 65.375 111.605 65.705 112.105 ;
        RECT 65.920 111.775 66.145 113.895 ;
        RECT 66.315 113.775 66.645 114.155 ;
        RECT 66.815 113.605 66.985 113.895 ;
        RECT 67.245 113.610 72.590 114.155 ;
        RECT 66.320 113.435 66.985 113.605 ;
        RECT 66.320 112.445 66.550 113.435 ;
        RECT 66.720 112.615 67.070 113.265 ;
        RECT 68.830 112.780 69.170 113.610 ;
        RECT 72.765 113.385 76.275 114.155 ;
        RECT 76.445 113.405 77.655 114.155 ;
        RECT 77.825 113.480 78.085 113.985 ;
        RECT 78.265 113.775 78.595 114.155 ;
        RECT 78.775 113.605 78.945 113.985 ;
        RECT 66.320 112.275 66.985 112.445 ;
        RECT 66.315 111.605 66.645 112.105 ;
        RECT 66.815 111.775 66.985 112.275 ;
        RECT 70.650 112.040 71.000 113.290 ;
        RECT 72.765 112.865 74.415 113.385 ;
        RECT 74.585 112.695 76.275 113.215 ;
        RECT 76.445 112.865 76.965 113.405 ;
        RECT 77.135 112.695 77.655 113.235 ;
        RECT 67.245 111.605 72.590 112.040 ;
        RECT 72.765 111.605 76.275 112.695 ;
        RECT 76.445 111.605 77.655 112.695 ;
        RECT 77.825 112.680 77.995 113.480 ;
        RECT 78.280 113.435 78.945 113.605 ;
        RECT 78.280 113.180 78.450 113.435 ;
        RECT 79.205 113.405 80.415 114.155 ;
        RECT 78.165 112.850 78.450 113.180 ;
        RECT 78.685 112.885 79.015 113.255 ;
        RECT 79.205 112.865 79.725 113.405 ;
        RECT 80.625 113.335 80.855 114.155 ;
        RECT 81.025 113.355 81.355 113.985 ;
        RECT 78.280 112.705 78.450 112.850 ;
        RECT 77.825 111.775 78.095 112.680 ;
        RECT 78.280 112.535 78.945 112.705 ;
        RECT 79.895 112.695 80.415 113.235 ;
        RECT 80.605 112.915 80.935 113.165 ;
        RECT 81.105 112.755 81.355 113.355 ;
        RECT 81.525 113.335 81.735 114.155 ;
        RECT 82.885 113.430 83.175 114.155 ;
        RECT 83.350 113.415 83.605 113.985 ;
        RECT 83.775 113.755 84.105 114.155 ;
        RECT 84.530 113.620 85.060 113.985 ;
        RECT 85.250 113.815 85.525 113.985 ;
        RECT 85.245 113.645 85.525 113.815 ;
        RECT 84.530 113.585 84.705 113.620 ;
        RECT 83.775 113.415 84.705 113.585 ;
        RECT 78.265 111.605 78.595 112.365 ;
        RECT 78.775 111.775 78.945 112.535 ;
        RECT 79.205 111.605 80.415 112.695 ;
        RECT 80.625 111.605 80.855 112.745 ;
        RECT 81.025 111.775 81.355 112.755 ;
        RECT 81.525 111.605 81.735 112.745 ;
        RECT 82.885 111.605 83.175 112.770 ;
        RECT 83.350 112.745 83.520 113.415 ;
        RECT 83.775 113.245 83.945 113.415 ;
        RECT 83.690 112.915 83.945 113.245 ;
        RECT 84.170 112.915 84.365 113.245 ;
        RECT 83.350 111.775 83.685 112.745 ;
        RECT 83.855 111.605 84.025 112.745 ;
        RECT 84.195 111.945 84.365 112.915 ;
        RECT 84.535 112.285 84.705 113.415 ;
        RECT 84.875 112.625 85.045 113.425 ;
        RECT 85.250 112.825 85.525 113.645 ;
        RECT 85.695 112.625 85.885 113.985 ;
        RECT 86.065 113.620 86.575 114.155 ;
        RECT 86.795 113.345 87.040 113.950 ;
        RECT 87.485 113.480 87.745 113.985 ;
        RECT 87.925 113.775 88.255 114.155 ;
        RECT 88.435 113.605 88.605 113.985 ;
        RECT 86.085 113.175 87.315 113.345 ;
        RECT 84.875 112.455 85.885 112.625 ;
        RECT 86.055 112.610 86.805 112.800 ;
        RECT 84.535 112.115 85.660 112.285 ;
        RECT 86.055 111.945 86.225 112.610 ;
        RECT 86.975 112.365 87.315 113.175 ;
        RECT 84.195 111.775 86.225 111.945 ;
        RECT 86.395 111.605 86.565 112.365 ;
        RECT 86.800 111.955 87.315 112.365 ;
        RECT 87.485 112.680 87.655 113.480 ;
        RECT 87.940 113.435 88.605 113.605 ;
        RECT 87.940 113.180 88.110 113.435 ;
        RECT 88.925 113.335 89.135 114.155 ;
        RECT 89.305 113.355 89.635 113.985 ;
        RECT 87.825 112.850 88.110 113.180 ;
        RECT 88.345 112.885 88.675 113.255 ;
        RECT 87.940 112.705 88.110 112.850 ;
        RECT 89.305 112.755 89.555 113.355 ;
        RECT 89.805 113.335 90.035 114.155 ;
        RECT 90.245 113.385 91.915 114.155 ;
        RECT 92.635 113.605 92.805 113.985 ;
        RECT 92.985 113.775 93.315 114.155 ;
        RECT 92.635 113.435 93.300 113.605 ;
        RECT 93.495 113.480 93.755 113.985 ;
        RECT 89.725 112.915 90.055 113.165 ;
        RECT 90.245 112.865 90.995 113.385 ;
        RECT 87.485 111.775 87.755 112.680 ;
        RECT 87.940 112.535 88.605 112.705 ;
        RECT 87.925 111.605 88.255 112.365 ;
        RECT 88.435 111.775 88.605 112.535 ;
        RECT 88.925 111.605 89.135 112.745 ;
        RECT 89.305 111.775 89.635 112.755 ;
        RECT 89.805 111.605 90.035 112.745 ;
        RECT 91.165 112.695 91.915 113.215 ;
        RECT 92.565 112.885 92.895 113.255 ;
        RECT 93.130 113.180 93.300 113.435 ;
        RECT 93.130 112.850 93.415 113.180 ;
        RECT 93.130 112.705 93.300 112.850 ;
        RECT 90.245 111.605 91.915 112.695 ;
        RECT 92.635 112.535 93.300 112.705 ;
        RECT 93.585 112.680 93.755 113.480 ;
        RECT 93.965 113.335 94.195 114.155 ;
        RECT 94.365 113.355 94.695 113.985 ;
        RECT 93.945 112.915 94.275 113.165 ;
        RECT 94.445 112.755 94.695 113.355 ;
        RECT 94.865 113.335 95.075 114.155 ;
        RECT 95.395 113.605 95.565 113.895 ;
        RECT 95.735 113.775 96.065 114.155 ;
        RECT 95.395 113.435 96.060 113.605 ;
        RECT 92.635 111.775 92.805 112.535 ;
        RECT 92.985 111.605 93.315 112.365 ;
        RECT 93.485 111.775 93.755 112.680 ;
        RECT 93.965 111.605 94.195 112.745 ;
        RECT 94.365 111.775 94.695 112.755 ;
        RECT 94.865 111.605 95.075 112.745 ;
        RECT 95.310 112.615 95.660 113.265 ;
        RECT 95.830 112.445 96.060 113.435 ;
        RECT 95.395 112.275 96.060 112.445 ;
        RECT 95.395 111.775 95.565 112.275 ;
        RECT 95.735 111.605 96.065 112.105 ;
        RECT 96.235 111.775 96.460 113.895 ;
        RECT 96.675 113.775 97.005 114.155 ;
        RECT 97.175 113.605 97.345 113.935 ;
        RECT 97.645 113.775 98.660 113.975 ;
        RECT 96.650 113.415 97.345 113.605 ;
        RECT 96.650 112.445 96.820 113.415 ;
        RECT 96.990 112.615 97.400 113.235 ;
        RECT 97.570 112.665 97.790 113.535 ;
        RECT 97.970 113.225 98.320 113.595 ;
        RECT 98.490 113.045 98.660 113.775 ;
        RECT 98.830 113.715 99.240 114.155 ;
        RECT 99.530 113.515 99.780 113.945 ;
        RECT 99.980 113.695 100.300 114.155 ;
        RECT 100.860 113.765 101.710 113.935 ;
        RECT 98.830 113.175 99.240 113.505 ;
        RECT 99.530 113.175 99.950 113.515 ;
        RECT 98.240 113.005 98.660 113.045 ;
        RECT 98.240 112.835 99.590 113.005 ;
        RECT 96.650 112.275 97.345 112.445 ;
        RECT 97.570 112.285 98.070 112.665 ;
        RECT 96.675 111.605 97.005 112.105 ;
        RECT 97.175 111.775 97.345 112.275 ;
        RECT 98.240 111.990 98.410 112.835 ;
        RECT 99.340 112.675 99.590 112.835 ;
        RECT 98.580 112.405 98.830 112.665 ;
        RECT 99.760 112.405 99.950 113.175 ;
        RECT 98.580 112.155 99.950 112.405 ;
        RECT 100.120 113.345 101.370 113.515 ;
        RECT 100.120 112.585 100.290 113.345 ;
        RECT 101.040 113.225 101.370 113.345 ;
        RECT 100.460 112.765 100.640 113.175 ;
        RECT 101.540 113.005 101.710 113.765 ;
        RECT 101.910 113.675 102.570 114.155 ;
        RECT 102.750 113.560 103.070 113.890 ;
        RECT 101.900 113.235 102.560 113.505 ;
        RECT 101.900 113.175 102.230 113.235 ;
        RECT 102.380 113.005 102.710 113.065 ;
        RECT 100.810 112.835 102.710 113.005 ;
        RECT 100.120 112.275 100.640 112.585 ;
        RECT 100.810 112.325 100.980 112.835 ;
        RECT 102.880 112.665 103.070 113.560 ;
        RECT 101.150 112.495 103.070 112.665 ;
        RECT 102.750 112.475 103.070 112.495 ;
        RECT 103.270 113.245 103.520 113.895 ;
        RECT 103.700 113.695 103.985 114.155 ;
        RECT 104.165 113.445 104.420 113.975 ;
        RECT 103.270 112.915 104.070 113.245 ;
        RECT 100.810 112.155 102.020 112.325 ;
        RECT 97.580 111.820 98.410 111.990 ;
        RECT 98.650 111.605 99.030 111.985 ;
        RECT 99.210 111.865 99.380 112.155 ;
        RECT 100.810 112.075 100.980 112.155 ;
        RECT 99.550 111.605 99.880 111.985 ;
        RECT 100.350 111.825 100.980 112.075 ;
        RECT 101.160 111.605 101.580 111.985 ;
        RECT 101.780 111.865 102.020 112.155 ;
        RECT 102.250 111.605 102.580 112.295 ;
        RECT 102.750 111.865 102.920 112.475 ;
        RECT 103.270 112.325 103.520 112.915 ;
        RECT 104.240 112.585 104.420 113.445 ;
        RECT 105.055 113.605 105.225 113.985 ;
        RECT 105.405 113.775 105.735 114.155 ;
        RECT 105.055 113.435 105.720 113.605 ;
        RECT 105.915 113.480 106.175 113.985 ;
        RECT 104.985 112.885 105.315 113.255 ;
        RECT 105.550 113.180 105.720 113.435 ;
        RECT 105.550 112.850 105.835 113.180 ;
        RECT 105.550 112.705 105.720 112.850 ;
        RECT 103.190 111.815 103.520 112.325 ;
        RECT 103.700 111.605 103.985 112.405 ;
        RECT 104.165 112.115 104.420 112.585 ;
        RECT 105.055 112.535 105.720 112.705 ;
        RECT 106.005 112.680 106.175 113.480 ;
        RECT 106.345 113.385 108.015 114.155 ;
        RECT 108.645 113.430 108.935 114.155 ;
        RECT 109.105 113.610 114.450 114.155 ;
        RECT 114.625 113.610 119.970 114.155 ;
        RECT 106.345 112.865 107.095 113.385 ;
        RECT 107.265 112.695 108.015 113.215 ;
        RECT 110.690 112.780 111.030 113.610 ;
        RECT 104.165 111.945 104.505 112.115 ;
        RECT 104.165 111.915 104.420 111.945 ;
        RECT 105.055 111.775 105.225 112.535 ;
        RECT 105.405 111.605 105.735 112.365 ;
        RECT 105.905 111.775 106.175 112.680 ;
        RECT 106.345 111.605 108.015 112.695 ;
        RECT 108.645 111.605 108.935 112.770 ;
        RECT 112.510 112.040 112.860 113.290 ;
        RECT 116.210 112.780 116.550 113.610 ;
        RECT 120.145 113.385 121.815 114.155 ;
        RECT 122.445 113.405 123.655 114.155 ;
        RECT 118.030 112.040 118.380 113.290 ;
        RECT 120.145 112.865 120.895 113.385 ;
        RECT 121.065 112.695 121.815 113.215 ;
        RECT 109.105 111.605 114.450 112.040 ;
        RECT 114.625 111.605 119.970 112.040 ;
        RECT 120.145 111.605 121.815 112.695 ;
        RECT 122.445 112.695 122.965 113.235 ;
        RECT 123.135 112.865 123.655 113.405 ;
        RECT 122.445 111.605 123.655 112.695 ;
        RECT 5.520 111.435 123.740 111.605 ;
        RECT 5.605 110.345 6.815 111.435 ;
        RECT 6.985 111.000 12.330 111.435 ;
        RECT 5.605 109.635 6.125 110.175 ;
        RECT 6.295 109.805 6.815 110.345 ;
        RECT 5.605 108.885 6.815 109.635 ;
        RECT 8.570 109.430 8.910 110.260 ;
        RECT 10.390 109.750 10.740 111.000 ;
        RECT 12.505 110.345 14.175 111.435 ;
        RECT 12.505 109.655 13.255 110.175 ;
        RECT 13.425 109.825 14.175 110.345 ;
        RECT 14.345 110.360 14.615 111.265 ;
        RECT 14.785 110.675 15.115 111.435 ;
        RECT 15.295 110.505 15.465 111.265 ;
        RECT 6.985 108.885 12.330 109.430 ;
        RECT 12.505 108.885 14.175 109.655 ;
        RECT 14.345 109.560 14.515 110.360 ;
        RECT 14.800 110.335 15.465 110.505 ;
        RECT 14.800 110.190 14.970 110.335 ;
        RECT 15.785 110.295 15.995 111.435 ;
        RECT 14.685 109.860 14.970 110.190 ;
        RECT 16.165 110.285 16.495 111.265 ;
        RECT 16.665 110.295 16.895 111.435 ;
        RECT 17.105 110.345 18.315 111.435 ;
        RECT 14.800 109.605 14.970 109.860 ;
        RECT 15.205 109.785 15.535 110.155 ;
        RECT 14.345 109.055 14.605 109.560 ;
        RECT 14.800 109.435 15.465 109.605 ;
        RECT 14.785 108.885 15.115 109.265 ;
        RECT 15.295 109.055 15.465 109.435 ;
        RECT 15.785 108.885 15.995 109.705 ;
        RECT 16.165 109.685 16.415 110.285 ;
        RECT 16.585 109.875 16.915 110.125 ;
        RECT 16.165 109.055 16.495 109.685 ;
        RECT 16.665 108.885 16.895 109.705 ;
        RECT 17.105 109.635 17.625 110.175 ;
        RECT 17.795 109.805 18.315 110.345 ;
        RECT 18.485 110.270 18.775 111.435 ;
        RECT 18.950 110.295 19.285 111.265 ;
        RECT 19.455 110.295 19.625 111.435 ;
        RECT 19.795 111.095 21.825 111.265 ;
        RECT 17.105 108.885 18.315 109.635 ;
        RECT 18.950 109.625 19.120 110.295 ;
        RECT 19.795 110.125 19.965 111.095 ;
        RECT 19.290 109.795 19.545 110.125 ;
        RECT 19.770 109.795 19.965 110.125 ;
        RECT 20.135 110.755 21.260 110.925 ;
        RECT 19.375 109.625 19.545 109.795 ;
        RECT 20.135 109.625 20.305 110.755 ;
        RECT 18.485 108.885 18.775 109.610 ;
        RECT 18.950 109.055 19.205 109.625 ;
        RECT 19.375 109.455 20.305 109.625 ;
        RECT 20.475 110.415 21.485 110.585 ;
        RECT 20.475 109.615 20.645 110.415 ;
        RECT 20.130 109.420 20.305 109.455 ;
        RECT 19.375 108.885 19.705 109.285 ;
        RECT 20.130 109.055 20.660 109.420 ;
        RECT 20.850 109.395 21.125 110.215 ;
        RECT 20.845 109.225 21.125 109.395 ;
        RECT 20.850 109.055 21.125 109.225 ;
        RECT 21.295 109.055 21.485 110.415 ;
        RECT 21.655 110.430 21.825 111.095 ;
        RECT 21.995 110.675 22.165 111.435 ;
        RECT 22.400 110.675 22.915 111.085 ;
        RECT 21.655 110.240 22.405 110.430 ;
        RECT 22.575 109.865 22.915 110.675 ;
        RECT 23.085 110.345 24.755 111.435 ;
        RECT 21.685 109.695 22.915 109.865 ;
        RECT 21.665 108.885 22.175 109.420 ;
        RECT 22.395 109.090 22.640 109.695 ;
        RECT 23.085 109.655 23.835 110.175 ;
        RECT 24.005 109.825 24.755 110.345 ;
        RECT 24.965 110.295 25.195 111.435 ;
        RECT 25.365 110.285 25.695 111.265 ;
        RECT 25.865 110.295 26.075 111.435 ;
        RECT 26.395 110.765 26.565 111.265 ;
        RECT 26.735 110.935 27.065 111.435 ;
        RECT 26.395 110.595 27.060 110.765 ;
        RECT 24.945 109.875 25.275 110.125 ;
        RECT 23.085 108.885 24.755 109.655 ;
        RECT 24.965 108.885 25.195 109.705 ;
        RECT 25.445 109.685 25.695 110.285 ;
        RECT 26.310 109.775 26.660 110.425 ;
        RECT 25.365 109.055 25.695 109.685 ;
        RECT 25.865 108.885 26.075 109.705 ;
        RECT 26.830 109.605 27.060 110.595 ;
        RECT 26.395 109.435 27.060 109.605 ;
        RECT 26.395 109.145 26.565 109.435 ;
        RECT 26.735 108.885 27.065 109.265 ;
        RECT 27.235 109.145 27.460 111.265 ;
        RECT 27.675 110.935 28.005 111.435 ;
        RECT 28.175 110.765 28.345 111.265 ;
        RECT 28.580 111.050 29.410 111.220 ;
        RECT 29.650 111.055 30.030 111.435 ;
        RECT 27.650 110.595 28.345 110.765 ;
        RECT 27.650 109.625 27.820 110.595 ;
        RECT 27.990 109.805 28.400 110.425 ;
        RECT 28.570 110.375 29.070 110.755 ;
        RECT 27.650 109.435 28.345 109.625 ;
        RECT 28.570 109.505 28.790 110.375 ;
        RECT 29.240 110.205 29.410 111.050 ;
        RECT 30.210 110.885 30.380 111.175 ;
        RECT 30.550 111.055 30.880 111.435 ;
        RECT 31.350 110.965 31.980 111.215 ;
        RECT 32.160 111.055 32.580 111.435 ;
        RECT 31.810 110.885 31.980 110.965 ;
        RECT 32.780 110.885 33.020 111.175 ;
        RECT 29.580 110.635 30.950 110.885 ;
        RECT 29.580 110.375 29.830 110.635 ;
        RECT 30.340 110.205 30.590 110.365 ;
        RECT 29.240 110.035 30.590 110.205 ;
        RECT 29.240 109.995 29.660 110.035 ;
        RECT 28.970 109.445 29.320 109.815 ;
        RECT 27.675 108.885 28.005 109.265 ;
        RECT 28.175 109.105 28.345 109.435 ;
        RECT 29.490 109.265 29.660 109.995 ;
        RECT 30.760 109.865 30.950 110.635 ;
        RECT 29.830 109.535 30.240 109.865 ;
        RECT 30.530 109.525 30.950 109.865 ;
        RECT 31.120 110.455 31.640 110.765 ;
        RECT 31.810 110.715 33.020 110.885 ;
        RECT 33.250 110.745 33.580 111.435 ;
        RECT 31.120 109.695 31.290 110.455 ;
        RECT 31.460 109.865 31.640 110.275 ;
        RECT 31.810 110.205 31.980 110.715 ;
        RECT 33.750 110.565 33.920 111.175 ;
        RECT 34.190 110.715 34.520 111.225 ;
        RECT 33.750 110.545 34.070 110.565 ;
        RECT 32.150 110.375 34.070 110.545 ;
        RECT 31.810 110.035 33.710 110.205 ;
        RECT 32.040 109.695 32.370 109.815 ;
        RECT 31.120 109.525 32.370 109.695 ;
        RECT 28.645 109.065 29.660 109.265 ;
        RECT 29.830 108.885 30.240 109.325 ;
        RECT 30.530 109.095 30.780 109.525 ;
        RECT 30.980 108.885 31.300 109.345 ;
        RECT 32.540 109.275 32.710 110.035 ;
        RECT 33.380 109.975 33.710 110.035 ;
        RECT 32.900 109.805 33.230 109.865 ;
        RECT 32.900 109.535 33.560 109.805 ;
        RECT 33.880 109.480 34.070 110.375 ;
        RECT 31.860 109.105 32.710 109.275 ;
        RECT 32.910 108.885 33.570 109.365 ;
        RECT 33.750 109.150 34.070 109.480 ;
        RECT 34.270 110.125 34.520 110.715 ;
        RECT 34.700 110.635 34.985 111.435 ;
        RECT 35.165 110.455 35.420 111.125 ;
        RECT 35.965 111.000 41.310 111.435 ;
        RECT 34.270 109.795 35.070 110.125 ;
        RECT 34.270 109.145 34.520 109.795 ;
        RECT 35.240 109.595 35.420 110.455 ;
        RECT 35.165 109.395 35.420 109.595 ;
        RECT 37.550 109.430 37.890 110.260 ;
        RECT 39.370 109.750 39.720 111.000 ;
        RECT 41.485 110.360 41.755 111.265 ;
        RECT 41.925 110.675 42.255 111.435 ;
        RECT 42.435 110.505 42.605 111.265 ;
        RECT 41.485 109.560 41.655 110.360 ;
        RECT 41.940 110.335 42.605 110.505 ;
        RECT 42.865 110.345 44.075 111.435 ;
        RECT 41.940 110.190 42.110 110.335 ;
        RECT 41.825 109.860 42.110 110.190 ;
        RECT 41.940 109.605 42.110 109.860 ;
        RECT 42.345 109.785 42.675 110.155 ;
        RECT 42.865 109.635 43.385 110.175 ;
        RECT 43.555 109.805 44.075 110.345 ;
        RECT 44.245 110.270 44.535 111.435 ;
        RECT 44.765 110.295 44.975 111.435 ;
        RECT 45.145 110.285 45.475 111.265 ;
        RECT 45.645 110.295 45.875 111.435 ;
        RECT 46.085 110.345 47.755 111.435 ;
        RECT 34.700 108.885 34.985 109.345 ;
        RECT 35.165 109.225 35.505 109.395 ;
        RECT 35.165 109.065 35.420 109.225 ;
        RECT 35.965 108.885 41.310 109.430 ;
        RECT 41.485 109.055 41.745 109.560 ;
        RECT 41.940 109.435 42.605 109.605 ;
        RECT 41.925 108.885 42.255 109.265 ;
        RECT 42.435 109.055 42.605 109.435 ;
        RECT 42.865 108.885 44.075 109.635 ;
        RECT 44.245 108.885 44.535 109.610 ;
        RECT 44.765 108.885 44.975 109.705 ;
        RECT 45.145 109.685 45.395 110.285 ;
        RECT 45.565 109.875 45.895 110.125 ;
        RECT 45.145 109.055 45.475 109.685 ;
        RECT 45.645 108.885 45.875 109.705 ;
        RECT 46.085 109.655 46.835 110.175 ;
        RECT 47.005 109.825 47.755 110.345 ;
        RECT 48.385 110.360 48.655 111.265 ;
        RECT 48.825 110.675 49.155 111.435 ;
        RECT 49.335 110.505 49.505 111.265 ;
        RECT 46.085 108.885 47.755 109.655 ;
        RECT 48.385 109.560 48.555 110.360 ;
        RECT 48.840 110.335 49.505 110.505 ;
        RECT 48.840 110.190 49.010 110.335 ;
        RECT 50.265 110.295 50.495 111.435 ;
        RECT 50.665 110.285 50.995 111.265 ;
        RECT 51.165 110.295 51.375 111.435 ;
        RECT 52.615 110.505 52.785 111.265 ;
        RECT 52.965 110.675 53.295 111.435 ;
        RECT 52.615 110.335 53.280 110.505 ;
        RECT 53.465 110.360 53.735 111.265 ;
        RECT 48.725 109.860 49.010 110.190 ;
        RECT 48.840 109.605 49.010 109.860 ;
        RECT 49.245 109.785 49.575 110.155 ;
        RECT 50.245 109.875 50.575 110.125 ;
        RECT 48.385 109.055 48.645 109.560 ;
        RECT 48.840 109.435 49.505 109.605 ;
        RECT 48.825 108.885 49.155 109.265 ;
        RECT 49.335 109.055 49.505 109.435 ;
        RECT 50.265 108.885 50.495 109.705 ;
        RECT 50.745 109.685 50.995 110.285 ;
        RECT 53.110 110.190 53.280 110.335 ;
        RECT 52.545 109.785 52.875 110.155 ;
        RECT 53.110 109.860 53.395 110.190 ;
        RECT 50.665 109.055 50.995 109.685 ;
        RECT 51.165 108.885 51.375 109.705 ;
        RECT 53.110 109.605 53.280 109.860 ;
        RECT 52.615 109.435 53.280 109.605 ;
        RECT 53.565 109.560 53.735 110.360 ;
        RECT 52.615 109.055 52.785 109.435 ;
        RECT 52.965 108.885 53.295 109.265 ;
        RECT 53.475 109.055 53.735 109.560 ;
        RECT 53.910 110.295 54.245 111.265 ;
        RECT 54.415 110.295 54.585 111.435 ;
        RECT 54.755 111.095 56.785 111.265 ;
        RECT 53.910 109.625 54.080 110.295 ;
        RECT 54.755 110.125 54.925 111.095 ;
        RECT 54.250 109.795 54.505 110.125 ;
        RECT 54.730 109.795 54.925 110.125 ;
        RECT 55.095 110.755 56.220 110.925 ;
        RECT 54.335 109.625 54.505 109.795 ;
        RECT 55.095 109.625 55.265 110.755 ;
        RECT 53.910 109.055 54.165 109.625 ;
        RECT 54.335 109.455 55.265 109.625 ;
        RECT 55.435 110.415 56.445 110.585 ;
        RECT 55.435 109.615 55.605 110.415 ;
        RECT 55.810 110.075 56.085 110.215 ;
        RECT 55.805 109.905 56.085 110.075 ;
        RECT 55.090 109.420 55.265 109.455 ;
        RECT 54.335 108.885 54.665 109.285 ;
        RECT 55.090 109.055 55.620 109.420 ;
        RECT 55.810 109.055 56.085 109.905 ;
        RECT 56.255 109.055 56.445 110.415 ;
        RECT 56.615 110.430 56.785 111.095 ;
        RECT 56.955 110.675 57.125 111.435 ;
        RECT 57.360 110.675 57.875 111.085 ;
        RECT 56.615 110.240 57.365 110.430 ;
        RECT 57.535 109.865 57.875 110.675 ;
        RECT 58.135 110.505 58.305 111.265 ;
        RECT 58.485 110.675 58.815 111.435 ;
        RECT 58.135 110.335 58.800 110.505 ;
        RECT 58.985 110.360 59.255 111.265 ;
        RECT 59.515 110.765 59.685 111.265 ;
        RECT 59.855 110.935 60.185 111.435 ;
        RECT 59.515 110.595 60.180 110.765 ;
        RECT 58.630 110.190 58.800 110.335 ;
        RECT 56.645 109.695 57.875 109.865 ;
        RECT 58.065 109.785 58.395 110.155 ;
        RECT 58.630 109.860 58.915 110.190 ;
        RECT 56.625 108.885 57.135 109.420 ;
        RECT 57.355 109.090 57.600 109.695 ;
        RECT 58.630 109.605 58.800 109.860 ;
        RECT 58.135 109.435 58.800 109.605 ;
        RECT 59.085 109.560 59.255 110.360 ;
        RECT 59.430 109.775 59.780 110.425 ;
        RECT 59.950 109.605 60.180 110.595 ;
        RECT 58.135 109.055 58.305 109.435 ;
        RECT 58.485 108.885 58.815 109.265 ;
        RECT 58.995 109.055 59.255 109.560 ;
        RECT 59.515 109.435 60.180 109.605 ;
        RECT 59.515 109.145 59.685 109.435 ;
        RECT 59.855 108.885 60.185 109.265 ;
        RECT 60.355 109.145 60.580 111.265 ;
        RECT 60.795 110.935 61.125 111.435 ;
        RECT 61.295 110.765 61.465 111.265 ;
        RECT 61.700 111.050 62.530 111.220 ;
        RECT 62.770 111.055 63.150 111.435 ;
        RECT 60.770 110.595 61.465 110.765 ;
        RECT 60.770 109.625 60.940 110.595 ;
        RECT 61.110 109.805 61.520 110.425 ;
        RECT 61.690 110.375 62.190 110.755 ;
        RECT 60.770 109.435 61.465 109.625 ;
        RECT 61.690 109.505 61.910 110.375 ;
        RECT 62.360 110.205 62.530 111.050 ;
        RECT 63.330 110.885 63.500 111.175 ;
        RECT 63.670 111.055 64.000 111.435 ;
        RECT 64.470 110.965 65.100 111.215 ;
        RECT 65.280 111.055 65.700 111.435 ;
        RECT 64.930 110.885 65.100 110.965 ;
        RECT 65.900 110.885 66.140 111.175 ;
        RECT 62.700 110.635 64.070 110.885 ;
        RECT 62.700 110.375 62.950 110.635 ;
        RECT 63.460 110.205 63.710 110.365 ;
        RECT 62.360 110.035 63.710 110.205 ;
        RECT 62.360 109.995 62.780 110.035 ;
        RECT 62.090 109.445 62.440 109.815 ;
        RECT 60.795 108.885 61.125 109.265 ;
        RECT 61.295 109.105 61.465 109.435 ;
        RECT 62.610 109.265 62.780 109.995 ;
        RECT 63.880 109.865 64.070 110.635 ;
        RECT 62.950 109.535 63.360 109.865 ;
        RECT 63.650 109.525 64.070 109.865 ;
        RECT 64.240 110.455 64.760 110.765 ;
        RECT 64.930 110.715 66.140 110.885 ;
        RECT 66.370 110.745 66.700 111.435 ;
        RECT 64.240 109.695 64.410 110.455 ;
        RECT 64.580 109.865 64.760 110.275 ;
        RECT 64.930 110.205 65.100 110.715 ;
        RECT 66.870 110.565 67.040 111.175 ;
        RECT 67.310 110.715 67.640 111.225 ;
        RECT 66.870 110.545 67.190 110.565 ;
        RECT 65.270 110.375 67.190 110.545 ;
        RECT 64.930 110.035 66.830 110.205 ;
        RECT 65.160 109.695 65.490 109.815 ;
        RECT 64.240 109.525 65.490 109.695 ;
        RECT 61.765 109.065 62.780 109.265 ;
        RECT 62.950 108.885 63.360 109.325 ;
        RECT 63.650 109.095 63.900 109.525 ;
        RECT 64.100 108.885 64.420 109.345 ;
        RECT 65.660 109.275 65.830 110.035 ;
        RECT 66.500 109.975 66.830 110.035 ;
        RECT 66.020 109.805 66.350 109.865 ;
        RECT 66.020 109.535 66.680 109.805 ;
        RECT 67.000 109.480 67.190 110.375 ;
        RECT 64.980 109.105 65.830 109.275 ;
        RECT 66.030 108.885 66.690 109.365 ;
        RECT 66.870 109.150 67.190 109.480 ;
        RECT 67.390 110.125 67.640 110.715 ;
        RECT 67.820 110.635 68.105 111.435 ;
        RECT 68.285 110.455 68.540 111.125 ;
        RECT 67.390 109.795 68.190 110.125 ;
        RECT 67.390 109.145 67.640 109.795 ;
        RECT 68.360 109.595 68.540 110.455 ;
        RECT 70.005 110.270 70.295 111.435 ;
        RECT 71.015 110.765 71.185 111.265 ;
        RECT 71.355 110.935 71.685 111.435 ;
        RECT 71.015 110.595 71.680 110.765 ;
        RECT 70.930 109.775 71.280 110.425 ;
        RECT 68.285 109.395 68.540 109.595 ;
        RECT 67.820 108.885 68.105 109.345 ;
        RECT 68.285 109.225 68.625 109.395 ;
        RECT 68.285 109.065 68.540 109.225 ;
        RECT 70.005 108.885 70.295 109.610 ;
        RECT 71.450 109.605 71.680 110.595 ;
        RECT 71.015 109.435 71.680 109.605 ;
        RECT 71.015 109.145 71.185 109.435 ;
        RECT 71.355 108.885 71.685 109.265 ;
        RECT 71.855 109.145 72.080 111.265 ;
        RECT 72.295 110.935 72.625 111.435 ;
        RECT 72.795 110.765 72.965 111.265 ;
        RECT 73.200 111.050 74.030 111.220 ;
        RECT 74.270 111.055 74.650 111.435 ;
        RECT 72.270 110.595 72.965 110.765 ;
        RECT 72.270 109.625 72.440 110.595 ;
        RECT 72.610 109.805 73.020 110.425 ;
        RECT 73.190 110.375 73.690 110.755 ;
        RECT 72.270 109.435 72.965 109.625 ;
        RECT 73.190 109.505 73.410 110.375 ;
        RECT 73.860 110.205 74.030 111.050 ;
        RECT 74.830 110.885 75.000 111.175 ;
        RECT 75.170 111.055 75.500 111.435 ;
        RECT 75.970 110.965 76.600 111.215 ;
        RECT 76.780 111.055 77.200 111.435 ;
        RECT 76.430 110.885 76.600 110.965 ;
        RECT 77.400 110.885 77.640 111.175 ;
        RECT 74.200 110.635 75.570 110.885 ;
        RECT 74.200 110.375 74.450 110.635 ;
        RECT 74.960 110.205 75.210 110.365 ;
        RECT 73.860 110.035 75.210 110.205 ;
        RECT 73.860 109.995 74.280 110.035 ;
        RECT 73.590 109.445 73.940 109.815 ;
        RECT 72.295 108.885 72.625 109.265 ;
        RECT 72.795 109.105 72.965 109.435 ;
        RECT 74.110 109.265 74.280 109.995 ;
        RECT 75.380 109.865 75.570 110.635 ;
        RECT 74.450 109.535 74.860 109.865 ;
        RECT 75.150 109.525 75.570 109.865 ;
        RECT 75.740 110.455 76.260 110.765 ;
        RECT 76.430 110.715 77.640 110.885 ;
        RECT 77.870 110.745 78.200 111.435 ;
        RECT 75.740 109.695 75.910 110.455 ;
        RECT 76.080 109.865 76.260 110.275 ;
        RECT 76.430 110.205 76.600 110.715 ;
        RECT 78.370 110.565 78.540 111.175 ;
        RECT 78.810 110.715 79.140 111.225 ;
        RECT 78.370 110.545 78.690 110.565 ;
        RECT 76.770 110.375 78.690 110.545 ;
        RECT 76.430 110.035 78.330 110.205 ;
        RECT 76.660 109.695 76.990 109.815 ;
        RECT 75.740 109.525 76.990 109.695 ;
        RECT 73.265 109.065 74.280 109.265 ;
        RECT 74.450 108.885 74.860 109.325 ;
        RECT 75.150 109.095 75.400 109.525 ;
        RECT 75.600 108.885 75.920 109.345 ;
        RECT 77.160 109.275 77.330 110.035 ;
        RECT 78.000 109.975 78.330 110.035 ;
        RECT 77.520 109.805 77.850 109.865 ;
        RECT 77.520 109.535 78.180 109.805 ;
        RECT 78.500 109.480 78.690 110.375 ;
        RECT 76.480 109.105 77.330 109.275 ;
        RECT 77.530 108.885 78.190 109.365 ;
        RECT 78.370 109.150 78.690 109.480 ;
        RECT 78.890 110.125 79.140 110.715 ;
        RECT 79.320 110.635 79.605 111.435 ;
        RECT 79.785 110.455 80.040 111.125 ;
        RECT 81.595 110.690 81.865 111.435 ;
        RECT 82.495 111.430 88.770 111.435 ;
        RECT 82.035 110.520 82.325 111.260 ;
        RECT 82.495 110.705 82.750 111.430 ;
        RECT 82.935 110.535 83.195 111.260 ;
        RECT 83.365 110.705 83.610 111.430 ;
        RECT 83.795 110.535 84.055 111.260 ;
        RECT 84.225 110.705 84.470 111.430 ;
        RECT 84.655 110.535 84.915 111.260 ;
        RECT 85.085 110.705 85.330 111.430 ;
        RECT 85.500 110.535 85.760 111.260 ;
        RECT 85.930 110.705 86.190 111.430 ;
        RECT 86.360 110.535 86.620 111.260 ;
        RECT 86.790 110.705 87.050 111.430 ;
        RECT 87.220 110.535 87.480 111.260 ;
        RECT 87.650 110.705 87.910 111.430 ;
        RECT 88.080 110.535 88.340 111.260 ;
        RECT 88.510 110.635 88.770 111.430 ;
        RECT 82.935 110.520 88.340 110.535 ;
        RECT 79.860 110.415 80.040 110.455 ;
        RECT 79.860 110.245 80.125 110.415 ;
        RECT 81.595 110.295 88.340 110.520 ;
        RECT 78.890 109.795 79.690 110.125 ;
        RECT 78.890 109.145 79.140 109.795 ;
        RECT 79.860 109.595 80.040 110.245 ;
        RECT 79.320 108.885 79.605 109.345 ;
        RECT 79.785 109.065 80.040 109.595 ;
        RECT 81.595 109.705 82.760 110.295 ;
        RECT 88.940 110.125 89.190 111.260 ;
        RECT 89.370 110.625 89.630 111.435 ;
        RECT 89.805 110.125 90.050 111.265 ;
        RECT 90.230 110.625 90.525 111.435 ;
        RECT 90.705 110.675 91.220 111.085 ;
        RECT 91.455 110.675 91.625 111.435 ;
        RECT 91.795 111.095 93.825 111.265 ;
        RECT 82.930 109.875 90.050 110.125 ;
        RECT 81.595 109.535 88.340 109.705 ;
        RECT 81.595 108.885 81.895 109.365 ;
        RECT 82.065 109.080 82.325 109.535 ;
        RECT 82.495 108.885 82.755 109.365 ;
        RECT 82.935 109.080 83.195 109.535 ;
        RECT 83.365 108.885 83.615 109.365 ;
        RECT 83.795 109.080 84.055 109.535 ;
        RECT 84.225 108.885 84.475 109.365 ;
        RECT 84.655 109.080 84.915 109.535 ;
        RECT 85.085 108.885 85.330 109.365 ;
        RECT 85.500 109.080 85.775 109.535 ;
        RECT 85.945 108.885 86.190 109.365 ;
        RECT 86.360 109.080 86.620 109.535 ;
        RECT 86.790 108.885 87.050 109.365 ;
        RECT 87.220 109.080 87.480 109.535 ;
        RECT 87.650 108.885 87.910 109.365 ;
        RECT 88.080 109.080 88.340 109.535 ;
        RECT 88.510 108.885 88.770 109.445 ;
        RECT 88.940 109.065 89.190 109.875 ;
        RECT 89.370 108.885 89.630 109.410 ;
        RECT 89.800 109.065 90.050 109.875 ;
        RECT 90.220 109.565 90.535 110.125 ;
        RECT 90.705 109.865 91.045 110.675 ;
        RECT 91.795 110.430 91.965 111.095 ;
        RECT 92.360 110.755 93.485 110.925 ;
        RECT 91.215 110.240 91.965 110.430 ;
        RECT 92.135 110.415 93.145 110.585 ;
        RECT 90.705 109.695 91.935 109.865 ;
        RECT 90.230 108.885 90.535 109.395 ;
        RECT 90.980 109.090 91.225 109.695 ;
        RECT 91.445 108.885 91.955 109.420 ;
        RECT 92.135 109.055 92.325 110.415 ;
        RECT 92.495 109.395 92.770 110.215 ;
        RECT 92.975 109.615 93.145 110.415 ;
        RECT 93.315 109.625 93.485 110.755 ;
        RECT 93.655 110.125 93.825 111.095 ;
        RECT 93.995 110.295 94.165 111.435 ;
        RECT 94.335 110.295 94.670 111.265 ;
        RECT 93.655 109.795 93.850 110.125 ;
        RECT 94.075 109.795 94.330 110.125 ;
        RECT 94.075 109.625 94.245 109.795 ;
        RECT 94.500 109.625 94.670 110.295 ;
        RECT 95.765 110.270 96.055 111.435 ;
        RECT 96.225 110.675 96.740 111.085 ;
        RECT 96.975 110.675 97.145 111.435 ;
        RECT 97.315 111.095 99.345 111.265 ;
        RECT 96.225 109.865 96.565 110.675 ;
        RECT 97.315 110.430 97.485 111.095 ;
        RECT 97.880 110.755 99.005 110.925 ;
        RECT 96.735 110.240 97.485 110.430 ;
        RECT 97.655 110.415 98.665 110.585 ;
        RECT 96.225 109.695 97.455 109.865 ;
        RECT 93.315 109.455 94.245 109.625 ;
        RECT 93.315 109.420 93.490 109.455 ;
        RECT 92.495 109.225 92.775 109.395 ;
        RECT 92.495 109.055 92.770 109.225 ;
        RECT 92.960 109.055 93.490 109.420 ;
        RECT 93.915 108.885 94.245 109.285 ;
        RECT 94.415 109.055 94.670 109.625 ;
        RECT 95.765 108.885 96.055 109.610 ;
        RECT 96.500 109.090 96.745 109.695 ;
        RECT 96.965 108.885 97.475 109.420 ;
        RECT 97.655 109.055 97.845 110.415 ;
        RECT 98.015 109.395 98.290 110.215 ;
        RECT 98.495 109.615 98.665 110.415 ;
        RECT 98.835 109.625 99.005 110.755 ;
        RECT 99.175 110.125 99.345 111.095 ;
        RECT 99.515 110.295 99.685 111.435 ;
        RECT 99.855 110.295 100.190 111.265 ;
        RECT 99.175 109.795 99.370 110.125 ;
        RECT 99.595 109.795 99.850 110.125 ;
        RECT 99.595 109.625 99.765 109.795 ;
        RECT 100.020 109.625 100.190 110.295 ;
        RECT 98.835 109.455 99.765 109.625 ;
        RECT 98.835 109.420 99.010 109.455 ;
        RECT 98.015 109.225 98.295 109.395 ;
        RECT 98.015 109.055 98.290 109.225 ;
        RECT 98.480 109.055 99.010 109.420 ;
        RECT 99.435 108.885 99.765 109.285 ;
        RECT 99.935 109.055 100.190 109.625 ;
        RECT 100.365 110.360 100.635 111.265 ;
        RECT 100.805 110.675 101.135 111.435 ;
        RECT 101.315 110.505 101.485 111.265 ;
        RECT 100.365 109.560 100.535 110.360 ;
        RECT 100.820 110.335 101.485 110.505 ;
        RECT 100.820 110.190 100.990 110.335 ;
        RECT 101.805 110.295 102.015 111.435 ;
        RECT 100.705 109.860 100.990 110.190 ;
        RECT 102.185 110.285 102.515 111.265 ;
        RECT 102.685 110.295 102.915 111.435 ;
        RECT 103.585 110.675 104.100 111.085 ;
        RECT 104.335 110.675 104.505 111.435 ;
        RECT 104.675 111.095 106.705 111.265 ;
        RECT 100.820 109.605 100.990 109.860 ;
        RECT 101.225 109.785 101.555 110.155 ;
        RECT 100.365 109.055 100.625 109.560 ;
        RECT 100.820 109.435 101.485 109.605 ;
        RECT 100.805 108.885 101.135 109.265 ;
        RECT 101.315 109.055 101.485 109.435 ;
        RECT 101.805 108.885 102.015 109.705 ;
        RECT 102.185 109.685 102.435 110.285 ;
        RECT 102.605 109.875 102.935 110.125 ;
        RECT 103.585 109.865 103.925 110.675 ;
        RECT 104.675 110.430 104.845 111.095 ;
        RECT 105.240 110.755 106.365 110.925 ;
        RECT 104.095 110.240 104.845 110.430 ;
        RECT 105.015 110.415 106.025 110.585 ;
        RECT 102.185 109.055 102.515 109.685 ;
        RECT 102.685 108.885 102.915 109.705 ;
        RECT 103.585 109.695 104.815 109.865 ;
        RECT 103.860 109.090 104.105 109.695 ;
        RECT 104.325 108.885 104.835 109.420 ;
        RECT 105.015 109.055 105.205 110.415 ;
        RECT 105.375 109.395 105.650 110.215 ;
        RECT 105.855 109.615 106.025 110.415 ;
        RECT 106.195 109.625 106.365 110.755 ;
        RECT 106.535 110.125 106.705 111.095 ;
        RECT 106.875 110.295 107.045 111.435 ;
        RECT 107.215 110.295 107.550 111.265 ;
        RECT 107.815 110.765 107.985 111.265 ;
        RECT 108.155 110.935 108.485 111.435 ;
        RECT 107.815 110.595 108.480 110.765 ;
        RECT 106.535 109.795 106.730 110.125 ;
        RECT 106.955 109.795 107.210 110.125 ;
        RECT 106.955 109.625 107.125 109.795 ;
        RECT 107.380 109.625 107.550 110.295 ;
        RECT 107.730 109.775 108.080 110.425 ;
        RECT 106.195 109.455 107.125 109.625 ;
        RECT 106.195 109.420 106.370 109.455 ;
        RECT 105.375 109.225 105.655 109.395 ;
        RECT 105.375 109.055 105.650 109.225 ;
        RECT 105.840 109.055 106.370 109.420 ;
        RECT 106.795 108.885 107.125 109.285 ;
        RECT 107.295 109.055 107.550 109.625 ;
        RECT 108.250 109.605 108.480 110.595 ;
        RECT 107.815 109.435 108.480 109.605 ;
        RECT 107.815 109.145 107.985 109.435 ;
        RECT 108.155 108.885 108.485 109.265 ;
        RECT 108.655 109.145 108.880 111.265 ;
        RECT 109.095 110.935 109.425 111.435 ;
        RECT 109.595 110.765 109.765 111.265 ;
        RECT 110.000 111.050 110.830 111.220 ;
        RECT 111.070 111.055 111.450 111.435 ;
        RECT 109.070 110.595 109.765 110.765 ;
        RECT 109.070 109.625 109.240 110.595 ;
        RECT 109.410 109.805 109.820 110.425 ;
        RECT 109.990 110.375 110.490 110.755 ;
        RECT 109.070 109.435 109.765 109.625 ;
        RECT 109.990 109.505 110.210 110.375 ;
        RECT 110.660 110.205 110.830 111.050 ;
        RECT 111.630 110.885 111.800 111.175 ;
        RECT 111.970 111.055 112.300 111.435 ;
        RECT 112.770 110.965 113.400 111.215 ;
        RECT 113.580 111.055 114.000 111.435 ;
        RECT 113.230 110.885 113.400 110.965 ;
        RECT 114.200 110.885 114.440 111.175 ;
        RECT 111.000 110.635 112.370 110.885 ;
        RECT 111.000 110.375 111.250 110.635 ;
        RECT 111.760 110.205 112.010 110.365 ;
        RECT 110.660 110.035 112.010 110.205 ;
        RECT 110.660 109.995 111.080 110.035 ;
        RECT 110.390 109.445 110.740 109.815 ;
        RECT 109.095 108.885 109.425 109.265 ;
        RECT 109.595 109.105 109.765 109.435 ;
        RECT 110.910 109.265 111.080 109.995 ;
        RECT 112.180 109.865 112.370 110.635 ;
        RECT 111.250 109.535 111.660 109.865 ;
        RECT 111.950 109.525 112.370 109.865 ;
        RECT 112.540 110.455 113.060 110.765 ;
        RECT 113.230 110.715 114.440 110.885 ;
        RECT 114.670 110.745 115.000 111.435 ;
        RECT 112.540 109.695 112.710 110.455 ;
        RECT 112.880 109.865 113.060 110.275 ;
        RECT 113.230 110.205 113.400 110.715 ;
        RECT 115.170 110.565 115.340 111.175 ;
        RECT 115.610 110.715 115.940 111.225 ;
        RECT 115.170 110.545 115.490 110.565 ;
        RECT 113.570 110.375 115.490 110.545 ;
        RECT 113.230 110.035 115.130 110.205 ;
        RECT 113.460 109.695 113.790 109.815 ;
        RECT 112.540 109.525 113.790 109.695 ;
        RECT 110.065 109.065 111.080 109.265 ;
        RECT 111.250 108.885 111.660 109.325 ;
        RECT 111.950 109.095 112.200 109.525 ;
        RECT 112.400 108.885 112.720 109.345 ;
        RECT 113.960 109.275 114.130 110.035 ;
        RECT 114.800 109.975 115.130 110.035 ;
        RECT 114.320 109.805 114.650 109.865 ;
        RECT 114.320 109.535 114.980 109.805 ;
        RECT 115.300 109.480 115.490 110.375 ;
        RECT 113.280 109.105 114.130 109.275 ;
        RECT 114.330 108.885 114.990 109.365 ;
        RECT 115.170 109.150 115.490 109.480 ;
        RECT 115.690 110.125 115.940 110.715 ;
        RECT 116.120 110.635 116.405 111.435 ;
        RECT 116.585 110.455 116.840 111.125 ;
        RECT 115.690 109.795 116.490 110.125 ;
        RECT 115.690 109.145 115.940 109.795 ;
        RECT 116.660 109.595 116.840 110.455 ;
        RECT 117.425 110.295 117.655 111.435 ;
        RECT 117.825 110.285 118.155 111.265 ;
        RECT 118.325 110.295 118.535 111.435 ;
        RECT 118.765 110.345 121.355 111.435 ;
        RECT 117.405 109.875 117.735 110.125 ;
        RECT 116.585 109.395 116.840 109.595 ;
        RECT 116.120 108.885 116.405 109.345 ;
        RECT 116.585 109.225 116.925 109.395 ;
        RECT 116.585 109.065 116.840 109.225 ;
        RECT 117.425 108.885 117.655 109.705 ;
        RECT 117.905 109.685 118.155 110.285 ;
        RECT 117.825 109.055 118.155 109.685 ;
        RECT 118.325 108.885 118.535 109.705 ;
        RECT 118.765 109.655 119.975 110.175 ;
        RECT 120.145 109.825 121.355 110.345 ;
        RECT 121.525 110.270 121.815 111.435 ;
        RECT 122.445 110.345 123.655 111.435 ;
        RECT 122.445 109.805 122.965 110.345 ;
        RECT 118.765 108.885 121.355 109.655 ;
        RECT 123.135 109.635 123.655 110.175 ;
        RECT 121.525 108.885 121.815 109.610 ;
        RECT 122.445 108.885 123.655 109.635 ;
        RECT 5.520 108.715 123.740 108.885 ;
        RECT 5.605 107.965 6.815 108.715 ;
        RECT 6.985 108.170 12.330 108.715 ;
        RECT 12.505 108.170 17.850 108.715 ;
        RECT 5.605 107.425 6.125 107.965 ;
        RECT 6.295 107.255 6.815 107.795 ;
        RECT 8.570 107.340 8.910 108.170 ;
        RECT 5.605 106.165 6.815 107.255 ;
        RECT 10.390 106.600 10.740 107.850 ;
        RECT 14.090 107.340 14.430 108.170 ;
        RECT 19.035 108.165 19.205 108.545 ;
        RECT 19.385 108.335 19.715 108.715 ;
        RECT 19.035 107.995 19.700 108.165 ;
        RECT 19.895 108.040 20.155 108.545 ;
        RECT 15.910 106.600 16.260 107.850 ;
        RECT 18.965 107.445 19.295 107.815 ;
        RECT 19.530 107.740 19.700 107.995 ;
        RECT 19.530 107.410 19.815 107.740 ;
        RECT 19.530 107.265 19.700 107.410 ;
        RECT 19.035 107.095 19.700 107.265 ;
        RECT 19.985 107.240 20.155 108.040 ;
        RECT 20.415 108.165 20.585 108.455 ;
        RECT 20.755 108.335 21.085 108.715 ;
        RECT 20.415 107.995 21.080 108.165 ;
        RECT 6.985 106.165 12.330 106.600 ;
        RECT 12.505 106.165 17.850 106.600 ;
        RECT 19.035 106.335 19.205 107.095 ;
        RECT 19.385 106.165 19.715 106.925 ;
        RECT 19.885 106.335 20.155 107.240 ;
        RECT 20.330 107.175 20.680 107.825 ;
        RECT 20.850 107.005 21.080 107.995 ;
        RECT 20.415 106.835 21.080 107.005 ;
        RECT 20.415 106.335 20.585 106.835 ;
        RECT 20.755 106.165 21.085 106.665 ;
        RECT 21.255 106.335 21.480 108.455 ;
        RECT 21.695 108.335 22.025 108.715 ;
        RECT 22.195 108.165 22.365 108.495 ;
        RECT 22.665 108.335 23.680 108.535 ;
        RECT 21.670 107.975 22.365 108.165 ;
        RECT 21.670 107.005 21.840 107.975 ;
        RECT 22.010 107.175 22.420 107.795 ;
        RECT 22.590 107.225 22.810 108.095 ;
        RECT 22.990 107.785 23.340 108.155 ;
        RECT 23.510 107.605 23.680 108.335 ;
        RECT 23.850 108.275 24.260 108.715 ;
        RECT 24.550 108.075 24.800 108.505 ;
        RECT 25.000 108.255 25.320 108.715 ;
        RECT 25.880 108.325 26.730 108.495 ;
        RECT 23.850 107.735 24.260 108.065 ;
        RECT 24.550 107.735 24.970 108.075 ;
        RECT 23.260 107.565 23.680 107.605 ;
        RECT 23.260 107.395 24.610 107.565 ;
        RECT 21.670 106.835 22.365 107.005 ;
        RECT 22.590 106.845 23.090 107.225 ;
        RECT 21.695 106.165 22.025 106.665 ;
        RECT 22.195 106.335 22.365 106.835 ;
        RECT 23.260 106.550 23.430 107.395 ;
        RECT 24.360 107.235 24.610 107.395 ;
        RECT 23.600 106.965 23.850 107.225 ;
        RECT 24.780 106.965 24.970 107.735 ;
        RECT 23.600 106.715 24.970 106.965 ;
        RECT 25.140 107.905 26.390 108.075 ;
        RECT 25.140 107.145 25.310 107.905 ;
        RECT 26.060 107.785 26.390 107.905 ;
        RECT 25.480 107.325 25.660 107.735 ;
        RECT 26.560 107.565 26.730 108.325 ;
        RECT 26.930 108.235 27.590 108.715 ;
        RECT 27.770 108.120 28.090 108.450 ;
        RECT 26.920 107.795 27.580 108.065 ;
        RECT 26.920 107.735 27.250 107.795 ;
        RECT 27.400 107.565 27.730 107.625 ;
        RECT 25.830 107.395 27.730 107.565 ;
        RECT 25.140 106.835 25.660 107.145 ;
        RECT 25.830 106.885 26.000 107.395 ;
        RECT 27.900 107.225 28.090 108.120 ;
        RECT 26.170 107.055 28.090 107.225 ;
        RECT 27.770 107.035 28.090 107.055 ;
        RECT 28.290 107.805 28.540 108.455 ;
        RECT 28.720 108.255 29.005 108.715 ;
        RECT 29.185 108.005 29.440 108.535 ;
        RECT 28.290 107.475 29.090 107.805 ;
        RECT 25.830 106.715 27.040 106.885 ;
        RECT 22.600 106.380 23.430 106.550 ;
        RECT 23.670 106.165 24.050 106.545 ;
        RECT 24.230 106.425 24.400 106.715 ;
        RECT 25.830 106.635 26.000 106.715 ;
        RECT 24.570 106.165 24.900 106.545 ;
        RECT 25.370 106.385 26.000 106.635 ;
        RECT 26.180 106.165 26.600 106.545 ;
        RECT 26.800 106.425 27.040 106.715 ;
        RECT 27.270 106.165 27.600 106.855 ;
        RECT 27.770 106.425 27.940 107.035 ;
        RECT 28.290 106.885 28.540 107.475 ;
        RECT 29.260 107.145 29.440 108.005 ;
        RECT 29.985 107.965 31.195 108.715 ;
        RECT 31.365 107.990 31.655 108.715 ;
        RECT 32.835 108.165 33.005 108.545 ;
        RECT 33.185 108.335 33.515 108.715 ;
        RECT 32.835 107.995 33.500 108.165 ;
        RECT 33.695 108.040 33.955 108.545 ;
        RECT 29.985 107.425 30.505 107.965 ;
        RECT 30.675 107.255 31.195 107.795 ;
        RECT 32.765 107.445 33.095 107.815 ;
        RECT 33.330 107.740 33.500 107.995 ;
        RECT 33.330 107.410 33.615 107.740 ;
        RECT 28.210 106.375 28.540 106.885 ;
        RECT 28.720 106.165 29.005 106.965 ;
        RECT 29.185 106.675 29.440 107.145 ;
        RECT 29.185 106.505 29.525 106.675 ;
        RECT 29.185 106.475 29.440 106.505 ;
        RECT 29.985 106.165 31.195 107.255 ;
        RECT 31.365 106.165 31.655 107.330 ;
        RECT 33.330 107.265 33.500 107.410 ;
        RECT 32.835 107.095 33.500 107.265 ;
        RECT 33.785 107.240 33.955 108.040 ;
        RECT 34.215 108.165 34.385 108.455 ;
        RECT 34.555 108.335 34.885 108.715 ;
        RECT 34.215 107.995 34.880 108.165 ;
        RECT 32.835 106.335 33.005 107.095 ;
        RECT 33.185 106.165 33.515 106.925 ;
        RECT 33.685 106.335 33.955 107.240 ;
        RECT 34.130 107.175 34.480 107.825 ;
        RECT 34.650 107.005 34.880 107.995 ;
        RECT 34.215 106.835 34.880 107.005 ;
        RECT 34.215 106.335 34.385 106.835 ;
        RECT 34.555 106.165 34.885 106.665 ;
        RECT 35.055 106.335 35.280 108.455 ;
        RECT 35.495 108.335 35.825 108.715 ;
        RECT 35.995 108.165 36.165 108.495 ;
        RECT 36.465 108.335 37.480 108.535 ;
        RECT 35.470 107.975 36.165 108.165 ;
        RECT 35.470 107.005 35.640 107.975 ;
        RECT 35.810 107.175 36.220 107.795 ;
        RECT 36.390 107.225 36.610 108.095 ;
        RECT 36.790 107.785 37.140 108.155 ;
        RECT 37.310 107.605 37.480 108.335 ;
        RECT 37.650 108.275 38.060 108.715 ;
        RECT 38.350 108.075 38.600 108.505 ;
        RECT 38.800 108.255 39.120 108.715 ;
        RECT 39.680 108.325 40.530 108.495 ;
        RECT 37.650 107.735 38.060 108.065 ;
        RECT 38.350 107.735 38.770 108.075 ;
        RECT 37.060 107.565 37.480 107.605 ;
        RECT 37.060 107.395 38.410 107.565 ;
        RECT 35.470 106.835 36.165 107.005 ;
        RECT 36.390 106.845 36.890 107.225 ;
        RECT 35.495 106.165 35.825 106.665 ;
        RECT 35.995 106.335 36.165 106.835 ;
        RECT 37.060 106.550 37.230 107.395 ;
        RECT 38.160 107.235 38.410 107.395 ;
        RECT 37.400 106.965 37.650 107.225 ;
        RECT 38.580 106.965 38.770 107.735 ;
        RECT 37.400 106.715 38.770 106.965 ;
        RECT 38.940 107.905 40.190 108.075 ;
        RECT 38.940 107.145 39.110 107.905 ;
        RECT 39.860 107.785 40.190 107.905 ;
        RECT 39.280 107.325 39.460 107.735 ;
        RECT 40.360 107.565 40.530 108.325 ;
        RECT 40.730 108.235 41.390 108.715 ;
        RECT 41.570 108.120 41.890 108.450 ;
        RECT 40.720 107.795 41.380 108.065 ;
        RECT 40.720 107.735 41.050 107.795 ;
        RECT 41.200 107.565 41.530 107.625 ;
        RECT 39.630 107.395 41.530 107.565 ;
        RECT 38.940 106.835 39.460 107.145 ;
        RECT 39.630 106.885 39.800 107.395 ;
        RECT 41.700 107.225 41.890 108.120 ;
        RECT 39.970 107.055 41.890 107.225 ;
        RECT 41.570 107.035 41.890 107.055 ;
        RECT 42.090 107.805 42.340 108.455 ;
        RECT 42.520 108.255 42.805 108.715 ;
        RECT 42.985 108.005 43.240 108.535 ;
        RECT 42.090 107.475 42.890 107.805 ;
        RECT 39.630 106.715 40.840 106.885 ;
        RECT 36.400 106.380 37.230 106.550 ;
        RECT 37.470 106.165 37.850 106.545 ;
        RECT 38.030 106.425 38.200 106.715 ;
        RECT 39.630 106.635 39.800 106.715 ;
        RECT 38.370 106.165 38.700 106.545 ;
        RECT 39.170 106.385 39.800 106.635 ;
        RECT 39.980 106.165 40.400 106.545 ;
        RECT 40.600 106.425 40.840 106.715 ;
        RECT 41.070 106.165 41.400 106.855 ;
        RECT 41.570 106.425 41.740 107.035 ;
        RECT 42.090 106.885 42.340 107.475 ;
        RECT 43.060 107.145 43.240 108.005 ;
        RECT 43.845 107.895 44.055 108.715 ;
        RECT 44.225 107.915 44.555 108.545 ;
        RECT 44.225 107.315 44.475 107.915 ;
        RECT 44.725 107.895 44.955 108.715 ;
        RECT 45.715 108.165 45.885 108.455 ;
        RECT 46.055 108.335 46.385 108.715 ;
        RECT 45.715 107.995 46.380 108.165 ;
        RECT 44.645 107.475 44.975 107.725 ;
        RECT 42.010 106.375 42.340 106.885 ;
        RECT 42.520 106.165 42.805 106.965 ;
        RECT 42.985 106.675 43.240 107.145 ;
        RECT 42.985 106.505 43.325 106.675 ;
        RECT 42.985 106.475 43.240 106.505 ;
        RECT 43.845 106.165 44.055 107.305 ;
        RECT 44.225 106.335 44.555 107.315 ;
        RECT 44.725 106.165 44.955 107.305 ;
        RECT 45.630 107.175 45.980 107.825 ;
        RECT 46.150 107.005 46.380 107.995 ;
        RECT 45.715 106.835 46.380 107.005 ;
        RECT 45.715 106.335 45.885 106.835 ;
        RECT 46.055 106.165 46.385 106.665 ;
        RECT 46.555 106.335 46.780 108.455 ;
        RECT 46.995 108.335 47.325 108.715 ;
        RECT 47.495 108.165 47.665 108.495 ;
        RECT 47.965 108.335 48.980 108.535 ;
        RECT 46.970 107.975 47.665 108.165 ;
        RECT 46.970 107.005 47.140 107.975 ;
        RECT 47.310 107.175 47.720 107.795 ;
        RECT 47.890 107.225 48.110 108.095 ;
        RECT 48.290 107.785 48.640 108.155 ;
        RECT 48.810 107.605 48.980 108.335 ;
        RECT 49.150 108.275 49.560 108.715 ;
        RECT 49.850 108.075 50.100 108.505 ;
        RECT 50.300 108.255 50.620 108.715 ;
        RECT 51.180 108.325 52.030 108.495 ;
        RECT 49.150 107.735 49.560 108.065 ;
        RECT 49.850 107.735 50.270 108.075 ;
        RECT 48.560 107.565 48.980 107.605 ;
        RECT 48.560 107.395 49.910 107.565 ;
        RECT 46.970 106.835 47.665 107.005 ;
        RECT 47.890 106.845 48.390 107.225 ;
        RECT 46.995 106.165 47.325 106.665 ;
        RECT 47.495 106.335 47.665 106.835 ;
        RECT 48.560 106.550 48.730 107.395 ;
        RECT 49.660 107.235 49.910 107.395 ;
        RECT 48.900 106.965 49.150 107.225 ;
        RECT 50.080 106.965 50.270 107.735 ;
        RECT 48.900 106.715 50.270 106.965 ;
        RECT 50.440 107.905 51.690 108.075 ;
        RECT 50.440 107.145 50.610 107.905 ;
        RECT 51.360 107.785 51.690 107.905 ;
        RECT 50.780 107.325 50.960 107.735 ;
        RECT 51.860 107.565 52.030 108.325 ;
        RECT 52.230 108.235 52.890 108.715 ;
        RECT 53.070 108.120 53.390 108.450 ;
        RECT 52.220 107.795 52.880 108.065 ;
        RECT 52.220 107.735 52.550 107.795 ;
        RECT 52.700 107.565 53.030 107.625 ;
        RECT 51.130 107.395 53.030 107.565 ;
        RECT 50.440 106.835 50.960 107.145 ;
        RECT 51.130 106.885 51.300 107.395 ;
        RECT 53.200 107.225 53.390 108.120 ;
        RECT 51.470 107.055 53.390 107.225 ;
        RECT 53.070 107.035 53.390 107.055 ;
        RECT 53.590 107.805 53.840 108.455 ;
        RECT 54.020 108.255 54.305 108.715 ;
        RECT 54.485 108.005 54.740 108.535 ;
        RECT 53.590 107.475 54.390 107.805 ;
        RECT 51.130 106.715 52.340 106.885 ;
        RECT 47.900 106.380 48.730 106.550 ;
        RECT 48.970 106.165 49.350 106.545 ;
        RECT 49.530 106.425 49.700 106.715 ;
        RECT 51.130 106.635 51.300 106.715 ;
        RECT 49.870 106.165 50.200 106.545 ;
        RECT 50.670 106.385 51.300 106.635 ;
        RECT 51.480 106.165 51.900 106.545 ;
        RECT 52.100 106.425 52.340 106.715 ;
        RECT 52.570 106.165 52.900 106.855 ;
        RECT 53.070 106.425 53.240 107.035 ;
        RECT 53.590 106.885 53.840 107.475 ;
        RECT 54.560 107.145 54.740 108.005 ;
        RECT 55.285 107.945 56.955 108.715 ;
        RECT 57.125 107.990 57.415 108.715 ;
        RECT 55.285 107.425 56.035 107.945 ;
        RECT 58.545 107.895 58.775 108.715 ;
        RECT 58.945 107.915 59.275 108.545 ;
        RECT 56.205 107.255 56.955 107.775 ;
        RECT 58.525 107.475 58.855 107.725 ;
        RECT 53.510 106.375 53.840 106.885 ;
        RECT 54.020 106.165 54.305 106.965 ;
        RECT 54.485 106.675 54.740 107.145 ;
        RECT 54.485 106.505 54.825 106.675 ;
        RECT 54.485 106.475 54.740 106.505 ;
        RECT 55.285 106.165 56.955 107.255 ;
        RECT 57.125 106.165 57.415 107.330 ;
        RECT 59.025 107.315 59.275 107.915 ;
        RECT 59.445 107.895 59.655 108.715 ;
        RECT 59.890 107.975 60.145 108.545 ;
        RECT 60.315 108.315 60.645 108.715 ;
        RECT 61.070 108.180 61.600 108.545 ;
        RECT 61.790 108.375 62.065 108.545 ;
        RECT 61.785 108.205 62.065 108.375 ;
        RECT 61.070 108.145 61.245 108.180 ;
        RECT 60.315 107.975 61.245 108.145 ;
        RECT 58.545 106.165 58.775 107.305 ;
        RECT 58.945 106.335 59.275 107.315 ;
        RECT 59.890 107.305 60.060 107.975 ;
        RECT 60.315 107.805 60.485 107.975 ;
        RECT 60.230 107.475 60.485 107.805 ;
        RECT 60.710 107.475 60.905 107.805 ;
        RECT 59.445 106.165 59.655 107.305 ;
        RECT 59.890 106.335 60.225 107.305 ;
        RECT 60.395 106.165 60.565 107.305 ;
        RECT 60.735 106.505 60.905 107.475 ;
        RECT 61.075 106.845 61.245 107.975 ;
        RECT 61.415 107.185 61.585 107.985 ;
        RECT 61.790 107.385 62.065 108.205 ;
        RECT 62.235 107.185 62.425 108.545 ;
        RECT 62.605 108.180 63.115 108.715 ;
        RECT 63.335 107.905 63.580 108.510 ;
        RECT 62.625 107.735 63.855 107.905 ;
        RECT 64.545 107.895 64.755 108.715 ;
        RECT 64.925 107.915 65.255 108.545 ;
        RECT 61.415 107.015 62.425 107.185 ;
        RECT 62.595 107.170 63.345 107.360 ;
        RECT 61.075 106.675 62.200 106.845 ;
        RECT 62.595 106.505 62.765 107.170 ;
        RECT 63.515 106.925 63.855 107.735 ;
        RECT 64.925 107.315 65.175 107.915 ;
        RECT 65.425 107.895 65.655 108.715 ;
        RECT 65.865 108.170 71.210 108.715 ;
        RECT 65.345 107.475 65.675 107.725 ;
        RECT 67.450 107.340 67.790 108.170 ;
        RECT 71.385 107.965 72.595 108.715 ;
        RECT 72.765 108.040 73.025 108.545 ;
        RECT 73.205 108.335 73.535 108.715 ;
        RECT 73.715 108.165 73.885 108.545 ;
        RECT 60.735 106.335 62.765 106.505 ;
        RECT 62.935 106.165 63.105 106.925 ;
        RECT 63.340 106.515 63.855 106.925 ;
        RECT 64.545 106.165 64.755 107.305 ;
        RECT 64.925 106.335 65.255 107.315 ;
        RECT 65.425 106.165 65.655 107.305 ;
        RECT 69.270 106.600 69.620 107.850 ;
        RECT 71.385 107.425 71.905 107.965 ;
        RECT 72.075 107.255 72.595 107.795 ;
        RECT 65.865 106.165 71.210 106.600 ;
        RECT 71.385 106.165 72.595 107.255 ;
        RECT 72.765 107.240 72.935 108.040 ;
        RECT 73.220 107.995 73.885 108.165 ;
        RECT 74.235 108.065 74.405 108.545 ;
        RECT 74.585 108.235 74.825 108.715 ;
        RECT 75.075 108.065 75.245 108.545 ;
        RECT 75.415 108.235 75.745 108.715 ;
        RECT 75.915 108.065 76.085 108.545 ;
        RECT 73.220 107.740 73.390 107.995 ;
        RECT 74.235 107.895 74.870 108.065 ;
        RECT 75.075 107.895 76.085 108.065 ;
        RECT 76.255 107.915 76.585 108.715 ;
        RECT 77.830 107.975 78.085 108.545 ;
        RECT 78.255 108.315 78.585 108.715 ;
        RECT 79.010 108.180 79.540 108.545 ;
        RECT 79.730 108.375 80.005 108.545 ;
        RECT 79.725 108.205 80.005 108.375 ;
        RECT 79.010 108.145 79.185 108.180 ;
        RECT 78.255 107.975 79.185 108.145 ;
        RECT 73.105 107.410 73.390 107.740 ;
        RECT 73.625 107.445 73.955 107.815 ;
        RECT 74.700 107.725 74.870 107.895 ;
        RECT 74.150 107.485 74.530 107.725 ;
        RECT 74.700 107.555 75.200 107.725 ;
        RECT 73.220 107.265 73.390 107.410 ;
        RECT 74.700 107.315 74.870 107.555 ;
        RECT 75.590 107.355 76.085 107.895 ;
        RECT 72.765 106.335 73.035 107.240 ;
        RECT 73.220 107.095 73.885 107.265 ;
        RECT 73.205 106.165 73.535 106.925 ;
        RECT 73.715 106.335 73.885 107.095 ;
        RECT 74.155 107.145 74.870 107.315 ;
        RECT 75.075 107.185 76.085 107.355 ;
        RECT 74.155 106.335 74.485 107.145 ;
        RECT 74.655 106.165 74.895 106.965 ;
        RECT 75.075 106.335 75.245 107.185 ;
        RECT 75.415 106.165 75.745 106.965 ;
        RECT 75.915 106.335 76.085 107.185 ;
        RECT 76.255 106.165 76.585 107.315 ;
        RECT 77.830 107.305 78.000 107.975 ;
        RECT 78.255 107.805 78.425 107.975 ;
        RECT 78.170 107.475 78.425 107.805 ;
        RECT 78.650 107.475 78.845 107.805 ;
        RECT 77.830 106.335 78.165 107.305 ;
        RECT 78.335 106.165 78.505 107.305 ;
        RECT 78.675 106.505 78.845 107.475 ;
        RECT 79.015 106.845 79.185 107.975 ;
        RECT 79.355 107.185 79.525 107.985 ;
        RECT 79.730 107.385 80.005 108.205 ;
        RECT 80.175 107.185 80.365 108.545 ;
        RECT 80.545 108.180 81.055 108.715 ;
        RECT 81.275 107.905 81.520 108.510 ;
        RECT 82.885 107.990 83.175 108.715 ;
        RECT 83.355 108.065 83.685 108.540 ;
        RECT 83.855 108.235 84.025 108.715 ;
        RECT 84.195 108.065 84.525 108.540 ;
        RECT 84.695 108.235 84.865 108.715 ;
        RECT 85.035 108.065 85.365 108.540 ;
        RECT 85.535 108.235 85.705 108.715 ;
        RECT 85.875 108.065 86.205 108.540 ;
        RECT 86.375 108.235 86.545 108.715 ;
        RECT 86.715 108.065 87.045 108.540 ;
        RECT 87.215 108.235 87.385 108.715 ;
        RECT 87.555 108.540 87.805 108.545 ;
        RECT 87.555 108.065 87.885 108.540 ;
        RECT 88.055 108.235 88.225 108.715 ;
        RECT 88.475 108.540 88.645 108.545 ;
        RECT 88.395 108.065 88.725 108.540 ;
        RECT 88.895 108.235 89.065 108.715 ;
        RECT 89.315 108.540 89.485 108.545 ;
        RECT 89.235 108.065 89.565 108.540 ;
        RECT 89.735 108.235 89.905 108.715 ;
        RECT 90.075 108.065 90.405 108.540 ;
        RECT 90.575 108.235 90.745 108.715 ;
        RECT 90.915 108.065 91.245 108.540 ;
        RECT 91.415 108.235 91.585 108.715 ;
        RECT 91.755 108.065 92.085 108.540 ;
        RECT 92.255 108.235 92.425 108.715 ;
        RECT 92.595 108.065 92.925 108.540 ;
        RECT 93.095 108.235 93.265 108.715 ;
        RECT 93.435 108.065 93.765 108.540 ;
        RECT 93.935 108.235 94.105 108.715 ;
        RECT 80.565 107.735 81.795 107.905 ;
        RECT 83.355 107.895 84.865 108.065 ;
        RECT 85.035 107.895 87.385 108.065 ;
        RECT 87.555 107.895 94.215 108.065 ;
        RECT 79.355 107.015 80.365 107.185 ;
        RECT 80.535 107.170 81.285 107.360 ;
        RECT 79.015 106.675 80.140 106.845 ;
        RECT 80.535 106.505 80.705 107.170 ;
        RECT 81.455 106.925 81.795 107.735 ;
        RECT 84.695 107.725 84.865 107.895 ;
        RECT 87.210 107.725 87.385 107.895 ;
        RECT 83.350 107.525 84.525 107.725 ;
        RECT 84.695 107.525 87.005 107.725 ;
        RECT 87.210 107.525 93.770 107.725 ;
        RECT 84.695 107.355 84.865 107.525 ;
        RECT 87.210 107.355 87.385 107.525 ;
        RECT 93.940 107.355 94.215 107.895 ;
        RECT 78.675 106.335 80.705 106.505 ;
        RECT 80.875 106.165 81.045 106.925 ;
        RECT 81.280 106.515 81.795 106.925 ;
        RECT 82.885 106.165 83.175 107.330 ;
        RECT 83.355 107.185 84.865 107.355 ;
        RECT 85.035 107.185 87.385 107.355 ;
        RECT 87.555 107.185 94.215 107.355 ;
        RECT 94.760 108.005 95.015 108.535 ;
        RECT 95.195 108.255 95.480 108.715 ;
        RECT 83.355 106.335 83.685 107.185 ;
        RECT 83.855 106.165 84.025 107.015 ;
        RECT 84.195 106.335 84.525 107.185 ;
        RECT 84.695 106.165 84.865 107.015 ;
        RECT 85.035 106.335 85.365 107.185 ;
        RECT 85.535 106.165 85.705 106.965 ;
        RECT 85.875 106.335 86.205 107.185 ;
        RECT 86.375 106.165 86.545 106.965 ;
        RECT 86.715 106.335 87.045 107.185 ;
        RECT 87.215 106.165 87.385 106.965 ;
        RECT 87.555 106.335 87.885 107.185 ;
        RECT 88.055 106.165 88.225 106.965 ;
        RECT 88.395 106.335 88.725 107.185 ;
        RECT 88.895 106.165 89.065 106.965 ;
        RECT 89.235 106.335 89.565 107.185 ;
        RECT 89.735 106.165 89.905 106.965 ;
        RECT 90.075 106.335 90.405 107.185 ;
        RECT 90.575 106.165 90.745 106.965 ;
        RECT 90.915 106.335 91.245 107.185 ;
        RECT 91.415 106.165 91.585 106.965 ;
        RECT 91.755 106.335 92.085 107.185 ;
        RECT 92.255 106.165 92.425 106.965 ;
        RECT 92.595 106.335 92.925 107.185 ;
        RECT 93.095 106.165 93.265 106.965 ;
        RECT 93.435 106.335 93.765 107.185 ;
        RECT 94.760 107.145 94.940 108.005 ;
        RECT 95.660 107.805 95.910 108.455 ;
        RECT 95.110 107.475 95.910 107.805 ;
        RECT 94.760 107.015 95.015 107.145 ;
        RECT 93.935 106.165 94.105 106.965 ;
        RECT 94.675 106.845 95.015 107.015 ;
        RECT 94.760 106.475 95.015 106.845 ;
        RECT 95.195 106.165 95.480 106.965 ;
        RECT 95.660 106.885 95.910 107.475 ;
        RECT 96.110 108.120 96.430 108.450 ;
        RECT 96.610 108.235 97.270 108.715 ;
        RECT 97.470 108.325 98.320 108.495 ;
        RECT 96.110 107.225 96.300 108.120 ;
        RECT 96.620 107.795 97.280 108.065 ;
        RECT 96.950 107.735 97.280 107.795 ;
        RECT 96.470 107.565 96.800 107.625 ;
        RECT 97.470 107.565 97.640 108.325 ;
        RECT 98.880 108.255 99.200 108.715 ;
        RECT 99.400 108.075 99.650 108.505 ;
        RECT 99.940 108.275 100.350 108.715 ;
        RECT 100.520 108.335 101.535 108.535 ;
        RECT 97.810 107.905 99.060 108.075 ;
        RECT 97.810 107.785 98.140 107.905 ;
        RECT 96.470 107.395 98.370 107.565 ;
        RECT 96.110 107.055 98.030 107.225 ;
        RECT 96.110 107.035 96.430 107.055 ;
        RECT 95.660 106.375 95.990 106.885 ;
        RECT 96.260 106.425 96.430 107.035 ;
        RECT 98.200 106.885 98.370 107.395 ;
        RECT 98.540 107.325 98.720 107.735 ;
        RECT 98.890 107.145 99.060 107.905 ;
        RECT 96.600 106.165 96.930 106.855 ;
        RECT 97.160 106.715 98.370 106.885 ;
        RECT 98.540 106.835 99.060 107.145 ;
        RECT 99.230 107.735 99.650 108.075 ;
        RECT 99.940 107.735 100.350 108.065 ;
        RECT 99.230 106.965 99.420 107.735 ;
        RECT 100.520 107.605 100.690 108.335 ;
        RECT 101.835 108.165 102.005 108.495 ;
        RECT 102.175 108.335 102.505 108.715 ;
        RECT 100.860 107.785 101.210 108.155 ;
        RECT 100.520 107.565 100.940 107.605 ;
        RECT 99.590 107.395 100.940 107.565 ;
        RECT 99.590 107.235 99.840 107.395 ;
        RECT 100.350 106.965 100.600 107.225 ;
        RECT 99.230 106.715 100.600 106.965 ;
        RECT 97.160 106.425 97.400 106.715 ;
        RECT 98.200 106.635 98.370 106.715 ;
        RECT 97.600 106.165 98.020 106.545 ;
        RECT 98.200 106.385 98.830 106.635 ;
        RECT 99.300 106.165 99.630 106.545 ;
        RECT 99.800 106.425 99.970 106.715 ;
        RECT 100.770 106.550 100.940 107.395 ;
        RECT 101.390 107.225 101.610 108.095 ;
        RECT 101.835 107.975 102.530 108.165 ;
        RECT 101.110 106.845 101.610 107.225 ;
        RECT 101.780 107.175 102.190 107.795 ;
        RECT 102.360 107.005 102.530 107.975 ;
        RECT 101.835 106.835 102.530 107.005 ;
        RECT 100.150 106.165 100.530 106.545 ;
        RECT 100.770 106.380 101.600 106.550 ;
        RECT 101.835 106.335 102.005 106.835 ;
        RECT 102.175 106.165 102.505 106.665 ;
        RECT 102.720 106.335 102.945 108.455 ;
        RECT 103.115 108.335 103.445 108.715 ;
        RECT 103.615 108.165 103.785 108.455 ;
        RECT 103.120 107.995 103.785 108.165 ;
        RECT 103.120 107.005 103.350 107.995 ;
        RECT 104.045 107.945 106.635 108.715 ;
        RECT 106.895 108.165 107.065 108.545 ;
        RECT 107.245 108.335 107.575 108.715 ;
        RECT 106.895 107.995 107.560 108.165 ;
        RECT 107.755 108.040 108.015 108.545 ;
        RECT 103.520 107.175 103.870 107.825 ;
        RECT 104.045 107.425 105.255 107.945 ;
        RECT 105.425 107.255 106.635 107.775 ;
        RECT 106.825 107.445 107.155 107.815 ;
        RECT 107.390 107.740 107.560 107.995 ;
        RECT 107.390 107.410 107.675 107.740 ;
        RECT 107.390 107.265 107.560 107.410 ;
        RECT 103.120 106.835 103.785 107.005 ;
        RECT 103.115 106.165 103.445 106.665 ;
        RECT 103.615 106.335 103.785 106.835 ;
        RECT 104.045 106.165 106.635 107.255 ;
        RECT 106.895 107.095 107.560 107.265 ;
        RECT 107.845 107.240 108.015 108.040 ;
        RECT 108.645 107.990 108.935 108.715 ;
        RECT 109.105 107.965 110.315 108.715 ;
        RECT 110.575 108.165 110.745 108.545 ;
        RECT 110.925 108.335 111.255 108.715 ;
        RECT 110.575 107.995 111.240 108.165 ;
        RECT 111.435 108.040 111.695 108.545 ;
        RECT 109.105 107.425 109.625 107.965 ;
        RECT 106.895 106.335 107.065 107.095 ;
        RECT 107.245 106.165 107.575 106.925 ;
        RECT 107.745 106.335 108.015 107.240 ;
        RECT 108.645 106.165 108.935 107.330 ;
        RECT 109.795 107.255 110.315 107.795 ;
        RECT 110.505 107.445 110.835 107.815 ;
        RECT 111.070 107.740 111.240 107.995 ;
        RECT 111.070 107.410 111.355 107.740 ;
        RECT 111.070 107.265 111.240 107.410 ;
        RECT 109.105 106.165 110.315 107.255 ;
        RECT 110.575 107.095 111.240 107.265 ;
        RECT 111.525 107.240 111.695 108.040 ;
        RECT 111.955 108.165 112.125 108.455 ;
        RECT 112.295 108.335 112.625 108.715 ;
        RECT 111.955 107.995 112.620 108.165 ;
        RECT 110.575 106.335 110.745 107.095 ;
        RECT 110.925 106.165 111.255 106.925 ;
        RECT 111.425 106.335 111.695 107.240 ;
        RECT 111.870 107.175 112.220 107.825 ;
        RECT 112.390 107.005 112.620 107.995 ;
        RECT 111.955 106.835 112.620 107.005 ;
        RECT 111.955 106.335 112.125 106.835 ;
        RECT 112.295 106.165 112.625 106.665 ;
        RECT 112.795 106.335 113.020 108.455 ;
        RECT 113.235 108.335 113.565 108.715 ;
        RECT 113.735 108.165 113.905 108.495 ;
        RECT 114.205 108.335 115.220 108.535 ;
        RECT 113.210 107.975 113.905 108.165 ;
        RECT 113.210 107.005 113.380 107.975 ;
        RECT 113.550 107.175 113.960 107.795 ;
        RECT 114.130 107.225 114.350 108.095 ;
        RECT 114.530 107.785 114.880 108.155 ;
        RECT 115.050 107.605 115.220 108.335 ;
        RECT 115.390 108.275 115.800 108.715 ;
        RECT 116.090 108.075 116.340 108.505 ;
        RECT 116.540 108.255 116.860 108.715 ;
        RECT 117.420 108.325 118.270 108.495 ;
        RECT 115.390 107.735 115.800 108.065 ;
        RECT 116.090 107.735 116.510 108.075 ;
        RECT 114.800 107.565 115.220 107.605 ;
        RECT 114.800 107.395 116.150 107.565 ;
        RECT 113.210 106.835 113.905 107.005 ;
        RECT 114.130 106.845 114.630 107.225 ;
        RECT 113.235 106.165 113.565 106.665 ;
        RECT 113.735 106.335 113.905 106.835 ;
        RECT 114.800 106.550 114.970 107.395 ;
        RECT 115.900 107.235 116.150 107.395 ;
        RECT 115.140 106.965 115.390 107.225 ;
        RECT 116.320 106.965 116.510 107.735 ;
        RECT 115.140 106.715 116.510 106.965 ;
        RECT 116.680 107.905 117.930 108.075 ;
        RECT 116.680 107.145 116.850 107.905 ;
        RECT 117.600 107.785 117.930 107.905 ;
        RECT 117.020 107.325 117.200 107.735 ;
        RECT 118.100 107.565 118.270 108.325 ;
        RECT 118.470 108.235 119.130 108.715 ;
        RECT 119.310 108.120 119.630 108.450 ;
        RECT 118.460 107.795 119.120 108.065 ;
        RECT 118.460 107.735 118.790 107.795 ;
        RECT 118.940 107.565 119.270 107.625 ;
        RECT 117.370 107.395 119.270 107.565 ;
        RECT 116.680 106.835 117.200 107.145 ;
        RECT 117.370 106.885 117.540 107.395 ;
        RECT 119.440 107.225 119.630 108.120 ;
        RECT 117.710 107.055 119.630 107.225 ;
        RECT 119.310 107.035 119.630 107.055 ;
        RECT 119.830 107.805 120.080 108.455 ;
        RECT 120.260 108.255 120.545 108.715 ;
        RECT 120.725 108.005 120.980 108.535 ;
        RECT 119.830 107.475 120.630 107.805 ;
        RECT 117.370 106.715 118.580 106.885 ;
        RECT 114.140 106.380 114.970 106.550 ;
        RECT 115.210 106.165 115.590 106.545 ;
        RECT 115.770 106.425 115.940 106.715 ;
        RECT 117.370 106.635 117.540 106.715 ;
        RECT 116.110 106.165 116.440 106.545 ;
        RECT 116.910 106.385 117.540 106.635 ;
        RECT 117.720 106.165 118.140 106.545 ;
        RECT 118.340 106.425 118.580 106.715 ;
        RECT 118.810 106.165 119.140 106.855 ;
        RECT 119.310 106.425 119.480 107.035 ;
        RECT 119.830 106.885 120.080 107.475 ;
        RECT 120.800 107.145 120.980 108.005 ;
        RECT 122.445 107.965 123.655 108.715 ;
        RECT 119.750 106.375 120.080 106.885 ;
        RECT 120.260 106.165 120.545 106.965 ;
        RECT 120.725 106.675 120.980 107.145 ;
        RECT 122.445 107.255 122.965 107.795 ;
        RECT 123.135 107.425 123.655 107.965 ;
        RECT 120.725 106.505 121.065 106.675 ;
        RECT 120.725 106.475 120.980 106.505 ;
        RECT 122.445 106.165 123.655 107.255 ;
        RECT 5.520 105.995 123.740 106.165 ;
        RECT 5.605 104.905 6.815 105.995 ;
        RECT 6.985 104.905 10.495 105.995 ;
        RECT 5.605 104.195 6.125 104.735 ;
        RECT 6.295 104.365 6.815 104.905 ;
        RECT 6.985 104.215 8.635 104.735 ;
        RECT 8.805 104.385 10.495 104.905 ;
        RECT 11.585 104.920 11.855 105.825 ;
        RECT 12.025 105.235 12.355 105.995 ;
        RECT 12.535 105.065 12.705 105.825 ;
        RECT 5.605 103.445 6.815 104.195 ;
        RECT 6.985 103.445 10.495 104.215 ;
        RECT 11.585 104.120 11.755 104.920 ;
        RECT 12.040 104.895 12.705 105.065 ;
        RECT 12.040 104.750 12.210 104.895 ;
        RECT 13.025 104.855 13.235 105.995 ;
        RECT 11.925 104.420 12.210 104.750 ;
        RECT 13.405 104.845 13.735 105.825 ;
        RECT 13.905 104.855 14.135 105.995 ;
        RECT 14.350 104.855 14.685 105.825 ;
        RECT 14.855 104.855 15.025 105.995 ;
        RECT 15.195 105.655 17.225 105.825 ;
        RECT 12.040 104.165 12.210 104.420 ;
        RECT 12.445 104.345 12.775 104.715 ;
        RECT 11.585 103.615 11.845 104.120 ;
        RECT 12.040 103.995 12.705 104.165 ;
        RECT 12.025 103.445 12.355 103.825 ;
        RECT 12.535 103.615 12.705 103.995 ;
        RECT 13.025 103.445 13.235 104.265 ;
        RECT 13.405 104.245 13.655 104.845 ;
        RECT 13.825 104.435 14.155 104.685 ;
        RECT 13.405 103.615 13.735 104.245 ;
        RECT 13.905 103.445 14.135 104.265 ;
        RECT 14.350 104.185 14.520 104.855 ;
        RECT 15.195 104.685 15.365 105.655 ;
        RECT 14.690 104.355 14.945 104.685 ;
        RECT 15.170 104.355 15.365 104.685 ;
        RECT 15.535 105.315 16.660 105.485 ;
        RECT 14.775 104.185 14.945 104.355 ;
        RECT 15.535 104.185 15.705 105.315 ;
        RECT 14.350 103.615 14.605 104.185 ;
        RECT 14.775 104.015 15.705 104.185 ;
        RECT 15.875 104.975 16.885 105.145 ;
        RECT 15.875 104.175 16.045 104.975 ;
        RECT 15.530 103.980 15.705 104.015 ;
        RECT 14.775 103.445 15.105 103.845 ;
        RECT 15.530 103.615 16.060 103.980 ;
        RECT 16.250 103.955 16.525 104.775 ;
        RECT 16.245 103.785 16.525 103.955 ;
        RECT 16.250 103.615 16.525 103.785 ;
        RECT 16.695 103.615 16.885 104.975 ;
        RECT 17.055 104.990 17.225 105.655 ;
        RECT 17.395 105.235 17.565 105.995 ;
        RECT 17.800 105.235 18.315 105.645 ;
        RECT 17.055 104.800 17.805 104.990 ;
        RECT 17.975 104.425 18.315 105.235 ;
        RECT 18.485 104.830 18.775 105.995 ;
        RECT 18.945 104.905 20.615 105.995 ;
        RECT 17.085 104.255 18.315 104.425 ;
        RECT 17.065 103.445 17.575 103.980 ;
        RECT 17.795 103.650 18.040 104.255 ;
        RECT 18.945 104.215 19.695 104.735 ;
        RECT 19.865 104.385 20.615 104.905 ;
        RECT 21.250 104.855 21.585 105.825 ;
        RECT 21.755 104.855 21.925 105.995 ;
        RECT 22.095 105.655 24.125 105.825 ;
        RECT 18.485 103.445 18.775 104.170 ;
        RECT 18.945 103.445 20.615 104.215 ;
        RECT 21.250 104.185 21.420 104.855 ;
        RECT 22.095 104.685 22.265 105.655 ;
        RECT 21.590 104.355 21.845 104.685 ;
        RECT 22.070 104.355 22.265 104.685 ;
        RECT 22.435 105.315 23.560 105.485 ;
        RECT 21.675 104.185 21.845 104.355 ;
        RECT 22.435 104.185 22.605 105.315 ;
        RECT 21.250 103.615 21.505 104.185 ;
        RECT 21.675 104.015 22.605 104.185 ;
        RECT 22.775 104.975 23.785 105.145 ;
        RECT 22.775 104.175 22.945 104.975 ;
        RECT 23.150 104.635 23.425 104.775 ;
        RECT 23.145 104.465 23.425 104.635 ;
        RECT 22.430 103.980 22.605 104.015 ;
        RECT 21.675 103.445 22.005 103.845 ;
        RECT 22.430 103.615 22.960 103.980 ;
        RECT 23.150 103.615 23.425 104.465 ;
        RECT 23.595 103.615 23.785 104.975 ;
        RECT 23.955 104.990 24.125 105.655 ;
        RECT 24.295 105.235 24.465 105.995 ;
        RECT 24.700 105.235 25.215 105.645 ;
        RECT 23.955 104.800 24.705 104.990 ;
        RECT 24.875 104.425 25.215 105.235 ;
        RECT 25.395 105.185 25.690 105.995 ;
        RECT 25.870 104.685 26.115 105.825 ;
        RECT 26.290 105.185 26.550 105.995 ;
        RECT 27.150 105.990 33.425 105.995 ;
        RECT 26.730 104.685 26.980 105.820 ;
        RECT 27.150 105.195 27.410 105.990 ;
        RECT 27.580 105.095 27.840 105.820 ;
        RECT 28.010 105.265 28.270 105.990 ;
        RECT 28.440 105.095 28.700 105.820 ;
        RECT 28.870 105.265 29.130 105.990 ;
        RECT 29.300 105.095 29.560 105.820 ;
        RECT 29.730 105.265 29.990 105.990 ;
        RECT 30.160 105.095 30.420 105.820 ;
        RECT 30.590 105.265 30.835 105.990 ;
        RECT 31.005 105.095 31.265 105.820 ;
        RECT 31.450 105.265 31.695 105.990 ;
        RECT 31.865 105.095 32.125 105.820 ;
        RECT 32.310 105.265 32.555 105.990 ;
        RECT 32.725 105.095 32.985 105.820 ;
        RECT 33.170 105.265 33.425 105.990 ;
        RECT 27.580 105.080 32.985 105.095 ;
        RECT 33.595 105.080 33.885 105.820 ;
        RECT 34.055 105.250 34.325 105.995 ;
        RECT 27.580 104.855 34.325 105.080 ;
        RECT 34.585 104.905 35.795 105.995 ;
        RECT 23.985 104.255 25.215 104.425 ;
        RECT 23.965 103.445 24.475 103.980 ;
        RECT 24.695 103.650 24.940 104.255 ;
        RECT 25.385 104.125 25.700 104.685 ;
        RECT 25.870 104.435 32.990 104.685 ;
        RECT 25.385 103.445 25.690 103.955 ;
        RECT 25.870 103.625 26.120 104.435 ;
        RECT 26.290 103.445 26.550 103.970 ;
        RECT 26.730 103.625 26.980 104.435 ;
        RECT 33.160 104.265 34.325 104.855 ;
        RECT 27.580 104.095 34.325 104.265 ;
        RECT 34.585 104.195 35.105 104.735 ;
        RECT 35.275 104.365 35.795 104.905 ;
        RECT 35.970 104.855 36.305 105.825 ;
        RECT 36.475 104.855 36.645 105.995 ;
        RECT 36.815 105.655 38.845 105.825 ;
        RECT 27.150 103.445 27.410 104.005 ;
        RECT 27.580 103.640 27.840 104.095 ;
        RECT 28.010 103.445 28.270 103.925 ;
        RECT 28.440 103.640 28.700 104.095 ;
        RECT 28.870 103.445 29.130 103.925 ;
        RECT 29.300 103.640 29.560 104.095 ;
        RECT 29.730 103.445 29.975 103.925 ;
        RECT 30.145 103.640 30.420 104.095 ;
        RECT 30.590 103.445 30.835 103.925 ;
        RECT 31.005 103.640 31.265 104.095 ;
        RECT 31.445 103.445 31.695 103.925 ;
        RECT 31.865 103.640 32.125 104.095 ;
        RECT 32.305 103.445 32.555 103.925 ;
        RECT 32.725 103.640 32.985 104.095 ;
        RECT 33.165 103.445 33.425 103.925 ;
        RECT 33.595 103.640 33.855 104.095 ;
        RECT 34.025 103.445 34.325 103.925 ;
        RECT 34.585 103.445 35.795 104.195 ;
        RECT 35.970 104.185 36.140 104.855 ;
        RECT 36.815 104.685 36.985 105.655 ;
        RECT 36.310 104.355 36.565 104.685 ;
        RECT 36.790 104.355 36.985 104.685 ;
        RECT 37.155 105.315 38.280 105.485 ;
        RECT 36.395 104.185 36.565 104.355 ;
        RECT 37.155 104.185 37.325 105.315 ;
        RECT 35.970 103.615 36.225 104.185 ;
        RECT 36.395 104.015 37.325 104.185 ;
        RECT 37.495 104.975 38.505 105.145 ;
        RECT 37.495 104.175 37.665 104.975 ;
        RECT 37.870 104.295 38.145 104.775 ;
        RECT 37.865 104.125 38.145 104.295 ;
        RECT 37.150 103.980 37.325 104.015 ;
        RECT 36.395 103.445 36.725 103.845 ;
        RECT 37.150 103.615 37.680 103.980 ;
        RECT 37.870 103.615 38.145 104.125 ;
        RECT 38.315 103.615 38.505 104.975 ;
        RECT 38.675 104.990 38.845 105.655 ;
        RECT 39.015 105.235 39.185 105.995 ;
        RECT 39.420 105.235 39.935 105.645 ;
        RECT 38.675 104.800 39.425 104.990 ;
        RECT 39.595 104.425 39.935 105.235 ;
        RECT 40.105 104.905 41.315 105.995 ;
        RECT 38.705 104.255 39.935 104.425 ;
        RECT 38.685 103.445 39.195 103.980 ;
        RECT 39.415 103.650 39.660 104.255 ;
        RECT 40.105 104.195 40.625 104.735 ;
        RECT 40.795 104.365 41.315 104.905 ;
        RECT 41.485 105.025 41.795 105.825 ;
        RECT 41.965 105.195 42.275 105.995 ;
        RECT 42.445 105.365 42.705 105.825 ;
        RECT 42.875 105.535 43.130 105.995 ;
        RECT 43.305 105.365 43.565 105.825 ;
        RECT 42.445 105.195 43.565 105.365 ;
        RECT 41.485 104.855 42.515 105.025 ;
        RECT 40.105 103.445 41.315 104.195 ;
        RECT 41.485 103.945 41.655 104.855 ;
        RECT 41.825 104.115 42.175 104.685 ;
        RECT 42.345 104.605 42.515 104.855 ;
        RECT 43.305 104.945 43.565 105.195 ;
        RECT 43.735 105.125 44.020 105.995 ;
        RECT 43.305 104.775 44.060 104.945 ;
        RECT 44.245 104.830 44.535 105.995 ;
        RECT 44.715 105.185 45.010 105.995 ;
        RECT 42.345 104.435 43.485 104.605 ;
        RECT 43.655 104.265 44.060 104.775 ;
        RECT 45.190 104.685 45.435 105.825 ;
        RECT 45.610 105.185 45.870 105.995 ;
        RECT 46.470 105.990 52.745 105.995 ;
        RECT 46.050 104.685 46.300 105.820 ;
        RECT 46.470 105.195 46.730 105.990 ;
        RECT 46.900 105.095 47.160 105.820 ;
        RECT 47.330 105.265 47.590 105.990 ;
        RECT 47.760 105.095 48.020 105.820 ;
        RECT 48.190 105.265 48.450 105.990 ;
        RECT 48.620 105.095 48.880 105.820 ;
        RECT 49.050 105.265 49.310 105.990 ;
        RECT 49.480 105.095 49.740 105.820 ;
        RECT 49.910 105.265 50.155 105.990 ;
        RECT 50.325 105.095 50.585 105.820 ;
        RECT 50.770 105.265 51.015 105.990 ;
        RECT 51.185 105.095 51.445 105.820 ;
        RECT 51.630 105.265 51.875 105.990 ;
        RECT 52.045 105.095 52.305 105.820 ;
        RECT 52.490 105.265 52.745 105.990 ;
        RECT 46.900 105.080 52.305 105.095 ;
        RECT 52.915 105.080 53.205 105.820 ;
        RECT 53.375 105.250 53.645 105.995 ;
        RECT 46.900 104.855 53.645 105.080 ;
        RECT 42.410 104.095 44.060 104.265 ;
        RECT 41.485 103.615 41.785 103.945 ;
        RECT 41.955 103.445 42.230 103.925 ;
        RECT 42.410 103.705 42.705 104.095 ;
        RECT 42.875 103.445 43.130 103.925 ;
        RECT 43.305 103.705 43.565 104.095 ;
        RECT 43.735 103.445 44.015 103.925 ;
        RECT 44.245 103.445 44.535 104.170 ;
        RECT 44.705 104.125 45.020 104.685 ;
        RECT 45.190 104.435 52.310 104.685 ;
        RECT 44.705 103.445 45.010 103.955 ;
        RECT 45.190 103.625 45.440 104.435 ;
        RECT 45.610 103.445 45.870 103.970 ;
        RECT 46.050 103.625 46.300 104.435 ;
        RECT 52.480 104.265 53.645 104.855 ;
        RECT 46.900 104.095 53.645 104.265 ;
        RECT 53.910 104.855 54.245 105.825 ;
        RECT 54.415 104.855 54.585 105.995 ;
        RECT 54.755 105.655 56.785 105.825 ;
        RECT 53.910 104.185 54.080 104.855 ;
        RECT 54.755 104.685 54.925 105.655 ;
        RECT 54.250 104.355 54.505 104.685 ;
        RECT 54.730 104.355 54.925 104.685 ;
        RECT 55.095 105.315 56.220 105.485 ;
        RECT 54.335 104.185 54.505 104.355 ;
        RECT 55.095 104.185 55.265 105.315 ;
        RECT 46.470 103.445 46.730 104.005 ;
        RECT 46.900 103.640 47.160 104.095 ;
        RECT 47.330 103.445 47.590 103.925 ;
        RECT 47.760 103.640 48.020 104.095 ;
        RECT 48.190 103.445 48.450 103.925 ;
        RECT 48.620 103.640 48.880 104.095 ;
        RECT 49.050 103.445 49.295 103.925 ;
        RECT 49.465 103.640 49.740 104.095 ;
        RECT 49.910 103.445 50.155 103.925 ;
        RECT 50.325 103.640 50.585 104.095 ;
        RECT 50.765 103.445 51.015 103.925 ;
        RECT 51.185 103.640 51.445 104.095 ;
        RECT 51.625 103.445 51.875 103.925 ;
        RECT 52.045 103.640 52.305 104.095 ;
        RECT 52.485 103.445 52.745 103.925 ;
        RECT 52.915 103.640 53.175 104.095 ;
        RECT 53.345 103.445 53.645 103.925 ;
        RECT 53.910 103.615 54.165 104.185 ;
        RECT 54.335 104.015 55.265 104.185 ;
        RECT 55.435 104.975 56.445 105.145 ;
        RECT 55.435 104.175 55.605 104.975 ;
        RECT 55.810 104.635 56.085 104.775 ;
        RECT 55.805 104.465 56.085 104.635 ;
        RECT 55.090 103.980 55.265 104.015 ;
        RECT 54.335 103.445 54.665 103.845 ;
        RECT 55.090 103.615 55.620 103.980 ;
        RECT 55.810 103.615 56.085 104.465 ;
        RECT 56.255 103.615 56.445 104.975 ;
        RECT 56.615 104.990 56.785 105.655 ;
        RECT 56.955 105.235 57.125 105.995 ;
        RECT 57.360 105.235 57.875 105.645 ;
        RECT 56.615 104.800 57.365 104.990 ;
        RECT 57.535 104.425 57.875 105.235 ;
        RECT 56.645 104.255 57.875 104.425 ;
        RECT 58.045 105.275 58.505 105.825 ;
        RECT 58.695 105.275 59.025 105.995 ;
        RECT 56.625 103.445 57.135 103.980 ;
        RECT 57.355 103.650 57.600 104.255 ;
        RECT 58.045 103.905 58.295 105.275 ;
        RECT 59.225 105.105 59.525 105.655 ;
        RECT 59.695 105.325 59.975 105.995 ;
        RECT 60.345 105.560 65.690 105.995 ;
        RECT 58.585 104.935 59.525 105.105 ;
        RECT 58.585 104.685 58.755 104.935 ;
        RECT 59.895 104.685 60.160 105.045 ;
        RECT 58.465 104.355 58.755 104.685 ;
        RECT 58.925 104.435 59.265 104.685 ;
        RECT 59.485 104.435 60.160 104.685 ;
        RECT 58.585 104.265 58.755 104.355 ;
        RECT 58.585 104.075 59.975 104.265 ;
        RECT 58.045 103.615 58.605 103.905 ;
        RECT 58.775 103.445 59.025 103.905 ;
        RECT 59.645 103.715 59.975 104.075 ;
        RECT 61.930 103.990 62.270 104.820 ;
        RECT 63.750 104.310 64.100 105.560 ;
        RECT 65.920 105.125 66.205 105.995 ;
        RECT 66.375 105.365 66.635 105.825 ;
        RECT 66.810 105.535 67.065 105.995 ;
        RECT 67.235 105.365 67.495 105.825 ;
        RECT 66.375 105.195 67.495 105.365 ;
        RECT 67.665 105.195 67.975 105.995 ;
        RECT 66.375 104.945 66.635 105.195 ;
        RECT 68.145 105.025 68.455 105.825 ;
        RECT 65.880 104.775 66.635 104.945 ;
        RECT 67.425 104.855 68.455 105.025 ;
        RECT 68.625 104.905 69.835 105.995 ;
        RECT 65.880 104.265 66.285 104.775 ;
        RECT 67.425 104.605 67.595 104.855 ;
        RECT 66.455 104.435 67.595 104.605 ;
        RECT 65.880 104.095 67.530 104.265 ;
        RECT 67.765 104.115 68.115 104.685 ;
        RECT 60.345 103.445 65.690 103.990 ;
        RECT 65.925 103.445 66.205 103.925 ;
        RECT 66.375 103.705 66.635 104.095 ;
        RECT 66.810 103.445 67.065 103.925 ;
        RECT 67.235 103.705 67.530 104.095 ;
        RECT 68.285 103.945 68.455 104.855 ;
        RECT 67.710 103.445 67.985 103.925 ;
        RECT 68.155 103.615 68.455 103.945 ;
        RECT 68.625 104.195 69.145 104.735 ;
        RECT 69.315 104.365 69.835 104.905 ;
        RECT 70.005 104.830 70.295 105.995 ;
        RECT 70.465 104.905 71.675 105.995 ;
        RECT 70.465 104.195 70.985 104.735 ;
        RECT 71.155 104.365 71.675 104.905 ;
        RECT 71.845 105.025 72.155 105.825 ;
        RECT 72.325 105.195 72.635 105.995 ;
        RECT 72.805 105.365 73.065 105.825 ;
        RECT 73.235 105.535 73.490 105.995 ;
        RECT 73.665 105.365 73.925 105.825 ;
        RECT 72.805 105.195 73.925 105.365 ;
        RECT 71.845 104.855 72.875 105.025 ;
        RECT 68.625 103.445 69.835 104.195 ;
        RECT 70.005 103.445 70.295 104.170 ;
        RECT 70.465 103.445 71.675 104.195 ;
        RECT 71.845 103.945 72.015 104.855 ;
        RECT 72.185 104.115 72.535 104.685 ;
        RECT 72.705 104.605 72.875 104.855 ;
        RECT 73.665 104.945 73.925 105.195 ;
        RECT 74.095 105.125 74.380 105.995 ;
        RECT 73.665 104.775 74.420 104.945 ;
        RECT 74.605 104.905 75.815 105.995 ;
        RECT 72.705 104.435 73.845 104.605 ;
        RECT 74.015 104.265 74.420 104.775 ;
        RECT 72.770 104.095 74.420 104.265 ;
        RECT 74.605 104.195 75.125 104.735 ;
        RECT 75.295 104.365 75.815 104.905 ;
        RECT 76.045 104.855 76.255 105.995 ;
        RECT 76.425 104.845 76.755 105.825 ;
        RECT 76.925 104.855 77.155 105.995 ;
        RECT 77.365 104.905 78.575 105.995 ;
        RECT 78.945 105.325 79.225 105.995 ;
        RECT 79.395 105.105 79.695 105.655 ;
        RECT 79.895 105.275 80.225 105.995 ;
        RECT 80.415 105.275 80.875 105.825 ;
        RECT 71.845 103.615 72.145 103.945 ;
        RECT 72.315 103.445 72.590 103.925 ;
        RECT 72.770 103.705 73.065 104.095 ;
        RECT 73.235 103.445 73.490 103.925 ;
        RECT 73.665 103.705 73.925 104.095 ;
        RECT 74.095 103.445 74.375 103.925 ;
        RECT 74.605 103.445 75.815 104.195 ;
        RECT 76.045 103.445 76.255 104.265 ;
        RECT 76.425 104.245 76.675 104.845 ;
        RECT 76.845 104.435 77.175 104.685 ;
        RECT 76.425 103.615 76.755 104.245 ;
        RECT 76.925 103.445 77.155 104.265 ;
        RECT 77.365 104.195 77.885 104.735 ;
        RECT 78.055 104.365 78.575 104.905 ;
        RECT 78.760 104.685 79.025 105.045 ;
        RECT 79.395 104.935 80.335 105.105 ;
        RECT 80.165 104.685 80.335 104.935 ;
        RECT 78.760 104.435 79.435 104.685 ;
        RECT 79.655 104.435 79.995 104.685 ;
        RECT 80.165 104.355 80.455 104.685 ;
        RECT 80.165 104.265 80.335 104.355 ;
        RECT 77.365 103.445 78.575 104.195 ;
        RECT 78.945 104.075 80.335 104.265 ;
        RECT 78.945 103.715 79.275 104.075 ;
        RECT 80.625 103.905 80.875 105.275 ;
        RECT 81.135 105.325 81.305 105.825 ;
        RECT 81.475 105.495 81.805 105.995 ;
        RECT 81.135 105.155 81.800 105.325 ;
        RECT 81.050 104.335 81.400 104.985 ;
        RECT 81.570 104.165 81.800 105.155 ;
        RECT 79.895 103.445 80.145 103.905 ;
        RECT 80.315 103.615 80.875 103.905 ;
        RECT 81.135 103.995 81.800 104.165 ;
        RECT 81.135 103.705 81.305 103.995 ;
        RECT 81.475 103.445 81.805 103.825 ;
        RECT 81.975 103.705 82.200 105.825 ;
        RECT 82.415 105.495 82.745 105.995 ;
        RECT 82.915 105.325 83.085 105.825 ;
        RECT 83.320 105.610 84.150 105.780 ;
        RECT 84.390 105.615 84.770 105.995 ;
        RECT 82.390 105.155 83.085 105.325 ;
        RECT 82.390 104.185 82.560 105.155 ;
        RECT 82.730 104.365 83.140 104.985 ;
        RECT 83.310 104.935 83.810 105.315 ;
        RECT 82.390 103.995 83.085 104.185 ;
        RECT 83.310 104.065 83.530 104.935 ;
        RECT 83.980 104.765 84.150 105.610 ;
        RECT 84.950 105.445 85.120 105.735 ;
        RECT 85.290 105.615 85.620 105.995 ;
        RECT 86.090 105.525 86.720 105.775 ;
        RECT 86.900 105.615 87.320 105.995 ;
        RECT 86.550 105.445 86.720 105.525 ;
        RECT 87.520 105.445 87.760 105.735 ;
        RECT 84.320 105.195 85.690 105.445 ;
        RECT 84.320 104.935 84.570 105.195 ;
        RECT 85.080 104.765 85.330 104.925 ;
        RECT 83.980 104.595 85.330 104.765 ;
        RECT 83.980 104.555 84.400 104.595 ;
        RECT 83.710 104.005 84.060 104.375 ;
        RECT 82.415 103.445 82.745 103.825 ;
        RECT 82.915 103.665 83.085 103.995 ;
        RECT 84.230 103.825 84.400 104.555 ;
        RECT 85.500 104.425 85.690 105.195 ;
        RECT 84.570 104.095 84.980 104.425 ;
        RECT 85.270 104.085 85.690 104.425 ;
        RECT 85.860 105.015 86.380 105.325 ;
        RECT 86.550 105.275 87.760 105.445 ;
        RECT 87.990 105.305 88.320 105.995 ;
        RECT 85.860 104.255 86.030 105.015 ;
        RECT 86.200 104.425 86.380 104.835 ;
        RECT 86.550 104.765 86.720 105.275 ;
        RECT 88.490 105.125 88.660 105.735 ;
        RECT 88.930 105.275 89.260 105.785 ;
        RECT 88.490 105.105 88.810 105.125 ;
        RECT 86.890 104.935 88.810 105.105 ;
        RECT 86.550 104.595 88.450 104.765 ;
        RECT 86.780 104.255 87.110 104.375 ;
        RECT 85.860 104.085 87.110 104.255 ;
        RECT 83.385 103.625 84.400 103.825 ;
        RECT 84.570 103.445 84.980 103.885 ;
        RECT 85.270 103.655 85.520 104.085 ;
        RECT 85.720 103.445 86.040 103.905 ;
        RECT 87.280 103.835 87.450 104.595 ;
        RECT 88.120 104.535 88.450 104.595 ;
        RECT 87.640 104.365 87.970 104.425 ;
        RECT 87.640 104.095 88.300 104.365 ;
        RECT 88.620 104.040 88.810 104.935 ;
        RECT 86.600 103.665 87.450 103.835 ;
        RECT 87.650 103.445 88.310 103.925 ;
        RECT 88.490 103.710 88.810 104.040 ;
        RECT 89.010 104.685 89.260 105.275 ;
        RECT 89.440 105.195 89.725 105.995 ;
        RECT 89.905 105.015 90.160 105.685 ;
        RECT 89.010 104.355 89.810 104.685 ;
        RECT 89.010 103.705 89.260 104.355 ;
        RECT 89.980 104.155 90.160 105.015 ;
        RECT 89.905 103.955 90.160 104.155 ;
        RECT 90.705 105.275 91.165 105.825 ;
        RECT 91.355 105.275 91.685 105.995 ;
        RECT 89.440 103.445 89.725 103.905 ;
        RECT 89.905 103.785 90.245 103.955 ;
        RECT 90.705 103.905 90.955 105.275 ;
        RECT 91.885 105.105 92.185 105.655 ;
        RECT 92.355 105.325 92.635 105.995 ;
        RECT 91.245 104.935 92.185 105.105 ;
        RECT 91.245 104.685 91.415 104.935 ;
        RECT 92.555 104.685 92.820 105.045 ;
        RECT 93.005 104.905 95.595 105.995 ;
        RECT 91.125 104.355 91.415 104.685 ;
        RECT 91.585 104.435 91.925 104.685 ;
        RECT 92.145 104.435 92.820 104.685 ;
        RECT 91.245 104.265 91.415 104.355 ;
        RECT 91.245 104.075 92.635 104.265 ;
        RECT 89.905 103.625 90.160 103.785 ;
        RECT 90.705 103.615 91.265 103.905 ;
        RECT 91.435 103.445 91.685 103.905 ;
        RECT 92.305 103.715 92.635 104.075 ;
        RECT 93.005 104.215 94.215 104.735 ;
        RECT 94.385 104.385 95.595 104.905 ;
        RECT 95.765 104.830 96.055 105.995 ;
        RECT 96.225 104.905 98.815 105.995 ;
        RECT 96.225 104.215 97.435 104.735 ;
        RECT 97.605 104.385 98.815 104.905 ;
        RECT 99.025 104.855 99.255 105.995 ;
        RECT 99.425 104.845 99.755 105.825 ;
        RECT 99.925 104.855 100.135 105.995 ;
        RECT 100.375 105.185 100.670 105.995 ;
        RECT 99.005 104.435 99.335 104.685 ;
        RECT 93.005 103.445 95.595 104.215 ;
        RECT 95.765 103.445 96.055 104.170 ;
        RECT 96.225 103.445 98.815 104.215 ;
        RECT 99.025 103.445 99.255 104.265 ;
        RECT 99.505 104.245 99.755 104.845 ;
        RECT 100.850 104.685 101.095 105.825 ;
        RECT 101.270 105.185 101.530 105.995 ;
        RECT 102.130 105.990 108.405 105.995 ;
        RECT 101.710 104.685 101.960 105.820 ;
        RECT 102.130 105.195 102.390 105.990 ;
        RECT 102.560 105.095 102.820 105.820 ;
        RECT 102.990 105.265 103.250 105.990 ;
        RECT 103.420 105.095 103.680 105.820 ;
        RECT 103.850 105.265 104.110 105.990 ;
        RECT 104.280 105.095 104.540 105.820 ;
        RECT 104.710 105.265 104.970 105.990 ;
        RECT 105.140 105.095 105.400 105.820 ;
        RECT 105.570 105.265 105.815 105.990 ;
        RECT 105.985 105.095 106.245 105.820 ;
        RECT 106.430 105.265 106.675 105.990 ;
        RECT 106.845 105.095 107.105 105.820 ;
        RECT 107.290 105.265 107.535 105.990 ;
        RECT 107.705 105.095 107.965 105.820 ;
        RECT 108.150 105.265 108.405 105.990 ;
        RECT 102.560 105.080 107.965 105.095 ;
        RECT 108.575 105.080 108.865 105.820 ;
        RECT 109.035 105.250 109.305 105.995 ;
        RECT 102.560 104.855 109.305 105.080 ;
        RECT 109.565 104.905 112.155 105.995 ;
        RECT 99.425 103.615 99.755 104.245 ;
        RECT 99.925 103.445 100.135 104.265 ;
        RECT 100.365 104.125 100.680 104.685 ;
        RECT 100.850 104.435 107.970 104.685 ;
        RECT 100.365 103.445 100.670 103.955 ;
        RECT 100.850 103.625 101.100 104.435 ;
        RECT 101.270 103.445 101.530 103.970 ;
        RECT 101.710 103.625 101.960 104.435 ;
        RECT 108.140 104.295 109.305 104.855 ;
        RECT 108.140 104.265 109.335 104.295 ;
        RECT 102.560 104.125 109.335 104.265 ;
        RECT 109.565 104.215 110.775 104.735 ;
        RECT 110.945 104.385 112.155 104.905 ;
        RECT 112.330 104.855 112.665 105.825 ;
        RECT 112.835 104.855 113.005 105.995 ;
        RECT 113.175 105.655 115.205 105.825 ;
        RECT 102.560 104.095 109.305 104.125 ;
        RECT 102.130 103.445 102.390 104.005 ;
        RECT 102.560 103.640 102.820 104.095 ;
        RECT 102.990 103.445 103.250 103.925 ;
        RECT 103.420 103.640 103.680 104.095 ;
        RECT 103.850 103.445 104.110 103.925 ;
        RECT 104.280 103.640 104.540 104.095 ;
        RECT 104.710 103.445 104.955 103.925 ;
        RECT 105.125 103.640 105.400 104.095 ;
        RECT 105.570 103.445 105.815 103.925 ;
        RECT 105.985 103.640 106.245 104.095 ;
        RECT 106.425 103.445 106.675 103.925 ;
        RECT 106.845 103.640 107.105 104.095 ;
        RECT 107.285 103.445 107.535 103.925 ;
        RECT 107.705 103.640 107.965 104.095 ;
        RECT 108.145 103.445 108.405 103.925 ;
        RECT 108.575 103.640 108.835 104.095 ;
        RECT 109.005 103.445 109.305 103.925 ;
        RECT 109.565 103.445 112.155 104.215 ;
        RECT 112.330 104.185 112.500 104.855 ;
        RECT 113.175 104.685 113.345 105.655 ;
        RECT 112.670 104.355 112.925 104.685 ;
        RECT 113.150 104.355 113.345 104.685 ;
        RECT 113.515 105.315 114.640 105.485 ;
        RECT 112.755 104.185 112.925 104.355 ;
        RECT 113.515 104.185 113.685 105.315 ;
        RECT 112.330 103.615 112.585 104.185 ;
        RECT 112.755 104.015 113.685 104.185 ;
        RECT 113.855 104.975 114.865 105.145 ;
        RECT 113.855 104.175 114.025 104.975 ;
        RECT 114.230 104.635 114.505 104.775 ;
        RECT 114.225 104.465 114.505 104.635 ;
        RECT 113.510 103.980 113.685 104.015 ;
        RECT 112.755 103.445 113.085 103.845 ;
        RECT 113.510 103.615 114.040 103.980 ;
        RECT 114.230 103.615 114.505 104.465 ;
        RECT 114.675 103.615 114.865 104.975 ;
        RECT 115.035 104.990 115.205 105.655 ;
        RECT 115.375 105.235 115.545 105.995 ;
        RECT 115.780 105.235 116.295 105.645 ;
        RECT 115.035 104.800 115.785 104.990 ;
        RECT 115.955 104.425 116.295 105.235 ;
        RECT 116.505 104.855 116.735 105.995 ;
        RECT 116.905 104.845 117.235 105.825 ;
        RECT 117.405 104.855 117.615 105.995 ;
        RECT 117.845 104.905 121.355 105.995 ;
        RECT 116.485 104.435 116.815 104.685 ;
        RECT 115.065 104.255 116.295 104.425 ;
        RECT 115.045 103.445 115.555 103.980 ;
        RECT 115.775 103.650 116.020 104.255 ;
        RECT 116.505 103.445 116.735 104.265 ;
        RECT 116.985 104.245 117.235 104.845 ;
        RECT 116.905 103.615 117.235 104.245 ;
        RECT 117.405 103.445 117.615 104.265 ;
        RECT 117.845 104.215 119.495 104.735 ;
        RECT 119.665 104.385 121.355 104.905 ;
        RECT 121.525 104.830 121.815 105.995 ;
        RECT 122.445 104.905 123.655 105.995 ;
        RECT 122.445 104.365 122.965 104.905 ;
        RECT 117.845 103.445 121.355 104.215 ;
        RECT 123.135 104.195 123.655 104.735 ;
        RECT 121.525 103.445 121.815 104.170 ;
        RECT 122.445 103.445 123.655 104.195 ;
        RECT 5.520 103.275 123.740 103.445 ;
        RECT 5.605 102.525 6.815 103.275 ;
        RECT 7.075 102.725 7.245 103.105 ;
        RECT 7.425 102.895 7.755 103.275 ;
        RECT 7.075 102.555 7.740 102.725 ;
        RECT 7.935 102.600 8.195 103.105 ;
        RECT 5.605 101.985 6.125 102.525 ;
        RECT 6.295 101.815 6.815 102.355 ;
        RECT 7.005 102.005 7.335 102.375 ;
        RECT 7.570 102.300 7.740 102.555 ;
        RECT 7.570 101.970 7.855 102.300 ;
        RECT 7.570 101.825 7.740 101.970 ;
        RECT 5.605 100.725 6.815 101.815 ;
        RECT 7.075 101.655 7.740 101.825 ;
        RECT 8.025 101.800 8.195 102.600 ;
        RECT 8.455 102.725 8.625 103.015 ;
        RECT 8.795 102.895 9.125 103.275 ;
        RECT 8.455 102.555 9.120 102.725 ;
        RECT 7.075 100.895 7.245 101.655 ;
        RECT 7.425 100.725 7.755 101.485 ;
        RECT 7.925 100.895 8.195 101.800 ;
        RECT 8.370 101.735 8.720 102.385 ;
        RECT 8.890 101.565 9.120 102.555 ;
        RECT 8.455 101.395 9.120 101.565 ;
        RECT 8.455 100.895 8.625 101.395 ;
        RECT 8.795 100.725 9.125 101.225 ;
        RECT 9.295 100.895 9.520 103.015 ;
        RECT 9.735 102.895 10.065 103.275 ;
        RECT 10.235 102.725 10.405 103.055 ;
        RECT 10.705 102.895 11.720 103.095 ;
        RECT 9.710 102.535 10.405 102.725 ;
        RECT 9.710 101.565 9.880 102.535 ;
        RECT 10.050 101.735 10.460 102.355 ;
        RECT 10.630 101.785 10.850 102.655 ;
        RECT 11.030 102.345 11.380 102.715 ;
        RECT 11.550 102.165 11.720 102.895 ;
        RECT 11.890 102.835 12.300 103.275 ;
        RECT 12.590 102.635 12.840 103.065 ;
        RECT 13.040 102.815 13.360 103.275 ;
        RECT 13.920 102.885 14.770 103.055 ;
        RECT 11.890 102.295 12.300 102.625 ;
        RECT 12.590 102.295 13.010 102.635 ;
        RECT 11.300 102.125 11.720 102.165 ;
        RECT 11.300 101.955 12.650 102.125 ;
        RECT 9.710 101.395 10.405 101.565 ;
        RECT 10.630 101.405 11.130 101.785 ;
        RECT 9.735 100.725 10.065 101.225 ;
        RECT 10.235 100.895 10.405 101.395 ;
        RECT 11.300 101.110 11.470 101.955 ;
        RECT 12.400 101.795 12.650 101.955 ;
        RECT 11.640 101.525 11.890 101.785 ;
        RECT 12.820 101.525 13.010 102.295 ;
        RECT 11.640 101.275 13.010 101.525 ;
        RECT 13.180 102.465 14.430 102.635 ;
        RECT 13.180 101.705 13.350 102.465 ;
        RECT 14.100 102.345 14.430 102.465 ;
        RECT 13.520 101.885 13.700 102.295 ;
        RECT 14.600 102.125 14.770 102.885 ;
        RECT 14.970 102.795 15.630 103.275 ;
        RECT 15.810 102.680 16.130 103.010 ;
        RECT 14.960 102.355 15.620 102.625 ;
        RECT 14.960 102.295 15.290 102.355 ;
        RECT 15.440 102.125 15.770 102.185 ;
        RECT 13.870 101.955 15.770 102.125 ;
        RECT 13.180 101.395 13.700 101.705 ;
        RECT 13.870 101.445 14.040 101.955 ;
        RECT 15.940 101.785 16.130 102.680 ;
        RECT 14.210 101.615 16.130 101.785 ;
        RECT 15.810 101.595 16.130 101.615 ;
        RECT 16.330 102.365 16.580 103.015 ;
        RECT 16.760 102.815 17.045 103.275 ;
        RECT 17.225 102.565 17.480 103.095 ;
        RECT 16.330 102.035 17.130 102.365 ;
        RECT 13.870 101.275 15.080 101.445 ;
        RECT 10.640 100.940 11.470 101.110 ;
        RECT 11.710 100.725 12.090 101.105 ;
        RECT 12.270 100.985 12.440 101.275 ;
        RECT 13.870 101.195 14.040 101.275 ;
        RECT 12.610 100.725 12.940 101.105 ;
        RECT 13.410 100.945 14.040 101.195 ;
        RECT 14.220 100.725 14.640 101.105 ;
        RECT 14.840 100.985 15.080 101.275 ;
        RECT 15.310 100.725 15.640 101.415 ;
        RECT 15.810 100.985 15.980 101.595 ;
        RECT 16.330 101.445 16.580 102.035 ;
        RECT 17.300 101.705 17.480 102.565 ;
        RECT 17.225 101.575 17.480 101.705 ;
        RECT 18.030 102.535 18.285 103.105 ;
        RECT 18.455 102.875 18.785 103.275 ;
        RECT 19.210 102.740 19.740 103.105 ;
        RECT 19.210 102.705 19.385 102.740 ;
        RECT 18.455 102.535 19.385 102.705 ;
        RECT 18.030 101.865 18.200 102.535 ;
        RECT 18.455 102.365 18.625 102.535 ;
        RECT 18.370 102.035 18.625 102.365 ;
        RECT 18.850 102.035 19.045 102.365 ;
        RECT 16.250 100.935 16.580 101.445 ;
        RECT 16.760 100.725 17.045 101.525 ;
        RECT 17.225 101.405 17.565 101.575 ;
        RECT 17.225 101.035 17.480 101.405 ;
        RECT 18.030 100.895 18.365 101.865 ;
        RECT 18.535 100.725 18.705 101.865 ;
        RECT 18.875 101.065 19.045 102.035 ;
        RECT 19.215 101.405 19.385 102.535 ;
        RECT 19.555 101.745 19.725 102.545 ;
        RECT 19.930 102.255 20.205 103.105 ;
        RECT 19.925 102.085 20.205 102.255 ;
        RECT 19.930 101.945 20.205 102.085 ;
        RECT 20.375 101.745 20.565 103.105 ;
        RECT 20.745 102.740 21.255 103.275 ;
        RECT 21.475 102.465 21.720 103.070 ;
        RECT 20.765 102.295 21.995 102.465 ;
        RECT 22.225 102.455 22.435 103.275 ;
        RECT 22.605 102.475 22.935 103.105 ;
        RECT 19.555 101.575 20.565 101.745 ;
        RECT 20.735 101.730 21.485 101.920 ;
        RECT 19.215 101.235 20.340 101.405 ;
        RECT 20.735 101.065 20.905 101.730 ;
        RECT 21.655 101.485 21.995 102.295 ;
        RECT 22.605 101.875 22.855 102.475 ;
        RECT 23.105 102.455 23.335 103.275 ;
        RECT 23.545 102.505 26.135 103.275 ;
        RECT 26.965 102.645 27.295 103.005 ;
        RECT 27.915 102.815 28.165 103.275 ;
        RECT 28.335 102.815 28.895 103.105 ;
        RECT 23.025 102.035 23.355 102.285 ;
        RECT 23.545 101.985 24.755 102.505 ;
        RECT 26.965 102.455 28.355 102.645 ;
        RECT 28.185 102.365 28.355 102.455 ;
        RECT 18.875 100.895 20.905 101.065 ;
        RECT 21.075 100.725 21.245 101.485 ;
        RECT 21.480 101.075 21.995 101.485 ;
        RECT 22.225 100.725 22.435 101.865 ;
        RECT 22.605 100.895 22.935 101.875 ;
        RECT 23.105 100.725 23.335 101.865 ;
        RECT 24.925 101.815 26.135 102.335 ;
        RECT 23.545 100.725 26.135 101.815 ;
        RECT 26.780 102.035 27.455 102.285 ;
        RECT 27.675 102.035 28.015 102.285 ;
        RECT 28.185 102.035 28.475 102.365 ;
        RECT 26.780 101.675 27.045 102.035 ;
        RECT 28.185 101.785 28.355 102.035 ;
        RECT 27.415 101.615 28.355 101.785 ;
        RECT 26.965 100.725 27.245 101.395 ;
        RECT 27.415 101.065 27.715 101.615 ;
        RECT 28.645 101.445 28.895 102.815 ;
        RECT 29.065 102.505 30.735 103.275 ;
        RECT 31.365 102.550 31.655 103.275 ;
        RECT 31.830 102.535 32.085 103.105 ;
        RECT 32.255 102.875 32.585 103.275 ;
        RECT 33.010 102.740 33.540 103.105 ;
        RECT 33.010 102.705 33.185 102.740 ;
        RECT 32.255 102.535 33.185 102.705 ;
        RECT 33.730 102.595 34.005 103.105 ;
        RECT 29.065 101.985 29.815 102.505 ;
        RECT 29.985 101.815 30.735 102.335 ;
        RECT 27.915 100.725 28.245 101.445 ;
        RECT 28.435 100.895 28.895 101.445 ;
        RECT 29.065 100.725 30.735 101.815 ;
        RECT 31.365 100.725 31.655 101.890 ;
        RECT 31.830 101.865 32.000 102.535 ;
        RECT 32.255 102.365 32.425 102.535 ;
        RECT 32.170 102.035 32.425 102.365 ;
        RECT 32.650 102.035 32.845 102.365 ;
        RECT 31.830 100.895 32.165 101.865 ;
        RECT 32.335 100.725 32.505 101.865 ;
        RECT 32.675 101.065 32.845 102.035 ;
        RECT 33.015 101.405 33.185 102.535 ;
        RECT 33.355 101.745 33.525 102.545 ;
        RECT 33.725 102.425 34.005 102.595 ;
        RECT 33.730 101.945 34.005 102.425 ;
        RECT 34.175 101.745 34.365 103.105 ;
        RECT 34.545 102.740 35.055 103.275 ;
        RECT 35.275 102.465 35.520 103.070 ;
        RECT 35.965 102.730 41.310 103.275 ;
        RECT 34.565 102.295 35.795 102.465 ;
        RECT 33.355 101.575 34.365 101.745 ;
        RECT 34.535 101.730 35.285 101.920 ;
        RECT 33.015 101.235 34.140 101.405 ;
        RECT 34.535 101.065 34.705 101.730 ;
        RECT 35.455 101.485 35.795 102.295 ;
        RECT 37.550 101.900 37.890 102.730 ;
        RECT 41.485 102.505 44.075 103.275 ;
        RECT 44.710 102.535 44.965 103.105 ;
        RECT 45.135 102.875 45.465 103.275 ;
        RECT 45.890 102.740 46.420 103.105 ;
        RECT 45.890 102.705 46.065 102.740 ;
        RECT 45.135 102.535 46.065 102.705 ;
        RECT 32.675 100.895 34.705 101.065 ;
        RECT 34.875 100.725 35.045 101.485 ;
        RECT 35.280 101.075 35.795 101.485 ;
        RECT 39.370 101.160 39.720 102.410 ;
        RECT 41.485 101.985 42.695 102.505 ;
        RECT 42.865 101.815 44.075 102.335 ;
        RECT 35.965 100.725 41.310 101.160 ;
        RECT 41.485 100.725 44.075 101.815 ;
        RECT 44.710 101.865 44.880 102.535 ;
        RECT 45.135 102.365 45.305 102.535 ;
        RECT 45.050 102.035 45.305 102.365 ;
        RECT 45.530 102.035 45.725 102.365 ;
        RECT 44.710 100.895 45.045 101.865 ;
        RECT 45.215 100.725 45.385 101.865 ;
        RECT 45.555 101.065 45.725 102.035 ;
        RECT 45.895 101.405 46.065 102.535 ;
        RECT 46.235 101.745 46.405 102.545 ;
        RECT 46.610 102.255 46.885 103.105 ;
        RECT 46.605 102.085 46.885 102.255 ;
        RECT 46.610 101.945 46.885 102.085 ;
        RECT 47.055 101.745 47.245 103.105 ;
        RECT 47.425 102.740 47.935 103.275 ;
        RECT 48.155 102.465 48.400 103.070 ;
        RECT 48.845 102.505 50.515 103.275 ;
        RECT 50.885 102.645 51.215 103.005 ;
        RECT 51.835 102.815 52.085 103.275 ;
        RECT 52.255 102.815 52.815 103.105 ;
        RECT 47.445 102.295 48.675 102.465 ;
        RECT 46.235 101.575 47.245 101.745 ;
        RECT 47.415 101.730 48.165 101.920 ;
        RECT 45.895 101.235 47.020 101.405 ;
        RECT 47.415 101.065 47.585 101.730 ;
        RECT 48.335 101.485 48.675 102.295 ;
        RECT 48.845 101.985 49.595 102.505 ;
        RECT 50.885 102.455 52.275 102.645 ;
        RECT 52.105 102.365 52.275 102.455 ;
        RECT 49.765 101.815 50.515 102.335 ;
        RECT 45.555 100.895 47.585 101.065 ;
        RECT 47.755 100.725 47.925 101.485 ;
        RECT 48.160 101.075 48.675 101.485 ;
        RECT 48.845 100.725 50.515 101.815 ;
        RECT 50.700 102.035 51.375 102.285 ;
        RECT 51.595 102.035 51.935 102.285 ;
        RECT 52.105 102.035 52.395 102.365 ;
        RECT 50.700 101.675 50.965 102.035 ;
        RECT 52.105 101.785 52.275 102.035 ;
        RECT 51.335 101.615 52.275 101.785 ;
        RECT 50.885 100.725 51.165 101.395 ;
        RECT 51.335 101.065 51.635 101.615 ;
        RECT 52.565 101.445 52.815 102.815 ;
        RECT 53.185 102.645 53.515 103.005 ;
        RECT 54.135 102.815 54.385 103.275 ;
        RECT 54.555 102.815 55.115 103.105 ;
        RECT 53.185 102.455 54.575 102.645 ;
        RECT 54.405 102.365 54.575 102.455 ;
        RECT 53.000 102.035 53.675 102.285 ;
        RECT 53.895 102.035 54.235 102.285 ;
        RECT 54.405 102.035 54.695 102.365 ;
        RECT 53.000 101.675 53.265 102.035 ;
        RECT 54.405 101.785 54.575 102.035 ;
        RECT 51.835 100.725 52.165 101.445 ;
        RECT 52.355 100.895 52.815 101.445 ;
        RECT 53.635 101.615 54.575 101.785 ;
        RECT 53.185 100.725 53.465 101.395 ;
        RECT 53.635 101.065 53.935 101.615 ;
        RECT 54.865 101.445 55.115 102.815 ;
        RECT 55.285 102.505 56.955 103.275 ;
        RECT 57.125 102.550 57.415 103.275 ;
        RECT 57.585 102.815 58.145 103.105 ;
        RECT 58.315 102.815 58.565 103.275 ;
        RECT 55.285 101.985 56.035 102.505 ;
        RECT 56.205 101.815 56.955 102.335 ;
        RECT 54.135 100.725 54.465 101.445 ;
        RECT 54.655 100.895 55.115 101.445 ;
        RECT 55.285 100.725 56.955 101.815 ;
        RECT 57.125 100.725 57.415 101.890 ;
        RECT 57.585 101.445 57.835 102.815 ;
        RECT 59.185 102.645 59.515 103.005 ;
        RECT 59.885 102.730 65.230 103.275 ;
        RECT 58.125 102.455 59.515 102.645 ;
        RECT 58.125 102.365 58.295 102.455 ;
        RECT 58.005 102.035 58.295 102.365 ;
        RECT 58.465 102.035 58.805 102.285 ;
        RECT 59.025 102.035 59.700 102.285 ;
        RECT 58.125 101.785 58.295 102.035 ;
        RECT 58.125 101.615 59.065 101.785 ;
        RECT 59.435 101.675 59.700 102.035 ;
        RECT 61.470 101.900 61.810 102.730 ;
        RECT 66.525 102.645 66.855 103.005 ;
        RECT 67.475 102.815 67.725 103.275 ;
        RECT 67.895 102.815 68.455 103.105 ;
        RECT 66.525 102.455 67.915 102.645 ;
        RECT 57.585 100.895 58.045 101.445 ;
        RECT 58.235 100.725 58.565 101.445 ;
        RECT 58.765 101.065 59.065 101.615 ;
        RECT 59.235 100.725 59.515 101.395 ;
        RECT 63.290 101.160 63.640 102.410 ;
        RECT 67.745 102.365 67.915 102.455 ;
        RECT 66.340 102.035 67.015 102.285 ;
        RECT 67.235 102.035 67.575 102.285 ;
        RECT 67.745 102.035 68.035 102.365 ;
        RECT 66.340 101.675 66.605 102.035 ;
        RECT 67.745 101.785 67.915 102.035 ;
        RECT 66.975 101.615 67.915 101.785 ;
        RECT 59.885 100.725 65.230 101.160 ;
        RECT 66.525 100.725 66.805 101.395 ;
        RECT 66.975 101.065 67.275 101.615 ;
        RECT 68.205 101.445 68.455 102.815 ;
        RECT 67.475 100.725 67.805 101.445 ;
        RECT 67.995 100.895 68.455 101.445 ;
        RECT 68.625 102.775 68.885 103.105 ;
        RECT 69.095 102.795 69.370 103.275 ;
        RECT 68.625 101.865 68.795 102.775 ;
        RECT 69.580 102.705 69.785 103.105 ;
        RECT 69.955 102.875 70.290 103.275 ;
        RECT 70.465 102.730 75.810 103.275 ;
        RECT 75.985 102.730 81.330 103.275 ;
        RECT 68.965 102.035 69.325 102.615 ;
        RECT 69.580 102.535 70.265 102.705 ;
        RECT 69.505 101.865 69.755 102.365 ;
        RECT 68.625 101.695 69.755 101.865 ;
        RECT 68.625 100.925 68.895 101.695 ;
        RECT 69.925 101.505 70.265 102.535 ;
        RECT 72.050 101.900 72.390 102.730 ;
        RECT 69.065 100.725 69.395 101.505 ;
        RECT 69.600 101.330 70.265 101.505 ;
        RECT 69.600 100.925 69.785 101.330 ;
        RECT 73.870 101.160 74.220 102.410 ;
        RECT 77.570 101.900 77.910 102.730 ;
        RECT 81.505 102.525 82.715 103.275 ;
        RECT 82.885 102.550 83.175 103.275 ;
        RECT 84.465 102.645 84.795 103.005 ;
        RECT 85.415 102.815 85.665 103.275 ;
        RECT 85.835 102.815 86.395 103.105 ;
        RECT 79.390 101.160 79.740 102.410 ;
        RECT 81.505 101.985 82.025 102.525 ;
        RECT 84.465 102.455 85.855 102.645 ;
        RECT 85.685 102.365 85.855 102.455 ;
        RECT 82.195 101.815 82.715 102.355 ;
        RECT 84.280 102.035 84.955 102.285 ;
        RECT 85.175 102.035 85.515 102.285 ;
        RECT 85.685 102.035 85.975 102.365 ;
        RECT 69.955 100.725 70.290 101.150 ;
        RECT 70.465 100.725 75.810 101.160 ;
        RECT 75.985 100.725 81.330 101.160 ;
        RECT 81.505 100.725 82.715 101.815 ;
        RECT 82.885 100.725 83.175 101.890 ;
        RECT 84.280 101.675 84.545 102.035 ;
        RECT 85.685 101.785 85.855 102.035 ;
        RECT 84.915 101.615 85.855 101.785 ;
        RECT 84.465 100.725 84.745 101.395 ;
        RECT 84.915 101.065 85.215 101.615 ;
        RECT 86.145 101.445 86.395 102.815 ;
        RECT 85.415 100.725 85.745 101.445 ;
        RECT 85.935 100.895 86.395 101.445 ;
        RECT 86.570 102.535 86.825 103.105 ;
        RECT 86.995 102.875 87.325 103.275 ;
        RECT 87.750 102.740 88.280 103.105 ;
        RECT 87.750 102.705 87.925 102.740 ;
        RECT 86.995 102.535 87.925 102.705 ;
        RECT 88.470 102.595 88.745 103.105 ;
        RECT 86.570 101.865 86.740 102.535 ;
        RECT 86.995 102.365 87.165 102.535 ;
        RECT 86.910 102.035 87.165 102.365 ;
        RECT 87.390 102.035 87.585 102.365 ;
        RECT 86.570 100.895 86.905 101.865 ;
        RECT 87.075 100.725 87.245 101.865 ;
        RECT 87.415 101.065 87.585 102.035 ;
        RECT 87.755 101.405 87.925 102.535 ;
        RECT 88.095 101.745 88.265 102.545 ;
        RECT 88.465 102.425 88.745 102.595 ;
        RECT 88.470 101.945 88.745 102.425 ;
        RECT 88.915 101.745 89.105 103.105 ;
        RECT 89.285 102.740 89.795 103.275 ;
        RECT 90.015 102.465 90.260 103.070 ;
        RECT 91.625 102.815 92.185 103.105 ;
        RECT 92.355 102.815 92.605 103.275 ;
        RECT 89.305 102.295 90.535 102.465 ;
        RECT 88.095 101.575 89.105 101.745 ;
        RECT 89.275 101.730 90.025 101.920 ;
        RECT 87.755 101.235 88.880 101.405 ;
        RECT 89.275 101.065 89.445 101.730 ;
        RECT 90.195 101.485 90.535 102.295 ;
        RECT 87.415 100.895 89.445 101.065 ;
        RECT 89.615 100.725 89.785 101.485 ;
        RECT 90.020 101.075 90.535 101.485 ;
        RECT 91.625 101.445 91.875 102.815 ;
        RECT 93.225 102.645 93.555 103.005 ;
        RECT 92.165 102.455 93.555 102.645 ;
        RECT 94.385 102.815 94.945 103.105 ;
        RECT 95.115 102.815 95.365 103.275 ;
        RECT 92.165 102.365 92.335 102.455 ;
        RECT 92.045 102.035 92.335 102.365 ;
        RECT 92.505 102.035 92.845 102.285 ;
        RECT 93.065 102.035 93.740 102.285 ;
        RECT 92.165 101.785 92.335 102.035 ;
        RECT 92.165 101.615 93.105 101.785 ;
        RECT 93.475 101.675 93.740 102.035 ;
        RECT 91.625 100.895 92.085 101.445 ;
        RECT 92.275 100.725 92.605 101.445 ;
        RECT 92.805 101.065 93.105 101.615 ;
        RECT 94.385 101.445 94.635 102.815 ;
        RECT 95.985 102.645 96.315 103.005 ;
        RECT 94.925 102.455 96.315 102.645 ;
        RECT 97.235 102.725 97.405 103.015 ;
        RECT 97.575 102.895 97.905 103.275 ;
        RECT 97.235 102.555 97.900 102.725 ;
        RECT 94.925 102.365 95.095 102.455 ;
        RECT 94.805 102.035 95.095 102.365 ;
        RECT 95.265 102.035 95.605 102.285 ;
        RECT 95.825 102.035 96.500 102.285 ;
        RECT 94.925 101.785 95.095 102.035 ;
        RECT 94.925 101.615 95.865 101.785 ;
        RECT 96.235 101.675 96.500 102.035 ;
        RECT 97.150 101.735 97.500 102.385 ;
        RECT 93.275 100.725 93.555 101.395 ;
        RECT 94.385 100.895 94.845 101.445 ;
        RECT 95.035 100.725 95.365 101.445 ;
        RECT 95.565 101.065 95.865 101.615 ;
        RECT 97.670 101.565 97.900 102.555 ;
        RECT 97.235 101.395 97.900 101.565 ;
        RECT 96.035 100.725 96.315 101.395 ;
        RECT 97.235 100.895 97.405 101.395 ;
        RECT 97.575 100.725 97.905 101.225 ;
        RECT 98.075 100.895 98.300 103.015 ;
        RECT 98.515 102.895 98.845 103.275 ;
        RECT 99.015 102.725 99.185 103.055 ;
        RECT 99.485 102.895 100.500 103.095 ;
        RECT 98.490 102.535 99.185 102.725 ;
        RECT 98.490 101.565 98.660 102.535 ;
        RECT 98.830 101.735 99.240 102.355 ;
        RECT 99.410 101.785 99.630 102.655 ;
        RECT 99.810 102.345 100.160 102.715 ;
        RECT 100.330 102.165 100.500 102.895 ;
        RECT 100.670 102.835 101.080 103.275 ;
        RECT 101.370 102.635 101.620 103.065 ;
        RECT 101.820 102.815 102.140 103.275 ;
        RECT 102.700 102.885 103.550 103.055 ;
        RECT 100.670 102.295 101.080 102.625 ;
        RECT 101.370 102.295 101.790 102.635 ;
        RECT 100.080 102.125 100.500 102.165 ;
        RECT 100.080 101.955 101.430 102.125 ;
        RECT 98.490 101.395 99.185 101.565 ;
        RECT 99.410 101.405 99.910 101.785 ;
        RECT 98.515 100.725 98.845 101.225 ;
        RECT 99.015 100.895 99.185 101.395 ;
        RECT 100.080 101.110 100.250 101.955 ;
        RECT 101.180 101.795 101.430 101.955 ;
        RECT 100.420 101.525 100.670 101.785 ;
        RECT 101.600 101.525 101.790 102.295 ;
        RECT 100.420 101.275 101.790 101.525 ;
        RECT 101.960 102.465 103.210 102.635 ;
        RECT 101.960 101.705 102.130 102.465 ;
        RECT 102.880 102.345 103.210 102.465 ;
        RECT 102.300 101.885 102.480 102.295 ;
        RECT 103.380 102.125 103.550 102.885 ;
        RECT 103.750 102.795 104.410 103.275 ;
        RECT 104.590 102.680 104.910 103.010 ;
        RECT 103.740 102.355 104.400 102.625 ;
        RECT 103.740 102.295 104.070 102.355 ;
        RECT 104.220 102.125 104.550 102.185 ;
        RECT 102.650 101.955 104.550 102.125 ;
        RECT 101.960 101.395 102.480 101.705 ;
        RECT 102.650 101.445 102.820 101.955 ;
        RECT 104.720 101.785 104.910 102.680 ;
        RECT 102.990 101.615 104.910 101.785 ;
        RECT 104.590 101.595 104.910 101.615 ;
        RECT 105.110 102.365 105.360 103.015 ;
        RECT 105.540 102.815 105.825 103.275 ;
        RECT 106.005 102.565 106.260 103.095 ;
        RECT 105.110 102.035 105.910 102.365 ;
        RECT 102.650 101.275 103.860 101.445 ;
        RECT 99.420 100.940 100.250 101.110 ;
        RECT 100.490 100.725 100.870 101.105 ;
        RECT 101.050 100.985 101.220 101.275 ;
        RECT 102.650 101.195 102.820 101.275 ;
        RECT 101.390 100.725 101.720 101.105 ;
        RECT 102.190 100.945 102.820 101.195 ;
        RECT 103.000 100.725 103.420 101.105 ;
        RECT 103.620 100.985 103.860 101.275 ;
        RECT 104.090 100.725 104.420 101.415 ;
        RECT 104.590 100.985 104.760 101.595 ;
        RECT 105.110 101.445 105.360 102.035 ;
        RECT 106.080 101.705 106.260 102.565 ;
        RECT 106.805 102.505 108.475 103.275 ;
        RECT 108.645 102.550 108.935 103.275 ;
        RECT 109.570 102.535 109.825 103.105 ;
        RECT 109.995 102.875 110.325 103.275 ;
        RECT 110.750 102.740 111.280 103.105 ;
        RECT 111.470 102.935 111.745 103.105 ;
        RECT 111.465 102.765 111.745 102.935 ;
        RECT 110.750 102.705 110.925 102.740 ;
        RECT 109.995 102.535 110.925 102.705 ;
        RECT 106.805 101.985 107.555 102.505 ;
        RECT 107.725 101.815 108.475 102.335 ;
        RECT 105.030 100.935 105.360 101.445 ;
        RECT 105.540 100.725 105.825 101.525 ;
        RECT 106.005 101.235 106.260 101.705 ;
        RECT 106.005 101.065 106.345 101.235 ;
        RECT 106.005 101.035 106.260 101.065 ;
        RECT 106.805 100.725 108.475 101.815 ;
        RECT 108.645 100.725 108.935 101.890 ;
        RECT 109.570 101.865 109.740 102.535 ;
        RECT 109.995 102.365 110.165 102.535 ;
        RECT 109.910 102.035 110.165 102.365 ;
        RECT 110.390 102.035 110.585 102.365 ;
        RECT 109.570 100.895 109.905 101.865 ;
        RECT 110.075 100.725 110.245 101.865 ;
        RECT 110.415 101.065 110.585 102.035 ;
        RECT 110.755 101.405 110.925 102.535 ;
        RECT 111.095 101.745 111.265 102.545 ;
        RECT 111.470 101.945 111.745 102.765 ;
        RECT 111.915 101.745 112.105 103.105 ;
        RECT 112.285 102.740 112.795 103.275 ;
        RECT 113.015 102.465 113.260 103.070 ;
        RECT 112.305 102.295 113.535 102.465 ;
        RECT 113.765 102.455 113.975 103.275 ;
        RECT 114.145 102.475 114.475 103.105 ;
        RECT 111.095 101.575 112.105 101.745 ;
        RECT 112.275 101.730 113.025 101.920 ;
        RECT 110.755 101.235 111.880 101.405 ;
        RECT 112.275 101.065 112.445 101.730 ;
        RECT 113.195 101.485 113.535 102.295 ;
        RECT 114.145 101.875 114.395 102.475 ;
        RECT 114.645 102.455 114.875 103.275 ;
        RECT 115.085 102.730 120.430 103.275 ;
        RECT 114.565 102.035 114.895 102.285 ;
        RECT 116.670 101.900 117.010 102.730 ;
        RECT 120.605 102.505 122.275 103.275 ;
        RECT 122.445 102.525 123.655 103.275 ;
        RECT 110.415 100.895 112.445 101.065 ;
        RECT 112.615 100.725 112.785 101.485 ;
        RECT 113.020 101.075 113.535 101.485 ;
        RECT 113.765 100.725 113.975 101.865 ;
        RECT 114.145 100.895 114.475 101.875 ;
        RECT 114.645 100.725 114.875 101.865 ;
        RECT 118.490 101.160 118.840 102.410 ;
        RECT 120.605 101.985 121.355 102.505 ;
        RECT 121.525 101.815 122.275 102.335 ;
        RECT 115.085 100.725 120.430 101.160 ;
        RECT 120.605 100.725 122.275 101.815 ;
        RECT 122.445 101.815 122.965 102.355 ;
        RECT 123.135 101.985 123.655 102.525 ;
        RECT 122.445 100.725 123.655 101.815 ;
        RECT 5.520 100.555 123.740 100.725 ;
        RECT 5.605 99.465 6.815 100.555 ;
        RECT 7.995 99.885 8.165 100.385 ;
        RECT 8.335 100.055 8.665 100.555 ;
        RECT 7.995 99.715 8.660 99.885 ;
        RECT 5.605 98.755 6.125 99.295 ;
        RECT 6.295 98.925 6.815 99.465 ;
        RECT 7.910 98.895 8.260 99.545 ;
        RECT 5.605 98.005 6.815 98.755 ;
        RECT 8.430 98.725 8.660 99.715 ;
        RECT 7.995 98.555 8.660 98.725 ;
        RECT 7.995 98.265 8.165 98.555 ;
        RECT 8.335 98.005 8.665 98.385 ;
        RECT 8.835 98.265 9.060 100.385 ;
        RECT 9.275 100.055 9.605 100.555 ;
        RECT 9.775 99.885 9.945 100.385 ;
        RECT 10.180 100.170 11.010 100.340 ;
        RECT 11.250 100.175 11.630 100.555 ;
        RECT 9.250 99.715 9.945 99.885 ;
        RECT 9.250 98.745 9.420 99.715 ;
        RECT 9.590 98.925 10.000 99.545 ;
        RECT 10.170 99.495 10.670 99.875 ;
        RECT 9.250 98.555 9.945 98.745 ;
        RECT 10.170 98.625 10.390 99.495 ;
        RECT 10.840 99.325 11.010 100.170 ;
        RECT 11.810 100.005 11.980 100.295 ;
        RECT 12.150 100.175 12.480 100.555 ;
        RECT 12.950 100.085 13.580 100.335 ;
        RECT 13.760 100.175 14.180 100.555 ;
        RECT 13.410 100.005 13.580 100.085 ;
        RECT 14.380 100.005 14.620 100.295 ;
        RECT 11.180 99.755 12.550 100.005 ;
        RECT 11.180 99.495 11.430 99.755 ;
        RECT 11.940 99.325 12.190 99.485 ;
        RECT 10.840 99.155 12.190 99.325 ;
        RECT 10.840 99.115 11.260 99.155 ;
        RECT 10.570 98.565 10.920 98.935 ;
        RECT 9.275 98.005 9.605 98.385 ;
        RECT 9.775 98.225 9.945 98.555 ;
        RECT 11.090 98.385 11.260 99.115 ;
        RECT 12.360 98.985 12.550 99.755 ;
        RECT 11.430 98.655 11.840 98.985 ;
        RECT 12.130 98.645 12.550 98.985 ;
        RECT 12.720 99.575 13.240 99.885 ;
        RECT 13.410 99.835 14.620 100.005 ;
        RECT 14.850 99.865 15.180 100.555 ;
        RECT 12.720 98.815 12.890 99.575 ;
        RECT 13.060 98.985 13.240 99.395 ;
        RECT 13.410 99.325 13.580 99.835 ;
        RECT 15.350 99.685 15.520 100.295 ;
        RECT 15.790 99.835 16.120 100.345 ;
        RECT 15.350 99.665 15.670 99.685 ;
        RECT 13.750 99.495 15.670 99.665 ;
        RECT 13.410 99.155 15.310 99.325 ;
        RECT 13.640 98.815 13.970 98.935 ;
        RECT 12.720 98.645 13.970 98.815 ;
        RECT 10.245 98.185 11.260 98.385 ;
        RECT 11.430 98.005 11.840 98.445 ;
        RECT 12.130 98.215 12.380 98.645 ;
        RECT 12.580 98.005 12.900 98.465 ;
        RECT 14.140 98.395 14.310 99.155 ;
        RECT 14.980 99.095 15.310 99.155 ;
        RECT 14.500 98.925 14.830 98.985 ;
        RECT 14.500 98.655 15.160 98.925 ;
        RECT 15.480 98.600 15.670 99.495 ;
        RECT 13.460 98.225 14.310 98.395 ;
        RECT 14.510 98.005 15.170 98.485 ;
        RECT 15.350 98.270 15.670 98.600 ;
        RECT 15.870 99.245 16.120 99.835 ;
        RECT 16.300 99.755 16.585 100.555 ;
        RECT 16.765 100.215 17.020 100.245 ;
        RECT 16.765 100.045 17.105 100.215 ;
        RECT 16.765 99.575 17.020 100.045 ;
        RECT 15.870 98.915 16.670 99.245 ;
        RECT 15.870 98.265 16.120 98.915 ;
        RECT 16.840 98.715 17.020 99.575 ;
        RECT 18.485 99.390 18.775 100.555 ;
        RECT 18.945 99.465 22.455 100.555 ;
        RECT 22.825 99.885 23.105 100.555 ;
        RECT 23.275 99.665 23.575 100.215 ;
        RECT 23.775 99.835 24.105 100.555 ;
        RECT 24.295 99.835 24.755 100.385 ;
        RECT 18.945 98.775 20.595 99.295 ;
        RECT 20.765 98.945 22.455 99.465 ;
        RECT 22.640 99.245 22.905 99.605 ;
        RECT 23.275 99.495 24.215 99.665 ;
        RECT 24.045 99.245 24.215 99.495 ;
        RECT 22.640 98.995 23.315 99.245 ;
        RECT 23.535 98.995 23.875 99.245 ;
        RECT 24.045 98.915 24.335 99.245 ;
        RECT 24.045 98.825 24.215 98.915 ;
        RECT 16.300 98.005 16.585 98.465 ;
        RECT 16.765 98.185 17.020 98.715 ;
        RECT 18.485 98.005 18.775 98.730 ;
        RECT 18.945 98.005 22.455 98.775 ;
        RECT 22.825 98.635 24.215 98.825 ;
        RECT 22.825 98.275 23.155 98.635 ;
        RECT 24.505 98.465 24.755 99.835 ;
        RECT 23.775 98.005 24.025 98.465 ;
        RECT 24.195 98.175 24.755 98.465 ;
        RECT 24.925 99.835 25.385 100.385 ;
        RECT 25.575 99.835 25.905 100.555 ;
        RECT 24.925 98.465 25.175 99.835 ;
        RECT 26.105 99.665 26.405 100.215 ;
        RECT 26.575 99.885 26.855 100.555 ;
        RECT 27.425 99.885 27.705 100.555 ;
        RECT 25.465 99.495 26.405 99.665 ;
        RECT 27.875 99.665 28.175 100.215 ;
        RECT 28.375 99.835 28.705 100.555 ;
        RECT 28.895 99.835 29.355 100.385 ;
        RECT 25.465 99.245 25.635 99.495 ;
        RECT 26.775 99.245 27.040 99.605 ;
        RECT 25.345 98.915 25.635 99.245 ;
        RECT 25.805 98.995 26.145 99.245 ;
        RECT 26.365 98.995 27.040 99.245 ;
        RECT 27.240 99.245 27.505 99.605 ;
        RECT 27.875 99.495 28.815 99.665 ;
        RECT 28.645 99.245 28.815 99.495 ;
        RECT 27.240 98.995 27.915 99.245 ;
        RECT 28.135 98.995 28.475 99.245 ;
        RECT 25.465 98.825 25.635 98.915 ;
        RECT 28.645 98.915 28.935 99.245 ;
        RECT 28.645 98.825 28.815 98.915 ;
        RECT 25.465 98.635 26.855 98.825 ;
        RECT 24.925 98.175 25.485 98.465 ;
        RECT 25.655 98.005 25.905 98.465 ;
        RECT 26.525 98.275 26.855 98.635 ;
        RECT 27.425 98.635 28.815 98.825 ;
        RECT 27.425 98.275 27.755 98.635 ;
        RECT 29.105 98.465 29.355 99.835 ;
        RECT 29.525 99.465 33.035 100.555 ;
        RECT 33.205 99.465 34.415 100.555 ;
        RECT 28.375 98.005 28.625 98.465 ;
        RECT 28.795 98.175 29.355 98.465 ;
        RECT 29.525 98.775 31.175 99.295 ;
        RECT 31.345 98.945 33.035 99.465 ;
        RECT 29.525 98.005 33.035 98.775 ;
        RECT 33.205 98.755 33.725 99.295 ;
        RECT 33.895 98.925 34.415 99.465 ;
        RECT 34.585 99.835 35.045 100.385 ;
        RECT 35.235 99.835 35.565 100.555 ;
        RECT 33.205 98.005 34.415 98.755 ;
        RECT 34.585 98.465 34.835 99.835 ;
        RECT 35.765 99.665 36.065 100.215 ;
        RECT 36.235 99.885 36.515 100.555 ;
        RECT 36.885 100.120 42.230 100.555 ;
        RECT 35.125 99.495 36.065 99.665 ;
        RECT 35.125 99.245 35.295 99.495 ;
        RECT 36.435 99.245 36.700 99.605 ;
        RECT 35.005 98.915 35.295 99.245 ;
        RECT 35.465 98.995 35.805 99.245 ;
        RECT 36.025 98.995 36.700 99.245 ;
        RECT 35.125 98.825 35.295 98.915 ;
        RECT 35.125 98.635 36.515 98.825 ;
        RECT 34.585 98.175 35.145 98.465 ;
        RECT 35.315 98.005 35.565 98.465 ;
        RECT 36.185 98.275 36.515 98.635 ;
        RECT 38.470 98.550 38.810 99.380 ;
        RECT 40.290 98.870 40.640 100.120 ;
        RECT 42.405 99.465 44.075 100.555 ;
        RECT 42.405 98.775 43.155 99.295 ;
        RECT 43.325 98.945 44.075 99.465 ;
        RECT 44.245 99.390 44.535 100.555 ;
        RECT 44.745 99.415 44.975 100.555 ;
        RECT 45.145 99.405 45.475 100.385 ;
        RECT 45.645 99.415 45.855 100.555 ;
        RECT 46.085 100.120 51.430 100.555 ;
        RECT 51.605 100.120 56.950 100.555 ;
        RECT 57.125 100.120 62.470 100.555 ;
        RECT 44.725 98.995 45.055 99.245 ;
        RECT 36.885 98.005 42.230 98.550 ;
        RECT 42.405 98.005 44.075 98.775 ;
        RECT 44.245 98.005 44.535 98.730 ;
        RECT 44.745 98.005 44.975 98.825 ;
        RECT 45.225 98.805 45.475 99.405 ;
        RECT 45.145 98.175 45.475 98.805 ;
        RECT 45.645 98.005 45.855 98.825 ;
        RECT 47.670 98.550 48.010 99.380 ;
        RECT 49.490 98.870 49.840 100.120 ;
        RECT 53.190 98.550 53.530 99.380 ;
        RECT 55.010 98.870 55.360 100.120 ;
        RECT 58.710 98.550 59.050 99.380 ;
        RECT 60.530 98.870 60.880 100.120 ;
        RECT 62.645 99.465 66.155 100.555 ;
        RECT 62.645 98.775 64.295 99.295 ;
        RECT 64.465 98.945 66.155 99.465 ;
        RECT 66.785 99.585 67.055 100.355 ;
        RECT 67.225 99.775 67.555 100.555 ;
        RECT 67.760 99.950 67.945 100.355 ;
        RECT 68.115 100.130 68.450 100.555 ;
        RECT 67.760 99.775 68.425 99.950 ;
        RECT 66.785 99.415 67.915 99.585 ;
        RECT 46.085 98.005 51.430 98.550 ;
        RECT 51.605 98.005 56.950 98.550 ;
        RECT 57.125 98.005 62.470 98.550 ;
        RECT 62.645 98.005 66.155 98.775 ;
        RECT 66.785 98.505 66.955 99.415 ;
        RECT 67.125 98.665 67.485 99.245 ;
        RECT 67.665 98.915 67.915 99.415 ;
        RECT 68.085 98.745 68.425 99.775 ;
        RECT 68.625 99.465 69.835 100.555 ;
        RECT 67.740 98.575 68.425 98.745 ;
        RECT 68.625 98.755 69.145 99.295 ;
        RECT 69.315 98.925 69.835 99.465 ;
        RECT 70.005 99.390 70.295 100.555 ;
        RECT 70.525 99.415 70.735 100.555 ;
        RECT 70.905 99.405 71.235 100.385 ;
        RECT 71.405 99.415 71.635 100.555 ;
        RECT 71.845 99.465 73.515 100.555 ;
        RECT 66.785 98.175 67.045 98.505 ;
        RECT 67.255 98.005 67.530 98.485 ;
        RECT 67.740 98.175 67.945 98.575 ;
        RECT 68.115 98.005 68.450 98.405 ;
        RECT 68.625 98.005 69.835 98.755 ;
        RECT 70.005 98.005 70.295 98.730 ;
        RECT 70.525 98.005 70.735 98.825 ;
        RECT 70.905 98.805 71.155 99.405 ;
        RECT 71.325 98.995 71.655 99.245 ;
        RECT 70.905 98.175 71.235 98.805 ;
        RECT 71.405 98.005 71.635 98.825 ;
        RECT 71.845 98.775 72.595 99.295 ;
        RECT 72.765 98.945 73.515 99.465 ;
        RECT 73.685 99.480 73.955 100.385 ;
        RECT 74.125 99.795 74.455 100.555 ;
        RECT 74.635 99.625 74.805 100.385 ;
        RECT 75.065 100.120 80.410 100.555 ;
        RECT 80.585 100.120 85.930 100.555 ;
        RECT 86.105 100.120 91.450 100.555 ;
        RECT 71.845 98.005 73.515 98.775 ;
        RECT 73.685 98.680 73.855 99.480 ;
        RECT 74.140 99.455 74.805 99.625 ;
        RECT 74.140 99.310 74.310 99.455 ;
        RECT 74.025 98.980 74.310 99.310 ;
        RECT 74.140 98.725 74.310 98.980 ;
        RECT 74.545 98.905 74.875 99.275 ;
        RECT 73.685 98.175 73.945 98.680 ;
        RECT 74.140 98.555 74.805 98.725 ;
        RECT 74.125 98.005 74.455 98.385 ;
        RECT 74.635 98.175 74.805 98.555 ;
        RECT 76.650 98.550 76.990 99.380 ;
        RECT 78.470 98.870 78.820 100.120 ;
        RECT 82.170 98.550 82.510 99.380 ;
        RECT 83.990 98.870 84.340 100.120 ;
        RECT 87.690 98.550 88.030 99.380 ;
        RECT 89.510 98.870 89.860 100.120 ;
        RECT 91.625 99.465 95.135 100.555 ;
        RECT 91.625 98.775 93.275 99.295 ;
        RECT 93.445 98.945 95.135 99.465 ;
        RECT 95.765 99.390 96.055 100.555 ;
        RECT 96.225 99.835 96.685 100.385 ;
        RECT 96.875 99.835 97.205 100.555 ;
        RECT 75.065 98.005 80.410 98.550 ;
        RECT 80.585 98.005 85.930 98.550 ;
        RECT 86.105 98.005 91.450 98.550 ;
        RECT 91.625 98.005 95.135 98.775 ;
        RECT 95.765 98.005 96.055 98.730 ;
        RECT 96.225 98.465 96.475 99.835 ;
        RECT 97.405 99.665 97.705 100.215 ;
        RECT 97.875 99.885 98.155 100.555 ;
        RECT 96.765 99.495 97.705 99.665 ;
        RECT 96.765 99.245 96.935 99.495 ;
        RECT 98.075 99.245 98.340 99.605 ;
        RECT 96.645 98.915 96.935 99.245 ;
        RECT 97.105 98.995 97.445 99.245 ;
        RECT 97.665 98.995 98.340 99.245 ;
        RECT 98.985 99.480 99.255 100.385 ;
        RECT 99.425 99.795 99.755 100.555 ;
        RECT 99.935 99.625 100.105 100.385 ;
        RECT 96.765 98.825 96.935 98.915 ;
        RECT 96.765 98.635 98.155 98.825 ;
        RECT 96.225 98.175 96.785 98.465 ;
        RECT 96.955 98.005 97.205 98.465 ;
        RECT 97.825 98.275 98.155 98.635 ;
        RECT 98.985 98.680 99.155 99.480 ;
        RECT 99.440 99.455 100.105 99.625 ;
        RECT 99.440 99.310 99.610 99.455 ;
        RECT 99.325 98.980 99.610 99.310 ;
        RECT 100.370 99.415 100.705 100.385 ;
        RECT 100.875 99.415 101.045 100.555 ;
        RECT 101.215 100.215 103.245 100.385 ;
        RECT 99.440 98.725 99.610 98.980 ;
        RECT 99.845 98.905 100.175 99.275 ;
        RECT 100.370 98.745 100.540 99.415 ;
        RECT 101.215 99.245 101.385 100.215 ;
        RECT 100.710 98.915 100.965 99.245 ;
        RECT 101.190 98.915 101.385 99.245 ;
        RECT 101.555 99.875 102.680 100.045 ;
        RECT 100.795 98.745 100.965 98.915 ;
        RECT 101.555 98.745 101.725 99.875 ;
        RECT 98.985 98.175 99.245 98.680 ;
        RECT 99.440 98.555 100.105 98.725 ;
        RECT 99.425 98.005 99.755 98.385 ;
        RECT 99.935 98.175 100.105 98.555 ;
        RECT 100.370 98.175 100.625 98.745 ;
        RECT 100.795 98.575 101.725 98.745 ;
        RECT 101.895 99.535 102.905 99.705 ;
        RECT 101.895 98.735 102.065 99.535 ;
        RECT 101.550 98.540 101.725 98.575 ;
        RECT 100.795 98.005 101.125 98.405 ;
        RECT 101.550 98.175 102.080 98.540 ;
        RECT 102.270 98.515 102.545 99.335 ;
        RECT 102.265 98.345 102.545 98.515 ;
        RECT 102.270 98.175 102.545 98.345 ;
        RECT 102.715 98.175 102.905 99.535 ;
        RECT 103.075 99.550 103.245 100.215 ;
        RECT 103.415 99.795 103.585 100.555 ;
        RECT 103.820 99.795 104.335 100.205 ;
        RECT 103.075 99.360 103.825 99.550 ;
        RECT 103.995 98.985 104.335 99.795 ;
        RECT 104.505 99.465 107.095 100.555 ;
        RECT 107.815 99.885 107.985 100.385 ;
        RECT 108.155 100.055 108.485 100.555 ;
        RECT 107.815 99.715 108.480 99.885 ;
        RECT 103.105 98.815 104.335 98.985 ;
        RECT 103.085 98.005 103.595 98.540 ;
        RECT 103.815 98.210 104.060 98.815 ;
        RECT 104.505 98.775 105.715 99.295 ;
        RECT 105.885 98.945 107.095 99.465 ;
        RECT 107.730 98.895 108.080 99.545 ;
        RECT 104.505 98.005 107.095 98.775 ;
        RECT 108.250 98.725 108.480 99.715 ;
        RECT 107.815 98.555 108.480 98.725 ;
        RECT 107.815 98.265 107.985 98.555 ;
        RECT 108.155 98.005 108.485 98.385 ;
        RECT 108.655 98.265 108.880 100.385 ;
        RECT 109.095 100.055 109.425 100.555 ;
        RECT 109.595 99.885 109.765 100.385 ;
        RECT 110.000 100.170 110.830 100.340 ;
        RECT 111.070 100.175 111.450 100.555 ;
        RECT 109.070 99.715 109.765 99.885 ;
        RECT 109.070 98.745 109.240 99.715 ;
        RECT 109.410 98.925 109.820 99.545 ;
        RECT 109.990 99.495 110.490 99.875 ;
        RECT 109.070 98.555 109.765 98.745 ;
        RECT 109.990 98.625 110.210 99.495 ;
        RECT 110.660 99.325 110.830 100.170 ;
        RECT 111.630 100.005 111.800 100.295 ;
        RECT 111.970 100.175 112.300 100.555 ;
        RECT 112.770 100.085 113.400 100.335 ;
        RECT 113.580 100.175 114.000 100.555 ;
        RECT 113.230 100.005 113.400 100.085 ;
        RECT 114.200 100.005 114.440 100.295 ;
        RECT 111.000 99.755 112.370 100.005 ;
        RECT 111.000 99.495 111.250 99.755 ;
        RECT 111.760 99.325 112.010 99.485 ;
        RECT 110.660 99.155 112.010 99.325 ;
        RECT 110.660 99.115 111.080 99.155 ;
        RECT 110.390 98.565 110.740 98.935 ;
        RECT 109.095 98.005 109.425 98.385 ;
        RECT 109.595 98.225 109.765 98.555 ;
        RECT 110.910 98.385 111.080 99.115 ;
        RECT 112.180 98.985 112.370 99.755 ;
        RECT 111.250 98.655 111.660 98.985 ;
        RECT 111.950 98.645 112.370 98.985 ;
        RECT 112.540 99.575 113.060 99.885 ;
        RECT 113.230 99.835 114.440 100.005 ;
        RECT 114.670 99.865 115.000 100.555 ;
        RECT 112.540 98.815 112.710 99.575 ;
        RECT 112.880 98.985 113.060 99.395 ;
        RECT 113.230 99.325 113.400 99.835 ;
        RECT 115.170 99.685 115.340 100.295 ;
        RECT 115.610 99.835 115.940 100.345 ;
        RECT 115.170 99.665 115.490 99.685 ;
        RECT 113.570 99.495 115.490 99.665 ;
        RECT 113.230 99.155 115.130 99.325 ;
        RECT 113.460 98.815 113.790 98.935 ;
        RECT 112.540 98.645 113.790 98.815 ;
        RECT 110.065 98.185 111.080 98.385 ;
        RECT 111.250 98.005 111.660 98.445 ;
        RECT 111.950 98.215 112.200 98.645 ;
        RECT 112.400 98.005 112.720 98.465 ;
        RECT 113.960 98.395 114.130 99.155 ;
        RECT 114.800 99.095 115.130 99.155 ;
        RECT 114.320 98.925 114.650 98.985 ;
        RECT 114.320 98.655 114.980 98.925 ;
        RECT 115.300 98.600 115.490 99.495 ;
        RECT 113.280 98.225 114.130 98.395 ;
        RECT 114.330 98.005 114.990 98.485 ;
        RECT 115.170 98.270 115.490 98.600 ;
        RECT 115.690 99.245 115.940 99.835 ;
        RECT 116.120 99.755 116.405 100.555 ;
        RECT 116.585 99.575 116.840 100.245 ;
        RECT 115.690 98.915 116.490 99.245 ;
        RECT 115.690 98.265 115.940 98.915 ;
        RECT 116.660 98.715 116.840 99.575 ;
        RECT 117.425 99.415 117.655 100.555 ;
        RECT 117.825 99.405 118.155 100.385 ;
        RECT 118.325 99.415 118.535 100.555 ;
        RECT 118.765 99.465 121.355 100.555 ;
        RECT 117.405 98.995 117.735 99.245 ;
        RECT 116.585 98.515 116.840 98.715 ;
        RECT 116.120 98.005 116.405 98.465 ;
        RECT 116.585 98.345 116.925 98.515 ;
        RECT 116.585 98.185 116.840 98.345 ;
        RECT 117.425 98.005 117.655 98.825 ;
        RECT 117.905 98.805 118.155 99.405 ;
        RECT 117.825 98.175 118.155 98.805 ;
        RECT 118.325 98.005 118.535 98.825 ;
        RECT 118.765 98.775 119.975 99.295 ;
        RECT 120.145 98.945 121.355 99.465 ;
        RECT 121.525 99.390 121.815 100.555 ;
        RECT 122.445 99.465 123.655 100.555 ;
        RECT 122.445 98.925 122.965 99.465 ;
        RECT 118.765 98.005 121.355 98.775 ;
        RECT 123.135 98.755 123.655 99.295 ;
        RECT 121.525 98.005 121.815 98.730 ;
        RECT 122.445 98.005 123.655 98.755 ;
        RECT 5.520 97.835 123.740 98.005 ;
        RECT 5.605 97.085 6.815 97.835 ;
        RECT 6.985 97.290 12.330 97.835 ;
        RECT 12.505 97.290 17.850 97.835 ;
        RECT 5.605 96.545 6.125 97.085 ;
        RECT 6.295 96.375 6.815 96.915 ;
        RECT 8.570 96.460 8.910 97.290 ;
        RECT 5.605 95.285 6.815 96.375 ;
        RECT 10.390 95.720 10.740 96.970 ;
        RECT 14.090 96.460 14.430 97.290 ;
        RECT 18.025 97.065 20.615 97.835 ;
        RECT 20.785 97.375 21.345 97.665 ;
        RECT 21.515 97.375 21.765 97.835 ;
        RECT 15.910 95.720 16.260 96.970 ;
        RECT 18.025 96.545 19.235 97.065 ;
        RECT 19.405 96.375 20.615 96.895 ;
        RECT 6.985 95.285 12.330 95.720 ;
        RECT 12.505 95.285 17.850 95.720 ;
        RECT 18.025 95.285 20.615 96.375 ;
        RECT 20.785 96.005 21.035 97.375 ;
        RECT 22.385 97.205 22.715 97.565 ;
        RECT 21.325 97.015 22.715 97.205 ;
        RECT 23.085 97.160 23.345 97.665 ;
        RECT 23.525 97.455 23.855 97.835 ;
        RECT 24.035 97.285 24.205 97.665 ;
        RECT 21.325 96.925 21.495 97.015 ;
        RECT 21.205 96.595 21.495 96.925 ;
        RECT 21.665 96.595 22.005 96.845 ;
        RECT 22.225 96.595 22.900 96.845 ;
        RECT 21.325 96.345 21.495 96.595 ;
        RECT 21.325 96.175 22.265 96.345 ;
        RECT 22.635 96.235 22.900 96.595 ;
        RECT 23.085 96.360 23.255 97.160 ;
        RECT 23.540 97.115 24.205 97.285 ;
        RECT 23.540 96.860 23.710 97.115 ;
        RECT 24.465 97.065 26.135 97.835 ;
        RECT 23.425 96.530 23.710 96.860 ;
        RECT 23.945 96.565 24.275 96.935 ;
        RECT 24.465 96.545 25.215 97.065 ;
        RECT 26.345 97.015 26.575 97.835 ;
        RECT 26.745 97.035 27.075 97.665 ;
        RECT 23.540 96.385 23.710 96.530 ;
        RECT 20.785 95.455 21.245 96.005 ;
        RECT 21.435 95.285 21.765 96.005 ;
        RECT 21.965 95.625 22.265 96.175 ;
        RECT 22.435 95.285 22.715 95.955 ;
        RECT 23.085 95.455 23.355 96.360 ;
        RECT 23.540 96.215 24.205 96.385 ;
        RECT 25.385 96.375 26.135 96.895 ;
        RECT 26.325 96.595 26.655 96.845 ;
        RECT 26.825 96.435 27.075 97.035 ;
        RECT 27.245 97.015 27.455 97.835 ;
        RECT 27.685 97.065 31.195 97.835 ;
        RECT 31.365 97.110 31.655 97.835 ;
        RECT 32.835 97.285 33.005 97.665 ;
        RECT 33.185 97.455 33.515 97.835 ;
        RECT 32.835 97.115 33.500 97.285 ;
        RECT 33.695 97.160 33.955 97.665 ;
        RECT 27.685 96.545 29.335 97.065 ;
        RECT 23.525 95.285 23.855 96.045 ;
        RECT 24.035 95.455 24.205 96.215 ;
        RECT 24.465 95.285 26.135 96.375 ;
        RECT 26.345 95.285 26.575 96.425 ;
        RECT 26.745 95.455 27.075 96.435 ;
        RECT 27.245 95.285 27.455 96.425 ;
        RECT 29.505 96.375 31.195 96.895 ;
        RECT 32.765 96.565 33.095 96.935 ;
        RECT 33.330 96.860 33.500 97.115 ;
        RECT 33.330 96.530 33.615 96.860 ;
        RECT 27.685 95.285 31.195 96.375 ;
        RECT 31.365 95.285 31.655 96.450 ;
        RECT 33.330 96.385 33.500 96.530 ;
        RECT 32.835 96.215 33.500 96.385 ;
        RECT 33.785 96.360 33.955 97.160 ;
        RECT 34.125 97.065 35.795 97.835 ;
        RECT 34.125 96.545 34.875 97.065 ;
        RECT 36.485 97.015 36.695 97.835 ;
        RECT 36.865 97.035 37.195 97.665 ;
        RECT 35.045 96.375 35.795 96.895 ;
        RECT 36.865 96.435 37.115 97.035 ;
        RECT 37.365 97.015 37.595 97.835 ;
        RECT 37.805 97.085 39.015 97.835 ;
        RECT 39.275 97.285 39.445 97.665 ;
        RECT 39.625 97.455 39.955 97.835 ;
        RECT 39.275 97.115 39.940 97.285 ;
        RECT 40.135 97.160 40.395 97.665 ;
        RECT 37.285 96.595 37.615 96.845 ;
        RECT 37.805 96.545 38.325 97.085 ;
        RECT 32.835 95.455 33.005 96.215 ;
        RECT 33.185 95.285 33.515 96.045 ;
        RECT 33.685 95.455 33.955 96.360 ;
        RECT 34.125 95.285 35.795 96.375 ;
        RECT 36.485 95.285 36.695 96.425 ;
        RECT 36.865 95.455 37.195 96.435 ;
        RECT 37.365 95.285 37.595 96.425 ;
        RECT 38.495 96.375 39.015 96.915 ;
        RECT 39.205 96.565 39.535 96.935 ;
        RECT 39.770 96.860 39.940 97.115 ;
        RECT 39.770 96.530 40.055 96.860 ;
        RECT 39.770 96.385 39.940 96.530 ;
        RECT 37.805 95.285 39.015 96.375 ;
        RECT 39.275 96.215 39.940 96.385 ;
        RECT 40.225 96.360 40.395 97.160 ;
        RECT 40.655 97.285 40.825 97.575 ;
        RECT 40.995 97.455 41.325 97.835 ;
        RECT 40.655 97.115 41.320 97.285 ;
        RECT 39.275 95.455 39.445 96.215 ;
        RECT 39.625 95.285 39.955 96.045 ;
        RECT 40.125 95.455 40.395 96.360 ;
        RECT 40.570 96.295 40.920 96.945 ;
        RECT 41.090 96.125 41.320 97.115 ;
        RECT 40.655 95.955 41.320 96.125 ;
        RECT 40.655 95.455 40.825 95.955 ;
        RECT 40.995 95.285 41.325 95.785 ;
        RECT 41.495 95.455 41.720 97.575 ;
        RECT 41.935 97.455 42.265 97.835 ;
        RECT 42.435 97.285 42.605 97.615 ;
        RECT 42.905 97.455 43.920 97.655 ;
        RECT 41.910 97.095 42.605 97.285 ;
        RECT 41.910 96.125 42.080 97.095 ;
        RECT 42.250 96.295 42.660 96.915 ;
        RECT 42.830 96.345 43.050 97.215 ;
        RECT 43.230 96.905 43.580 97.275 ;
        RECT 43.750 96.725 43.920 97.455 ;
        RECT 44.090 97.395 44.500 97.835 ;
        RECT 44.790 97.195 45.040 97.625 ;
        RECT 45.240 97.375 45.560 97.835 ;
        RECT 46.120 97.445 46.970 97.615 ;
        RECT 44.090 96.855 44.500 97.185 ;
        RECT 44.790 96.855 45.210 97.195 ;
        RECT 43.500 96.685 43.920 96.725 ;
        RECT 43.500 96.515 44.850 96.685 ;
        RECT 41.910 95.955 42.605 96.125 ;
        RECT 42.830 95.965 43.330 96.345 ;
        RECT 41.935 95.285 42.265 95.785 ;
        RECT 42.435 95.455 42.605 95.955 ;
        RECT 43.500 95.670 43.670 96.515 ;
        RECT 44.600 96.355 44.850 96.515 ;
        RECT 43.840 96.085 44.090 96.345 ;
        RECT 45.020 96.085 45.210 96.855 ;
        RECT 43.840 95.835 45.210 96.085 ;
        RECT 45.380 97.025 46.630 97.195 ;
        RECT 45.380 96.265 45.550 97.025 ;
        RECT 46.300 96.905 46.630 97.025 ;
        RECT 45.720 96.445 45.900 96.855 ;
        RECT 46.800 96.685 46.970 97.445 ;
        RECT 47.170 97.355 47.830 97.835 ;
        RECT 48.010 97.240 48.330 97.570 ;
        RECT 47.160 96.915 47.820 97.185 ;
        RECT 47.160 96.855 47.490 96.915 ;
        RECT 47.640 96.685 47.970 96.745 ;
        RECT 46.070 96.515 47.970 96.685 ;
        RECT 45.380 95.955 45.900 96.265 ;
        RECT 46.070 96.005 46.240 96.515 ;
        RECT 48.140 96.345 48.330 97.240 ;
        RECT 46.410 96.175 48.330 96.345 ;
        RECT 48.010 96.155 48.330 96.175 ;
        RECT 48.530 96.925 48.780 97.575 ;
        RECT 48.960 97.375 49.245 97.835 ;
        RECT 49.425 97.125 49.680 97.655 ;
        RECT 48.530 96.595 49.330 96.925 ;
        RECT 46.070 95.835 47.280 96.005 ;
        RECT 42.840 95.500 43.670 95.670 ;
        RECT 43.910 95.285 44.290 95.665 ;
        RECT 44.470 95.545 44.640 95.835 ;
        RECT 46.070 95.755 46.240 95.835 ;
        RECT 44.810 95.285 45.140 95.665 ;
        RECT 45.610 95.505 46.240 95.755 ;
        RECT 46.420 95.285 46.840 95.665 ;
        RECT 47.040 95.545 47.280 95.835 ;
        RECT 47.510 95.285 47.840 95.975 ;
        RECT 48.010 95.545 48.180 96.155 ;
        RECT 48.530 96.005 48.780 96.595 ;
        RECT 49.500 96.265 49.680 97.125 ;
        RECT 50.225 97.065 52.815 97.835 ;
        RECT 53.445 97.160 53.715 97.505 ;
        RECT 53.905 97.435 54.285 97.835 ;
        RECT 54.455 97.265 54.625 97.615 ;
        RECT 54.795 97.435 55.125 97.835 ;
        RECT 55.325 97.265 55.495 97.615 ;
        RECT 55.695 97.335 56.025 97.835 ;
        RECT 50.225 96.545 51.435 97.065 ;
        RECT 51.605 96.375 52.815 96.895 ;
        RECT 48.450 95.495 48.780 96.005 ;
        RECT 48.960 95.285 49.245 96.085 ;
        RECT 49.425 95.795 49.680 96.265 ;
        RECT 49.425 95.625 49.765 95.795 ;
        RECT 49.425 95.595 49.680 95.625 ;
        RECT 50.225 95.285 52.815 96.375 ;
        RECT 53.445 96.425 53.615 97.160 ;
        RECT 53.885 97.095 55.495 97.265 ;
        RECT 53.885 96.925 54.055 97.095 ;
        RECT 53.785 96.595 54.055 96.925 ;
        RECT 54.225 96.595 54.630 96.925 ;
        RECT 53.885 96.425 54.055 96.595 ;
        RECT 53.445 95.455 53.715 96.425 ;
        RECT 53.885 96.255 54.610 96.425 ;
        RECT 54.800 96.305 55.510 96.925 ;
        RECT 55.680 96.595 56.030 97.165 ;
        RECT 57.125 97.110 57.415 97.835 ;
        RECT 57.585 97.065 60.175 97.835 ;
        RECT 60.435 97.285 60.605 97.575 ;
        RECT 60.775 97.455 61.105 97.835 ;
        RECT 60.435 97.115 61.100 97.285 ;
        RECT 57.585 96.545 58.795 97.065 ;
        RECT 54.440 96.135 54.610 96.255 ;
        RECT 55.710 96.135 56.030 96.425 ;
        RECT 53.925 95.285 54.205 96.085 ;
        RECT 54.440 95.965 56.030 96.135 ;
        RECT 54.375 95.505 56.030 95.795 ;
        RECT 57.125 95.285 57.415 96.450 ;
        RECT 58.965 96.375 60.175 96.895 ;
        RECT 57.585 95.285 60.175 96.375 ;
        RECT 60.350 96.295 60.700 96.945 ;
        RECT 60.870 96.125 61.100 97.115 ;
        RECT 60.435 95.955 61.100 96.125 ;
        RECT 60.435 95.455 60.605 95.955 ;
        RECT 60.775 95.285 61.105 95.785 ;
        RECT 61.275 95.455 61.500 97.575 ;
        RECT 61.715 97.455 62.045 97.835 ;
        RECT 62.215 97.285 62.385 97.615 ;
        RECT 62.685 97.455 63.700 97.655 ;
        RECT 61.690 97.095 62.385 97.285 ;
        RECT 61.690 96.125 61.860 97.095 ;
        RECT 62.030 96.295 62.440 96.915 ;
        RECT 62.610 96.345 62.830 97.215 ;
        RECT 63.010 96.905 63.360 97.275 ;
        RECT 63.530 96.725 63.700 97.455 ;
        RECT 63.870 97.395 64.280 97.835 ;
        RECT 64.570 97.195 64.820 97.625 ;
        RECT 65.020 97.375 65.340 97.835 ;
        RECT 65.900 97.445 66.750 97.615 ;
        RECT 63.870 96.855 64.280 97.185 ;
        RECT 64.570 96.855 64.990 97.195 ;
        RECT 63.280 96.685 63.700 96.725 ;
        RECT 63.280 96.515 64.630 96.685 ;
        RECT 61.690 95.955 62.385 96.125 ;
        RECT 62.610 95.965 63.110 96.345 ;
        RECT 61.715 95.285 62.045 95.785 ;
        RECT 62.215 95.455 62.385 95.955 ;
        RECT 63.280 95.670 63.450 96.515 ;
        RECT 64.380 96.355 64.630 96.515 ;
        RECT 63.620 96.085 63.870 96.345 ;
        RECT 64.800 96.085 64.990 96.855 ;
        RECT 63.620 95.835 64.990 96.085 ;
        RECT 65.160 97.025 66.410 97.195 ;
        RECT 65.160 96.265 65.330 97.025 ;
        RECT 66.080 96.905 66.410 97.025 ;
        RECT 65.500 96.445 65.680 96.855 ;
        RECT 66.580 96.685 66.750 97.445 ;
        RECT 66.950 97.355 67.610 97.835 ;
        RECT 67.790 97.240 68.110 97.570 ;
        RECT 66.940 96.915 67.600 97.185 ;
        RECT 66.940 96.855 67.270 96.915 ;
        RECT 67.420 96.685 67.750 96.745 ;
        RECT 65.850 96.515 67.750 96.685 ;
        RECT 65.160 95.955 65.680 96.265 ;
        RECT 65.850 96.005 66.020 96.515 ;
        RECT 67.920 96.345 68.110 97.240 ;
        RECT 66.190 96.175 68.110 96.345 ;
        RECT 67.790 96.155 68.110 96.175 ;
        RECT 68.310 96.925 68.560 97.575 ;
        RECT 68.740 97.375 69.025 97.835 ;
        RECT 69.205 97.125 69.460 97.655 ;
        RECT 68.310 96.595 69.110 96.925 ;
        RECT 65.850 95.835 67.060 96.005 ;
        RECT 62.620 95.500 63.450 95.670 ;
        RECT 63.690 95.285 64.070 95.665 ;
        RECT 64.250 95.545 64.420 95.835 ;
        RECT 65.850 95.755 66.020 95.835 ;
        RECT 64.590 95.285 64.920 95.665 ;
        RECT 65.390 95.505 66.020 95.755 ;
        RECT 66.200 95.285 66.620 95.665 ;
        RECT 66.820 95.545 67.060 95.835 ;
        RECT 67.290 95.285 67.620 95.975 ;
        RECT 67.790 95.545 67.960 96.155 ;
        RECT 68.310 96.005 68.560 96.595 ;
        RECT 69.280 96.265 69.460 97.125 ;
        RECT 70.095 97.285 70.265 97.575 ;
        RECT 70.435 97.455 70.765 97.835 ;
        RECT 70.095 97.115 70.760 97.285 ;
        RECT 70.010 96.295 70.360 96.945 ;
        RECT 68.230 95.495 68.560 96.005 ;
        RECT 68.740 95.285 69.025 96.085 ;
        RECT 69.205 95.795 69.460 96.265 ;
        RECT 70.530 96.125 70.760 97.115 ;
        RECT 70.095 95.955 70.760 96.125 ;
        RECT 69.205 95.625 69.545 95.795 ;
        RECT 69.205 95.595 69.460 95.625 ;
        RECT 70.095 95.455 70.265 95.955 ;
        RECT 70.435 95.285 70.765 95.785 ;
        RECT 70.935 95.455 71.160 97.575 ;
        RECT 71.375 97.455 71.705 97.835 ;
        RECT 71.875 97.285 72.045 97.615 ;
        RECT 72.345 97.455 73.360 97.655 ;
        RECT 71.350 97.095 72.045 97.285 ;
        RECT 71.350 96.125 71.520 97.095 ;
        RECT 71.690 96.295 72.100 96.915 ;
        RECT 72.270 96.345 72.490 97.215 ;
        RECT 72.670 96.905 73.020 97.275 ;
        RECT 73.190 96.725 73.360 97.455 ;
        RECT 73.530 97.395 73.940 97.835 ;
        RECT 74.230 97.195 74.480 97.625 ;
        RECT 74.680 97.375 75.000 97.835 ;
        RECT 75.560 97.445 76.410 97.615 ;
        RECT 73.530 96.855 73.940 97.185 ;
        RECT 74.230 96.855 74.650 97.195 ;
        RECT 72.940 96.685 73.360 96.725 ;
        RECT 72.940 96.515 74.290 96.685 ;
        RECT 71.350 95.955 72.045 96.125 ;
        RECT 72.270 95.965 72.770 96.345 ;
        RECT 71.375 95.285 71.705 95.785 ;
        RECT 71.875 95.455 72.045 95.955 ;
        RECT 72.940 95.670 73.110 96.515 ;
        RECT 74.040 96.355 74.290 96.515 ;
        RECT 73.280 96.085 73.530 96.345 ;
        RECT 74.460 96.085 74.650 96.855 ;
        RECT 73.280 95.835 74.650 96.085 ;
        RECT 74.820 97.025 76.070 97.195 ;
        RECT 74.820 96.265 74.990 97.025 ;
        RECT 75.740 96.905 76.070 97.025 ;
        RECT 75.160 96.445 75.340 96.855 ;
        RECT 76.240 96.685 76.410 97.445 ;
        RECT 76.610 97.355 77.270 97.835 ;
        RECT 77.450 97.240 77.770 97.570 ;
        RECT 76.600 96.915 77.260 97.185 ;
        RECT 76.600 96.855 76.930 96.915 ;
        RECT 77.080 96.685 77.410 96.745 ;
        RECT 75.510 96.515 77.410 96.685 ;
        RECT 74.820 95.955 75.340 96.265 ;
        RECT 75.510 96.005 75.680 96.515 ;
        RECT 77.580 96.345 77.770 97.240 ;
        RECT 75.850 96.175 77.770 96.345 ;
        RECT 77.450 96.155 77.770 96.175 ;
        RECT 77.970 96.925 78.220 97.575 ;
        RECT 78.400 97.375 78.685 97.835 ;
        RECT 78.865 97.125 79.120 97.655 ;
        RECT 77.970 96.595 78.770 96.925 ;
        RECT 75.510 95.835 76.720 96.005 ;
        RECT 72.280 95.500 73.110 95.670 ;
        RECT 73.350 95.285 73.730 95.665 ;
        RECT 73.910 95.545 74.080 95.835 ;
        RECT 75.510 95.755 75.680 95.835 ;
        RECT 74.250 95.285 74.580 95.665 ;
        RECT 75.050 95.505 75.680 95.755 ;
        RECT 75.860 95.285 76.280 95.665 ;
        RECT 76.480 95.545 76.720 95.835 ;
        RECT 76.950 95.285 77.280 95.975 ;
        RECT 77.450 95.545 77.620 96.155 ;
        RECT 77.970 96.005 78.220 96.595 ;
        RECT 78.940 96.265 79.120 97.125 ;
        RECT 79.665 97.065 82.255 97.835 ;
        RECT 82.885 97.110 83.175 97.835 ;
        RECT 83.345 97.290 88.690 97.835 ;
        RECT 88.865 97.290 94.210 97.835 ;
        RECT 79.665 96.545 80.875 97.065 ;
        RECT 81.045 96.375 82.255 96.895 ;
        RECT 84.930 96.460 85.270 97.290 ;
        RECT 77.890 95.495 78.220 96.005 ;
        RECT 78.400 95.285 78.685 96.085 ;
        RECT 78.865 95.795 79.120 96.265 ;
        RECT 78.865 95.625 79.205 95.795 ;
        RECT 78.865 95.595 79.120 95.625 ;
        RECT 79.665 95.285 82.255 96.375 ;
        RECT 82.885 95.285 83.175 96.450 ;
        RECT 86.750 95.720 87.100 96.970 ;
        RECT 90.450 96.460 90.790 97.290 ;
        RECT 94.385 97.065 97.895 97.835 ;
        RECT 98.065 97.085 99.275 97.835 ;
        RECT 99.645 97.205 99.975 97.565 ;
        RECT 100.595 97.375 100.845 97.835 ;
        RECT 101.015 97.375 101.575 97.665 ;
        RECT 92.270 95.720 92.620 96.970 ;
        RECT 94.385 96.545 96.035 97.065 ;
        RECT 96.205 96.375 97.895 96.895 ;
        RECT 98.065 96.545 98.585 97.085 ;
        RECT 99.645 97.015 101.035 97.205 ;
        RECT 100.865 96.925 101.035 97.015 ;
        RECT 98.755 96.375 99.275 96.915 ;
        RECT 83.345 95.285 88.690 95.720 ;
        RECT 88.865 95.285 94.210 95.720 ;
        RECT 94.385 95.285 97.895 96.375 ;
        RECT 98.065 95.285 99.275 96.375 ;
        RECT 99.460 96.595 100.135 96.845 ;
        RECT 100.355 96.595 100.695 96.845 ;
        RECT 100.865 96.595 101.155 96.925 ;
        RECT 99.460 96.235 99.725 96.595 ;
        RECT 100.865 96.345 101.035 96.595 ;
        RECT 100.095 96.175 101.035 96.345 ;
        RECT 99.645 95.285 99.925 95.955 ;
        RECT 100.095 95.625 100.395 96.175 ;
        RECT 101.325 96.005 101.575 97.375 ;
        RECT 101.745 97.290 107.090 97.835 ;
        RECT 103.330 96.460 103.670 97.290 ;
        RECT 107.265 97.085 108.475 97.835 ;
        RECT 108.645 97.110 108.935 97.835 ;
        RECT 109.105 97.160 109.365 97.665 ;
        RECT 109.545 97.455 109.875 97.835 ;
        RECT 110.055 97.285 110.225 97.665 ;
        RECT 100.595 95.285 100.925 96.005 ;
        RECT 101.115 95.455 101.575 96.005 ;
        RECT 105.150 95.720 105.500 96.970 ;
        RECT 107.265 96.545 107.785 97.085 ;
        RECT 107.955 96.375 108.475 96.915 ;
        RECT 101.745 95.285 107.090 95.720 ;
        RECT 107.265 95.285 108.475 96.375 ;
        RECT 108.645 95.285 108.935 96.450 ;
        RECT 109.105 96.360 109.275 97.160 ;
        RECT 109.560 97.115 110.225 97.285 ;
        RECT 110.575 97.285 110.745 97.665 ;
        RECT 110.925 97.455 111.255 97.835 ;
        RECT 110.575 97.115 111.240 97.285 ;
        RECT 111.435 97.160 111.695 97.665 ;
        RECT 109.560 96.860 109.730 97.115 ;
        RECT 109.445 96.530 109.730 96.860 ;
        RECT 109.965 96.565 110.295 96.935 ;
        RECT 110.505 96.565 110.835 96.935 ;
        RECT 111.070 96.860 111.240 97.115 ;
        RECT 109.560 96.385 109.730 96.530 ;
        RECT 111.070 96.530 111.355 96.860 ;
        RECT 111.070 96.385 111.240 96.530 ;
        RECT 109.105 95.455 109.375 96.360 ;
        RECT 109.560 96.215 110.225 96.385 ;
        RECT 109.545 95.285 109.875 96.045 ;
        RECT 110.055 95.455 110.225 96.215 ;
        RECT 110.575 96.215 111.240 96.385 ;
        RECT 111.525 96.360 111.695 97.160 ;
        RECT 111.955 97.285 112.125 97.575 ;
        RECT 112.295 97.455 112.625 97.835 ;
        RECT 111.955 97.115 112.620 97.285 ;
        RECT 110.575 95.455 110.745 96.215 ;
        RECT 110.925 95.285 111.255 96.045 ;
        RECT 111.425 95.455 111.695 96.360 ;
        RECT 111.870 96.295 112.220 96.945 ;
        RECT 112.390 96.125 112.620 97.115 ;
        RECT 111.955 95.955 112.620 96.125 ;
        RECT 111.955 95.455 112.125 95.955 ;
        RECT 112.295 95.285 112.625 95.785 ;
        RECT 112.795 95.455 113.020 97.575 ;
        RECT 113.235 97.455 113.565 97.835 ;
        RECT 113.735 97.285 113.905 97.615 ;
        RECT 114.205 97.455 115.220 97.655 ;
        RECT 113.210 97.095 113.905 97.285 ;
        RECT 113.210 96.125 113.380 97.095 ;
        RECT 113.550 96.295 113.960 96.915 ;
        RECT 114.130 96.345 114.350 97.215 ;
        RECT 114.530 96.905 114.880 97.275 ;
        RECT 115.050 96.725 115.220 97.455 ;
        RECT 115.390 97.395 115.800 97.835 ;
        RECT 116.090 97.195 116.340 97.625 ;
        RECT 116.540 97.375 116.860 97.835 ;
        RECT 117.420 97.445 118.270 97.615 ;
        RECT 115.390 96.855 115.800 97.185 ;
        RECT 116.090 96.855 116.510 97.195 ;
        RECT 114.800 96.685 115.220 96.725 ;
        RECT 114.800 96.515 116.150 96.685 ;
        RECT 113.210 95.955 113.905 96.125 ;
        RECT 114.130 95.965 114.630 96.345 ;
        RECT 113.235 95.285 113.565 95.785 ;
        RECT 113.735 95.455 113.905 95.955 ;
        RECT 114.800 95.670 114.970 96.515 ;
        RECT 115.900 96.355 116.150 96.515 ;
        RECT 115.140 96.085 115.390 96.345 ;
        RECT 116.320 96.085 116.510 96.855 ;
        RECT 115.140 95.835 116.510 96.085 ;
        RECT 116.680 97.025 117.930 97.195 ;
        RECT 116.680 96.265 116.850 97.025 ;
        RECT 117.600 96.905 117.930 97.025 ;
        RECT 117.020 96.445 117.200 96.855 ;
        RECT 118.100 96.685 118.270 97.445 ;
        RECT 118.470 97.355 119.130 97.835 ;
        RECT 119.310 97.240 119.630 97.570 ;
        RECT 118.460 96.915 119.120 97.185 ;
        RECT 118.460 96.855 118.790 96.915 ;
        RECT 118.940 96.685 119.270 96.745 ;
        RECT 117.370 96.515 119.270 96.685 ;
        RECT 116.680 95.955 117.200 96.265 ;
        RECT 117.370 96.005 117.540 96.515 ;
        RECT 119.440 96.345 119.630 97.240 ;
        RECT 117.710 96.175 119.630 96.345 ;
        RECT 119.310 96.155 119.630 96.175 ;
        RECT 119.830 96.925 120.080 97.575 ;
        RECT 120.260 97.375 120.545 97.835 ;
        RECT 120.725 97.125 120.980 97.655 ;
        RECT 119.830 96.595 120.630 96.925 ;
        RECT 120.800 96.815 120.980 97.125 ;
        RECT 122.445 97.085 123.655 97.835 ;
        RECT 120.800 96.645 121.065 96.815 ;
        RECT 117.370 95.835 118.580 96.005 ;
        RECT 114.140 95.500 114.970 95.670 ;
        RECT 115.210 95.285 115.590 95.665 ;
        RECT 115.770 95.545 115.940 95.835 ;
        RECT 117.370 95.755 117.540 95.835 ;
        RECT 116.110 95.285 116.440 95.665 ;
        RECT 116.910 95.505 117.540 95.755 ;
        RECT 117.720 95.285 118.140 95.665 ;
        RECT 118.340 95.545 118.580 95.835 ;
        RECT 118.810 95.285 119.140 95.975 ;
        RECT 119.310 95.545 119.480 96.155 ;
        RECT 119.830 96.005 120.080 96.595 ;
        RECT 120.800 96.265 120.980 96.645 ;
        RECT 119.750 95.495 120.080 96.005 ;
        RECT 120.260 95.285 120.545 96.085 ;
        RECT 120.725 95.595 120.980 96.265 ;
        RECT 122.445 96.375 122.965 96.915 ;
        RECT 123.135 96.545 123.655 97.085 ;
        RECT 122.445 95.285 123.655 96.375 ;
        RECT 5.520 95.115 123.740 95.285 ;
        RECT 5.605 94.025 6.815 95.115 ;
        RECT 6.985 94.680 12.330 95.115 ;
        RECT 12.505 94.680 17.850 95.115 ;
        RECT 5.605 93.315 6.125 93.855 ;
        RECT 6.295 93.485 6.815 94.025 ;
        RECT 5.605 92.565 6.815 93.315 ;
        RECT 8.570 93.110 8.910 93.940 ;
        RECT 10.390 93.430 10.740 94.680 ;
        RECT 14.090 93.110 14.430 93.940 ;
        RECT 15.910 93.430 16.260 94.680 ;
        RECT 18.485 93.950 18.775 95.115 ;
        RECT 18.945 94.025 21.535 95.115 ;
        RECT 21.795 94.445 21.965 94.945 ;
        RECT 22.135 94.615 22.465 95.115 ;
        RECT 21.795 94.275 22.460 94.445 ;
        RECT 18.945 93.335 20.155 93.855 ;
        RECT 20.325 93.505 21.535 94.025 ;
        RECT 21.710 93.455 22.060 94.105 ;
        RECT 6.985 92.565 12.330 93.110 ;
        RECT 12.505 92.565 17.850 93.110 ;
        RECT 18.485 92.565 18.775 93.290 ;
        RECT 18.945 92.565 21.535 93.335 ;
        RECT 22.230 93.285 22.460 94.275 ;
        RECT 21.795 93.115 22.460 93.285 ;
        RECT 21.795 92.825 21.965 93.115 ;
        RECT 22.135 92.565 22.465 92.945 ;
        RECT 22.635 92.825 22.860 94.945 ;
        RECT 23.075 94.615 23.405 95.115 ;
        RECT 23.575 94.445 23.745 94.945 ;
        RECT 23.980 94.730 24.810 94.900 ;
        RECT 25.050 94.735 25.430 95.115 ;
        RECT 23.050 94.275 23.745 94.445 ;
        RECT 23.050 93.305 23.220 94.275 ;
        RECT 23.390 93.485 23.800 94.105 ;
        RECT 23.970 94.055 24.470 94.435 ;
        RECT 23.050 93.115 23.745 93.305 ;
        RECT 23.970 93.185 24.190 94.055 ;
        RECT 24.640 93.885 24.810 94.730 ;
        RECT 25.610 94.565 25.780 94.855 ;
        RECT 25.950 94.735 26.280 95.115 ;
        RECT 26.750 94.645 27.380 94.895 ;
        RECT 27.560 94.735 27.980 95.115 ;
        RECT 27.210 94.565 27.380 94.645 ;
        RECT 28.180 94.565 28.420 94.855 ;
        RECT 24.980 94.315 26.350 94.565 ;
        RECT 24.980 94.055 25.230 94.315 ;
        RECT 25.740 93.885 25.990 94.045 ;
        RECT 24.640 93.715 25.990 93.885 ;
        RECT 24.640 93.675 25.060 93.715 ;
        RECT 24.370 93.125 24.720 93.495 ;
        RECT 23.075 92.565 23.405 92.945 ;
        RECT 23.575 92.785 23.745 93.115 ;
        RECT 24.890 92.945 25.060 93.675 ;
        RECT 26.160 93.545 26.350 94.315 ;
        RECT 25.230 93.215 25.640 93.545 ;
        RECT 25.930 93.205 26.350 93.545 ;
        RECT 26.520 94.135 27.040 94.445 ;
        RECT 27.210 94.395 28.420 94.565 ;
        RECT 28.650 94.425 28.980 95.115 ;
        RECT 26.520 93.375 26.690 94.135 ;
        RECT 26.860 93.545 27.040 93.955 ;
        RECT 27.210 93.885 27.380 94.395 ;
        RECT 29.150 94.245 29.320 94.855 ;
        RECT 29.590 94.395 29.920 94.905 ;
        RECT 29.150 94.225 29.470 94.245 ;
        RECT 27.550 94.055 29.470 94.225 ;
        RECT 27.210 93.715 29.110 93.885 ;
        RECT 27.440 93.375 27.770 93.495 ;
        RECT 26.520 93.205 27.770 93.375 ;
        RECT 24.045 92.745 25.060 92.945 ;
        RECT 25.230 92.565 25.640 93.005 ;
        RECT 25.930 92.775 26.180 93.205 ;
        RECT 26.380 92.565 26.700 93.025 ;
        RECT 27.940 92.955 28.110 93.715 ;
        RECT 28.780 93.655 29.110 93.715 ;
        RECT 28.300 93.485 28.630 93.545 ;
        RECT 28.300 93.215 28.960 93.485 ;
        RECT 29.280 93.160 29.470 94.055 ;
        RECT 27.260 92.785 28.110 92.955 ;
        RECT 28.310 92.565 28.970 93.045 ;
        RECT 29.150 92.830 29.470 93.160 ;
        RECT 29.670 93.805 29.920 94.395 ;
        RECT 30.100 94.315 30.385 95.115 ;
        RECT 30.565 94.775 30.820 94.805 ;
        RECT 30.565 94.605 30.905 94.775 ;
        RECT 30.565 94.135 30.820 94.605 ;
        RECT 31.455 94.445 31.625 94.945 ;
        RECT 31.795 94.615 32.125 95.115 ;
        RECT 31.455 94.275 32.120 94.445 ;
        RECT 29.670 93.475 30.470 93.805 ;
        RECT 29.670 92.825 29.920 93.475 ;
        RECT 30.640 93.275 30.820 94.135 ;
        RECT 31.370 93.455 31.720 94.105 ;
        RECT 31.890 93.285 32.120 94.275 ;
        RECT 30.100 92.565 30.385 93.025 ;
        RECT 30.565 92.745 30.820 93.275 ;
        RECT 31.455 93.115 32.120 93.285 ;
        RECT 31.455 92.825 31.625 93.115 ;
        RECT 31.795 92.565 32.125 92.945 ;
        RECT 32.295 92.825 32.520 94.945 ;
        RECT 32.735 94.615 33.065 95.115 ;
        RECT 33.235 94.445 33.405 94.945 ;
        RECT 33.640 94.730 34.470 94.900 ;
        RECT 34.710 94.735 35.090 95.115 ;
        RECT 32.710 94.275 33.405 94.445 ;
        RECT 32.710 93.305 32.880 94.275 ;
        RECT 33.050 93.485 33.460 94.105 ;
        RECT 33.630 94.055 34.130 94.435 ;
        RECT 32.710 93.115 33.405 93.305 ;
        RECT 33.630 93.185 33.850 94.055 ;
        RECT 34.300 93.885 34.470 94.730 ;
        RECT 35.270 94.565 35.440 94.855 ;
        RECT 35.610 94.735 35.940 95.115 ;
        RECT 36.410 94.645 37.040 94.895 ;
        RECT 37.220 94.735 37.640 95.115 ;
        RECT 36.870 94.565 37.040 94.645 ;
        RECT 37.840 94.565 38.080 94.855 ;
        RECT 34.640 94.315 36.010 94.565 ;
        RECT 34.640 94.055 34.890 94.315 ;
        RECT 35.400 93.885 35.650 94.045 ;
        RECT 34.300 93.715 35.650 93.885 ;
        RECT 34.300 93.675 34.720 93.715 ;
        RECT 34.030 93.125 34.380 93.495 ;
        RECT 32.735 92.565 33.065 92.945 ;
        RECT 33.235 92.785 33.405 93.115 ;
        RECT 34.550 92.945 34.720 93.675 ;
        RECT 35.820 93.545 36.010 94.315 ;
        RECT 34.890 93.215 35.300 93.545 ;
        RECT 35.590 93.205 36.010 93.545 ;
        RECT 36.180 94.135 36.700 94.445 ;
        RECT 36.870 94.395 38.080 94.565 ;
        RECT 38.310 94.425 38.640 95.115 ;
        RECT 36.180 93.375 36.350 94.135 ;
        RECT 36.520 93.545 36.700 93.955 ;
        RECT 36.870 93.885 37.040 94.395 ;
        RECT 38.810 94.245 38.980 94.855 ;
        RECT 39.250 94.395 39.580 94.905 ;
        RECT 38.810 94.225 39.130 94.245 ;
        RECT 37.210 94.055 39.130 94.225 ;
        RECT 36.870 93.715 38.770 93.885 ;
        RECT 37.100 93.375 37.430 93.495 ;
        RECT 36.180 93.205 37.430 93.375 ;
        RECT 33.705 92.745 34.720 92.945 ;
        RECT 34.890 92.565 35.300 93.005 ;
        RECT 35.590 92.775 35.840 93.205 ;
        RECT 36.040 92.565 36.360 93.025 ;
        RECT 37.600 92.955 37.770 93.715 ;
        RECT 38.440 93.655 38.770 93.715 ;
        RECT 37.960 93.485 38.290 93.545 ;
        RECT 37.960 93.215 38.620 93.485 ;
        RECT 38.940 93.160 39.130 94.055 ;
        RECT 36.920 92.785 37.770 92.955 ;
        RECT 37.970 92.565 38.630 93.045 ;
        RECT 38.810 92.830 39.130 93.160 ;
        RECT 39.330 93.805 39.580 94.395 ;
        RECT 39.760 94.315 40.045 95.115 ;
        RECT 40.225 94.135 40.480 94.805 ;
        RECT 39.330 93.475 40.130 93.805 ;
        RECT 39.330 92.825 39.580 93.475 ;
        RECT 40.300 93.275 40.480 94.135 ;
        RECT 41.025 94.025 43.615 95.115 ;
        RECT 40.225 93.075 40.480 93.275 ;
        RECT 41.025 93.335 42.235 93.855 ;
        RECT 42.405 93.505 43.615 94.025 ;
        RECT 44.245 93.950 44.535 95.115 ;
        RECT 44.710 93.975 45.045 94.945 ;
        RECT 45.215 93.975 45.385 95.115 ;
        RECT 45.555 94.775 47.585 94.945 ;
        RECT 39.760 92.565 40.045 93.025 ;
        RECT 40.225 92.905 40.565 93.075 ;
        RECT 40.225 92.745 40.480 92.905 ;
        RECT 41.025 92.565 43.615 93.335 ;
        RECT 44.710 93.305 44.880 93.975 ;
        RECT 45.555 93.805 45.725 94.775 ;
        RECT 45.050 93.475 45.305 93.805 ;
        RECT 45.530 93.475 45.725 93.805 ;
        RECT 45.895 94.435 47.020 94.605 ;
        RECT 45.135 93.305 45.305 93.475 ;
        RECT 45.895 93.305 46.065 94.435 ;
        RECT 44.245 92.565 44.535 93.290 ;
        RECT 44.710 92.735 44.965 93.305 ;
        RECT 45.135 93.135 46.065 93.305 ;
        RECT 46.235 94.095 47.245 94.265 ;
        RECT 46.235 93.295 46.405 94.095 ;
        RECT 45.890 93.100 46.065 93.135 ;
        RECT 45.135 92.565 45.465 92.965 ;
        RECT 45.890 92.735 46.420 93.100 ;
        RECT 46.610 93.075 46.885 93.895 ;
        RECT 46.605 92.905 46.885 93.075 ;
        RECT 46.610 92.735 46.885 92.905 ;
        RECT 47.055 92.735 47.245 94.095 ;
        RECT 47.415 94.110 47.585 94.775 ;
        RECT 47.755 94.355 47.925 95.115 ;
        RECT 48.160 94.355 48.675 94.765 ;
        RECT 47.415 93.920 48.165 94.110 ;
        RECT 48.335 93.545 48.675 94.355 ;
        RECT 48.845 94.025 50.515 95.115 ;
        RECT 47.445 93.375 48.675 93.545 ;
        RECT 47.425 92.565 47.935 93.100 ;
        RECT 48.155 92.770 48.400 93.375 ;
        RECT 48.845 93.335 49.595 93.855 ;
        RECT 49.765 93.505 50.515 94.025 ;
        RECT 51.350 94.145 51.680 94.945 ;
        RECT 51.850 94.315 52.180 95.115 ;
        RECT 52.480 94.145 52.810 94.945 ;
        RECT 53.455 94.315 53.705 95.115 ;
        RECT 51.350 93.975 53.785 94.145 ;
        RECT 53.975 93.975 54.145 95.115 ;
        RECT 54.315 93.975 54.655 94.945 ;
        RECT 54.825 94.025 56.495 95.115 ;
        RECT 56.755 94.445 56.925 94.945 ;
        RECT 57.095 94.615 57.425 95.115 ;
        RECT 56.755 94.275 57.420 94.445 ;
        RECT 51.145 93.555 51.495 93.805 ;
        RECT 51.680 93.345 51.850 93.975 ;
        RECT 52.020 93.555 52.350 93.755 ;
        RECT 52.520 93.555 52.850 93.755 ;
        RECT 53.020 93.555 53.440 93.755 ;
        RECT 53.615 93.725 53.785 93.975 ;
        RECT 53.615 93.555 54.310 93.725 ;
        RECT 48.845 92.565 50.515 93.335 ;
        RECT 51.350 92.735 51.850 93.345 ;
        RECT 52.480 93.215 53.705 93.385 ;
        RECT 54.480 93.365 54.655 93.975 ;
        RECT 52.480 92.735 52.810 93.215 ;
        RECT 52.980 92.565 53.205 93.025 ;
        RECT 53.375 92.735 53.705 93.215 ;
        RECT 53.895 92.565 54.145 93.365 ;
        RECT 54.315 92.735 54.655 93.365 ;
        RECT 54.825 93.335 55.575 93.855 ;
        RECT 55.745 93.505 56.495 94.025 ;
        RECT 56.670 93.455 57.020 94.105 ;
        RECT 54.825 92.565 56.495 93.335 ;
        RECT 57.190 93.285 57.420 94.275 ;
        RECT 56.755 93.115 57.420 93.285 ;
        RECT 56.755 92.825 56.925 93.115 ;
        RECT 57.095 92.565 57.425 92.945 ;
        RECT 57.595 92.825 57.820 94.945 ;
        RECT 58.035 94.615 58.365 95.115 ;
        RECT 58.535 94.445 58.705 94.945 ;
        RECT 58.940 94.730 59.770 94.900 ;
        RECT 60.010 94.735 60.390 95.115 ;
        RECT 58.010 94.275 58.705 94.445 ;
        RECT 58.010 93.305 58.180 94.275 ;
        RECT 58.350 93.485 58.760 94.105 ;
        RECT 58.930 94.055 59.430 94.435 ;
        RECT 58.010 93.115 58.705 93.305 ;
        RECT 58.930 93.185 59.150 94.055 ;
        RECT 59.600 93.885 59.770 94.730 ;
        RECT 60.570 94.565 60.740 94.855 ;
        RECT 60.910 94.735 61.240 95.115 ;
        RECT 61.710 94.645 62.340 94.895 ;
        RECT 62.520 94.735 62.940 95.115 ;
        RECT 62.170 94.565 62.340 94.645 ;
        RECT 63.140 94.565 63.380 94.855 ;
        RECT 59.940 94.315 61.310 94.565 ;
        RECT 59.940 94.055 60.190 94.315 ;
        RECT 60.700 93.885 60.950 94.045 ;
        RECT 59.600 93.715 60.950 93.885 ;
        RECT 59.600 93.675 60.020 93.715 ;
        RECT 59.330 93.125 59.680 93.495 ;
        RECT 58.035 92.565 58.365 92.945 ;
        RECT 58.535 92.785 58.705 93.115 ;
        RECT 59.850 92.945 60.020 93.675 ;
        RECT 61.120 93.545 61.310 94.315 ;
        RECT 60.190 93.215 60.600 93.545 ;
        RECT 60.890 93.205 61.310 93.545 ;
        RECT 61.480 94.135 62.000 94.445 ;
        RECT 62.170 94.395 63.380 94.565 ;
        RECT 63.610 94.425 63.940 95.115 ;
        RECT 61.480 93.375 61.650 94.135 ;
        RECT 61.820 93.545 62.000 93.955 ;
        RECT 62.170 93.885 62.340 94.395 ;
        RECT 64.110 94.245 64.280 94.855 ;
        RECT 64.550 94.395 64.880 94.905 ;
        RECT 64.110 94.225 64.430 94.245 ;
        RECT 62.510 94.055 64.430 94.225 ;
        RECT 62.170 93.715 64.070 93.885 ;
        RECT 62.400 93.375 62.730 93.495 ;
        RECT 61.480 93.205 62.730 93.375 ;
        RECT 59.005 92.745 60.020 92.945 ;
        RECT 60.190 92.565 60.600 93.005 ;
        RECT 60.890 92.775 61.140 93.205 ;
        RECT 61.340 92.565 61.660 93.025 ;
        RECT 62.900 92.955 63.070 93.715 ;
        RECT 63.740 93.655 64.070 93.715 ;
        RECT 63.260 93.485 63.590 93.545 ;
        RECT 63.260 93.215 63.920 93.485 ;
        RECT 64.240 93.160 64.430 94.055 ;
        RECT 62.220 92.785 63.070 92.955 ;
        RECT 63.270 92.565 63.930 93.045 ;
        RECT 64.110 92.830 64.430 93.160 ;
        RECT 64.630 93.805 64.880 94.395 ;
        RECT 65.060 94.315 65.345 95.115 ;
        RECT 65.525 94.135 65.780 94.805 ;
        RECT 64.630 93.475 65.430 93.805 ;
        RECT 64.630 92.825 64.880 93.475 ;
        RECT 65.600 93.275 65.780 94.135 ;
        RECT 65.525 93.075 65.780 93.275 ;
        RECT 66.325 94.040 66.595 94.945 ;
        RECT 66.765 94.355 67.095 95.115 ;
        RECT 67.275 94.185 67.445 94.945 ;
        RECT 66.325 93.240 66.495 94.040 ;
        RECT 66.780 94.015 67.445 94.185 ;
        RECT 67.705 94.040 67.975 94.945 ;
        RECT 68.145 94.355 68.475 95.115 ;
        RECT 68.655 94.185 68.825 94.945 ;
        RECT 66.780 93.870 66.950 94.015 ;
        RECT 66.665 93.540 66.950 93.870 ;
        RECT 66.780 93.285 66.950 93.540 ;
        RECT 67.185 93.465 67.515 93.835 ;
        RECT 65.060 92.565 65.345 93.025 ;
        RECT 65.525 92.905 65.865 93.075 ;
        RECT 65.525 92.745 65.780 92.905 ;
        RECT 66.325 92.735 66.585 93.240 ;
        RECT 66.780 93.115 67.445 93.285 ;
        RECT 66.765 92.565 67.095 92.945 ;
        RECT 67.275 92.735 67.445 93.115 ;
        RECT 67.705 93.240 67.875 94.040 ;
        RECT 68.160 94.015 68.825 94.185 ;
        RECT 68.160 93.870 68.330 94.015 ;
        RECT 70.005 93.950 70.295 95.115 ;
        RECT 70.470 93.975 70.805 94.945 ;
        RECT 70.975 93.975 71.145 95.115 ;
        RECT 71.315 94.775 73.345 94.945 ;
        RECT 68.045 93.540 68.330 93.870 ;
        RECT 68.160 93.285 68.330 93.540 ;
        RECT 68.565 93.465 68.895 93.835 ;
        RECT 70.470 93.305 70.640 93.975 ;
        RECT 71.315 93.805 71.485 94.775 ;
        RECT 70.810 93.475 71.065 93.805 ;
        RECT 71.290 93.475 71.485 93.805 ;
        RECT 71.655 94.435 72.780 94.605 ;
        RECT 70.895 93.305 71.065 93.475 ;
        RECT 71.655 93.305 71.825 94.435 ;
        RECT 67.705 92.735 67.965 93.240 ;
        RECT 68.160 93.115 68.825 93.285 ;
        RECT 68.145 92.565 68.475 92.945 ;
        RECT 68.655 92.735 68.825 93.115 ;
        RECT 70.005 92.565 70.295 93.290 ;
        RECT 70.470 92.735 70.725 93.305 ;
        RECT 70.895 93.135 71.825 93.305 ;
        RECT 71.995 94.095 73.005 94.265 ;
        RECT 71.995 93.295 72.165 94.095 ;
        RECT 72.370 93.415 72.645 93.895 ;
        RECT 72.365 93.245 72.645 93.415 ;
        RECT 71.650 93.100 71.825 93.135 ;
        RECT 70.895 92.565 71.225 92.965 ;
        RECT 71.650 92.735 72.180 93.100 ;
        RECT 72.370 92.735 72.645 93.245 ;
        RECT 72.815 92.735 73.005 94.095 ;
        RECT 73.175 94.110 73.345 94.775 ;
        RECT 73.515 94.355 73.685 95.115 ;
        RECT 73.920 94.355 74.435 94.765 ;
        RECT 73.175 93.920 73.925 94.110 ;
        RECT 74.095 93.545 74.435 94.355 ;
        RECT 74.645 93.975 74.875 95.115 ;
        RECT 75.045 93.965 75.375 94.945 ;
        RECT 75.545 93.975 75.755 95.115 ;
        RECT 76.910 93.975 77.245 94.945 ;
        RECT 77.415 93.975 77.585 95.115 ;
        RECT 77.755 94.775 79.785 94.945 ;
        RECT 74.625 93.555 74.955 93.805 ;
        RECT 73.205 93.375 74.435 93.545 ;
        RECT 73.185 92.565 73.695 93.100 ;
        RECT 73.915 92.770 74.160 93.375 ;
        RECT 74.645 92.565 74.875 93.385 ;
        RECT 75.125 93.365 75.375 93.965 ;
        RECT 75.045 92.735 75.375 93.365 ;
        RECT 75.545 92.565 75.755 93.385 ;
        RECT 76.910 93.305 77.080 93.975 ;
        RECT 77.755 93.805 77.925 94.775 ;
        RECT 77.250 93.475 77.505 93.805 ;
        RECT 77.730 93.475 77.925 93.805 ;
        RECT 78.095 94.435 79.220 94.605 ;
        RECT 77.335 93.305 77.505 93.475 ;
        RECT 78.095 93.305 78.265 94.435 ;
        RECT 76.910 92.735 77.165 93.305 ;
        RECT 77.335 93.135 78.265 93.305 ;
        RECT 78.435 94.095 79.445 94.265 ;
        RECT 78.435 93.295 78.605 94.095 ;
        RECT 78.090 93.100 78.265 93.135 ;
        RECT 77.335 92.565 77.665 92.965 ;
        RECT 78.090 92.735 78.620 93.100 ;
        RECT 78.810 93.075 79.085 93.895 ;
        RECT 78.805 92.905 79.085 93.075 ;
        RECT 78.810 92.735 79.085 92.905 ;
        RECT 79.255 92.735 79.445 94.095 ;
        RECT 79.615 94.110 79.785 94.775 ;
        RECT 79.955 94.355 80.125 95.115 ;
        RECT 80.360 94.355 80.875 94.765 ;
        RECT 79.615 93.920 80.365 94.110 ;
        RECT 80.535 93.545 80.875 94.355 ;
        RECT 81.045 94.025 82.715 95.115 ;
        RECT 79.645 93.375 80.875 93.545 ;
        RECT 79.625 92.565 80.135 93.100 ;
        RECT 80.355 92.770 80.600 93.375 ;
        RECT 81.045 93.335 81.795 93.855 ;
        RECT 81.965 93.505 82.715 94.025 ;
        RECT 83.090 94.145 83.420 94.945 ;
        RECT 83.590 94.315 83.920 95.115 ;
        RECT 84.220 94.145 84.550 94.945 ;
        RECT 85.195 94.315 85.445 95.115 ;
        RECT 83.090 93.975 85.525 94.145 ;
        RECT 85.715 93.975 85.885 95.115 ;
        RECT 86.055 93.975 86.395 94.945 ;
        RECT 86.770 94.145 87.100 94.945 ;
        RECT 87.270 94.315 87.600 95.115 ;
        RECT 87.900 94.145 88.230 94.945 ;
        RECT 88.875 94.315 89.125 95.115 ;
        RECT 86.770 93.975 89.205 94.145 ;
        RECT 89.395 93.975 89.565 95.115 ;
        RECT 89.735 93.975 90.075 94.945 ;
        RECT 90.245 94.025 91.915 95.115 ;
        RECT 82.885 93.555 83.235 93.805 ;
        RECT 83.420 93.345 83.590 93.975 ;
        RECT 83.760 93.555 84.090 93.755 ;
        RECT 84.260 93.555 84.590 93.755 ;
        RECT 84.760 93.555 85.180 93.755 ;
        RECT 85.355 93.725 85.525 93.975 ;
        RECT 85.355 93.555 86.050 93.725 ;
        RECT 81.045 92.565 82.715 93.335 ;
        RECT 83.090 92.735 83.590 93.345 ;
        RECT 84.220 93.215 85.445 93.385 ;
        RECT 86.220 93.365 86.395 93.975 ;
        RECT 86.565 93.555 86.915 93.805 ;
        RECT 84.220 92.735 84.550 93.215 ;
        RECT 84.720 92.565 84.945 93.025 ;
        RECT 85.115 92.735 85.445 93.215 ;
        RECT 85.635 92.565 85.885 93.365 ;
        RECT 86.055 92.735 86.395 93.365 ;
        RECT 87.100 93.345 87.270 93.975 ;
        RECT 87.440 93.555 87.770 93.755 ;
        RECT 87.940 93.555 88.270 93.755 ;
        RECT 88.440 93.555 88.860 93.755 ;
        RECT 89.035 93.725 89.205 93.975 ;
        RECT 89.035 93.555 89.730 93.725 ;
        RECT 89.900 93.415 90.075 93.975 ;
        RECT 86.770 92.735 87.270 93.345 ;
        RECT 87.900 93.215 89.125 93.385 ;
        RECT 89.845 93.365 90.075 93.415 ;
        RECT 87.900 92.735 88.230 93.215 ;
        RECT 88.400 92.565 88.625 93.025 ;
        RECT 88.795 92.735 89.125 93.215 ;
        RECT 89.315 92.565 89.565 93.365 ;
        RECT 89.735 92.735 90.075 93.365 ;
        RECT 90.245 93.335 90.995 93.855 ;
        RECT 91.165 93.505 91.915 94.025 ;
        RECT 92.545 93.975 92.815 94.945 ;
        RECT 93.025 94.315 93.305 95.115 ;
        RECT 93.475 94.605 95.130 94.895 ;
        RECT 93.540 94.265 95.130 94.435 ;
        RECT 93.540 94.145 93.710 94.265 ;
        RECT 92.985 93.975 93.710 94.145 ;
        RECT 90.245 92.565 91.915 93.335 ;
        RECT 92.545 93.240 92.715 93.975 ;
        RECT 92.985 93.805 93.155 93.975 ;
        RECT 92.885 93.475 93.155 93.805 ;
        RECT 93.325 93.475 93.730 93.805 ;
        RECT 93.900 93.475 94.610 94.095 ;
        RECT 94.810 93.975 95.130 94.265 ;
        RECT 95.765 93.950 96.055 95.115 ;
        RECT 96.230 94.605 97.885 94.895 ;
        RECT 96.230 94.265 97.820 94.435 ;
        RECT 98.055 94.315 98.335 95.115 ;
        RECT 96.230 93.975 96.550 94.265 ;
        RECT 97.650 94.145 97.820 94.265 ;
        RECT 92.985 93.305 93.155 93.475 ;
        RECT 92.545 92.895 92.815 93.240 ;
        RECT 92.985 93.135 94.595 93.305 ;
        RECT 94.780 93.235 95.130 93.805 ;
        RECT 93.005 92.565 93.385 92.965 ;
        RECT 93.555 92.785 93.725 93.135 ;
        RECT 93.895 92.565 94.225 92.965 ;
        RECT 94.425 92.785 94.595 93.135 ;
        RECT 94.795 92.565 95.125 93.065 ;
        RECT 95.765 92.565 96.055 93.290 ;
        RECT 96.230 93.235 96.580 93.805 ;
        RECT 96.750 93.475 97.460 94.095 ;
        RECT 97.650 93.975 98.375 94.145 ;
        RECT 98.545 93.975 98.815 94.945 ;
        RECT 98.985 94.025 100.655 95.115 ;
        RECT 101.025 94.445 101.305 95.115 ;
        RECT 101.475 94.225 101.775 94.775 ;
        RECT 101.975 94.395 102.305 95.115 ;
        RECT 102.495 94.395 102.955 94.945 ;
        RECT 98.205 93.805 98.375 93.975 ;
        RECT 97.630 93.475 98.035 93.805 ;
        RECT 98.205 93.475 98.475 93.805 ;
        RECT 98.205 93.305 98.375 93.475 ;
        RECT 96.765 93.135 98.375 93.305 ;
        RECT 98.645 93.240 98.815 93.975 ;
        RECT 96.235 92.565 96.565 93.065 ;
        RECT 96.765 92.785 96.935 93.135 ;
        RECT 97.135 92.565 97.465 92.965 ;
        RECT 97.635 92.785 97.805 93.135 ;
        RECT 97.975 92.565 98.355 92.965 ;
        RECT 98.545 92.895 98.815 93.240 ;
        RECT 98.985 93.335 99.735 93.855 ;
        RECT 99.905 93.505 100.655 94.025 ;
        RECT 100.840 93.805 101.105 94.165 ;
        RECT 101.475 94.055 102.415 94.225 ;
        RECT 102.245 93.805 102.415 94.055 ;
        RECT 100.840 93.555 101.515 93.805 ;
        RECT 101.735 93.555 102.075 93.805 ;
        RECT 102.245 93.475 102.535 93.805 ;
        RECT 102.245 93.385 102.415 93.475 ;
        RECT 98.985 92.565 100.655 93.335 ;
        RECT 101.025 93.195 102.415 93.385 ;
        RECT 101.025 92.835 101.355 93.195 ;
        RECT 102.705 93.025 102.955 94.395 ;
        RECT 101.975 92.565 102.225 93.025 ;
        RECT 102.395 92.735 102.955 93.025 ;
        RECT 103.125 94.395 103.585 94.945 ;
        RECT 103.775 94.395 104.105 95.115 ;
        RECT 103.125 93.025 103.375 94.395 ;
        RECT 104.305 94.225 104.605 94.775 ;
        RECT 104.775 94.445 105.055 95.115 ;
        RECT 103.665 94.055 104.605 94.225 ;
        RECT 105.425 94.395 105.885 94.945 ;
        RECT 106.075 94.395 106.405 95.115 ;
        RECT 103.665 93.805 103.835 94.055 ;
        RECT 104.975 93.805 105.240 94.165 ;
        RECT 103.545 93.475 103.835 93.805 ;
        RECT 104.005 93.555 104.345 93.805 ;
        RECT 104.565 93.555 105.240 93.805 ;
        RECT 103.665 93.385 103.835 93.475 ;
        RECT 103.665 93.195 105.055 93.385 ;
        RECT 103.125 92.735 103.685 93.025 ;
        RECT 103.855 92.565 104.105 93.025 ;
        RECT 104.725 92.835 105.055 93.195 ;
        RECT 105.425 93.025 105.675 94.395 ;
        RECT 106.605 94.225 106.905 94.775 ;
        RECT 107.075 94.445 107.355 95.115 ;
        RECT 105.965 94.055 106.905 94.225 ;
        RECT 105.965 93.805 106.135 94.055 ;
        RECT 107.275 93.805 107.540 94.165 ;
        RECT 107.725 94.025 111.235 95.115 ;
        RECT 111.405 94.025 112.615 95.115 ;
        RECT 105.845 93.475 106.135 93.805 ;
        RECT 106.305 93.555 106.645 93.805 ;
        RECT 106.865 93.555 107.540 93.805 ;
        RECT 105.965 93.385 106.135 93.475 ;
        RECT 105.965 93.195 107.355 93.385 ;
        RECT 105.425 92.735 105.985 93.025 ;
        RECT 106.155 92.565 106.405 93.025 ;
        RECT 107.025 92.835 107.355 93.195 ;
        RECT 107.725 93.335 109.375 93.855 ;
        RECT 109.545 93.505 111.235 94.025 ;
        RECT 107.725 92.565 111.235 93.335 ;
        RECT 111.405 93.315 111.925 93.855 ;
        RECT 112.095 93.485 112.615 94.025 ;
        RECT 112.790 93.975 113.125 94.945 ;
        RECT 113.295 93.975 113.465 95.115 ;
        RECT 113.635 94.775 115.665 94.945 ;
        RECT 111.405 92.565 112.615 93.315 ;
        RECT 112.790 93.305 112.960 93.975 ;
        RECT 113.635 93.805 113.805 94.775 ;
        RECT 113.130 93.475 113.385 93.805 ;
        RECT 113.610 93.475 113.805 93.805 ;
        RECT 113.975 94.435 115.100 94.605 ;
        RECT 113.215 93.305 113.385 93.475 ;
        RECT 113.975 93.305 114.145 94.435 ;
        RECT 112.790 92.735 113.045 93.305 ;
        RECT 113.215 93.135 114.145 93.305 ;
        RECT 114.315 94.095 115.325 94.265 ;
        RECT 114.315 93.295 114.485 94.095 ;
        RECT 114.690 93.755 114.965 93.895 ;
        RECT 114.685 93.585 114.965 93.755 ;
        RECT 113.970 93.100 114.145 93.135 ;
        RECT 113.215 92.565 113.545 92.965 ;
        RECT 113.970 92.735 114.500 93.100 ;
        RECT 114.690 92.735 114.965 93.585 ;
        RECT 115.135 92.735 115.325 94.095 ;
        RECT 115.495 94.110 115.665 94.775 ;
        RECT 115.835 94.355 116.005 95.115 ;
        RECT 116.240 94.355 116.755 94.765 ;
        RECT 115.495 93.920 116.245 94.110 ;
        RECT 116.415 93.545 116.755 94.355 ;
        RECT 116.925 94.025 120.435 95.115 ;
        RECT 115.525 93.375 116.755 93.545 ;
        RECT 115.505 92.565 116.015 93.100 ;
        RECT 116.235 92.770 116.480 93.375 ;
        RECT 116.925 93.335 118.575 93.855 ;
        RECT 118.745 93.505 120.435 94.025 ;
        RECT 121.525 93.950 121.815 95.115 ;
        RECT 122.445 94.025 123.655 95.115 ;
        RECT 122.445 93.485 122.965 94.025 ;
        RECT 116.925 92.565 120.435 93.335 ;
        RECT 123.135 93.315 123.655 93.855 ;
        RECT 121.525 92.565 121.815 93.290 ;
        RECT 122.445 92.565 123.655 93.315 ;
        RECT 5.520 92.395 123.740 92.565 ;
        RECT 5.605 91.645 6.815 92.395 ;
        RECT 5.605 91.105 6.125 91.645 ;
        RECT 6.985 91.625 10.495 92.395 ;
        RECT 11.585 91.720 11.845 92.225 ;
        RECT 12.025 92.015 12.355 92.395 ;
        RECT 12.535 91.845 12.705 92.225 ;
        RECT 6.295 90.935 6.815 91.475 ;
        RECT 6.985 91.105 8.635 91.625 ;
        RECT 8.805 90.935 10.495 91.455 ;
        RECT 5.605 89.845 6.815 90.935 ;
        RECT 6.985 89.845 10.495 90.935 ;
        RECT 11.585 90.920 11.755 91.720 ;
        RECT 12.040 91.675 12.705 91.845 ;
        RECT 12.040 91.420 12.210 91.675 ;
        RECT 12.965 91.645 14.175 92.395 ;
        RECT 14.350 91.655 14.605 92.225 ;
        RECT 14.775 91.995 15.105 92.395 ;
        RECT 15.530 91.860 16.060 92.225 ;
        RECT 15.530 91.825 15.705 91.860 ;
        RECT 14.775 91.655 15.705 91.825 ;
        RECT 11.925 91.090 12.210 91.420 ;
        RECT 12.445 91.125 12.775 91.495 ;
        RECT 12.965 91.105 13.485 91.645 ;
        RECT 12.040 90.945 12.210 91.090 ;
        RECT 11.585 90.015 11.855 90.920 ;
        RECT 12.040 90.775 12.705 90.945 ;
        RECT 13.655 90.935 14.175 91.475 ;
        RECT 12.025 89.845 12.355 90.605 ;
        RECT 12.535 90.015 12.705 90.775 ;
        RECT 12.965 89.845 14.175 90.935 ;
        RECT 14.350 90.985 14.520 91.655 ;
        RECT 14.775 91.485 14.945 91.655 ;
        RECT 14.690 91.155 14.945 91.485 ;
        RECT 15.170 91.155 15.365 91.485 ;
        RECT 14.350 90.015 14.685 90.985 ;
        RECT 14.855 89.845 15.025 90.985 ;
        RECT 15.195 90.185 15.365 91.155 ;
        RECT 15.535 90.525 15.705 91.655 ;
        RECT 15.875 90.865 16.045 91.665 ;
        RECT 16.250 91.375 16.525 92.225 ;
        RECT 16.245 91.205 16.525 91.375 ;
        RECT 16.250 91.065 16.525 91.205 ;
        RECT 16.695 90.865 16.885 92.225 ;
        RECT 17.065 91.860 17.575 92.395 ;
        RECT 17.795 91.585 18.040 92.190 ;
        RECT 18.485 91.625 21.995 92.395 ;
        RECT 22.165 91.645 23.375 92.395 ;
        RECT 23.550 91.655 23.805 92.225 ;
        RECT 23.975 91.995 24.305 92.395 ;
        RECT 24.730 91.860 25.260 92.225 ;
        RECT 24.730 91.825 24.905 91.860 ;
        RECT 23.975 91.655 24.905 91.825 ;
        RECT 17.085 91.415 18.315 91.585 ;
        RECT 15.875 90.695 16.885 90.865 ;
        RECT 17.055 90.850 17.805 91.040 ;
        RECT 15.535 90.355 16.660 90.525 ;
        RECT 17.055 90.185 17.225 90.850 ;
        RECT 17.975 90.605 18.315 91.415 ;
        RECT 18.485 91.105 20.135 91.625 ;
        RECT 20.305 90.935 21.995 91.455 ;
        RECT 22.165 91.105 22.685 91.645 ;
        RECT 22.855 90.935 23.375 91.475 ;
        RECT 15.195 90.015 17.225 90.185 ;
        RECT 17.395 89.845 17.565 90.605 ;
        RECT 17.800 90.195 18.315 90.605 ;
        RECT 18.485 89.845 21.995 90.935 ;
        RECT 22.165 89.845 23.375 90.935 ;
        RECT 23.550 90.985 23.720 91.655 ;
        RECT 23.975 91.485 24.145 91.655 ;
        RECT 23.890 91.155 24.145 91.485 ;
        RECT 24.370 91.155 24.565 91.485 ;
        RECT 23.550 90.015 23.885 90.985 ;
        RECT 24.055 89.845 24.225 90.985 ;
        RECT 24.395 90.185 24.565 91.155 ;
        RECT 24.735 90.525 24.905 91.655 ;
        RECT 25.075 90.865 25.245 91.665 ;
        RECT 25.450 91.375 25.725 92.225 ;
        RECT 25.445 91.205 25.725 91.375 ;
        RECT 25.450 91.065 25.725 91.205 ;
        RECT 25.895 90.865 26.085 92.225 ;
        RECT 26.265 91.860 26.775 92.395 ;
        RECT 26.995 91.585 27.240 92.190 ;
        RECT 27.685 91.625 31.195 92.395 ;
        RECT 31.365 91.670 31.655 92.395 ;
        RECT 32.750 91.655 33.005 92.225 ;
        RECT 33.175 91.995 33.505 92.395 ;
        RECT 33.930 91.860 34.460 92.225 ;
        RECT 33.930 91.825 34.105 91.860 ;
        RECT 33.175 91.655 34.105 91.825 ;
        RECT 34.650 91.715 34.925 92.225 ;
        RECT 26.285 91.415 27.515 91.585 ;
        RECT 25.075 90.695 26.085 90.865 ;
        RECT 26.255 90.850 27.005 91.040 ;
        RECT 24.735 90.355 25.860 90.525 ;
        RECT 26.255 90.185 26.425 90.850 ;
        RECT 27.175 90.605 27.515 91.415 ;
        RECT 27.685 91.105 29.335 91.625 ;
        RECT 29.505 90.935 31.195 91.455 ;
        RECT 24.395 90.015 26.425 90.185 ;
        RECT 26.595 89.845 26.765 90.605 ;
        RECT 27.000 90.195 27.515 90.605 ;
        RECT 27.685 89.845 31.195 90.935 ;
        RECT 31.365 89.845 31.655 91.010 ;
        RECT 32.750 90.985 32.920 91.655 ;
        RECT 33.175 91.485 33.345 91.655 ;
        RECT 33.090 91.155 33.345 91.485 ;
        RECT 33.570 91.155 33.765 91.485 ;
        RECT 32.750 90.015 33.085 90.985 ;
        RECT 33.255 89.845 33.425 90.985 ;
        RECT 33.595 90.185 33.765 91.155 ;
        RECT 33.935 90.525 34.105 91.655 ;
        RECT 34.275 90.865 34.445 91.665 ;
        RECT 34.645 91.545 34.925 91.715 ;
        RECT 34.650 91.065 34.925 91.545 ;
        RECT 35.095 90.865 35.285 92.225 ;
        RECT 35.465 91.860 35.975 92.395 ;
        RECT 36.195 91.585 36.440 92.190 ;
        RECT 36.885 91.625 38.555 92.395 ;
        RECT 39.275 91.845 39.445 92.225 ;
        RECT 39.625 92.015 39.955 92.395 ;
        RECT 39.275 91.675 39.940 91.845 ;
        RECT 40.135 91.720 40.395 92.225 ;
        RECT 35.485 91.415 36.715 91.585 ;
        RECT 34.275 90.695 35.285 90.865 ;
        RECT 35.455 90.850 36.205 91.040 ;
        RECT 33.935 90.355 35.060 90.525 ;
        RECT 35.455 90.185 35.625 90.850 ;
        RECT 36.375 90.605 36.715 91.415 ;
        RECT 36.885 91.105 37.635 91.625 ;
        RECT 37.805 90.935 38.555 91.455 ;
        RECT 39.205 91.125 39.535 91.495 ;
        RECT 39.770 91.420 39.940 91.675 ;
        RECT 39.770 91.090 40.055 91.420 ;
        RECT 39.770 90.945 39.940 91.090 ;
        RECT 33.595 90.015 35.625 90.185 ;
        RECT 35.795 89.845 35.965 90.605 ;
        RECT 36.200 90.195 36.715 90.605 ;
        RECT 36.885 89.845 38.555 90.935 ;
        RECT 39.275 90.775 39.940 90.945 ;
        RECT 40.225 90.920 40.395 91.720 ;
        RECT 40.655 91.845 40.825 92.135 ;
        RECT 40.995 92.015 41.325 92.395 ;
        RECT 40.655 91.675 41.320 91.845 ;
        RECT 39.275 90.015 39.445 90.775 ;
        RECT 39.625 89.845 39.955 90.605 ;
        RECT 40.125 90.015 40.395 90.920 ;
        RECT 40.570 90.855 40.920 91.505 ;
        RECT 41.090 90.685 41.320 91.675 ;
        RECT 40.655 90.515 41.320 90.685 ;
        RECT 40.655 90.015 40.825 90.515 ;
        RECT 40.995 89.845 41.325 90.345 ;
        RECT 41.495 90.015 41.720 92.135 ;
        RECT 41.935 92.015 42.265 92.395 ;
        RECT 42.435 91.845 42.605 92.175 ;
        RECT 42.905 92.015 43.920 92.215 ;
        RECT 41.910 91.655 42.605 91.845 ;
        RECT 41.910 90.685 42.080 91.655 ;
        RECT 42.250 90.855 42.660 91.475 ;
        RECT 42.830 90.905 43.050 91.775 ;
        RECT 43.230 91.465 43.580 91.835 ;
        RECT 43.750 91.285 43.920 92.015 ;
        RECT 44.090 91.955 44.500 92.395 ;
        RECT 44.790 91.755 45.040 92.185 ;
        RECT 45.240 91.935 45.560 92.395 ;
        RECT 46.120 92.005 46.970 92.175 ;
        RECT 44.090 91.415 44.500 91.745 ;
        RECT 44.790 91.415 45.210 91.755 ;
        RECT 43.500 91.245 43.920 91.285 ;
        RECT 43.500 91.075 44.850 91.245 ;
        RECT 41.910 90.515 42.605 90.685 ;
        RECT 42.830 90.525 43.330 90.905 ;
        RECT 41.935 89.845 42.265 90.345 ;
        RECT 42.435 90.015 42.605 90.515 ;
        RECT 43.500 90.230 43.670 91.075 ;
        RECT 44.600 90.915 44.850 91.075 ;
        RECT 43.840 90.645 44.090 90.905 ;
        RECT 45.020 90.645 45.210 91.415 ;
        RECT 43.840 90.395 45.210 90.645 ;
        RECT 45.380 91.585 46.630 91.755 ;
        RECT 45.380 90.825 45.550 91.585 ;
        RECT 46.300 91.465 46.630 91.585 ;
        RECT 45.720 91.005 45.900 91.415 ;
        RECT 46.800 91.245 46.970 92.005 ;
        RECT 47.170 91.915 47.830 92.395 ;
        RECT 48.010 91.800 48.330 92.130 ;
        RECT 47.160 91.475 47.820 91.745 ;
        RECT 47.160 91.415 47.490 91.475 ;
        RECT 47.640 91.245 47.970 91.305 ;
        RECT 46.070 91.075 47.970 91.245 ;
        RECT 45.380 90.515 45.900 90.825 ;
        RECT 46.070 90.565 46.240 91.075 ;
        RECT 48.140 90.905 48.330 91.800 ;
        RECT 46.410 90.735 48.330 90.905 ;
        RECT 48.010 90.715 48.330 90.735 ;
        RECT 48.530 91.485 48.780 92.135 ;
        RECT 48.960 91.935 49.245 92.395 ;
        RECT 49.425 91.685 49.680 92.215 ;
        RECT 48.530 91.155 49.330 91.485 ;
        RECT 46.070 90.395 47.280 90.565 ;
        RECT 42.840 90.060 43.670 90.230 ;
        RECT 43.910 89.845 44.290 90.225 ;
        RECT 44.470 90.105 44.640 90.395 ;
        RECT 46.070 90.315 46.240 90.395 ;
        RECT 44.810 89.845 45.140 90.225 ;
        RECT 45.610 90.065 46.240 90.315 ;
        RECT 46.420 89.845 46.840 90.225 ;
        RECT 47.040 90.105 47.280 90.395 ;
        RECT 47.510 89.845 47.840 90.535 ;
        RECT 48.010 90.105 48.180 90.715 ;
        RECT 48.530 90.565 48.780 91.155 ;
        RECT 49.500 90.825 49.680 91.685 ;
        RECT 50.430 91.615 50.930 92.225 ;
        RECT 50.225 91.155 50.575 91.405 ;
        RECT 50.760 90.985 50.930 91.615 ;
        RECT 51.560 91.745 51.890 92.225 ;
        RECT 52.060 91.935 52.285 92.395 ;
        RECT 52.455 91.745 52.785 92.225 ;
        RECT 51.560 91.575 52.785 91.745 ;
        RECT 52.975 91.595 53.225 92.395 ;
        RECT 53.395 91.595 53.735 92.225 ;
        RECT 53.915 91.895 54.245 92.395 ;
        RECT 54.445 91.825 54.615 92.175 ;
        RECT 54.815 91.995 55.145 92.395 ;
        RECT 55.315 91.825 55.485 92.175 ;
        RECT 55.655 91.995 56.035 92.395 ;
        RECT 53.505 91.545 53.735 91.595 ;
        RECT 51.100 91.205 51.430 91.405 ;
        RECT 51.600 91.205 51.930 91.405 ;
        RECT 52.100 91.205 52.520 91.405 ;
        RECT 52.695 91.235 53.390 91.405 ;
        RECT 52.695 90.985 52.865 91.235 ;
        RECT 53.560 90.985 53.735 91.545 ;
        RECT 53.910 91.155 54.260 91.725 ;
        RECT 54.445 91.655 56.055 91.825 ;
        RECT 56.225 91.720 56.495 92.065 ;
        RECT 55.885 91.485 56.055 91.655 ;
        RECT 48.450 90.055 48.780 90.565 ;
        RECT 48.960 89.845 49.245 90.645 ;
        RECT 49.425 90.355 49.680 90.825 ;
        RECT 50.430 90.815 52.865 90.985 ;
        RECT 49.425 90.185 49.765 90.355 ;
        RECT 49.425 90.155 49.680 90.185 ;
        RECT 50.430 90.015 50.760 90.815 ;
        RECT 50.930 89.845 51.260 90.645 ;
        RECT 51.560 90.015 51.890 90.815 ;
        RECT 52.535 89.845 52.785 90.645 ;
        RECT 53.055 89.845 53.225 90.985 ;
        RECT 53.395 90.015 53.735 90.985 ;
        RECT 53.910 90.695 54.230 90.985 ;
        RECT 54.430 90.865 55.140 91.485 ;
        RECT 55.310 91.155 55.715 91.485 ;
        RECT 55.885 91.155 56.155 91.485 ;
        RECT 55.885 90.985 56.055 91.155 ;
        RECT 56.325 90.985 56.495 91.720 ;
        RECT 57.125 91.670 57.415 92.395 ;
        RECT 57.585 91.625 61.095 92.395 ;
        RECT 57.585 91.105 59.235 91.625 ;
        RECT 61.305 91.575 61.535 92.395 ;
        RECT 61.705 91.595 62.035 92.225 ;
        RECT 55.330 90.815 56.055 90.985 ;
        RECT 55.330 90.695 55.500 90.815 ;
        RECT 53.910 90.525 55.500 90.695 ;
        RECT 53.910 90.065 55.565 90.355 ;
        RECT 55.735 89.845 56.015 90.645 ;
        RECT 56.225 90.015 56.495 90.985 ;
        RECT 57.125 89.845 57.415 91.010 ;
        RECT 59.405 90.935 61.095 91.455 ;
        RECT 61.285 91.155 61.615 91.405 ;
        RECT 61.785 90.995 62.035 91.595 ;
        RECT 62.205 91.575 62.415 92.395 ;
        RECT 63.380 91.585 63.625 92.190 ;
        RECT 63.845 91.860 64.355 92.395 ;
        RECT 57.585 89.845 61.095 90.935 ;
        RECT 61.305 89.845 61.535 90.985 ;
        RECT 61.705 90.015 62.035 90.995 ;
        RECT 63.105 91.415 64.335 91.585 ;
        RECT 62.205 89.845 62.415 90.985 ;
        RECT 63.105 90.605 63.445 91.415 ;
        RECT 63.615 90.850 64.365 91.040 ;
        RECT 63.105 90.195 63.620 90.605 ;
        RECT 63.855 89.845 64.025 90.605 ;
        RECT 64.195 90.185 64.365 90.850 ;
        RECT 64.535 90.865 64.725 92.225 ;
        RECT 64.895 92.055 65.170 92.225 ;
        RECT 64.895 91.885 65.175 92.055 ;
        RECT 64.895 91.065 65.170 91.885 ;
        RECT 65.360 91.860 65.890 92.225 ;
        RECT 66.315 91.995 66.645 92.395 ;
        RECT 65.715 91.825 65.890 91.860 ;
        RECT 65.375 90.865 65.545 91.665 ;
        RECT 64.535 90.695 65.545 90.865 ;
        RECT 65.715 91.655 66.645 91.825 ;
        RECT 66.815 91.655 67.070 92.225 ;
        RECT 67.245 91.850 72.590 92.395 ;
        RECT 72.765 91.850 78.110 92.395 ;
        RECT 65.715 90.525 65.885 91.655 ;
        RECT 66.475 91.485 66.645 91.655 ;
        RECT 64.760 90.355 65.885 90.525 ;
        RECT 66.055 91.155 66.250 91.485 ;
        RECT 66.475 91.155 66.730 91.485 ;
        RECT 66.055 90.185 66.225 91.155 ;
        RECT 66.900 90.985 67.070 91.655 ;
        RECT 68.830 91.020 69.170 91.850 ;
        RECT 64.195 90.015 66.225 90.185 ;
        RECT 66.395 89.845 66.565 90.985 ;
        RECT 66.735 90.015 67.070 90.985 ;
        RECT 70.650 90.280 71.000 91.530 ;
        RECT 74.350 91.020 74.690 91.850 ;
        RECT 78.285 91.625 79.955 92.395 ;
        RECT 80.585 91.720 80.845 92.225 ;
        RECT 81.025 92.015 81.355 92.395 ;
        RECT 81.535 91.845 81.705 92.225 ;
        RECT 76.170 90.280 76.520 91.530 ;
        RECT 78.285 91.105 79.035 91.625 ;
        RECT 79.205 90.935 79.955 91.455 ;
        RECT 67.245 89.845 72.590 90.280 ;
        RECT 72.765 89.845 78.110 90.280 ;
        RECT 78.285 89.845 79.955 90.935 ;
        RECT 80.585 90.920 80.755 91.720 ;
        RECT 81.040 91.675 81.705 91.845 ;
        RECT 81.040 91.420 81.210 91.675 ;
        RECT 82.885 91.670 83.175 92.395 ;
        RECT 83.350 91.655 83.605 92.225 ;
        RECT 83.775 91.995 84.105 92.395 ;
        RECT 84.530 91.860 85.060 92.225 ;
        RECT 84.530 91.825 84.705 91.860 ;
        RECT 83.775 91.655 84.705 91.825 ;
        RECT 80.925 91.090 81.210 91.420 ;
        RECT 81.445 91.125 81.775 91.495 ;
        RECT 81.040 90.945 81.210 91.090 ;
        RECT 80.585 90.015 80.855 90.920 ;
        RECT 81.040 90.775 81.705 90.945 ;
        RECT 81.025 89.845 81.355 90.605 ;
        RECT 81.535 90.015 81.705 90.775 ;
        RECT 82.885 89.845 83.175 91.010 ;
        RECT 83.350 90.985 83.520 91.655 ;
        RECT 83.775 91.485 83.945 91.655 ;
        RECT 83.690 91.155 83.945 91.485 ;
        RECT 84.170 91.155 84.365 91.485 ;
        RECT 83.350 90.015 83.685 90.985 ;
        RECT 83.855 89.845 84.025 90.985 ;
        RECT 84.195 90.185 84.365 91.155 ;
        RECT 84.535 90.525 84.705 91.655 ;
        RECT 84.875 90.865 85.045 91.665 ;
        RECT 85.250 91.375 85.525 92.225 ;
        RECT 85.245 91.205 85.525 91.375 ;
        RECT 85.250 91.065 85.525 91.205 ;
        RECT 85.695 90.865 85.885 92.225 ;
        RECT 86.065 91.860 86.575 92.395 ;
        RECT 86.795 91.585 87.040 92.190 ;
        RECT 87.690 91.615 88.190 92.225 ;
        RECT 86.085 91.415 87.315 91.585 ;
        RECT 84.875 90.695 85.885 90.865 ;
        RECT 86.055 90.850 86.805 91.040 ;
        RECT 84.535 90.355 85.660 90.525 ;
        RECT 86.055 90.185 86.225 90.850 ;
        RECT 86.975 90.605 87.315 91.415 ;
        RECT 87.485 91.155 87.835 91.405 ;
        RECT 88.020 90.985 88.190 91.615 ;
        RECT 88.820 91.745 89.150 92.225 ;
        RECT 89.320 91.935 89.545 92.395 ;
        RECT 89.715 91.745 90.045 92.225 ;
        RECT 88.820 91.575 90.045 91.745 ;
        RECT 90.235 91.595 90.485 92.395 ;
        RECT 90.655 91.595 90.995 92.225 ;
        RECT 91.175 91.895 91.505 92.395 ;
        RECT 91.705 91.825 91.875 92.175 ;
        RECT 92.075 91.995 92.405 92.395 ;
        RECT 92.575 91.825 92.745 92.175 ;
        RECT 92.915 91.995 93.295 92.395 ;
        RECT 90.765 91.545 90.995 91.595 ;
        RECT 88.360 91.205 88.690 91.405 ;
        RECT 88.860 91.205 89.190 91.405 ;
        RECT 89.360 91.205 89.780 91.405 ;
        RECT 89.955 91.235 90.650 91.405 ;
        RECT 89.955 90.985 90.125 91.235 ;
        RECT 90.820 90.985 90.995 91.545 ;
        RECT 91.170 91.155 91.520 91.725 ;
        RECT 91.705 91.655 93.315 91.825 ;
        RECT 93.485 91.720 93.755 92.065 ;
        RECT 93.925 91.850 99.270 92.395 ;
        RECT 99.445 91.850 104.790 92.395 ;
        RECT 93.145 91.485 93.315 91.655 ;
        RECT 91.690 91.035 92.400 91.485 ;
        RECT 92.570 91.155 92.975 91.485 ;
        RECT 93.145 91.155 93.415 91.485 ;
        RECT 84.195 90.015 86.225 90.185 ;
        RECT 86.395 89.845 86.565 90.605 ;
        RECT 86.800 90.195 87.315 90.605 ;
        RECT 87.690 90.815 90.125 90.985 ;
        RECT 87.690 90.015 88.020 90.815 ;
        RECT 88.190 89.845 88.520 90.645 ;
        RECT 88.820 90.015 89.150 90.815 ;
        RECT 89.795 89.845 90.045 90.645 ;
        RECT 90.315 89.845 90.485 90.985 ;
        RECT 90.655 90.015 90.995 90.985 ;
        RECT 91.170 90.695 91.490 90.985 ;
        RECT 91.685 90.865 92.400 91.035 ;
        RECT 93.145 90.985 93.315 91.155 ;
        RECT 93.585 90.985 93.755 91.720 ;
        RECT 95.510 91.020 95.850 91.850 ;
        RECT 92.590 90.815 93.315 90.985 ;
        RECT 92.590 90.695 92.760 90.815 ;
        RECT 91.170 90.525 92.760 90.695 ;
        RECT 91.170 90.065 92.825 90.355 ;
        RECT 92.995 89.845 93.275 90.645 ;
        RECT 93.485 90.015 93.755 90.985 ;
        RECT 97.330 90.280 97.680 91.530 ;
        RECT 101.030 91.020 101.370 91.850 ;
        RECT 104.965 91.625 108.475 92.395 ;
        RECT 108.645 91.670 108.935 92.395 ;
        RECT 109.105 91.850 114.450 92.395 ;
        RECT 114.625 91.850 119.970 92.395 ;
        RECT 102.850 90.280 103.200 91.530 ;
        RECT 104.965 91.105 106.615 91.625 ;
        RECT 106.785 90.935 108.475 91.455 ;
        RECT 110.690 91.020 111.030 91.850 ;
        RECT 93.925 89.845 99.270 90.280 ;
        RECT 99.445 89.845 104.790 90.280 ;
        RECT 104.965 89.845 108.475 90.935 ;
        RECT 108.645 89.845 108.935 91.010 ;
        RECT 112.510 90.280 112.860 91.530 ;
        RECT 116.210 91.020 116.550 91.850 ;
        RECT 120.145 91.625 121.815 92.395 ;
        RECT 122.445 91.645 123.655 92.395 ;
        RECT 118.030 90.280 118.380 91.530 ;
        RECT 120.145 91.105 120.895 91.625 ;
        RECT 121.065 90.935 121.815 91.455 ;
        RECT 109.105 89.845 114.450 90.280 ;
        RECT 114.625 89.845 119.970 90.280 ;
        RECT 120.145 89.845 121.815 90.935 ;
        RECT 122.445 90.935 122.965 91.475 ;
        RECT 123.135 91.105 123.655 91.645 ;
        RECT 122.445 89.845 123.655 90.935 ;
        RECT 5.520 89.675 123.740 89.845 ;
        RECT 5.605 88.585 6.815 89.675 ;
        RECT 6.985 88.585 8.655 89.675 ;
        RECT 8.915 89.005 9.085 89.505 ;
        RECT 9.255 89.175 9.585 89.675 ;
        RECT 8.915 88.835 9.580 89.005 ;
        RECT 5.605 87.875 6.125 88.415 ;
        RECT 6.295 88.045 6.815 88.585 ;
        RECT 6.985 87.895 7.735 88.415 ;
        RECT 7.905 88.065 8.655 88.585 ;
        RECT 8.830 88.015 9.180 88.665 ;
        RECT 5.605 87.125 6.815 87.875 ;
        RECT 6.985 87.125 8.655 87.895 ;
        RECT 9.350 87.845 9.580 88.835 ;
        RECT 8.915 87.675 9.580 87.845 ;
        RECT 8.915 87.385 9.085 87.675 ;
        RECT 9.255 87.125 9.585 87.505 ;
        RECT 9.755 87.385 9.980 89.505 ;
        RECT 10.195 89.175 10.525 89.675 ;
        RECT 10.695 89.005 10.865 89.505 ;
        RECT 11.100 89.290 11.930 89.460 ;
        RECT 12.170 89.295 12.550 89.675 ;
        RECT 10.170 88.835 10.865 89.005 ;
        RECT 10.170 87.865 10.340 88.835 ;
        RECT 10.510 88.045 10.920 88.665 ;
        RECT 11.090 88.615 11.590 88.995 ;
        RECT 10.170 87.675 10.865 87.865 ;
        RECT 11.090 87.745 11.310 88.615 ;
        RECT 11.760 88.445 11.930 89.290 ;
        RECT 12.730 89.125 12.900 89.415 ;
        RECT 13.070 89.295 13.400 89.675 ;
        RECT 13.870 89.205 14.500 89.455 ;
        RECT 14.680 89.295 15.100 89.675 ;
        RECT 14.330 89.125 14.500 89.205 ;
        RECT 15.300 89.125 15.540 89.415 ;
        RECT 12.100 88.875 13.470 89.125 ;
        RECT 12.100 88.615 12.350 88.875 ;
        RECT 12.860 88.445 13.110 88.605 ;
        RECT 11.760 88.275 13.110 88.445 ;
        RECT 11.760 88.235 12.180 88.275 ;
        RECT 11.490 87.685 11.840 88.055 ;
        RECT 10.195 87.125 10.525 87.505 ;
        RECT 10.695 87.345 10.865 87.675 ;
        RECT 12.010 87.505 12.180 88.235 ;
        RECT 13.280 88.105 13.470 88.875 ;
        RECT 12.350 87.775 12.760 88.105 ;
        RECT 13.050 87.765 13.470 88.105 ;
        RECT 13.640 88.695 14.160 89.005 ;
        RECT 14.330 88.955 15.540 89.125 ;
        RECT 15.770 88.985 16.100 89.675 ;
        RECT 13.640 87.935 13.810 88.695 ;
        RECT 13.980 88.105 14.160 88.515 ;
        RECT 14.330 88.445 14.500 88.955 ;
        RECT 16.270 88.805 16.440 89.415 ;
        RECT 16.710 88.955 17.040 89.465 ;
        RECT 16.270 88.785 16.590 88.805 ;
        RECT 14.670 88.615 16.590 88.785 ;
        RECT 14.330 88.275 16.230 88.445 ;
        RECT 14.560 87.935 14.890 88.055 ;
        RECT 13.640 87.765 14.890 87.935 ;
        RECT 11.165 87.305 12.180 87.505 ;
        RECT 12.350 87.125 12.760 87.565 ;
        RECT 13.050 87.335 13.300 87.765 ;
        RECT 13.500 87.125 13.820 87.585 ;
        RECT 15.060 87.515 15.230 88.275 ;
        RECT 15.900 88.215 16.230 88.275 ;
        RECT 15.420 88.045 15.750 88.105 ;
        RECT 15.420 87.775 16.080 88.045 ;
        RECT 16.400 87.720 16.590 88.615 ;
        RECT 14.380 87.345 15.230 87.515 ;
        RECT 15.430 87.125 16.090 87.605 ;
        RECT 16.270 87.390 16.590 87.720 ;
        RECT 16.790 88.365 17.040 88.955 ;
        RECT 17.220 88.875 17.505 89.675 ;
        RECT 17.685 89.335 17.940 89.365 ;
        RECT 17.685 89.165 18.025 89.335 ;
        RECT 17.685 88.695 17.940 89.165 ;
        RECT 16.790 88.035 17.590 88.365 ;
        RECT 16.790 87.385 17.040 88.035 ;
        RECT 17.760 87.835 17.940 88.695 ;
        RECT 18.485 88.510 18.775 89.675 ;
        RECT 18.945 89.240 24.290 89.675 ;
        RECT 17.220 87.125 17.505 87.585 ;
        RECT 17.685 87.305 17.940 87.835 ;
        RECT 18.485 87.125 18.775 87.850 ;
        RECT 20.530 87.670 20.870 88.500 ;
        RECT 22.350 87.990 22.700 89.240 ;
        RECT 24.470 89.165 26.125 89.455 ;
        RECT 24.470 88.825 26.060 88.995 ;
        RECT 26.295 88.875 26.575 89.675 ;
        RECT 24.470 88.535 24.790 88.825 ;
        RECT 25.890 88.705 26.060 88.825 ;
        RECT 24.985 88.485 25.700 88.655 ;
        RECT 25.890 88.535 26.615 88.705 ;
        RECT 26.785 88.535 27.055 89.505 ;
        RECT 27.225 89.240 32.570 89.675 ;
        RECT 24.470 87.795 24.820 88.365 ;
        RECT 24.990 88.035 25.700 88.485 ;
        RECT 26.445 88.365 26.615 88.535 ;
        RECT 25.870 88.035 26.275 88.365 ;
        RECT 26.445 88.035 26.715 88.365 ;
        RECT 26.445 87.865 26.615 88.035 ;
        RECT 25.005 87.695 26.615 87.865 ;
        RECT 26.885 87.800 27.055 88.535 ;
        RECT 18.945 87.125 24.290 87.670 ;
        RECT 24.475 87.125 24.805 87.625 ;
        RECT 25.005 87.345 25.175 87.695 ;
        RECT 25.375 87.125 25.705 87.525 ;
        RECT 25.875 87.345 26.045 87.695 ;
        RECT 26.215 87.125 26.595 87.525 ;
        RECT 26.785 87.455 27.055 87.800 ;
        RECT 28.810 87.670 29.150 88.500 ;
        RECT 30.630 87.990 30.980 89.240 ;
        RECT 32.745 88.585 33.955 89.675 ;
        RECT 34.130 89.165 35.785 89.455 ;
        RECT 32.745 87.875 33.265 88.415 ;
        RECT 33.435 88.045 33.955 88.585 ;
        RECT 34.130 88.825 35.720 88.995 ;
        RECT 35.955 88.875 36.235 89.675 ;
        RECT 34.130 88.535 34.450 88.825 ;
        RECT 35.550 88.705 35.720 88.825 ;
        RECT 27.225 87.125 32.570 87.670 ;
        RECT 32.745 87.125 33.955 87.875 ;
        RECT 34.130 87.795 34.480 88.365 ;
        RECT 34.650 88.035 35.360 88.655 ;
        RECT 35.550 88.535 36.275 88.705 ;
        RECT 36.445 88.535 36.715 89.505 ;
        RECT 36.885 89.240 42.230 89.675 ;
        RECT 36.105 88.365 36.275 88.535 ;
        RECT 35.530 88.035 35.935 88.365 ;
        RECT 36.105 88.035 36.375 88.365 ;
        RECT 36.105 87.865 36.275 88.035 ;
        RECT 34.665 87.695 36.275 87.865 ;
        RECT 36.545 87.800 36.715 88.535 ;
        RECT 34.135 87.125 34.465 87.625 ;
        RECT 34.665 87.345 34.835 87.695 ;
        RECT 35.035 87.125 35.365 87.525 ;
        RECT 35.535 87.345 35.705 87.695 ;
        RECT 35.875 87.125 36.255 87.525 ;
        RECT 36.445 87.455 36.715 87.800 ;
        RECT 38.470 87.670 38.810 88.500 ;
        RECT 40.290 87.990 40.640 89.240 ;
        RECT 42.905 88.535 43.135 89.675 ;
        RECT 43.305 88.525 43.635 89.505 ;
        RECT 43.805 88.535 44.015 89.675 ;
        RECT 42.885 88.115 43.215 88.365 ;
        RECT 36.885 87.125 42.230 87.670 ;
        RECT 42.905 87.125 43.135 87.945 ;
        RECT 43.385 87.925 43.635 88.525 ;
        RECT 44.245 88.510 44.535 89.675 ;
        RECT 45.630 88.535 45.965 89.505 ;
        RECT 46.135 88.535 46.305 89.675 ;
        RECT 46.475 89.335 48.505 89.505 ;
        RECT 43.305 87.295 43.635 87.925 ;
        RECT 43.805 87.125 44.015 87.945 ;
        RECT 45.630 87.865 45.800 88.535 ;
        RECT 46.475 88.365 46.645 89.335 ;
        RECT 45.970 88.035 46.225 88.365 ;
        RECT 46.450 88.035 46.645 88.365 ;
        RECT 46.815 88.995 47.940 89.165 ;
        RECT 46.055 87.865 46.225 88.035 ;
        RECT 46.815 87.865 46.985 88.995 ;
        RECT 44.245 87.125 44.535 87.850 ;
        RECT 45.630 87.295 45.885 87.865 ;
        RECT 46.055 87.695 46.985 87.865 ;
        RECT 47.155 88.655 48.165 88.825 ;
        RECT 47.155 87.855 47.325 88.655 ;
        RECT 47.530 88.315 47.805 88.455 ;
        RECT 47.525 88.145 47.805 88.315 ;
        RECT 46.810 87.660 46.985 87.695 ;
        RECT 46.055 87.125 46.385 87.525 ;
        RECT 46.810 87.295 47.340 87.660 ;
        RECT 47.530 87.295 47.805 88.145 ;
        RECT 47.975 87.295 48.165 88.655 ;
        RECT 48.335 88.670 48.505 89.335 ;
        RECT 48.675 88.915 48.845 89.675 ;
        RECT 49.080 88.915 49.595 89.325 ;
        RECT 49.765 89.240 55.110 89.675 ;
        RECT 48.335 88.480 49.085 88.670 ;
        RECT 49.255 88.105 49.595 88.915 ;
        RECT 48.365 87.935 49.595 88.105 ;
        RECT 48.345 87.125 48.855 87.660 ;
        RECT 49.075 87.330 49.320 87.935 ;
        RECT 51.350 87.670 51.690 88.500 ;
        RECT 53.170 87.990 53.520 89.240 ;
        RECT 55.285 88.585 58.795 89.675 ;
        RECT 55.285 87.895 56.935 88.415 ;
        RECT 57.105 88.065 58.795 88.585 ;
        RECT 59.425 88.600 59.695 89.505 ;
        RECT 59.865 88.915 60.195 89.675 ;
        RECT 60.375 88.745 60.545 89.505 ;
        RECT 60.805 89.240 66.150 89.675 ;
        RECT 49.765 87.125 55.110 87.670 ;
        RECT 55.285 87.125 58.795 87.895 ;
        RECT 59.425 87.800 59.595 88.600 ;
        RECT 59.880 88.575 60.545 88.745 ;
        RECT 59.880 88.430 60.050 88.575 ;
        RECT 59.765 88.100 60.050 88.430 ;
        RECT 59.880 87.845 60.050 88.100 ;
        RECT 60.285 88.025 60.615 88.395 ;
        RECT 59.425 87.295 59.685 87.800 ;
        RECT 59.880 87.675 60.545 87.845 ;
        RECT 59.865 87.125 60.195 87.505 ;
        RECT 60.375 87.295 60.545 87.675 ;
        RECT 62.390 87.670 62.730 88.500 ;
        RECT 64.210 87.990 64.560 89.240 ;
        RECT 66.530 88.705 66.860 89.505 ;
        RECT 67.030 88.875 67.360 89.675 ;
        RECT 67.660 88.705 67.990 89.505 ;
        RECT 68.635 88.875 68.885 89.675 ;
        RECT 66.530 88.535 68.965 88.705 ;
        RECT 69.155 88.535 69.325 89.675 ;
        RECT 69.495 88.535 69.835 89.505 ;
        RECT 66.325 88.115 66.675 88.365 ;
        RECT 66.860 87.905 67.030 88.535 ;
        RECT 67.200 88.115 67.530 88.315 ;
        RECT 67.700 88.115 68.030 88.315 ;
        RECT 68.200 88.115 68.620 88.315 ;
        RECT 68.795 88.285 68.965 88.535 ;
        RECT 68.795 88.115 69.490 88.285 ;
        RECT 60.805 87.125 66.150 87.670 ;
        RECT 66.530 87.295 67.030 87.905 ;
        RECT 67.660 87.775 68.885 87.945 ;
        RECT 69.660 87.925 69.835 88.535 ;
        RECT 70.005 88.510 70.295 89.675 ;
        RECT 70.465 89.240 75.810 89.675 ;
        RECT 67.660 87.295 67.990 87.775 ;
        RECT 68.160 87.125 68.385 87.585 ;
        RECT 68.555 87.295 68.885 87.775 ;
        RECT 69.075 87.125 69.325 87.925 ;
        RECT 69.495 87.295 69.835 87.925 ;
        RECT 70.005 87.125 70.295 87.850 ;
        RECT 72.050 87.670 72.390 88.500 ;
        RECT 73.870 87.990 74.220 89.240 ;
        RECT 75.985 88.585 77.655 89.675 ;
        RECT 78.375 89.005 78.545 89.505 ;
        RECT 78.715 89.175 79.045 89.675 ;
        RECT 78.375 88.835 79.040 89.005 ;
        RECT 75.985 87.895 76.735 88.415 ;
        RECT 76.905 88.065 77.655 88.585 ;
        RECT 78.290 88.015 78.640 88.665 ;
        RECT 70.465 87.125 75.810 87.670 ;
        RECT 75.985 87.125 77.655 87.895 ;
        RECT 78.810 87.845 79.040 88.835 ;
        RECT 78.375 87.675 79.040 87.845 ;
        RECT 78.375 87.385 78.545 87.675 ;
        RECT 78.715 87.125 79.045 87.505 ;
        RECT 79.215 87.385 79.440 89.505 ;
        RECT 79.655 89.175 79.985 89.675 ;
        RECT 80.155 89.005 80.325 89.505 ;
        RECT 80.560 89.290 81.390 89.460 ;
        RECT 81.630 89.295 82.010 89.675 ;
        RECT 79.630 88.835 80.325 89.005 ;
        RECT 79.630 87.865 79.800 88.835 ;
        RECT 79.970 88.045 80.380 88.665 ;
        RECT 80.550 88.615 81.050 88.995 ;
        RECT 79.630 87.675 80.325 87.865 ;
        RECT 80.550 87.745 80.770 88.615 ;
        RECT 81.220 88.445 81.390 89.290 ;
        RECT 82.190 89.125 82.360 89.415 ;
        RECT 82.530 89.295 82.860 89.675 ;
        RECT 83.330 89.205 83.960 89.455 ;
        RECT 84.140 89.295 84.560 89.675 ;
        RECT 83.790 89.125 83.960 89.205 ;
        RECT 84.760 89.125 85.000 89.415 ;
        RECT 81.560 88.875 82.930 89.125 ;
        RECT 81.560 88.615 81.810 88.875 ;
        RECT 82.320 88.445 82.570 88.605 ;
        RECT 81.220 88.275 82.570 88.445 ;
        RECT 81.220 88.235 81.640 88.275 ;
        RECT 80.950 87.685 81.300 88.055 ;
        RECT 79.655 87.125 79.985 87.505 ;
        RECT 80.155 87.345 80.325 87.675 ;
        RECT 81.470 87.505 81.640 88.235 ;
        RECT 82.740 88.105 82.930 88.875 ;
        RECT 81.810 87.775 82.220 88.105 ;
        RECT 82.510 87.765 82.930 88.105 ;
        RECT 83.100 88.695 83.620 89.005 ;
        RECT 83.790 88.955 85.000 89.125 ;
        RECT 85.230 88.985 85.560 89.675 ;
        RECT 83.100 87.935 83.270 88.695 ;
        RECT 83.440 88.105 83.620 88.515 ;
        RECT 83.790 88.445 83.960 88.955 ;
        RECT 85.730 88.805 85.900 89.415 ;
        RECT 86.170 88.955 86.500 89.465 ;
        RECT 85.730 88.785 86.050 88.805 ;
        RECT 84.130 88.615 86.050 88.785 ;
        RECT 83.790 88.275 85.690 88.445 ;
        RECT 84.020 87.935 84.350 88.055 ;
        RECT 83.100 87.765 84.350 87.935 ;
        RECT 80.625 87.305 81.640 87.505 ;
        RECT 81.810 87.125 82.220 87.565 ;
        RECT 82.510 87.335 82.760 87.765 ;
        RECT 82.960 87.125 83.280 87.585 ;
        RECT 84.520 87.515 84.690 88.275 ;
        RECT 85.360 88.215 85.690 88.275 ;
        RECT 84.880 88.045 85.210 88.105 ;
        RECT 84.880 87.775 85.540 88.045 ;
        RECT 85.860 87.720 86.050 88.615 ;
        RECT 83.840 87.345 84.690 87.515 ;
        RECT 84.890 87.125 85.550 87.605 ;
        RECT 85.730 87.390 86.050 87.720 ;
        RECT 86.250 88.365 86.500 88.955 ;
        RECT 86.680 88.875 86.965 89.675 ;
        RECT 87.145 88.995 87.400 89.365 ;
        RECT 87.145 88.825 87.485 88.995 ;
        RECT 87.145 88.695 87.400 88.825 ;
        RECT 86.250 88.035 87.050 88.365 ;
        RECT 86.250 87.385 86.500 88.035 ;
        RECT 87.220 87.835 87.400 88.695 ;
        RECT 88.005 88.535 88.215 89.675 ;
        RECT 88.385 88.525 88.715 89.505 ;
        RECT 88.885 88.535 89.115 89.675 ;
        RECT 89.325 89.240 94.670 89.675 ;
        RECT 86.680 87.125 86.965 87.585 ;
        RECT 87.145 87.305 87.400 87.835 ;
        RECT 88.005 87.125 88.215 87.945 ;
        RECT 88.385 87.925 88.635 88.525 ;
        RECT 88.805 88.115 89.135 88.365 ;
        RECT 88.385 87.295 88.715 87.925 ;
        RECT 88.885 87.125 89.115 87.945 ;
        RECT 90.910 87.670 91.250 88.500 ;
        RECT 92.730 87.990 93.080 89.240 ;
        RECT 95.765 88.510 96.055 89.675 ;
        RECT 96.225 88.585 99.735 89.675 ;
        RECT 100.370 89.165 102.025 89.455 ;
        RECT 96.225 87.895 97.875 88.415 ;
        RECT 98.045 88.065 99.735 88.585 ;
        RECT 100.370 88.825 101.960 88.995 ;
        RECT 102.195 88.875 102.475 89.675 ;
        RECT 100.370 88.535 100.690 88.825 ;
        RECT 101.790 88.705 101.960 88.825 ;
        RECT 89.325 87.125 94.670 87.670 ;
        RECT 95.765 87.125 96.055 87.850 ;
        RECT 96.225 87.125 99.735 87.895 ;
        RECT 100.370 87.795 100.720 88.365 ;
        RECT 100.890 88.035 101.600 88.655 ;
        RECT 101.790 88.535 102.515 88.705 ;
        RECT 102.685 88.535 102.955 89.505 ;
        RECT 103.130 89.165 104.785 89.455 ;
        RECT 103.130 88.825 104.720 88.995 ;
        RECT 104.955 88.875 105.235 89.675 ;
        RECT 103.130 88.535 103.450 88.825 ;
        RECT 104.550 88.705 104.720 88.825 ;
        RECT 102.345 88.365 102.515 88.535 ;
        RECT 101.770 88.035 102.175 88.365 ;
        RECT 102.345 88.035 102.615 88.365 ;
        RECT 102.345 87.865 102.515 88.035 ;
        RECT 100.905 87.695 102.515 87.865 ;
        RECT 102.785 87.800 102.955 88.535 ;
        RECT 103.645 88.485 104.360 88.655 ;
        RECT 104.550 88.535 105.275 88.705 ;
        RECT 105.445 88.535 105.715 89.505 ;
        RECT 105.885 89.240 111.230 89.675 ;
        RECT 100.375 87.125 100.705 87.625 ;
        RECT 100.905 87.345 101.075 87.695 ;
        RECT 101.275 87.125 101.605 87.525 ;
        RECT 101.775 87.345 101.945 87.695 ;
        RECT 102.115 87.125 102.495 87.525 ;
        RECT 102.685 87.455 102.955 87.800 ;
        RECT 103.130 87.795 103.480 88.365 ;
        RECT 103.650 88.035 104.360 88.485 ;
        RECT 105.105 88.365 105.275 88.535 ;
        RECT 104.530 88.035 104.935 88.365 ;
        RECT 105.105 88.035 105.375 88.365 ;
        RECT 105.105 87.865 105.275 88.035 ;
        RECT 103.665 87.695 105.275 87.865 ;
        RECT 105.545 87.800 105.715 88.535 ;
        RECT 103.135 87.125 103.465 87.625 ;
        RECT 103.665 87.345 103.835 87.695 ;
        RECT 104.035 87.125 104.365 87.525 ;
        RECT 104.535 87.345 104.705 87.695 ;
        RECT 104.875 87.125 105.255 87.525 ;
        RECT 105.445 87.455 105.715 87.800 ;
        RECT 107.470 87.670 107.810 88.500 ;
        RECT 109.290 87.990 109.640 89.240 ;
        RECT 111.405 88.585 112.615 89.675 ;
        RECT 111.405 87.875 111.925 88.415 ;
        RECT 112.095 88.045 112.615 88.585 ;
        RECT 112.875 88.745 113.045 89.505 ;
        RECT 113.225 88.915 113.555 89.675 ;
        RECT 112.875 88.575 113.540 88.745 ;
        RECT 113.725 88.600 113.995 89.505 ;
        RECT 113.370 88.430 113.540 88.575 ;
        RECT 112.805 88.025 113.135 88.395 ;
        RECT 113.370 88.100 113.655 88.430 ;
        RECT 105.885 87.125 111.230 87.670 ;
        RECT 111.405 87.125 112.615 87.875 ;
        RECT 113.370 87.845 113.540 88.100 ;
        RECT 112.875 87.675 113.540 87.845 ;
        RECT 113.825 87.800 113.995 88.600 ;
        RECT 114.225 88.535 114.435 89.675 ;
        RECT 114.605 88.525 114.935 89.505 ;
        RECT 115.105 88.535 115.335 89.675 ;
        RECT 115.545 89.240 120.890 89.675 ;
        RECT 112.875 87.295 113.045 87.675 ;
        RECT 113.225 87.125 113.555 87.505 ;
        RECT 113.735 87.295 113.995 87.800 ;
        RECT 114.225 87.125 114.435 87.945 ;
        RECT 114.605 87.925 114.855 88.525 ;
        RECT 115.025 88.115 115.355 88.365 ;
        RECT 114.605 87.295 114.935 87.925 ;
        RECT 115.105 87.125 115.335 87.945 ;
        RECT 117.130 87.670 117.470 88.500 ;
        RECT 118.950 87.990 119.300 89.240 ;
        RECT 121.525 88.510 121.815 89.675 ;
        RECT 122.445 88.585 123.655 89.675 ;
        RECT 122.445 88.045 122.965 88.585 ;
        RECT 123.135 87.875 123.655 88.415 ;
        RECT 115.545 87.125 120.890 87.670 ;
        RECT 121.525 87.125 121.815 87.850 ;
        RECT 122.445 87.125 123.655 87.875 ;
        RECT 5.520 86.955 123.740 87.125 ;
        RECT 5.605 86.205 6.815 86.955 ;
        RECT 7.995 86.405 8.165 86.695 ;
        RECT 8.335 86.575 8.665 86.955 ;
        RECT 7.995 86.235 8.660 86.405 ;
        RECT 5.605 85.665 6.125 86.205 ;
        RECT 6.295 85.495 6.815 86.035 ;
        RECT 5.605 84.405 6.815 85.495 ;
        RECT 7.910 85.415 8.260 86.065 ;
        RECT 8.430 85.245 8.660 86.235 ;
        RECT 7.995 85.075 8.660 85.245 ;
        RECT 7.995 84.575 8.165 85.075 ;
        RECT 8.335 84.405 8.665 84.905 ;
        RECT 8.835 84.575 9.060 86.695 ;
        RECT 9.275 86.575 9.605 86.955 ;
        RECT 9.775 86.405 9.945 86.735 ;
        RECT 10.245 86.575 11.260 86.775 ;
        RECT 9.250 86.215 9.945 86.405 ;
        RECT 9.250 85.245 9.420 86.215 ;
        RECT 9.590 85.415 10.000 86.035 ;
        RECT 10.170 85.465 10.390 86.335 ;
        RECT 10.570 86.025 10.920 86.395 ;
        RECT 11.090 85.845 11.260 86.575 ;
        RECT 11.430 86.515 11.840 86.955 ;
        RECT 12.130 86.315 12.380 86.745 ;
        RECT 12.580 86.495 12.900 86.955 ;
        RECT 13.460 86.565 14.310 86.735 ;
        RECT 11.430 85.975 11.840 86.305 ;
        RECT 12.130 85.975 12.550 86.315 ;
        RECT 10.840 85.805 11.260 85.845 ;
        RECT 10.840 85.635 12.190 85.805 ;
        RECT 9.250 85.075 9.945 85.245 ;
        RECT 10.170 85.085 10.670 85.465 ;
        RECT 9.275 84.405 9.605 84.905 ;
        RECT 9.775 84.575 9.945 85.075 ;
        RECT 10.840 84.790 11.010 85.635 ;
        RECT 11.940 85.475 12.190 85.635 ;
        RECT 11.180 85.205 11.430 85.465 ;
        RECT 12.360 85.205 12.550 85.975 ;
        RECT 11.180 84.955 12.550 85.205 ;
        RECT 12.720 86.145 13.970 86.315 ;
        RECT 12.720 85.385 12.890 86.145 ;
        RECT 13.640 86.025 13.970 86.145 ;
        RECT 13.060 85.565 13.240 85.975 ;
        RECT 14.140 85.805 14.310 86.565 ;
        RECT 14.510 86.475 15.170 86.955 ;
        RECT 15.350 86.360 15.670 86.690 ;
        RECT 14.500 86.035 15.160 86.305 ;
        RECT 14.500 85.975 14.830 86.035 ;
        RECT 14.980 85.805 15.310 85.865 ;
        RECT 13.410 85.635 15.310 85.805 ;
        RECT 12.720 85.075 13.240 85.385 ;
        RECT 13.410 85.125 13.580 85.635 ;
        RECT 15.480 85.465 15.670 86.360 ;
        RECT 13.750 85.295 15.670 85.465 ;
        RECT 15.350 85.275 15.670 85.295 ;
        RECT 15.870 86.045 16.120 86.695 ;
        RECT 16.300 86.495 16.585 86.955 ;
        RECT 16.765 86.245 17.020 86.775 ;
        RECT 15.870 85.715 16.670 86.045 ;
        RECT 13.410 84.955 14.620 85.125 ;
        RECT 10.180 84.620 11.010 84.790 ;
        RECT 11.250 84.405 11.630 84.785 ;
        RECT 11.810 84.665 11.980 84.955 ;
        RECT 13.410 84.875 13.580 84.955 ;
        RECT 12.150 84.405 12.480 84.785 ;
        RECT 12.950 84.625 13.580 84.875 ;
        RECT 13.760 84.405 14.180 84.785 ;
        RECT 14.380 84.665 14.620 84.955 ;
        RECT 14.850 84.405 15.180 85.095 ;
        RECT 15.350 84.665 15.520 85.275 ;
        RECT 15.870 85.125 16.120 85.715 ;
        RECT 16.840 85.595 17.020 86.245 ;
        RECT 17.570 86.215 17.825 86.785 ;
        RECT 17.995 86.555 18.325 86.955 ;
        RECT 18.750 86.420 19.280 86.785 ;
        RECT 18.750 86.385 18.925 86.420 ;
        RECT 17.995 86.215 18.925 86.385 ;
        RECT 16.840 85.425 17.105 85.595 ;
        RECT 17.570 85.545 17.740 86.215 ;
        RECT 17.995 86.045 18.165 86.215 ;
        RECT 17.910 85.715 18.165 86.045 ;
        RECT 18.390 85.715 18.585 86.045 ;
        RECT 16.840 85.385 17.020 85.425 ;
        RECT 15.790 84.615 16.120 85.125 ;
        RECT 16.300 84.405 16.585 85.205 ;
        RECT 16.765 84.715 17.020 85.385 ;
        RECT 17.570 84.575 17.905 85.545 ;
        RECT 18.075 84.405 18.245 85.545 ;
        RECT 18.415 84.745 18.585 85.715 ;
        RECT 18.755 85.085 18.925 86.215 ;
        RECT 19.095 85.425 19.265 86.225 ;
        RECT 19.470 85.935 19.745 86.785 ;
        RECT 19.465 85.765 19.745 85.935 ;
        RECT 19.470 85.625 19.745 85.765 ;
        RECT 19.915 85.425 20.105 86.785 ;
        RECT 20.285 86.420 20.795 86.955 ;
        RECT 21.015 86.145 21.260 86.750 ;
        RECT 21.705 86.185 24.295 86.955 ;
        RECT 20.305 85.975 21.535 86.145 ;
        RECT 19.095 85.255 20.105 85.425 ;
        RECT 20.275 85.410 21.025 85.600 ;
        RECT 18.755 84.915 19.880 85.085 ;
        RECT 20.275 84.745 20.445 85.410 ;
        RECT 21.195 85.165 21.535 85.975 ;
        RECT 21.705 85.665 22.915 86.185 ;
        RECT 24.670 86.175 25.170 86.785 ;
        RECT 23.085 85.495 24.295 86.015 ;
        RECT 24.465 85.715 24.815 85.965 ;
        RECT 25.000 85.545 25.170 86.175 ;
        RECT 25.800 86.305 26.130 86.785 ;
        RECT 26.300 86.495 26.525 86.955 ;
        RECT 26.695 86.305 27.025 86.785 ;
        RECT 25.800 86.135 27.025 86.305 ;
        RECT 27.215 86.155 27.465 86.955 ;
        RECT 27.635 86.155 27.975 86.785 ;
        RECT 28.155 86.455 28.485 86.955 ;
        RECT 28.685 86.385 28.855 86.735 ;
        RECT 29.055 86.555 29.385 86.955 ;
        RECT 29.555 86.385 29.725 86.735 ;
        RECT 29.895 86.555 30.275 86.955 ;
        RECT 27.745 86.105 27.975 86.155 ;
        RECT 25.340 85.765 25.670 85.965 ;
        RECT 25.840 85.765 26.170 85.965 ;
        RECT 26.340 85.765 26.760 85.965 ;
        RECT 26.935 85.795 27.630 85.965 ;
        RECT 26.935 85.545 27.105 85.795 ;
        RECT 27.800 85.545 27.975 86.105 ;
        RECT 28.150 85.715 28.500 86.285 ;
        RECT 28.685 86.215 30.295 86.385 ;
        RECT 30.465 86.280 30.735 86.625 ;
        RECT 30.125 86.045 30.295 86.215 ;
        RECT 28.670 85.595 29.380 86.045 ;
        RECT 29.550 85.715 29.955 86.045 ;
        RECT 30.125 85.715 30.395 86.045 ;
        RECT 18.415 84.575 20.445 84.745 ;
        RECT 20.615 84.405 20.785 85.165 ;
        RECT 21.020 84.755 21.535 85.165 ;
        RECT 21.705 84.405 24.295 85.495 ;
        RECT 24.670 85.375 27.105 85.545 ;
        RECT 24.670 84.575 25.000 85.375 ;
        RECT 25.170 84.405 25.500 85.205 ;
        RECT 25.800 84.575 26.130 85.375 ;
        RECT 26.775 84.405 27.025 85.205 ;
        RECT 27.295 84.405 27.465 85.545 ;
        RECT 27.635 84.575 27.975 85.545 ;
        RECT 28.150 85.255 28.470 85.545 ;
        RECT 28.665 85.425 29.380 85.595 ;
        RECT 30.125 85.545 30.295 85.715 ;
        RECT 30.565 85.545 30.735 86.280 ;
        RECT 31.365 86.230 31.655 86.955 ;
        RECT 32.030 86.175 32.530 86.785 ;
        RECT 31.825 85.715 32.175 85.965 ;
        RECT 29.570 85.375 30.295 85.545 ;
        RECT 29.570 85.255 29.740 85.375 ;
        RECT 28.150 85.085 29.740 85.255 ;
        RECT 28.150 84.625 29.805 84.915 ;
        RECT 29.975 84.405 30.255 85.205 ;
        RECT 30.465 84.575 30.735 85.545 ;
        RECT 31.365 84.405 31.655 85.570 ;
        RECT 32.360 85.545 32.530 86.175 ;
        RECT 33.160 86.305 33.490 86.785 ;
        RECT 33.660 86.495 33.885 86.955 ;
        RECT 34.055 86.305 34.385 86.785 ;
        RECT 33.160 86.135 34.385 86.305 ;
        RECT 34.575 86.155 34.825 86.955 ;
        RECT 34.995 86.155 35.335 86.785 ;
        RECT 35.505 86.410 40.850 86.955 ;
        RECT 41.025 86.410 46.370 86.955 ;
        RECT 46.545 86.410 51.890 86.955 ;
        RECT 32.700 85.765 33.030 85.965 ;
        RECT 33.200 85.765 33.530 85.965 ;
        RECT 33.700 85.765 34.120 85.965 ;
        RECT 34.295 85.795 34.990 85.965 ;
        RECT 34.295 85.545 34.465 85.795 ;
        RECT 35.160 85.545 35.335 86.155 ;
        RECT 37.090 85.580 37.430 86.410 ;
        RECT 32.030 85.375 34.465 85.545 ;
        RECT 32.030 84.575 32.360 85.375 ;
        RECT 32.530 84.405 32.860 85.205 ;
        RECT 33.160 84.575 33.490 85.375 ;
        RECT 34.135 84.405 34.385 85.205 ;
        RECT 34.655 84.405 34.825 85.545 ;
        RECT 34.995 84.575 35.335 85.545 ;
        RECT 38.910 84.840 39.260 86.090 ;
        RECT 42.610 85.580 42.950 86.410 ;
        RECT 44.430 84.840 44.780 86.090 ;
        RECT 48.130 85.580 48.470 86.410 ;
        RECT 52.065 86.185 55.575 86.955 ;
        RECT 55.745 86.205 56.955 86.955 ;
        RECT 57.125 86.230 57.415 86.955 ;
        RECT 57.675 86.405 57.845 86.695 ;
        RECT 58.015 86.575 58.345 86.955 ;
        RECT 57.675 86.235 58.340 86.405 ;
        RECT 49.950 84.840 50.300 86.090 ;
        RECT 52.065 85.665 53.715 86.185 ;
        RECT 53.885 85.495 55.575 86.015 ;
        RECT 55.745 85.665 56.265 86.205 ;
        RECT 56.435 85.495 56.955 86.035 ;
        RECT 35.505 84.405 40.850 84.840 ;
        RECT 41.025 84.405 46.370 84.840 ;
        RECT 46.545 84.405 51.890 84.840 ;
        RECT 52.065 84.405 55.575 85.495 ;
        RECT 55.745 84.405 56.955 85.495 ;
        RECT 57.125 84.405 57.415 85.570 ;
        RECT 57.590 85.415 57.940 86.065 ;
        RECT 58.110 85.245 58.340 86.235 ;
        RECT 57.675 85.075 58.340 85.245 ;
        RECT 57.675 84.575 57.845 85.075 ;
        RECT 58.015 84.405 58.345 84.905 ;
        RECT 58.515 84.575 58.740 86.695 ;
        RECT 58.955 86.575 59.285 86.955 ;
        RECT 59.455 86.405 59.625 86.735 ;
        RECT 59.925 86.575 60.940 86.775 ;
        RECT 58.930 86.215 59.625 86.405 ;
        RECT 58.930 85.245 59.100 86.215 ;
        RECT 59.270 85.415 59.680 86.035 ;
        RECT 59.850 85.465 60.070 86.335 ;
        RECT 60.250 86.025 60.600 86.395 ;
        RECT 60.770 85.845 60.940 86.575 ;
        RECT 61.110 86.515 61.520 86.955 ;
        RECT 61.810 86.315 62.060 86.745 ;
        RECT 62.260 86.495 62.580 86.955 ;
        RECT 63.140 86.565 63.990 86.735 ;
        RECT 61.110 85.975 61.520 86.305 ;
        RECT 61.810 85.975 62.230 86.315 ;
        RECT 60.520 85.805 60.940 85.845 ;
        RECT 60.520 85.635 61.870 85.805 ;
        RECT 58.930 85.075 59.625 85.245 ;
        RECT 59.850 85.085 60.350 85.465 ;
        RECT 58.955 84.405 59.285 84.905 ;
        RECT 59.455 84.575 59.625 85.075 ;
        RECT 60.520 84.790 60.690 85.635 ;
        RECT 61.620 85.475 61.870 85.635 ;
        RECT 60.860 85.205 61.110 85.465 ;
        RECT 62.040 85.205 62.230 85.975 ;
        RECT 60.860 84.955 62.230 85.205 ;
        RECT 62.400 86.145 63.650 86.315 ;
        RECT 62.400 85.385 62.570 86.145 ;
        RECT 63.320 86.025 63.650 86.145 ;
        RECT 62.740 85.565 62.920 85.975 ;
        RECT 63.820 85.805 63.990 86.565 ;
        RECT 64.190 86.475 64.850 86.955 ;
        RECT 65.030 86.360 65.350 86.690 ;
        RECT 64.180 86.035 64.840 86.305 ;
        RECT 64.180 85.975 64.510 86.035 ;
        RECT 64.660 85.805 64.990 85.865 ;
        RECT 63.090 85.635 64.990 85.805 ;
        RECT 62.400 85.075 62.920 85.385 ;
        RECT 63.090 85.125 63.260 85.635 ;
        RECT 65.160 85.465 65.350 86.360 ;
        RECT 63.430 85.295 65.350 85.465 ;
        RECT 65.030 85.275 65.350 85.295 ;
        RECT 65.550 86.045 65.800 86.695 ;
        RECT 65.980 86.495 66.265 86.955 ;
        RECT 66.445 86.245 66.700 86.775 ;
        RECT 65.550 85.715 66.350 86.045 ;
        RECT 63.090 84.955 64.300 85.125 ;
        RECT 59.860 84.620 60.690 84.790 ;
        RECT 60.930 84.405 61.310 84.785 ;
        RECT 61.490 84.665 61.660 84.955 ;
        RECT 63.090 84.875 63.260 84.955 ;
        RECT 61.830 84.405 62.160 84.785 ;
        RECT 62.630 84.625 63.260 84.875 ;
        RECT 63.440 84.405 63.860 84.785 ;
        RECT 64.060 84.665 64.300 84.955 ;
        RECT 64.530 84.405 64.860 85.095 ;
        RECT 65.030 84.665 65.200 85.275 ;
        RECT 65.550 85.125 65.800 85.715 ;
        RECT 66.520 85.385 66.700 86.245 ;
        RECT 67.910 86.175 68.410 86.785 ;
        RECT 67.705 85.715 68.055 85.965 ;
        RECT 68.240 85.545 68.410 86.175 ;
        RECT 69.040 86.305 69.370 86.785 ;
        RECT 69.540 86.495 69.765 86.955 ;
        RECT 69.935 86.305 70.265 86.785 ;
        RECT 69.040 86.135 70.265 86.305 ;
        RECT 70.455 86.155 70.705 86.955 ;
        RECT 70.875 86.155 71.215 86.785 ;
        RECT 71.385 86.410 76.730 86.955 ;
        RECT 76.905 86.410 82.250 86.955 ;
        RECT 68.580 85.765 68.910 85.965 ;
        RECT 69.080 85.765 69.410 85.965 ;
        RECT 69.580 85.765 70.000 85.965 ;
        RECT 70.175 85.795 70.870 85.965 ;
        RECT 70.175 85.545 70.345 85.795 ;
        RECT 71.040 85.545 71.215 86.155 ;
        RECT 72.970 85.580 73.310 86.410 ;
        RECT 65.470 84.615 65.800 85.125 ;
        RECT 65.980 84.405 66.265 85.205 ;
        RECT 66.445 84.915 66.700 85.385 ;
        RECT 67.910 85.375 70.345 85.545 ;
        RECT 66.445 84.745 66.785 84.915 ;
        RECT 66.445 84.715 66.700 84.745 ;
        RECT 67.910 84.575 68.240 85.375 ;
        RECT 68.410 84.405 68.740 85.205 ;
        RECT 69.040 84.575 69.370 85.375 ;
        RECT 70.015 84.405 70.265 85.205 ;
        RECT 70.535 84.405 70.705 85.545 ;
        RECT 70.875 84.575 71.215 85.545 ;
        RECT 74.790 84.840 75.140 86.090 ;
        RECT 78.490 85.580 78.830 86.410 ;
        RECT 82.885 86.230 83.175 86.955 ;
        RECT 83.435 86.405 83.605 86.785 ;
        RECT 83.785 86.575 84.115 86.955 ;
        RECT 83.435 86.235 84.100 86.405 ;
        RECT 84.295 86.280 84.555 86.785 ;
        RECT 80.310 84.840 80.660 86.090 ;
        RECT 83.365 85.685 83.695 86.055 ;
        RECT 83.930 85.980 84.100 86.235 ;
        RECT 83.930 85.650 84.215 85.980 ;
        RECT 71.385 84.405 76.730 84.840 ;
        RECT 76.905 84.405 82.250 84.840 ;
        RECT 82.885 84.405 83.175 85.570 ;
        RECT 83.930 85.505 84.100 85.650 ;
        RECT 83.435 85.335 84.100 85.505 ;
        RECT 84.385 85.480 84.555 86.280 ;
        RECT 84.815 86.405 84.985 86.695 ;
        RECT 85.155 86.575 85.485 86.955 ;
        RECT 84.815 86.235 85.480 86.405 ;
        RECT 83.435 84.575 83.605 85.335 ;
        RECT 83.785 84.405 84.115 85.165 ;
        RECT 84.285 84.575 84.555 85.480 ;
        RECT 84.730 85.415 85.080 86.065 ;
        RECT 85.250 85.245 85.480 86.235 ;
        RECT 84.815 85.075 85.480 85.245 ;
        RECT 84.815 84.575 84.985 85.075 ;
        RECT 85.155 84.405 85.485 84.905 ;
        RECT 85.655 84.575 85.880 86.695 ;
        RECT 86.095 86.575 86.425 86.955 ;
        RECT 86.595 86.405 86.765 86.735 ;
        RECT 87.065 86.575 88.080 86.775 ;
        RECT 86.070 86.215 86.765 86.405 ;
        RECT 86.070 85.245 86.240 86.215 ;
        RECT 86.410 85.415 86.820 86.035 ;
        RECT 86.990 85.465 87.210 86.335 ;
        RECT 87.390 86.025 87.740 86.395 ;
        RECT 87.910 85.845 88.080 86.575 ;
        RECT 88.250 86.515 88.660 86.955 ;
        RECT 88.950 86.315 89.200 86.745 ;
        RECT 89.400 86.495 89.720 86.955 ;
        RECT 90.280 86.565 91.130 86.735 ;
        RECT 88.250 85.975 88.660 86.305 ;
        RECT 88.950 85.975 89.370 86.315 ;
        RECT 87.660 85.805 88.080 85.845 ;
        RECT 87.660 85.635 89.010 85.805 ;
        RECT 86.070 85.075 86.765 85.245 ;
        RECT 86.990 85.085 87.490 85.465 ;
        RECT 86.095 84.405 86.425 84.905 ;
        RECT 86.595 84.575 86.765 85.075 ;
        RECT 87.660 84.790 87.830 85.635 ;
        RECT 88.760 85.475 89.010 85.635 ;
        RECT 88.000 85.205 88.250 85.465 ;
        RECT 89.180 85.205 89.370 85.975 ;
        RECT 88.000 84.955 89.370 85.205 ;
        RECT 89.540 86.145 90.790 86.315 ;
        RECT 89.540 85.385 89.710 86.145 ;
        RECT 90.460 86.025 90.790 86.145 ;
        RECT 89.880 85.565 90.060 85.975 ;
        RECT 90.960 85.805 91.130 86.565 ;
        RECT 91.330 86.475 91.990 86.955 ;
        RECT 92.170 86.360 92.490 86.690 ;
        RECT 91.320 86.035 91.980 86.305 ;
        RECT 91.320 85.975 91.650 86.035 ;
        RECT 91.800 85.805 92.130 85.865 ;
        RECT 90.230 85.635 92.130 85.805 ;
        RECT 89.540 85.075 90.060 85.385 ;
        RECT 90.230 85.125 90.400 85.635 ;
        RECT 92.300 85.465 92.490 86.360 ;
        RECT 90.570 85.295 92.490 85.465 ;
        RECT 92.170 85.275 92.490 85.295 ;
        RECT 92.690 86.045 92.940 86.695 ;
        RECT 93.120 86.495 93.405 86.955 ;
        RECT 93.585 86.245 93.840 86.775 ;
        RECT 92.690 85.715 93.490 86.045 ;
        RECT 90.230 84.955 91.440 85.125 ;
        RECT 87.000 84.620 87.830 84.790 ;
        RECT 88.070 84.405 88.450 84.785 ;
        RECT 88.630 84.665 88.800 84.955 ;
        RECT 90.230 84.875 90.400 84.955 ;
        RECT 88.970 84.405 89.300 84.785 ;
        RECT 89.770 84.625 90.400 84.875 ;
        RECT 90.580 84.405 91.000 84.785 ;
        RECT 91.200 84.665 91.440 84.955 ;
        RECT 91.670 84.405 92.000 85.095 ;
        RECT 92.170 84.665 92.340 85.275 ;
        RECT 92.690 85.125 92.940 85.715 ;
        RECT 93.660 85.385 93.840 86.245 ;
        RECT 94.445 86.135 94.655 86.955 ;
        RECT 94.825 86.155 95.155 86.785 ;
        RECT 94.825 85.555 95.075 86.155 ;
        RECT 95.325 86.135 95.555 86.955 ;
        RECT 95.765 86.185 99.275 86.955 ;
        RECT 99.915 86.455 100.245 86.955 ;
        RECT 100.445 86.385 100.615 86.735 ;
        RECT 100.815 86.555 101.145 86.955 ;
        RECT 101.315 86.385 101.485 86.735 ;
        RECT 101.655 86.555 102.035 86.955 ;
        RECT 95.245 85.715 95.575 85.965 ;
        RECT 95.765 85.665 97.415 86.185 ;
        RECT 92.610 84.615 92.940 85.125 ;
        RECT 93.120 84.405 93.405 85.205 ;
        RECT 93.585 84.915 93.840 85.385 ;
        RECT 93.585 84.745 93.925 84.915 ;
        RECT 93.585 84.715 93.840 84.745 ;
        RECT 94.445 84.405 94.655 85.545 ;
        RECT 94.825 84.575 95.155 85.555 ;
        RECT 95.325 84.405 95.555 85.545 ;
        RECT 97.585 85.495 99.275 86.015 ;
        RECT 99.910 85.715 100.260 86.285 ;
        RECT 100.445 86.215 102.055 86.385 ;
        RECT 102.225 86.280 102.495 86.625 ;
        RECT 102.675 86.455 103.005 86.955 ;
        RECT 103.205 86.385 103.375 86.735 ;
        RECT 103.575 86.555 103.905 86.955 ;
        RECT 104.075 86.385 104.245 86.735 ;
        RECT 104.415 86.555 104.795 86.955 ;
        RECT 101.885 86.045 102.055 86.215 ;
        RECT 100.430 85.595 101.140 86.045 ;
        RECT 101.310 85.715 101.715 86.045 ;
        RECT 101.885 85.715 102.155 86.045 ;
        RECT 95.765 84.405 99.275 85.495 ;
        RECT 99.910 85.255 100.230 85.545 ;
        RECT 100.425 85.425 101.140 85.595 ;
        RECT 101.885 85.545 102.055 85.715 ;
        RECT 102.325 85.545 102.495 86.280 ;
        RECT 102.670 85.715 103.020 86.285 ;
        RECT 103.205 86.215 104.815 86.385 ;
        RECT 104.985 86.280 105.255 86.625 ;
        RECT 104.645 86.045 104.815 86.215 ;
        RECT 101.330 85.375 102.055 85.545 ;
        RECT 101.330 85.255 101.500 85.375 ;
        RECT 99.910 85.085 101.500 85.255 ;
        RECT 99.910 84.625 101.565 84.915 ;
        RECT 101.735 84.405 102.015 85.205 ;
        RECT 102.225 84.575 102.495 85.545 ;
        RECT 102.670 85.255 102.990 85.545 ;
        RECT 103.190 85.425 103.900 86.045 ;
        RECT 104.070 85.715 104.475 86.045 ;
        RECT 104.645 85.715 104.915 86.045 ;
        RECT 104.645 85.545 104.815 85.715 ;
        RECT 105.085 85.545 105.255 86.280 ;
        RECT 105.425 86.185 108.015 86.955 ;
        RECT 108.645 86.230 108.935 86.955 ;
        RECT 109.195 86.405 109.365 86.695 ;
        RECT 109.535 86.575 109.865 86.955 ;
        RECT 109.195 86.235 109.860 86.405 ;
        RECT 105.425 85.665 106.635 86.185 ;
        RECT 104.090 85.375 104.815 85.545 ;
        RECT 104.090 85.255 104.260 85.375 ;
        RECT 102.670 85.085 104.260 85.255 ;
        RECT 102.670 84.625 104.325 84.915 ;
        RECT 104.495 84.405 104.775 85.205 ;
        RECT 104.985 84.575 105.255 85.545 ;
        RECT 106.805 85.495 108.015 86.015 ;
        RECT 105.425 84.405 108.015 85.495 ;
        RECT 108.645 84.405 108.935 85.570 ;
        RECT 109.110 85.415 109.460 86.065 ;
        RECT 109.630 85.245 109.860 86.235 ;
        RECT 109.195 85.075 109.860 85.245 ;
        RECT 109.195 84.575 109.365 85.075 ;
        RECT 109.535 84.405 109.865 84.905 ;
        RECT 110.035 84.575 110.260 86.695 ;
        RECT 110.475 86.575 110.805 86.955 ;
        RECT 110.975 86.405 111.145 86.735 ;
        RECT 111.445 86.575 112.460 86.775 ;
        RECT 110.450 86.215 111.145 86.405 ;
        RECT 110.450 85.245 110.620 86.215 ;
        RECT 110.790 85.415 111.200 86.035 ;
        RECT 111.370 85.465 111.590 86.335 ;
        RECT 111.770 86.025 112.120 86.395 ;
        RECT 112.290 85.845 112.460 86.575 ;
        RECT 112.630 86.515 113.040 86.955 ;
        RECT 113.330 86.315 113.580 86.745 ;
        RECT 113.780 86.495 114.100 86.955 ;
        RECT 114.660 86.565 115.510 86.735 ;
        RECT 112.630 85.975 113.040 86.305 ;
        RECT 113.330 85.975 113.750 86.315 ;
        RECT 112.040 85.805 112.460 85.845 ;
        RECT 112.040 85.635 113.390 85.805 ;
        RECT 110.450 85.075 111.145 85.245 ;
        RECT 111.370 85.085 111.870 85.465 ;
        RECT 110.475 84.405 110.805 84.905 ;
        RECT 110.975 84.575 111.145 85.075 ;
        RECT 112.040 84.790 112.210 85.635 ;
        RECT 113.140 85.475 113.390 85.635 ;
        RECT 112.380 85.205 112.630 85.465 ;
        RECT 113.560 85.205 113.750 85.975 ;
        RECT 112.380 84.955 113.750 85.205 ;
        RECT 113.920 86.145 115.170 86.315 ;
        RECT 113.920 85.385 114.090 86.145 ;
        RECT 114.840 86.025 115.170 86.145 ;
        RECT 114.260 85.565 114.440 85.975 ;
        RECT 115.340 85.805 115.510 86.565 ;
        RECT 115.710 86.475 116.370 86.955 ;
        RECT 116.550 86.360 116.870 86.690 ;
        RECT 115.700 86.035 116.360 86.305 ;
        RECT 115.700 85.975 116.030 86.035 ;
        RECT 116.180 85.805 116.510 85.865 ;
        RECT 114.610 85.635 116.510 85.805 ;
        RECT 113.920 85.075 114.440 85.385 ;
        RECT 114.610 85.125 114.780 85.635 ;
        RECT 116.680 85.465 116.870 86.360 ;
        RECT 114.950 85.295 116.870 85.465 ;
        RECT 116.550 85.275 116.870 85.295 ;
        RECT 117.070 86.045 117.320 86.695 ;
        RECT 117.500 86.495 117.785 86.955 ;
        RECT 117.965 86.245 118.220 86.775 ;
        RECT 117.070 85.715 117.870 86.045 ;
        RECT 114.610 84.955 115.820 85.125 ;
        RECT 111.380 84.620 112.210 84.790 ;
        RECT 112.450 84.405 112.830 84.785 ;
        RECT 113.010 84.665 113.180 84.955 ;
        RECT 114.610 84.875 114.780 84.955 ;
        RECT 113.350 84.405 113.680 84.785 ;
        RECT 114.150 84.625 114.780 84.875 ;
        RECT 114.960 84.405 115.380 84.785 ;
        RECT 115.580 84.665 115.820 84.955 ;
        RECT 116.050 84.405 116.380 85.095 ;
        RECT 116.550 84.665 116.720 85.275 ;
        RECT 117.070 85.125 117.320 85.715 ;
        RECT 118.040 85.385 118.220 86.245 ;
        RECT 118.805 86.135 119.035 86.955 ;
        RECT 119.205 86.155 119.535 86.785 ;
        RECT 118.785 85.715 119.115 85.965 ;
        RECT 119.285 85.555 119.535 86.155 ;
        RECT 119.705 86.135 119.915 86.955 ;
        RECT 120.145 86.185 121.815 86.955 ;
        RECT 122.445 86.205 123.655 86.955 ;
        RECT 120.145 85.665 120.895 86.185 ;
        RECT 116.990 84.615 117.320 85.125 ;
        RECT 117.500 84.405 117.785 85.205 ;
        RECT 117.965 84.915 118.220 85.385 ;
        RECT 117.965 84.745 118.305 84.915 ;
        RECT 117.965 84.715 118.220 84.745 ;
        RECT 118.805 84.405 119.035 85.545 ;
        RECT 119.205 84.575 119.535 85.555 ;
        RECT 119.705 84.405 119.915 85.545 ;
        RECT 121.065 85.495 121.815 86.015 ;
        RECT 120.145 84.405 121.815 85.495 ;
        RECT 122.445 85.495 122.965 86.035 ;
        RECT 123.135 85.665 123.655 86.205 ;
        RECT 122.445 84.405 123.655 85.495 ;
        RECT 5.520 84.235 123.740 84.405 ;
        RECT 5.605 83.145 6.815 84.235 ;
        RECT 6.985 83.145 10.495 84.235 ;
        RECT 5.605 82.435 6.125 82.975 ;
        RECT 6.295 82.605 6.815 83.145 ;
        RECT 6.985 82.455 8.635 82.975 ;
        RECT 8.805 82.625 10.495 83.145 ;
        RECT 10.665 83.160 10.935 84.065 ;
        RECT 11.105 83.475 11.435 84.235 ;
        RECT 11.615 83.305 11.785 84.065 ;
        RECT 5.605 81.685 6.815 82.435 ;
        RECT 6.985 81.685 10.495 82.455 ;
        RECT 10.665 82.360 10.835 83.160 ;
        RECT 11.120 83.135 11.785 83.305 ;
        RECT 11.120 82.990 11.290 83.135 ;
        RECT 13.025 83.095 13.235 84.235 ;
        RECT 11.005 82.660 11.290 82.990 ;
        RECT 13.405 83.085 13.735 84.065 ;
        RECT 13.905 83.095 14.135 84.235 ;
        RECT 14.405 83.095 14.615 84.235 ;
        RECT 14.785 83.085 15.115 84.065 ;
        RECT 15.285 83.095 15.515 84.235 ;
        RECT 15.725 83.145 18.315 84.235 ;
        RECT 11.120 82.405 11.290 82.660 ;
        RECT 11.525 82.585 11.855 82.955 ;
        RECT 10.665 81.855 10.925 82.360 ;
        RECT 11.120 82.235 11.785 82.405 ;
        RECT 11.105 81.685 11.435 82.065 ;
        RECT 11.615 81.855 11.785 82.235 ;
        RECT 13.025 81.685 13.235 82.505 ;
        RECT 13.405 82.485 13.655 83.085 ;
        RECT 13.825 82.675 14.155 82.925 ;
        RECT 13.405 81.855 13.735 82.485 ;
        RECT 13.905 81.685 14.135 82.505 ;
        RECT 14.405 81.685 14.615 82.505 ;
        RECT 14.785 82.485 15.035 83.085 ;
        RECT 15.205 82.675 15.535 82.925 ;
        RECT 14.785 81.855 15.115 82.485 ;
        RECT 15.285 81.685 15.515 82.505 ;
        RECT 15.725 82.455 16.935 82.975 ;
        RECT 17.105 82.625 18.315 83.145 ;
        RECT 18.485 83.070 18.775 84.235 ;
        RECT 18.945 83.145 21.535 84.235 ;
        RECT 18.945 82.455 20.155 82.975 ;
        RECT 20.325 82.625 21.535 83.145 ;
        RECT 22.370 83.265 22.700 84.065 ;
        RECT 22.870 83.435 23.200 84.235 ;
        RECT 23.500 83.265 23.830 84.065 ;
        RECT 24.475 83.435 24.725 84.235 ;
        RECT 22.370 83.095 24.805 83.265 ;
        RECT 24.995 83.095 25.165 84.235 ;
        RECT 25.335 83.095 25.675 84.065 ;
        RECT 25.845 83.800 31.190 84.235 ;
        RECT 31.365 83.800 36.710 84.235 ;
        RECT 22.165 82.675 22.515 82.925 ;
        RECT 22.700 82.465 22.870 83.095 ;
        RECT 23.040 82.675 23.370 82.875 ;
        RECT 23.540 82.675 23.870 82.875 ;
        RECT 24.040 82.675 24.460 82.875 ;
        RECT 24.635 82.845 24.805 83.095 ;
        RECT 24.635 82.675 25.330 82.845 ;
        RECT 15.725 81.685 18.315 82.455 ;
        RECT 18.485 81.685 18.775 82.410 ;
        RECT 18.945 81.685 21.535 82.455 ;
        RECT 22.370 81.855 22.870 82.465 ;
        RECT 23.500 82.335 24.725 82.505 ;
        RECT 25.500 82.485 25.675 83.095 ;
        RECT 23.500 81.855 23.830 82.335 ;
        RECT 24.000 81.685 24.225 82.145 ;
        RECT 24.395 81.855 24.725 82.335 ;
        RECT 24.915 81.685 25.165 82.485 ;
        RECT 25.335 81.855 25.675 82.485 ;
        RECT 27.430 82.230 27.770 83.060 ;
        RECT 29.250 82.550 29.600 83.800 ;
        RECT 32.950 82.230 33.290 83.060 ;
        RECT 34.770 82.550 35.120 83.800 ;
        RECT 36.885 83.145 39.475 84.235 ;
        RECT 36.885 82.455 38.095 82.975 ;
        RECT 38.265 82.625 39.475 83.145 ;
        RECT 40.110 83.095 40.445 84.065 ;
        RECT 40.615 83.095 40.785 84.235 ;
        RECT 40.955 83.895 42.985 84.065 ;
        RECT 25.845 81.685 31.190 82.230 ;
        RECT 31.365 81.685 36.710 82.230 ;
        RECT 36.885 81.685 39.475 82.455 ;
        RECT 40.110 82.425 40.280 83.095 ;
        RECT 40.955 82.925 41.125 83.895 ;
        RECT 40.450 82.595 40.705 82.925 ;
        RECT 40.930 82.595 41.125 82.925 ;
        RECT 41.295 83.555 42.420 83.725 ;
        RECT 40.535 82.425 40.705 82.595 ;
        RECT 41.295 82.425 41.465 83.555 ;
        RECT 40.110 81.855 40.365 82.425 ;
        RECT 40.535 82.255 41.465 82.425 ;
        RECT 41.635 83.215 42.645 83.385 ;
        RECT 41.635 82.415 41.805 83.215 ;
        RECT 42.010 82.535 42.285 83.015 ;
        RECT 42.005 82.365 42.285 82.535 ;
        RECT 41.290 82.220 41.465 82.255 ;
        RECT 40.535 81.685 40.865 82.085 ;
        RECT 41.290 81.855 41.820 82.220 ;
        RECT 42.010 81.855 42.285 82.365 ;
        RECT 42.455 81.855 42.645 83.215 ;
        RECT 42.815 83.230 42.985 83.895 ;
        RECT 43.155 83.475 43.325 84.235 ;
        RECT 43.560 83.475 44.075 83.885 ;
        RECT 42.815 83.040 43.565 83.230 ;
        RECT 43.735 82.665 44.075 83.475 ;
        RECT 44.245 83.070 44.535 84.235 ;
        RECT 44.710 83.095 45.045 84.065 ;
        RECT 45.215 83.095 45.385 84.235 ;
        RECT 45.555 83.895 47.585 84.065 ;
        RECT 42.845 82.495 44.075 82.665 ;
        RECT 42.825 81.685 43.335 82.220 ;
        RECT 43.555 81.890 43.800 82.495 ;
        RECT 44.710 82.425 44.880 83.095 ;
        RECT 45.555 82.925 45.725 83.895 ;
        RECT 45.050 82.595 45.305 82.925 ;
        RECT 45.530 82.595 45.725 82.925 ;
        RECT 45.895 83.555 47.020 83.725 ;
        RECT 45.135 82.425 45.305 82.595 ;
        RECT 45.895 82.425 46.065 83.555 ;
        RECT 44.245 81.685 44.535 82.410 ;
        RECT 44.710 81.855 44.965 82.425 ;
        RECT 45.135 82.255 46.065 82.425 ;
        RECT 46.235 83.215 47.245 83.385 ;
        RECT 46.235 82.415 46.405 83.215 ;
        RECT 46.610 82.875 46.885 83.015 ;
        RECT 46.605 82.705 46.885 82.875 ;
        RECT 45.890 82.220 46.065 82.255 ;
        RECT 45.135 81.685 45.465 82.085 ;
        RECT 45.890 81.855 46.420 82.220 ;
        RECT 46.610 81.855 46.885 82.705 ;
        RECT 47.055 81.855 47.245 83.215 ;
        RECT 47.415 83.230 47.585 83.895 ;
        RECT 47.755 83.475 47.925 84.235 ;
        RECT 48.160 83.475 48.675 83.885 ;
        RECT 47.415 83.040 48.165 83.230 ;
        RECT 48.335 82.665 48.675 83.475 ;
        RECT 48.845 83.145 50.515 84.235 ;
        RECT 47.445 82.495 48.675 82.665 ;
        RECT 47.425 81.685 47.935 82.220 ;
        RECT 48.155 81.890 48.400 82.495 ;
        RECT 48.845 82.455 49.595 82.975 ;
        RECT 49.765 82.625 50.515 83.145 ;
        RECT 51.350 83.265 51.680 84.065 ;
        RECT 51.850 83.435 52.180 84.235 ;
        RECT 52.480 83.265 52.810 84.065 ;
        RECT 53.455 83.435 53.705 84.235 ;
        RECT 51.350 83.095 53.785 83.265 ;
        RECT 53.975 83.095 54.145 84.235 ;
        RECT 54.315 83.095 54.655 84.065 ;
        RECT 51.145 82.675 51.495 82.925 ;
        RECT 51.680 82.465 51.850 83.095 ;
        RECT 52.020 82.675 52.350 82.875 ;
        RECT 52.520 82.675 52.850 82.875 ;
        RECT 53.020 82.675 53.440 82.875 ;
        RECT 53.615 82.845 53.785 83.095 ;
        RECT 53.615 82.675 54.310 82.845 ;
        RECT 54.480 82.535 54.655 83.095 ;
        RECT 48.845 81.685 50.515 82.455 ;
        RECT 51.350 81.855 51.850 82.465 ;
        RECT 52.480 82.335 53.705 82.505 ;
        RECT 54.425 82.485 54.655 82.535 ;
        RECT 52.480 81.855 52.810 82.335 ;
        RECT 52.980 81.685 53.205 82.145 ;
        RECT 53.375 81.855 53.705 82.335 ;
        RECT 53.895 81.685 54.145 82.485 ;
        RECT 54.315 81.855 54.655 82.485 ;
        RECT 54.825 83.095 55.095 84.065 ;
        RECT 55.305 83.435 55.585 84.235 ;
        RECT 55.755 83.725 57.410 84.015 ;
        RECT 55.820 83.385 57.410 83.555 ;
        RECT 55.820 83.265 55.990 83.385 ;
        RECT 55.265 83.095 55.990 83.265 ;
        RECT 54.825 82.360 54.995 83.095 ;
        RECT 55.265 82.925 55.435 83.095 ;
        RECT 56.180 83.045 56.895 83.215 ;
        RECT 57.090 83.095 57.410 83.385 ;
        RECT 57.585 83.145 60.175 84.235 ;
        RECT 55.165 82.595 55.435 82.925 ;
        RECT 55.605 82.595 56.010 82.925 ;
        RECT 56.180 82.595 56.890 83.045 ;
        RECT 55.265 82.425 55.435 82.595 ;
        RECT 54.825 82.015 55.095 82.360 ;
        RECT 55.265 82.255 56.875 82.425 ;
        RECT 57.060 82.355 57.410 82.925 ;
        RECT 57.585 82.455 58.795 82.975 ;
        RECT 58.965 82.625 60.175 83.145 ;
        RECT 60.385 83.095 60.615 84.235 ;
        RECT 60.785 83.085 61.115 84.065 ;
        RECT 61.285 83.095 61.495 84.235 ;
        RECT 62.190 83.095 62.525 84.065 ;
        RECT 62.695 83.095 62.865 84.235 ;
        RECT 63.035 83.895 65.065 84.065 ;
        RECT 60.365 82.675 60.695 82.925 ;
        RECT 55.285 81.685 55.665 82.085 ;
        RECT 55.835 81.905 56.005 82.255 ;
        RECT 56.175 81.685 56.505 82.085 ;
        RECT 56.705 81.905 56.875 82.255 ;
        RECT 57.075 81.685 57.405 82.185 ;
        RECT 57.585 81.685 60.175 82.455 ;
        RECT 60.385 81.685 60.615 82.505 ;
        RECT 60.865 82.485 61.115 83.085 ;
        RECT 60.785 81.855 61.115 82.485 ;
        RECT 61.285 81.685 61.495 82.505 ;
        RECT 62.190 82.425 62.360 83.095 ;
        RECT 63.035 82.925 63.205 83.895 ;
        RECT 62.530 82.595 62.785 82.925 ;
        RECT 63.010 82.595 63.205 82.925 ;
        RECT 63.375 83.555 64.500 83.725 ;
        RECT 62.615 82.425 62.785 82.595 ;
        RECT 63.375 82.425 63.545 83.555 ;
        RECT 62.190 81.855 62.445 82.425 ;
        RECT 62.615 82.255 63.545 82.425 ;
        RECT 63.715 83.215 64.725 83.385 ;
        RECT 63.715 82.415 63.885 83.215 ;
        RECT 64.090 82.875 64.365 83.015 ;
        RECT 64.085 82.705 64.365 82.875 ;
        RECT 63.370 82.220 63.545 82.255 ;
        RECT 62.615 81.685 62.945 82.085 ;
        RECT 63.370 81.855 63.900 82.220 ;
        RECT 64.090 81.855 64.365 82.705 ;
        RECT 64.535 81.855 64.725 83.215 ;
        RECT 64.895 83.230 65.065 83.895 ;
        RECT 65.235 83.475 65.405 84.235 ;
        RECT 65.640 83.475 66.155 83.885 ;
        RECT 64.895 83.040 65.645 83.230 ;
        RECT 65.815 82.665 66.155 83.475 ;
        RECT 66.530 83.265 66.860 84.065 ;
        RECT 67.030 83.435 67.360 84.235 ;
        RECT 67.660 83.265 67.990 84.065 ;
        RECT 68.635 83.435 68.885 84.235 ;
        RECT 66.530 83.095 68.965 83.265 ;
        RECT 69.155 83.095 69.325 84.235 ;
        RECT 69.495 83.095 69.835 84.065 ;
        RECT 66.325 82.675 66.675 82.925 ;
        RECT 64.925 82.495 66.155 82.665 ;
        RECT 64.905 81.685 65.415 82.220 ;
        RECT 65.635 81.890 65.880 82.495 ;
        RECT 66.860 82.465 67.030 83.095 ;
        RECT 67.200 82.675 67.530 82.875 ;
        RECT 67.700 82.675 68.030 82.875 ;
        RECT 68.200 82.675 68.620 82.875 ;
        RECT 68.795 82.845 68.965 83.095 ;
        RECT 69.605 83.045 69.835 83.095 ;
        RECT 70.005 83.070 70.295 84.235 ;
        RECT 70.465 83.385 70.725 84.065 ;
        RECT 70.895 83.455 71.145 84.235 ;
        RECT 71.395 83.685 71.645 84.065 ;
        RECT 71.815 83.855 72.170 84.235 ;
        RECT 73.175 83.845 73.510 84.065 ;
        RECT 72.775 83.685 73.005 83.725 ;
        RECT 71.395 83.485 73.005 83.685 ;
        RECT 71.395 83.475 72.230 83.485 ;
        RECT 72.820 83.395 73.005 83.485 ;
        RECT 68.795 82.675 69.490 82.845 ;
        RECT 66.530 81.855 67.030 82.465 ;
        RECT 67.660 82.335 68.885 82.505 ;
        RECT 69.660 82.485 69.835 83.045 ;
        RECT 67.660 81.855 67.990 82.335 ;
        RECT 68.160 81.685 68.385 82.145 ;
        RECT 68.555 81.855 68.885 82.335 ;
        RECT 69.075 81.685 69.325 82.485 ;
        RECT 69.495 81.855 69.835 82.485 ;
        RECT 70.005 81.685 70.295 82.410 ;
        RECT 70.465 82.195 70.635 83.385 ;
        RECT 72.335 83.285 72.665 83.315 ;
        RECT 70.865 83.225 72.665 83.285 ;
        RECT 73.255 83.225 73.510 83.845 ;
        RECT 73.685 83.800 79.030 84.235 ;
        RECT 70.805 83.115 73.510 83.225 ;
        RECT 70.805 83.080 71.005 83.115 ;
        RECT 70.805 82.505 70.975 83.080 ;
        RECT 72.335 83.055 73.510 83.115 ;
        RECT 71.205 82.640 71.615 82.945 ;
        RECT 71.785 82.675 72.115 82.885 ;
        RECT 70.805 82.385 71.075 82.505 ;
        RECT 70.805 82.340 71.650 82.385 ;
        RECT 70.895 82.215 71.650 82.340 ;
        RECT 71.905 82.275 72.115 82.675 ;
        RECT 72.360 82.675 72.835 82.885 ;
        RECT 73.025 82.675 73.515 82.875 ;
        RECT 72.360 82.275 72.580 82.675 ;
        RECT 70.465 82.185 70.695 82.195 ;
        RECT 70.465 81.855 70.725 82.185 ;
        RECT 71.480 82.065 71.650 82.215 ;
        RECT 70.895 81.685 71.225 82.045 ;
        RECT 71.480 81.855 72.780 82.065 ;
        RECT 73.055 81.685 73.510 82.450 ;
        RECT 75.270 82.230 75.610 83.060 ;
        RECT 77.090 82.550 77.440 83.800 ;
        RECT 79.205 83.145 81.795 84.235 ;
        RECT 79.205 82.455 80.415 82.975 ;
        RECT 80.585 82.625 81.795 83.145 ;
        RECT 82.430 83.095 82.765 84.065 ;
        RECT 82.935 83.095 83.105 84.235 ;
        RECT 83.275 83.895 85.305 84.065 ;
        RECT 73.685 81.685 79.030 82.230 ;
        RECT 79.205 81.685 81.795 82.455 ;
        RECT 82.430 82.425 82.600 83.095 ;
        RECT 83.275 82.925 83.445 83.895 ;
        RECT 82.770 82.595 83.025 82.925 ;
        RECT 83.250 82.595 83.445 82.925 ;
        RECT 83.615 83.555 84.740 83.725 ;
        RECT 82.855 82.425 83.025 82.595 ;
        RECT 83.615 82.425 83.785 83.555 ;
        RECT 82.430 81.855 82.685 82.425 ;
        RECT 82.855 82.255 83.785 82.425 ;
        RECT 83.955 83.215 84.965 83.385 ;
        RECT 83.955 82.415 84.125 83.215 ;
        RECT 83.610 82.220 83.785 82.255 ;
        RECT 82.855 81.685 83.185 82.085 ;
        RECT 83.610 81.855 84.140 82.220 ;
        RECT 84.330 82.195 84.605 83.015 ;
        RECT 84.325 82.025 84.605 82.195 ;
        RECT 84.330 81.855 84.605 82.025 ;
        RECT 84.775 81.855 84.965 83.215 ;
        RECT 85.135 83.230 85.305 83.895 ;
        RECT 85.475 83.475 85.645 84.235 ;
        RECT 85.880 83.475 86.395 83.885 ;
        RECT 86.565 83.800 91.910 84.235 ;
        RECT 85.135 83.040 85.885 83.230 ;
        RECT 86.055 82.665 86.395 83.475 ;
        RECT 85.165 82.495 86.395 82.665 ;
        RECT 85.145 81.685 85.655 82.220 ;
        RECT 85.875 81.890 86.120 82.495 ;
        RECT 88.150 82.230 88.490 83.060 ;
        RECT 89.970 82.550 90.320 83.800 ;
        RECT 92.085 83.145 95.595 84.235 ;
        RECT 92.085 82.455 93.735 82.975 ;
        RECT 93.905 82.625 95.595 83.145 ;
        RECT 95.765 83.070 96.055 84.235 ;
        RECT 96.225 83.145 98.815 84.235 ;
        RECT 96.225 82.455 97.435 82.975 ;
        RECT 97.605 82.625 98.815 83.145 ;
        RECT 99.650 83.265 99.980 84.065 ;
        RECT 100.150 83.435 100.480 84.235 ;
        RECT 100.780 83.265 101.110 84.065 ;
        RECT 101.755 83.435 102.005 84.235 ;
        RECT 99.650 83.095 102.085 83.265 ;
        RECT 102.275 83.095 102.445 84.235 ;
        RECT 102.615 83.095 102.955 84.065 ;
        RECT 99.445 82.675 99.795 82.925 ;
        RECT 99.980 82.465 100.150 83.095 ;
        RECT 100.320 82.675 100.650 82.875 ;
        RECT 100.820 82.675 101.150 82.875 ;
        RECT 101.320 82.675 101.740 82.875 ;
        RECT 101.915 82.845 102.085 83.095 ;
        RECT 101.915 82.675 102.610 82.845 ;
        RECT 86.565 81.685 91.910 82.230 ;
        RECT 92.085 81.685 95.595 82.455 ;
        RECT 95.765 81.685 96.055 82.410 ;
        RECT 96.225 81.685 98.815 82.455 ;
        RECT 99.650 81.855 100.150 82.465 ;
        RECT 100.780 82.335 102.005 82.505 ;
        RECT 102.780 82.485 102.955 83.095 ;
        RECT 100.780 81.855 101.110 82.335 ;
        RECT 101.280 81.685 101.505 82.145 ;
        RECT 101.675 81.855 102.005 82.335 ;
        RECT 102.195 81.685 102.445 82.485 ;
        RECT 102.615 81.855 102.955 82.485 ;
        RECT 103.125 83.095 103.465 84.065 ;
        RECT 103.635 83.095 103.805 84.235 ;
        RECT 104.075 83.435 104.325 84.235 ;
        RECT 104.970 83.265 105.300 84.065 ;
        RECT 105.600 83.435 105.930 84.235 ;
        RECT 106.100 83.265 106.430 84.065 ;
        RECT 103.995 83.095 106.430 83.265 ;
        RECT 107.725 83.475 108.240 83.885 ;
        RECT 108.475 83.475 108.645 84.235 ;
        RECT 108.815 83.895 110.845 84.065 ;
        RECT 103.125 82.485 103.300 83.095 ;
        RECT 103.995 82.845 104.165 83.095 ;
        RECT 103.470 82.675 104.165 82.845 ;
        RECT 104.340 82.675 104.760 82.875 ;
        RECT 104.930 82.675 105.260 82.875 ;
        RECT 105.430 82.675 105.760 82.875 ;
        RECT 103.125 81.855 103.465 82.485 ;
        RECT 103.635 81.685 103.885 82.485 ;
        RECT 104.075 82.335 105.300 82.505 ;
        RECT 104.075 81.855 104.405 82.335 ;
        RECT 104.575 81.685 104.800 82.145 ;
        RECT 104.970 81.855 105.300 82.335 ;
        RECT 105.930 82.465 106.100 83.095 ;
        RECT 106.285 82.675 106.635 82.925 ;
        RECT 107.725 82.665 108.065 83.475 ;
        RECT 108.815 83.230 108.985 83.895 ;
        RECT 109.380 83.555 110.505 83.725 ;
        RECT 108.235 83.040 108.985 83.230 ;
        RECT 109.155 83.215 110.165 83.385 ;
        RECT 107.725 82.495 108.955 82.665 ;
        RECT 105.930 81.855 106.430 82.465 ;
        RECT 108.000 81.890 108.245 82.495 ;
        RECT 108.465 81.685 108.975 82.220 ;
        RECT 109.155 81.855 109.345 83.215 ;
        RECT 109.515 82.195 109.790 83.015 ;
        RECT 109.995 82.415 110.165 83.215 ;
        RECT 110.335 82.425 110.505 83.555 ;
        RECT 110.675 82.925 110.845 83.895 ;
        RECT 111.015 83.095 111.185 84.235 ;
        RECT 111.355 83.095 111.690 84.065 ;
        RECT 111.955 83.565 112.125 84.065 ;
        RECT 112.295 83.735 112.625 84.235 ;
        RECT 111.955 83.395 112.620 83.565 ;
        RECT 110.675 82.595 110.870 82.925 ;
        RECT 111.095 82.595 111.350 82.925 ;
        RECT 111.095 82.425 111.265 82.595 ;
        RECT 111.520 82.425 111.690 83.095 ;
        RECT 111.870 82.575 112.220 83.225 ;
        RECT 110.335 82.255 111.265 82.425 ;
        RECT 110.335 82.220 110.510 82.255 ;
        RECT 109.515 82.025 109.795 82.195 ;
        RECT 109.515 81.855 109.790 82.025 ;
        RECT 109.980 81.855 110.510 82.220 ;
        RECT 110.935 81.685 111.265 82.085 ;
        RECT 111.435 81.855 111.690 82.425 ;
        RECT 112.390 82.405 112.620 83.395 ;
        RECT 111.955 82.235 112.620 82.405 ;
        RECT 111.955 81.945 112.125 82.235 ;
        RECT 112.295 81.685 112.625 82.065 ;
        RECT 112.795 81.945 113.020 84.065 ;
        RECT 113.235 83.735 113.565 84.235 ;
        RECT 113.735 83.565 113.905 84.065 ;
        RECT 114.140 83.850 114.970 84.020 ;
        RECT 115.210 83.855 115.590 84.235 ;
        RECT 113.210 83.395 113.905 83.565 ;
        RECT 113.210 82.425 113.380 83.395 ;
        RECT 113.550 82.605 113.960 83.225 ;
        RECT 114.130 83.175 114.630 83.555 ;
        RECT 113.210 82.235 113.905 82.425 ;
        RECT 114.130 82.305 114.350 83.175 ;
        RECT 114.800 83.005 114.970 83.850 ;
        RECT 115.770 83.685 115.940 83.975 ;
        RECT 116.110 83.855 116.440 84.235 ;
        RECT 116.910 83.765 117.540 84.015 ;
        RECT 117.720 83.855 118.140 84.235 ;
        RECT 117.370 83.685 117.540 83.765 ;
        RECT 118.340 83.685 118.580 83.975 ;
        RECT 115.140 83.435 116.510 83.685 ;
        RECT 115.140 83.175 115.390 83.435 ;
        RECT 115.900 83.005 116.150 83.165 ;
        RECT 114.800 82.835 116.150 83.005 ;
        RECT 114.800 82.795 115.220 82.835 ;
        RECT 114.530 82.245 114.880 82.615 ;
        RECT 113.235 81.685 113.565 82.065 ;
        RECT 113.735 81.905 113.905 82.235 ;
        RECT 115.050 82.065 115.220 82.795 ;
        RECT 116.320 82.665 116.510 83.435 ;
        RECT 115.390 82.335 115.800 82.665 ;
        RECT 116.090 82.325 116.510 82.665 ;
        RECT 116.680 83.255 117.200 83.565 ;
        RECT 117.370 83.515 118.580 83.685 ;
        RECT 118.810 83.545 119.140 84.235 ;
        RECT 116.680 82.495 116.850 83.255 ;
        RECT 117.020 82.665 117.200 83.075 ;
        RECT 117.370 83.005 117.540 83.515 ;
        RECT 119.310 83.365 119.480 83.975 ;
        RECT 119.750 83.515 120.080 84.025 ;
        RECT 119.310 83.345 119.630 83.365 ;
        RECT 117.710 83.175 119.630 83.345 ;
        RECT 117.370 82.835 119.270 83.005 ;
        RECT 117.600 82.495 117.930 82.615 ;
        RECT 116.680 82.325 117.930 82.495 ;
        RECT 114.205 81.865 115.220 82.065 ;
        RECT 115.390 81.685 115.800 82.125 ;
        RECT 116.090 81.895 116.340 82.325 ;
        RECT 116.540 81.685 116.860 82.145 ;
        RECT 118.100 82.075 118.270 82.835 ;
        RECT 118.940 82.775 119.270 82.835 ;
        RECT 118.460 82.605 118.790 82.665 ;
        RECT 118.460 82.335 119.120 82.605 ;
        RECT 119.440 82.280 119.630 83.175 ;
        RECT 117.420 81.905 118.270 82.075 ;
        RECT 118.470 81.685 119.130 82.165 ;
        RECT 119.310 81.950 119.630 82.280 ;
        RECT 119.830 82.925 120.080 83.515 ;
        RECT 120.260 83.435 120.545 84.235 ;
        RECT 120.725 83.255 120.980 83.925 ;
        RECT 120.800 83.215 120.980 83.255 ;
        RECT 120.800 83.045 121.065 83.215 ;
        RECT 121.525 83.070 121.815 84.235 ;
        RECT 122.445 83.145 123.655 84.235 ;
        RECT 119.830 82.595 120.630 82.925 ;
        RECT 119.830 81.945 120.080 82.595 ;
        RECT 120.800 82.395 120.980 83.045 ;
        RECT 122.445 82.605 122.965 83.145 ;
        RECT 123.135 82.435 123.655 82.975 ;
        RECT 120.260 81.685 120.545 82.145 ;
        RECT 120.725 81.865 120.980 82.395 ;
        RECT 121.525 81.685 121.815 82.410 ;
        RECT 122.445 81.685 123.655 82.435 ;
        RECT 5.520 81.515 123.740 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 6.985 80.970 12.330 81.515 ;
        RECT 12.505 80.970 17.850 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 8.570 80.140 8.910 80.970 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 10.390 79.400 10.740 80.650 ;
        RECT 14.090 80.140 14.430 80.970 ;
        RECT 18.945 80.840 19.215 81.185 ;
        RECT 19.405 81.115 19.785 81.515 ;
        RECT 19.955 80.945 20.125 81.295 ;
        RECT 20.295 81.115 20.625 81.515 ;
        RECT 20.825 80.945 20.995 81.295 ;
        RECT 21.195 81.015 21.525 81.515 ;
        RECT 15.910 79.400 16.260 80.650 ;
        RECT 18.945 80.105 19.115 80.840 ;
        RECT 19.385 80.775 20.995 80.945 ;
        RECT 19.385 80.605 19.555 80.775 ;
        RECT 19.285 80.275 19.555 80.605 ;
        RECT 19.725 80.275 20.130 80.605 ;
        RECT 19.385 80.105 19.555 80.275 ;
        RECT 20.300 80.155 21.010 80.605 ;
        RECT 21.180 80.275 21.530 80.845 ;
        RECT 21.705 80.715 22.045 81.345 ;
        RECT 22.215 80.715 22.465 81.515 ;
        RECT 22.655 80.865 22.985 81.345 ;
        RECT 23.155 81.055 23.380 81.515 ;
        RECT 23.550 80.865 23.880 81.345 ;
        RECT 21.705 80.665 21.935 80.715 ;
        RECT 22.655 80.695 23.880 80.865 ;
        RECT 24.510 80.735 25.010 81.345 ;
        RECT 25.590 80.735 26.090 81.345 ;
        RECT 6.985 78.965 12.330 79.400 ;
        RECT 12.505 78.965 17.850 79.400 ;
        RECT 18.945 79.135 19.215 80.105 ;
        RECT 19.385 79.935 20.110 80.105 ;
        RECT 20.300 79.985 21.015 80.155 ;
        RECT 21.705 80.105 21.880 80.665 ;
        RECT 22.050 80.355 22.745 80.525 ;
        RECT 22.575 80.105 22.745 80.355 ;
        RECT 22.920 80.325 23.340 80.525 ;
        RECT 23.510 80.325 23.840 80.525 ;
        RECT 24.010 80.325 24.340 80.525 ;
        RECT 24.510 80.105 24.680 80.735 ;
        RECT 24.865 80.275 25.215 80.525 ;
        RECT 25.385 80.275 25.735 80.525 ;
        RECT 25.920 80.105 26.090 80.735 ;
        RECT 26.720 80.865 27.050 81.345 ;
        RECT 27.220 81.055 27.445 81.515 ;
        RECT 27.615 80.865 27.945 81.345 ;
        RECT 26.720 80.695 27.945 80.865 ;
        RECT 28.135 80.715 28.385 81.515 ;
        RECT 28.555 80.715 28.895 81.345 ;
        RECT 26.260 80.325 26.590 80.525 ;
        RECT 26.760 80.325 27.090 80.525 ;
        RECT 27.260 80.325 27.680 80.525 ;
        RECT 27.855 80.355 28.550 80.525 ;
        RECT 27.855 80.105 28.025 80.355 ;
        RECT 28.720 80.105 28.895 80.715 ;
        RECT 29.065 80.745 30.735 81.515 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 31.825 80.745 35.335 81.515 ;
        RECT 35.505 80.765 36.715 81.515 ;
        RECT 36.885 80.840 37.145 81.345 ;
        RECT 37.325 81.135 37.655 81.515 ;
        RECT 37.835 80.965 38.005 81.345 ;
        RECT 29.065 80.225 29.815 80.745 ;
        RECT 19.940 79.815 20.110 79.935 ;
        RECT 21.210 79.815 21.530 80.105 ;
        RECT 19.425 78.965 19.705 79.765 ;
        RECT 19.940 79.645 21.530 79.815 ;
        RECT 19.875 79.185 21.530 79.475 ;
        RECT 21.705 79.135 22.045 80.105 ;
        RECT 22.215 78.965 22.385 80.105 ;
        RECT 22.575 79.935 25.010 80.105 ;
        RECT 22.655 78.965 22.905 79.765 ;
        RECT 23.550 79.135 23.880 79.935 ;
        RECT 24.180 78.965 24.510 79.765 ;
        RECT 24.680 79.135 25.010 79.935 ;
        RECT 25.590 79.935 28.025 80.105 ;
        RECT 25.590 79.135 25.920 79.935 ;
        RECT 26.090 78.965 26.420 79.765 ;
        RECT 26.720 79.135 27.050 79.935 ;
        RECT 27.695 78.965 27.945 79.765 ;
        RECT 28.215 78.965 28.385 80.105 ;
        RECT 28.555 79.135 28.895 80.105 ;
        RECT 29.985 80.055 30.735 80.575 ;
        RECT 31.825 80.225 33.475 80.745 ;
        RECT 29.065 78.965 30.735 80.055 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 33.645 80.055 35.335 80.575 ;
        RECT 35.505 80.225 36.025 80.765 ;
        RECT 36.195 80.055 36.715 80.595 ;
        RECT 31.825 78.965 35.335 80.055 ;
        RECT 35.505 78.965 36.715 80.055 ;
        RECT 36.885 80.040 37.055 80.840 ;
        RECT 37.340 80.795 38.005 80.965 ;
        RECT 38.355 80.965 38.525 81.345 ;
        RECT 38.705 81.135 39.035 81.515 ;
        RECT 38.355 80.795 39.020 80.965 ;
        RECT 39.215 80.840 39.475 81.345 ;
        RECT 37.340 80.540 37.510 80.795 ;
        RECT 37.225 80.210 37.510 80.540 ;
        RECT 37.745 80.245 38.075 80.615 ;
        RECT 38.285 80.245 38.615 80.615 ;
        RECT 38.850 80.540 39.020 80.795 ;
        RECT 37.340 80.065 37.510 80.210 ;
        RECT 38.850 80.210 39.135 80.540 ;
        RECT 38.850 80.065 39.020 80.210 ;
        RECT 36.885 79.135 37.155 80.040 ;
        RECT 37.340 79.895 38.005 80.065 ;
        RECT 37.325 78.965 37.655 79.725 ;
        RECT 37.835 79.135 38.005 79.895 ;
        RECT 38.355 79.895 39.020 80.065 ;
        RECT 39.305 80.040 39.475 80.840 ;
        RECT 39.735 80.965 39.905 81.255 ;
        RECT 40.075 81.135 40.405 81.515 ;
        RECT 39.735 80.795 40.400 80.965 ;
        RECT 38.355 79.135 38.525 79.895 ;
        RECT 38.705 78.965 39.035 79.725 ;
        RECT 39.205 79.135 39.475 80.040 ;
        RECT 39.650 79.975 40.000 80.625 ;
        RECT 40.170 79.805 40.400 80.795 ;
        RECT 39.735 79.635 40.400 79.805 ;
        RECT 39.735 79.135 39.905 79.635 ;
        RECT 40.075 78.965 40.405 79.465 ;
        RECT 40.575 79.135 40.800 81.255 ;
        RECT 41.015 81.135 41.345 81.515 ;
        RECT 41.515 80.965 41.685 81.295 ;
        RECT 41.985 81.135 43.000 81.335 ;
        RECT 40.990 80.775 41.685 80.965 ;
        RECT 40.990 79.805 41.160 80.775 ;
        RECT 41.330 79.975 41.740 80.595 ;
        RECT 41.910 80.025 42.130 80.895 ;
        RECT 42.310 80.585 42.660 80.955 ;
        RECT 42.830 80.405 43.000 81.135 ;
        RECT 43.170 81.075 43.580 81.515 ;
        RECT 43.870 80.875 44.120 81.305 ;
        RECT 44.320 81.055 44.640 81.515 ;
        RECT 45.200 81.125 46.050 81.295 ;
        RECT 43.170 80.535 43.580 80.865 ;
        RECT 43.870 80.535 44.290 80.875 ;
        RECT 42.580 80.365 43.000 80.405 ;
        RECT 42.580 80.195 43.930 80.365 ;
        RECT 40.990 79.635 41.685 79.805 ;
        RECT 41.910 79.645 42.410 80.025 ;
        RECT 41.015 78.965 41.345 79.465 ;
        RECT 41.515 79.135 41.685 79.635 ;
        RECT 42.580 79.350 42.750 80.195 ;
        RECT 43.680 80.035 43.930 80.195 ;
        RECT 42.920 79.765 43.170 80.025 ;
        RECT 44.100 79.765 44.290 80.535 ;
        RECT 42.920 79.515 44.290 79.765 ;
        RECT 44.460 80.705 45.710 80.875 ;
        RECT 44.460 79.945 44.630 80.705 ;
        RECT 45.380 80.585 45.710 80.705 ;
        RECT 44.800 80.125 44.980 80.535 ;
        RECT 45.880 80.365 46.050 81.125 ;
        RECT 46.250 81.035 46.910 81.515 ;
        RECT 47.090 80.920 47.410 81.250 ;
        RECT 46.240 80.595 46.900 80.865 ;
        RECT 46.240 80.535 46.570 80.595 ;
        RECT 46.720 80.365 47.050 80.425 ;
        RECT 45.150 80.195 47.050 80.365 ;
        RECT 44.460 79.635 44.980 79.945 ;
        RECT 45.150 79.685 45.320 80.195 ;
        RECT 47.220 80.025 47.410 80.920 ;
        RECT 45.490 79.855 47.410 80.025 ;
        RECT 47.090 79.835 47.410 79.855 ;
        RECT 47.610 80.605 47.860 81.255 ;
        RECT 48.040 81.055 48.325 81.515 ;
        RECT 48.505 81.175 48.760 81.335 ;
        RECT 48.505 81.005 48.845 81.175 ;
        RECT 48.505 80.805 48.760 81.005 ;
        RECT 47.610 80.275 48.410 80.605 ;
        RECT 45.150 79.515 46.360 79.685 ;
        RECT 41.920 79.180 42.750 79.350 ;
        RECT 42.990 78.965 43.370 79.345 ;
        RECT 43.550 79.225 43.720 79.515 ;
        RECT 45.150 79.435 45.320 79.515 ;
        RECT 43.890 78.965 44.220 79.345 ;
        RECT 44.690 79.185 45.320 79.435 ;
        RECT 45.500 78.965 45.920 79.345 ;
        RECT 46.120 79.225 46.360 79.515 ;
        RECT 46.590 78.965 46.920 79.655 ;
        RECT 47.090 79.225 47.260 79.835 ;
        RECT 47.610 79.685 47.860 80.275 ;
        RECT 48.580 79.945 48.760 80.805 ;
        RECT 49.305 80.765 50.515 81.515 ;
        RECT 49.305 80.225 49.825 80.765 ;
        RECT 50.890 80.735 51.390 81.345 ;
        RECT 49.995 80.055 50.515 80.595 ;
        RECT 50.685 80.275 51.035 80.525 ;
        RECT 51.220 80.105 51.390 80.735 ;
        RECT 52.020 80.865 52.350 81.345 ;
        RECT 52.520 81.055 52.745 81.515 ;
        RECT 52.915 80.865 53.245 81.345 ;
        RECT 52.020 80.695 53.245 80.865 ;
        RECT 53.435 80.715 53.685 81.515 ;
        RECT 53.855 80.715 54.195 81.345 ;
        RECT 54.375 81.015 54.705 81.515 ;
        RECT 54.905 80.945 55.075 81.295 ;
        RECT 55.275 81.115 55.605 81.515 ;
        RECT 55.775 80.945 55.945 81.295 ;
        RECT 56.115 81.115 56.495 81.515 ;
        RECT 53.965 80.665 54.195 80.715 ;
        RECT 51.560 80.325 51.890 80.525 ;
        RECT 52.060 80.325 52.390 80.525 ;
        RECT 52.560 80.325 52.980 80.525 ;
        RECT 53.155 80.355 53.850 80.525 ;
        RECT 53.155 80.105 53.325 80.355 ;
        RECT 54.020 80.105 54.195 80.665 ;
        RECT 54.370 80.275 54.720 80.845 ;
        RECT 54.905 80.775 56.515 80.945 ;
        RECT 56.685 80.840 56.955 81.185 ;
        RECT 56.345 80.605 56.515 80.775 ;
        RECT 47.530 79.175 47.860 79.685 ;
        RECT 48.040 78.965 48.325 79.765 ;
        RECT 48.505 79.275 48.760 79.945 ;
        RECT 49.305 78.965 50.515 80.055 ;
        RECT 50.890 79.935 53.325 80.105 ;
        RECT 50.890 79.135 51.220 79.935 ;
        RECT 51.390 78.965 51.720 79.765 ;
        RECT 52.020 79.135 52.350 79.935 ;
        RECT 52.995 78.965 53.245 79.765 ;
        RECT 53.515 78.965 53.685 80.105 ;
        RECT 53.855 79.135 54.195 80.105 ;
        RECT 54.370 79.815 54.690 80.105 ;
        RECT 54.890 79.985 55.600 80.605 ;
        RECT 55.770 80.275 56.175 80.605 ;
        RECT 56.345 80.275 56.615 80.605 ;
        RECT 56.345 80.105 56.515 80.275 ;
        RECT 56.785 80.105 56.955 80.840 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 57.585 80.970 62.930 81.515 ;
        RECT 59.170 80.140 59.510 80.970 ;
        RECT 63.105 80.745 65.695 81.515 ;
        RECT 65.955 80.965 66.125 81.255 ;
        RECT 66.295 81.135 66.625 81.515 ;
        RECT 65.955 80.795 66.620 80.965 ;
        RECT 55.790 79.935 56.515 80.105 ;
        RECT 55.790 79.815 55.960 79.935 ;
        RECT 54.370 79.645 55.960 79.815 ;
        RECT 54.370 79.185 56.025 79.475 ;
        RECT 56.195 78.965 56.475 79.765 ;
        RECT 56.685 79.135 56.955 80.105 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 60.990 79.400 61.340 80.650 ;
        RECT 63.105 80.225 64.315 80.745 ;
        RECT 64.485 80.055 65.695 80.575 ;
        RECT 57.585 78.965 62.930 79.400 ;
        RECT 63.105 78.965 65.695 80.055 ;
        RECT 65.870 79.975 66.220 80.625 ;
        RECT 66.390 79.805 66.620 80.795 ;
        RECT 65.955 79.635 66.620 79.805 ;
        RECT 65.955 79.135 66.125 79.635 ;
        RECT 66.295 78.965 66.625 79.465 ;
        RECT 66.795 79.135 67.020 81.255 ;
        RECT 67.235 81.135 67.565 81.515 ;
        RECT 67.735 80.965 67.905 81.295 ;
        RECT 68.205 81.135 69.220 81.335 ;
        RECT 67.210 80.775 67.905 80.965 ;
        RECT 67.210 79.805 67.380 80.775 ;
        RECT 67.550 79.975 67.960 80.595 ;
        RECT 68.130 80.025 68.350 80.895 ;
        RECT 68.530 80.585 68.880 80.955 ;
        RECT 69.050 80.405 69.220 81.135 ;
        RECT 69.390 81.075 69.800 81.515 ;
        RECT 70.090 80.875 70.340 81.305 ;
        RECT 70.540 81.055 70.860 81.515 ;
        RECT 71.420 81.125 72.270 81.295 ;
        RECT 69.390 80.535 69.800 80.865 ;
        RECT 70.090 80.535 70.510 80.875 ;
        RECT 68.800 80.365 69.220 80.405 ;
        RECT 68.800 80.195 70.150 80.365 ;
        RECT 67.210 79.635 67.905 79.805 ;
        RECT 68.130 79.645 68.630 80.025 ;
        RECT 67.235 78.965 67.565 79.465 ;
        RECT 67.735 79.135 67.905 79.635 ;
        RECT 68.800 79.350 68.970 80.195 ;
        RECT 69.900 80.035 70.150 80.195 ;
        RECT 69.140 79.765 69.390 80.025 ;
        RECT 70.320 79.765 70.510 80.535 ;
        RECT 69.140 79.515 70.510 79.765 ;
        RECT 70.680 80.705 71.930 80.875 ;
        RECT 70.680 79.945 70.850 80.705 ;
        RECT 71.600 80.585 71.930 80.705 ;
        RECT 71.020 80.125 71.200 80.535 ;
        RECT 72.100 80.365 72.270 81.125 ;
        RECT 72.470 81.035 73.130 81.515 ;
        RECT 73.310 80.920 73.630 81.250 ;
        RECT 72.460 80.595 73.120 80.865 ;
        RECT 72.460 80.535 72.790 80.595 ;
        RECT 72.940 80.365 73.270 80.425 ;
        RECT 71.370 80.195 73.270 80.365 ;
        RECT 70.680 79.635 71.200 79.945 ;
        RECT 71.370 79.685 71.540 80.195 ;
        RECT 73.440 80.025 73.630 80.920 ;
        RECT 71.710 79.855 73.630 80.025 ;
        RECT 73.310 79.835 73.630 79.855 ;
        RECT 73.830 80.605 74.080 81.255 ;
        RECT 74.260 81.055 74.545 81.515 ;
        RECT 74.725 80.805 74.980 81.335 ;
        RECT 73.830 80.275 74.630 80.605 ;
        RECT 71.370 79.515 72.580 79.685 ;
        RECT 68.140 79.180 68.970 79.350 ;
        RECT 69.210 78.965 69.590 79.345 ;
        RECT 69.770 79.225 69.940 79.515 ;
        RECT 71.370 79.435 71.540 79.515 ;
        RECT 70.110 78.965 70.440 79.345 ;
        RECT 70.910 79.185 71.540 79.435 ;
        RECT 71.720 78.965 72.140 79.345 ;
        RECT 72.340 79.225 72.580 79.515 ;
        RECT 72.810 78.965 73.140 79.655 ;
        RECT 73.310 79.225 73.480 79.835 ;
        RECT 73.830 79.685 74.080 80.275 ;
        RECT 74.800 79.945 74.980 80.805 ;
        RECT 75.565 80.695 75.795 81.515 ;
        RECT 75.965 80.715 76.295 81.345 ;
        RECT 75.545 80.275 75.875 80.525 ;
        RECT 76.045 80.115 76.295 80.715 ;
        RECT 76.465 80.695 76.675 81.515 ;
        RECT 76.905 80.765 78.115 81.515 ;
        RECT 78.285 80.840 78.545 81.345 ;
        RECT 78.725 81.135 79.055 81.515 ;
        RECT 79.235 80.965 79.405 81.345 ;
        RECT 76.905 80.225 77.425 80.765 ;
        RECT 73.750 79.175 74.080 79.685 ;
        RECT 74.260 78.965 74.545 79.765 ;
        RECT 74.725 79.475 74.980 79.945 ;
        RECT 74.725 79.305 75.065 79.475 ;
        RECT 74.725 79.275 74.980 79.305 ;
        RECT 75.565 78.965 75.795 80.105 ;
        RECT 75.965 79.135 76.295 80.115 ;
        RECT 76.465 78.965 76.675 80.105 ;
        RECT 77.595 80.055 78.115 80.595 ;
        RECT 76.905 78.965 78.115 80.055 ;
        RECT 78.285 80.040 78.455 80.840 ;
        RECT 78.740 80.795 79.405 80.965 ;
        RECT 78.740 80.540 78.910 80.795 ;
        RECT 79.665 80.765 80.875 81.515 ;
        RECT 78.625 80.210 78.910 80.540 ;
        RECT 79.145 80.245 79.475 80.615 ;
        RECT 79.665 80.225 80.185 80.765 ;
        RECT 81.105 80.695 81.315 81.515 ;
        RECT 81.485 80.715 81.815 81.345 ;
        RECT 78.740 80.065 78.910 80.210 ;
        RECT 78.285 79.135 78.555 80.040 ;
        RECT 78.740 79.895 79.405 80.065 ;
        RECT 80.355 80.055 80.875 80.595 ;
        RECT 81.485 80.115 81.735 80.715 ;
        RECT 81.985 80.695 82.215 81.515 ;
        RECT 82.885 80.790 83.175 81.515 ;
        RECT 84.010 80.735 84.510 81.345 ;
        RECT 81.905 80.275 82.235 80.525 ;
        RECT 83.805 80.275 84.155 80.525 ;
        RECT 78.725 78.965 79.055 79.725 ;
        RECT 79.235 79.135 79.405 79.895 ;
        RECT 79.665 78.965 80.875 80.055 ;
        RECT 81.105 78.965 81.315 80.105 ;
        RECT 81.485 79.135 81.815 80.115 ;
        RECT 81.985 78.965 82.215 80.105 ;
        RECT 82.885 78.965 83.175 80.130 ;
        RECT 84.340 80.105 84.510 80.735 ;
        RECT 85.140 80.865 85.470 81.345 ;
        RECT 85.640 81.055 85.865 81.515 ;
        RECT 86.035 80.865 86.365 81.345 ;
        RECT 85.140 80.695 86.365 80.865 ;
        RECT 86.555 80.715 86.805 81.515 ;
        RECT 86.975 80.715 87.315 81.345 ;
        RECT 87.495 81.015 87.825 81.515 ;
        RECT 88.025 80.945 88.195 81.295 ;
        RECT 88.395 81.115 88.725 81.515 ;
        RECT 88.895 80.945 89.065 81.295 ;
        RECT 89.235 81.115 89.615 81.515 ;
        RECT 87.085 80.665 87.315 80.715 ;
        RECT 84.680 80.325 85.010 80.525 ;
        RECT 85.180 80.325 85.510 80.525 ;
        RECT 85.680 80.325 86.100 80.525 ;
        RECT 86.275 80.355 86.970 80.525 ;
        RECT 86.275 80.105 86.445 80.355 ;
        RECT 87.140 80.105 87.315 80.665 ;
        RECT 87.490 80.275 87.840 80.845 ;
        RECT 88.025 80.775 89.635 80.945 ;
        RECT 89.805 80.840 90.075 81.185 ;
        RECT 90.245 80.970 95.590 81.515 ;
        RECT 89.465 80.605 89.635 80.775 ;
        RECT 84.010 79.935 86.445 80.105 ;
        RECT 84.010 79.135 84.340 79.935 ;
        RECT 84.510 78.965 84.840 79.765 ;
        RECT 85.140 79.135 85.470 79.935 ;
        RECT 86.115 78.965 86.365 79.765 ;
        RECT 86.635 78.965 86.805 80.105 ;
        RECT 86.975 79.135 87.315 80.105 ;
        RECT 87.490 79.815 87.810 80.105 ;
        RECT 88.010 79.985 88.720 80.605 ;
        RECT 88.890 80.275 89.295 80.605 ;
        RECT 89.465 80.275 89.735 80.605 ;
        RECT 89.465 80.105 89.635 80.275 ;
        RECT 89.905 80.105 90.075 80.840 ;
        RECT 91.830 80.140 92.170 80.970 ;
        RECT 95.765 80.715 96.105 81.345 ;
        RECT 96.275 80.715 96.525 81.515 ;
        RECT 96.715 80.865 97.045 81.345 ;
        RECT 97.215 81.055 97.440 81.515 ;
        RECT 97.610 80.865 97.940 81.345 ;
        RECT 88.910 79.935 89.635 80.105 ;
        RECT 88.910 79.815 89.080 79.935 ;
        RECT 87.490 79.645 89.080 79.815 ;
        RECT 87.490 79.185 89.145 79.475 ;
        RECT 89.315 78.965 89.595 79.765 ;
        RECT 89.805 79.135 90.075 80.105 ;
        RECT 93.650 79.400 94.000 80.650 ;
        RECT 95.765 80.105 95.940 80.715 ;
        RECT 96.715 80.695 97.940 80.865 ;
        RECT 98.570 80.735 99.070 81.345 ;
        RECT 99.650 80.735 100.150 81.345 ;
        RECT 96.110 80.355 96.805 80.525 ;
        RECT 96.635 80.105 96.805 80.355 ;
        RECT 96.980 80.325 97.400 80.525 ;
        RECT 97.570 80.325 97.900 80.525 ;
        RECT 98.070 80.325 98.400 80.525 ;
        RECT 98.570 80.105 98.740 80.735 ;
        RECT 98.925 80.275 99.275 80.525 ;
        RECT 99.445 80.275 99.795 80.525 ;
        RECT 99.980 80.105 100.150 80.735 ;
        RECT 100.780 80.865 101.110 81.345 ;
        RECT 101.280 81.055 101.505 81.515 ;
        RECT 101.675 80.865 102.005 81.345 ;
        RECT 100.780 80.695 102.005 80.865 ;
        RECT 102.195 80.715 102.445 81.515 ;
        RECT 102.615 80.715 102.955 81.345 ;
        RECT 103.125 80.970 108.470 81.515 ;
        RECT 100.320 80.325 100.650 80.525 ;
        RECT 100.820 80.325 101.150 80.525 ;
        RECT 101.320 80.325 101.740 80.525 ;
        RECT 101.915 80.355 102.610 80.525 ;
        RECT 101.915 80.105 102.085 80.355 ;
        RECT 102.780 80.105 102.955 80.715 ;
        RECT 104.710 80.140 105.050 80.970 ;
        RECT 108.645 80.790 108.935 81.515 ;
        RECT 109.195 80.965 109.365 81.345 ;
        RECT 109.545 81.135 109.875 81.515 ;
        RECT 109.195 80.795 109.860 80.965 ;
        RECT 110.055 80.840 110.315 81.345 ;
        RECT 90.245 78.965 95.590 79.400 ;
        RECT 95.765 79.135 96.105 80.105 ;
        RECT 96.275 78.965 96.445 80.105 ;
        RECT 96.635 79.935 99.070 80.105 ;
        RECT 96.715 78.965 96.965 79.765 ;
        RECT 97.610 79.135 97.940 79.935 ;
        RECT 98.240 78.965 98.570 79.765 ;
        RECT 98.740 79.135 99.070 79.935 ;
        RECT 99.650 79.935 102.085 80.105 ;
        RECT 99.650 79.135 99.980 79.935 ;
        RECT 100.150 78.965 100.480 79.765 ;
        RECT 100.780 79.135 101.110 79.935 ;
        RECT 101.755 78.965 102.005 79.765 ;
        RECT 102.275 78.965 102.445 80.105 ;
        RECT 102.615 79.135 102.955 80.105 ;
        RECT 106.530 79.400 106.880 80.650 ;
        RECT 109.125 80.245 109.455 80.615 ;
        RECT 109.690 80.540 109.860 80.795 ;
        RECT 109.690 80.210 109.975 80.540 ;
        RECT 103.125 78.965 108.470 79.400 ;
        RECT 108.645 78.965 108.935 80.130 ;
        RECT 109.690 80.065 109.860 80.210 ;
        RECT 109.195 79.895 109.860 80.065 ;
        RECT 110.145 80.040 110.315 80.840 ;
        RECT 110.485 80.765 111.695 81.515 ;
        RECT 111.870 80.775 112.125 81.345 ;
        RECT 112.295 81.115 112.625 81.515 ;
        RECT 113.050 80.980 113.580 81.345 ;
        RECT 113.770 81.175 114.045 81.345 ;
        RECT 113.765 81.005 114.045 81.175 ;
        RECT 113.050 80.945 113.225 80.980 ;
        RECT 112.295 80.775 113.225 80.945 ;
        RECT 110.485 80.225 111.005 80.765 ;
        RECT 111.175 80.055 111.695 80.595 ;
        RECT 109.195 79.135 109.365 79.895 ;
        RECT 109.545 78.965 109.875 79.725 ;
        RECT 110.045 79.135 110.315 80.040 ;
        RECT 110.485 78.965 111.695 80.055 ;
        RECT 111.870 80.105 112.040 80.775 ;
        RECT 112.295 80.605 112.465 80.775 ;
        RECT 112.210 80.275 112.465 80.605 ;
        RECT 112.690 80.275 112.885 80.605 ;
        RECT 111.870 79.135 112.205 80.105 ;
        RECT 112.375 78.965 112.545 80.105 ;
        RECT 112.715 79.305 112.885 80.275 ;
        RECT 113.055 79.645 113.225 80.775 ;
        RECT 113.395 79.985 113.565 80.785 ;
        RECT 113.770 80.185 114.045 81.005 ;
        RECT 114.215 79.985 114.405 81.345 ;
        RECT 114.585 80.980 115.095 81.515 ;
        RECT 115.315 80.705 115.560 81.310 ;
        RECT 114.605 80.535 115.835 80.705 ;
        RECT 116.065 80.695 116.275 81.515 ;
        RECT 116.445 80.715 116.775 81.345 ;
        RECT 113.395 79.815 114.405 79.985 ;
        RECT 114.575 79.970 115.325 80.160 ;
        RECT 113.055 79.475 114.180 79.645 ;
        RECT 114.575 79.305 114.745 79.970 ;
        RECT 115.495 79.725 115.835 80.535 ;
        RECT 116.445 80.115 116.695 80.715 ;
        RECT 116.945 80.695 117.175 81.515 ;
        RECT 117.385 80.745 120.895 81.515 ;
        RECT 121.065 80.765 122.275 81.515 ;
        RECT 122.445 80.765 123.655 81.515 ;
        RECT 116.865 80.275 117.195 80.525 ;
        RECT 117.385 80.225 119.035 80.745 ;
        RECT 112.715 79.135 114.745 79.305 ;
        RECT 114.915 78.965 115.085 79.725 ;
        RECT 115.320 79.315 115.835 79.725 ;
        RECT 116.065 78.965 116.275 80.105 ;
        RECT 116.445 79.135 116.775 80.115 ;
        RECT 116.945 78.965 117.175 80.105 ;
        RECT 119.205 80.055 120.895 80.575 ;
        RECT 121.065 80.225 121.585 80.765 ;
        RECT 121.755 80.055 122.275 80.595 ;
        RECT 117.385 78.965 120.895 80.055 ;
        RECT 121.065 78.965 122.275 80.055 ;
        RECT 122.445 80.055 122.965 80.595 ;
        RECT 123.135 80.225 123.655 80.765 ;
        RECT 122.445 78.965 123.655 80.055 ;
        RECT 5.520 78.795 123.740 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 6.985 78.360 12.330 78.795 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 8.570 76.790 8.910 77.620 ;
        RECT 10.390 77.110 10.740 78.360 ;
        RECT 13.430 77.655 13.765 78.625 ;
        RECT 13.935 77.655 14.105 78.795 ;
        RECT 14.275 78.455 16.305 78.625 ;
        RECT 13.430 76.985 13.600 77.655 ;
        RECT 14.275 77.485 14.445 78.455 ;
        RECT 13.770 77.155 14.025 77.485 ;
        RECT 14.250 77.155 14.445 77.485 ;
        RECT 14.615 78.115 15.740 78.285 ;
        RECT 13.855 76.985 14.025 77.155 ;
        RECT 14.615 76.985 14.785 78.115 ;
        RECT 6.985 76.245 12.330 76.790 ;
        RECT 13.430 76.415 13.685 76.985 ;
        RECT 13.855 76.815 14.785 76.985 ;
        RECT 14.955 77.775 15.965 77.945 ;
        RECT 14.955 76.975 15.125 77.775 ;
        RECT 14.610 76.780 14.785 76.815 ;
        RECT 13.855 76.245 14.185 76.645 ;
        RECT 14.610 76.415 15.140 76.780 ;
        RECT 15.330 76.755 15.605 77.575 ;
        RECT 15.325 76.585 15.605 76.755 ;
        RECT 15.330 76.415 15.605 76.585 ;
        RECT 15.775 76.415 15.965 77.775 ;
        RECT 16.135 77.790 16.305 78.455 ;
        RECT 16.475 78.035 16.645 78.795 ;
        RECT 16.880 78.035 17.395 78.445 ;
        RECT 16.135 77.600 16.885 77.790 ;
        RECT 17.055 77.225 17.395 78.035 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 19.405 77.655 19.675 78.625 ;
        RECT 19.885 77.995 20.165 78.795 ;
        RECT 20.335 78.285 21.990 78.575 ;
        RECT 20.400 77.945 21.990 78.115 ;
        RECT 20.400 77.825 20.570 77.945 ;
        RECT 19.845 77.655 20.570 77.825 ;
        RECT 16.165 77.055 17.395 77.225 ;
        RECT 16.145 76.245 16.655 76.780 ;
        RECT 16.875 76.450 17.120 77.055 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 19.405 76.920 19.575 77.655 ;
        RECT 19.845 77.485 20.015 77.655 ;
        RECT 19.745 77.155 20.015 77.485 ;
        RECT 20.185 77.155 20.590 77.485 ;
        RECT 20.760 77.155 21.470 77.775 ;
        RECT 21.670 77.655 21.990 77.945 ;
        RECT 22.165 77.655 22.505 78.625 ;
        RECT 22.675 77.655 22.845 78.795 ;
        RECT 23.115 77.995 23.365 78.795 ;
        RECT 24.010 77.825 24.340 78.625 ;
        RECT 24.640 77.995 24.970 78.795 ;
        RECT 25.140 77.825 25.470 78.625 ;
        RECT 23.035 77.655 25.470 77.825 ;
        RECT 25.845 77.705 27.055 78.795 ;
        RECT 19.845 76.985 20.015 77.155 ;
        RECT 19.405 76.575 19.675 76.920 ;
        RECT 19.845 76.815 21.455 76.985 ;
        RECT 21.640 76.915 21.990 77.485 ;
        RECT 22.165 77.095 22.340 77.655 ;
        RECT 23.035 77.405 23.205 77.655 ;
        RECT 22.510 77.235 23.205 77.405 ;
        RECT 23.380 77.235 23.800 77.435 ;
        RECT 23.970 77.235 24.300 77.435 ;
        RECT 24.470 77.235 24.800 77.435 ;
        RECT 22.165 77.045 22.395 77.095 ;
        RECT 19.865 76.245 20.245 76.645 ;
        RECT 20.415 76.465 20.585 76.815 ;
        RECT 20.755 76.245 21.085 76.645 ;
        RECT 21.285 76.465 21.455 76.815 ;
        RECT 21.655 76.245 21.985 76.745 ;
        RECT 22.165 76.415 22.505 77.045 ;
        RECT 22.675 76.245 22.925 77.045 ;
        RECT 23.115 76.895 24.340 77.065 ;
        RECT 23.115 76.415 23.445 76.895 ;
        RECT 23.615 76.245 23.840 76.705 ;
        RECT 24.010 76.415 24.340 76.895 ;
        RECT 24.970 77.025 25.140 77.655 ;
        RECT 25.325 77.235 25.675 77.485 ;
        RECT 24.970 76.415 25.470 77.025 ;
        RECT 25.845 76.995 26.365 77.535 ;
        RECT 26.535 77.165 27.055 77.705 ;
        RECT 27.225 77.655 27.495 78.625 ;
        RECT 27.705 77.995 27.985 78.795 ;
        RECT 28.155 78.285 29.810 78.575 ;
        RECT 28.220 77.945 29.810 78.115 ;
        RECT 28.220 77.825 28.390 77.945 ;
        RECT 27.665 77.655 28.390 77.825 ;
        RECT 25.845 76.245 27.055 76.995 ;
        RECT 27.225 76.920 27.395 77.655 ;
        RECT 27.665 77.485 27.835 77.655 ;
        RECT 27.565 77.155 27.835 77.485 ;
        RECT 28.005 77.155 28.410 77.485 ;
        RECT 28.580 77.155 29.290 77.775 ;
        RECT 29.490 77.655 29.810 77.945 ;
        RECT 29.985 77.705 33.495 78.795 ;
        RECT 33.665 77.705 34.875 78.795 ;
        RECT 35.050 78.125 35.305 78.625 ;
        RECT 35.475 78.295 35.805 78.795 ;
        RECT 35.050 77.955 35.800 78.125 ;
        RECT 27.665 76.985 27.835 77.155 ;
        RECT 27.225 76.575 27.495 76.920 ;
        RECT 27.665 76.815 29.275 76.985 ;
        RECT 29.460 76.915 29.810 77.485 ;
        RECT 29.985 77.015 31.635 77.535 ;
        RECT 31.805 77.185 33.495 77.705 ;
        RECT 27.685 76.245 28.065 76.645 ;
        RECT 28.235 76.465 28.405 76.815 ;
        RECT 28.575 76.245 28.905 76.645 ;
        RECT 29.105 76.465 29.275 76.815 ;
        RECT 29.475 76.245 29.805 76.745 ;
        RECT 29.985 76.245 33.495 77.015 ;
        RECT 33.665 76.995 34.185 77.535 ;
        RECT 34.355 77.165 34.875 77.705 ;
        RECT 35.050 77.135 35.400 77.785 ;
        RECT 33.665 76.245 34.875 76.995 ;
        RECT 35.570 76.965 35.800 77.955 ;
        RECT 35.050 76.795 35.800 76.965 ;
        RECT 35.050 76.505 35.305 76.795 ;
        RECT 35.475 76.245 35.805 76.625 ;
        RECT 35.975 76.505 36.145 78.625 ;
        RECT 36.315 77.825 36.640 78.610 ;
        RECT 36.810 78.335 37.060 78.795 ;
        RECT 37.230 78.295 37.480 78.625 ;
        RECT 37.695 78.295 38.375 78.625 ;
        RECT 37.230 78.165 37.400 78.295 ;
        RECT 37.005 77.995 37.400 78.165 ;
        RECT 36.375 76.775 36.835 77.825 ;
        RECT 37.005 76.635 37.175 77.995 ;
        RECT 37.570 77.735 38.035 78.125 ;
        RECT 37.345 76.925 37.695 77.545 ;
        RECT 37.865 77.145 38.035 77.735 ;
        RECT 38.205 77.515 38.375 78.295 ;
        RECT 38.545 78.195 38.715 78.535 ;
        RECT 38.950 78.365 39.280 78.795 ;
        RECT 39.450 78.195 39.620 78.535 ;
        RECT 39.915 78.335 40.285 78.795 ;
        RECT 38.545 78.025 39.620 78.195 ;
        RECT 40.455 78.165 40.625 78.625 ;
        RECT 40.860 78.285 41.730 78.625 ;
        RECT 41.900 78.335 42.150 78.795 ;
        RECT 40.065 77.995 40.625 78.165 ;
        RECT 40.065 77.855 40.235 77.995 ;
        RECT 38.735 77.685 40.235 77.855 ;
        RECT 40.930 77.825 41.390 78.115 ;
        RECT 38.205 77.345 39.895 77.515 ;
        RECT 37.865 76.925 38.220 77.145 ;
        RECT 38.390 76.635 38.560 77.345 ;
        RECT 38.765 76.925 39.555 77.175 ;
        RECT 39.725 77.165 39.895 77.345 ;
        RECT 40.065 76.995 40.235 77.685 ;
        RECT 36.505 76.245 36.835 76.605 ;
        RECT 37.005 76.465 37.500 76.635 ;
        RECT 37.705 76.465 38.560 76.635 ;
        RECT 39.435 76.245 39.765 76.705 ;
        RECT 39.975 76.605 40.235 76.995 ;
        RECT 40.425 77.815 41.390 77.825 ;
        RECT 41.560 77.905 41.730 78.285 ;
        RECT 42.320 78.245 42.490 78.535 ;
        RECT 42.670 78.415 43.000 78.795 ;
        RECT 42.320 78.075 43.120 78.245 ;
        RECT 40.425 77.655 41.100 77.815 ;
        RECT 41.560 77.735 42.780 77.905 ;
        RECT 40.425 76.865 40.635 77.655 ;
        RECT 41.560 77.645 41.730 77.735 ;
        RECT 40.805 76.865 41.155 77.485 ;
        RECT 41.325 77.475 41.730 77.645 ;
        RECT 41.325 76.695 41.495 77.475 ;
        RECT 41.665 77.025 41.885 77.305 ;
        RECT 42.065 77.195 42.605 77.565 ;
        RECT 42.950 77.485 43.120 78.075 ;
        RECT 43.340 77.655 43.645 78.795 ;
        RECT 43.815 77.605 44.070 78.485 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.745 77.655 44.975 78.795 ;
        RECT 45.145 77.645 45.475 78.625 ;
        RECT 45.645 77.655 45.855 78.795 ;
        RECT 46.085 78.360 51.430 78.795 ;
        RECT 51.605 78.360 56.950 78.795 ;
        RECT 57.125 78.360 62.470 78.795 ;
        RECT 42.950 77.455 43.690 77.485 ;
        RECT 41.665 76.855 42.195 77.025 ;
        RECT 39.975 76.435 40.325 76.605 ;
        RECT 40.545 76.415 41.495 76.695 ;
        RECT 41.665 76.245 41.855 76.685 ;
        RECT 42.025 76.625 42.195 76.855 ;
        RECT 42.365 76.795 42.605 77.195 ;
        RECT 42.775 77.155 43.690 77.455 ;
        RECT 42.775 76.980 43.100 77.155 ;
        RECT 42.775 76.625 43.095 76.980 ;
        RECT 43.860 76.955 44.070 77.605 ;
        RECT 44.725 77.235 45.055 77.485 ;
        RECT 42.025 76.455 43.095 76.625 ;
        RECT 43.340 76.245 43.645 76.705 ;
        RECT 43.815 76.425 44.070 76.955 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 44.745 76.245 44.975 77.065 ;
        RECT 45.225 77.045 45.475 77.645 ;
        RECT 45.145 76.415 45.475 77.045 ;
        RECT 45.645 76.245 45.855 77.065 ;
        RECT 47.670 76.790 48.010 77.620 ;
        RECT 49.490 77.110 49.840 78.360 ;
        RECT 53.190 76.790 53.530 77.620 ;
        RECT 55.010 77.110 55.360 78.360 ;
        RECT 58.710 76.790 59.050 77.620 ;
        RECT 60.530 77.110 60.880 78.360 ;
        RECT 62.645 77.705 65.235 78.795 ;
        RECT 62.645 77.015 63.855 77.535 ;
        RECT 64.025 77.185 65.235 77.705 ;
        RECT 65.410 77.645 65.670 78.795 ;
        RECT 65.845 77.720 66.100 78.625 ;
        RECT 66.270 78.035 66.600 78.795 ;
        RECT 66.815 77.865 66.985 78.625 ;
        RECT 46.085 76.245 51.430 76.790 ;
        RECT 51.605 76.245 56.950 76.790 ;
        RECT 57.125 76.245 62.470 76.790 ;
        RECT 62.645 76.245 65.235 77.015 ;
        RECT 65.410 76.245 65.670 77.085 ;
        RECT 65.845 76.990 66.015 77.720 ;
        RECT 66.270 77.695 66.985 77.865 ;
        RECT 67.245 77.705 69.835 78.795 ;
        RECT 66.270 77.485 66.440 77.695 ;
        RECT 66.185 77.155 66.440 77.485 ;
        RECT 65.845 76.415 66.100 76.990 ;
        RECT 66.270 76.965 66.440 77.155 ;
        RECT 66.720 77.145 67.075 77.515 ;
        RECT 67.245 77.015 68.455 77.535 ;
        RECT 68.625 77.185 69.835 77.705 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.670 77.825 71.000 78.625 ;
        RECT 71.170 77.995 71.500 78.795 ;
        RECT 71.800 77.825 72.130 78.625 ;
        RECT 72.775 77.995 73.025 78.795 ;
        RECT 70.670 77.655 73.105 77.825 ;
        RECT 73.295 77.655 73.465 78.795 ;
        RECT 73.635 77.655 73.975 78.625 ;
        RECT 74.145 77.705 75.815 78.795 ;
        RECT 76.075 78.125 76.245 78.625 ;
        RECT 76.415 78.295 76.745 78.795 ;
        RECT 76.075 77.955 76.740 78.125 ;
        RECT 70.465 77.235 70.815 77.485 ;
        RECT 71.000 77.025 71.170 77.655 ;
        RECT 71.340 77.235 71.670 77.435 ;
        RECT 71.840 77.235 72.170 77.435 ;
        RECT 72.340 77.235 72.760 77.435 ;
        RECT 72.935 77.405 73.105 77.655 ;
        RECT 72.935 77.235 73.630 77.405 ;
        RECT 66.270 76.795 66.985 76.965 ;
        RECT 66.270 76.245 66.600 76.625 ;
        RECT 66.815 76.415 66.985 76.795 ;
        RECT 67.245 76.245 69.835 77.015 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 70.670 76.415 71.170 77.025 ;
        RECT 71.800 76.895 73.025 77.065 ;
        RECT 73.800 77.045 73.975 77.655 ;
        RECT 71.800 76.415 72.130 76.895 ;
        RECT 72.300 76.245 72.525 76.705 ;
        RECT 72.695 76.415 73.025 76.895 ;
        RECT 73.215 76.245 73.465 77.045 ;
        RECT 73.635 76.415 73.975 77.045 ;
        RECT 74.145 77.015 74.895 77.535 ;
        RECT 75.065 77.185 75.815 77.705 ;
        RECT 75.990 77.135 76.340 77.785 ;
        RECT 74.145 76.245 75.815 77.015 ;
        RECT 76.510 76.965 76.740 77.955 ;
        RECT 76.075 76.795 76.740 76.965 ;
        RECT 76.075 76.505 76.245 76.795 ;
        RECT 76.415 76.245 76.745 76.625 ;
        RECT 76.915 76.505 77.140 78.625 ;
        RECT 77.355 78.295 77.685 78.795 ;
        RECT 77.855 78.125 78.025 78.625 ;
        RECT 78.260 78.410 79.090 78.580 ;
        RECT 79.330 78.415 79.710 78.795 ;
        RECT 77.330 77.955 78.025 78.125 ;
        RECT 77.330 76.985 77.500 77.955 ;
        RECT 77.670 77.165 78.080 77.785 ;
        RECT 78.250 77.735 78.750 78.115 ;
        RECT 77.330 76.795 78.025 76.985 ;
        RECT 78.250 76.865 78.470 77.735 ;
        RECT 78.920 77.565 79.090 78.410 ;
        RECT 79.890 78.245 80.060 78.535 ;
        RECT 80.230 78.415 80.560 78.795 ;
        RECT 81.030 78.325 81.660 78.575 ;
        RECT 81.840 78.415 82.260 78.795 ;
        RECT 81.490 78.245 81.660 78.325 ;
        RECT 82.460 78.245 82.700 78.535 ;
        RECT 79.260 77.995 80.630 78.245 ;
        RECT 79.260 77.735 79.510 77.995 ;
        RECT 80.020 77.565 80.270 77.725 ;
        RECT 78.920 77.395 80.270 77.565 ;
        RECT 78.920 77.355 79.340 77.395 ;
        RECT 78.650 76.805 79.000 77.175 ;
        RECT 77.355 76.245 77.685 76.625 ;
        RECT 77.855 76.465 78.025 76.795 ;
        RECT 79.170 76.625 79.340 77.355 ;
        RECT 80.440 77.225 80.630 77.995 ;
        RECT 79.510 76.895 79.920 77.225 ;
        RECT 80.210 76.885 80.630 77.225 ;
        RECT 80.800 77.815 81.320 78.125 ;
        RECT 81.490 78.075 82.700 78.245 ;
        RECT 82.930 78.105 83.260 78.795 ;
        RECT 80.800 77.055 80.970 77.815 ;
        RECT 81.140 77.225 81.320 77.635 ;
        RECT 81.490 77.565 81.660 78.075 ;
        RECT 83.430 77.925 83.600 78.535 ;
        RECT 83.870 78.075 84.200 78.585 ;
        RECT 83.430 77.905 83.750 77.925 ;
        RECT 81.830 77.735 83.750 77.905 ;
        RECT 81.490 77.395 83.390 77.565 ;
        RECT 81.720 77.055 82.050 77.175 ;
        RECT 80.800 76.885 82.050 77.055 ;
        RECT 78.325 76.425 79.340 76.625 ;
        RECT 79.510 76.245 79.920 76.685 ;
        RECT 80.210 76.455 80.460 76.885 ;
        RECT 80.660 76.245 80.980 76.705 ;
        RECT 82.220 76.635 82.390 77.395 ;
        RECT 83.060 77.335 83.390 77.395 ;
        RECT 82.580 77.165 82.910 77.225 ;
        RECT 82.580 76.895 83.240 77.165 ;
        RECT 83.560 76.840 83.750 77.735 ;
        RECT 81.540 76.465 82.390 76.635 ;
        RECT 82.590 76.245 83.250 76.725 ;
        RECT 83.430 76.510 83.750 76.840 ;
        RECT 83.950 77.485 84.200 78.075 ;
        RECT 84.380 77.995 84.665 78.795 ;
        RECT 84.845 78.115 85.100 78.485 ;
        RECT 84.845 77.945 85.185 78.115 ;
        RECT 84.845 77.815 85.100 77.945 ;
        RECT 83.950 77.155 84.750 77.485 ;
        RECT 83.950 76.505 84.200 77.155 ;
        RECT 84.920 76.955 85.100 77.815 ;
        RECT 84.380 76.245 84.665 76.705 ;
        RECT 84.845 76.425 85.100 76.955 ;
        RECT 85.650 77.655 85.985 78.625 ;
        RECT 86.155 77.655 86.325 78.795 ;
        RECT 86.495 78.455 88.525 78.625 ;
        RECT 85.650 76.985 85.820 77.655 ;
        RECT 86.495 77.485 86.665 78.455 ;
        RECT 85.990 77.155 86.245 77.485 ;
        RECT 86.470 77.155 86.665 77.485 ;
        RECT 86.835 78.115 87.960 78.285 ;
        RECT 86.075 76.985 86.245 77.155 ;
        RECT 86.835 76.985 87.005 78.115 ;
        RECT 85.650 76.415 85.905 76.985 ;
        RECT 86.075 76.815 87.005 76.985 ;
        RECT 87.175 77.775 88.185 77.945 ;
        RECT 87.175 76.975 87.345 77.775 ;
        RECT 86.830 76.780 87.005 76.815 ;
        RECT 86.075 76.245 86.405 76.645 ;
        RECT 86.830 76.415 87.360 76.780 ;
        RECT 87.550 76.755 87.825 77.575 ;
        RECT 87.545 76.585 87.825 76.755 ;
        RECT 87.550 76.415 87.825 76.585 ;
        RECT 87.995 76.415 88.185 77.775 ;
        RECT 88.355 77.790 88.525 78.455 ;
        RECT 88.695 78.035 88.865 78.795 ;
        RECT 89.100 78.035 89.615 78.445 ;
        RECT 89.785 78.360 95.130 78.795 ;
        RECT 88.355 77.600 89.105 77.790 ;
        RECT 89.275 77.225 89.615 78.035 ;
        RECT 88.385 77.055 89.615 77.225 ;
        RECT 88.365 76.245 88.875 76.780 ;
        RECT 89.095 76.450 89.340 77.055 ;
        RECT 91.370 76.790 91.710 77.620 ;
        RECT 93.190 77.110 93.540 78.360 ;
        RECT 95.765 77.630 96.055 78.795 ;
        RECT 96.225 78.360 101.570 78.795 ;
        RECT 101.745 78.360 107.090 78.795 ;
        RECT 89.785 76.245 95.130 76.790 ;
        RECT 95.765 76.245 96.055 76.970 ;
        RECT 97.810 76.790 98.150 77.620 ;
        RECT 99.630 77.110 99.980 78.360 ;
        RECT 103.330 76.790 103.670 77.620 ;
        RECT 105.150 77.110 105.500 78.360 ;
        RECT 107.265 77.705 108.935 78.795 ;
        RECT 107.265 77.015 108.015 77.535 ;
        RECT 108.185 77.185 108.935 77.705 ;
        RECT 109.655 77.865 109.825 78.625 ;
        RECT 110.005 78.035 110.335 78.795 ;
        RECT 109.655 77.695 110.320 77.865 ;
        RECT 110.505 77.720 110.775 78.625 ;
        RECT 111.035 78.125 111.205 78.625 ;
        RECT 111.375 78.295 111.705 78.795 ;
        RECT 111.035 77.955 111.700 78.125 ;
        RECT 110.150 77.550 110.320 77.695 ;
        RECT 109.585 77.145 109.915 77.515 ;
        RECT 110.150 77.220 110.435 77.550 ;
        RECT 96.225 76.245 101.570 76.790 ;
        RECT 101.745 76.245 107.090 76.790 ;
        RECT 107.265 76.245 108.935 77.015 ;
        RECT 110.150 76.965 110.320 77.220 ;
        RECT 109.655 76.795 110.320 76.965 ;
        RECT 110.605 76.920 110.775 77.720 ;
        RECT 110.950 77.135 111.300 77.785 ;
        RECT 111.470 76.965 111.700 77.955 ;
        RECT 109.655 76.415 109.825 76.795 ;
        RECT 110.005 76.245 110.335 76.625 ;
        RECT 110.515 76.415 110.775 76.920 ;
        RECT 111.035 76.795 111.700 76.965 ;
        RECT 111.035 76.505 111.205 76.795 ;
        RECT 111.375 76.245 111.705 76.625 ;
        RECT 111.875 76.505 112.100 78.625 ;
        RECT 112.315 78.295 112.645 78.795 ;
        RECT 112.815 78.125 112.985 78.625 ;
        RECT 113.220 78.410 114.050 78.580 ;
        RECT 114.290 78.415 114.670 78.795 ;
        RECT 112.290 77.955 112.985 78.125 ;
        RECT 112.290 76.985 112.460 77.955 ;
        RECT 112.630 77.165 113.040 77.785 ;
        RECT 113.210 77.735 113.710 78.115 ;
        RECT 112.290 76.795 112.985 76.985 ;
        RECT 113.210 76.865 113.430 77.735 ;
        RECT 113.880 77.565 114.050 78.410 ;
        RECT 114.850 78.245 115.020 78.535 ;
        RECT 115.190 78.415 115.520 78.795 ;
        RECT 115.990 78.325 116.620 78.575 ;
        RECT 116.800 78.415 117.220 78.795 ;
        RECT 116.450 78.245 116.620 78.325 ;
        RECT 117.420 78.245 117.660 78.535 ;
        RECT 114.220 77.995 115.590 78.245 ;
        RECT 114.220 77.735 114.470 77.995 ;
        RECT 114.980 77.565 115.230 77.725 ;
        RECT 113.880 77.395 115.230 77.565 ;
        RECT 113.880 77.355 114.300 77.395 ;
        RECT 113.610 76.805 113.960 77.175 ;
        RECT 112.315 76.245 112.645 76.625 ;
        RECT 112.815 76.465 112.985 76.795 ;
        RECT 114.130 76.625 114.300 77.355 ;
        RECT 115.400 77.225 115.590 77.995 ;
        RECT 114.470 76.895 114.880 77.225 ;
        RECT 115.170 76.885 115.590 77.225 ;
        RECT 115.760 77.815 116.280 78.125 ;
        RECT 116.450 78.075 117.660 78.245 ;
        RECT 117.890 78.105 118.220 78.795 ;
        RECT 115.760 77.055 115.930 77.815 ;
        RECT 116.100 77.225 116.280 77.635 ;
        RECT 116.450 77.565 116.620 78.075 ;
        RECT 118.390 77.925 118.560 78.535 ;
        RECT 118.830 78.075 119.160 78.585 ;
        RECT 118.390 77.905 118.710 77.925 ;
        RECT 116.790 77.735 118.710 77.905 ;
        RECT 116.450 77.395 118.350 77.565 ;
        RECT 116.680 77.055 117.010 77.175 ;
        RECT 115.760 76.885 117.010 77.055 ;
        RECT 113.285 76.425 114.300 76.625 ;
        RECT 114.470 76.245 114.880 76.685 ;
        RECT 115.170 76.455 115.420 76.885 ;
        RECT 115.620 76.245 115.940 76.705 ;
        RECT 117.180 76.635 117.350 77.395 ;
        RECT 118.020 77.335 118.350 77.395 ;
        RECT 117.540 77.165 117.870 77.225 ;
        RECT 117.540 76.895 118.200 77.165 ;
        RECT 118.520 76.840 118.710 77.735 ;
        RECT 116.500 76.465 117.350 76.635 ;
        RECT 117.550 76.245 118.210 76.725 ;
        RECT 118.390 76.510 118.710 76.840 ;
        RECT 118.910 77.485 119.160 78.075 ;
        RECT 119.340 77.995 119.625 78.795 ;
        RECT 119.805 77.815 120.060 78.485 ;
        RECT 118.910 77.155 119.710 77.485 ;
        RECT 118.910 76.505 119.160 77.155 ;
        RECT 119.880 76.955 120.060 77.815 ;
        RECT 121.525 77.630 121.815 78.795 ;
        RECT 122.445 77.705 123.655 78.795 ;
        RECT 122.445 77.165 122.965 77.705 ;
        RECT 123.135 76.995 123.655 77.535 ;
        RECT 119.805 76.755 120.060 76.955 ;
        RECT 119.340 76.245 119.625 76.705 ;
        RECT 119.805 76.585 120.145 76.755 ;
        RECT 119.805 76.425 120.060 76.585 ;
        RECT 121.525 76.245 121.815 76.970 ;
        RECT 122.445 76.245 123.655 76.995 ;
        RECT 5.520 76.075 123.740 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 6.985 75.305 9.575 76.075 ;
        RECT 10.205 75.400 10.465 75.905 ;
        RECT 10.645 75.695 10.975 76.075 ;
        RECT 11.155 75.525 11.325 75.905 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 6.985 74.785 8.195 75.305 ;
        RECT 8.365 74.615 9.575 75.135 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 6.985 73.525 9.575 74.615 ;
        RECT 10.205 74.600 10.375 75.400 ;
        RECT 10.660 75.355 11.325 75.525 ;
        RECT 11.585 75.400 11.845 75.905 ;
        RECT 12.025 75.695 12.355 76.075 ;
        RECT 12.535 75.525 12.705 75.905 ;
        RECT 10.660 75.100 10.830 75.355 ;
        RECT 10.545 74.770 10.830 75.100 ;
        RECT 11.065 74.805 11.395 75.175 ;
        RECT 10.660 74.625 10.830 74.770 ;
        RECT 10.205 73.695 10.475 74.600 ;
        RECT 10.660 74.455 11.325 74.625 ;
        RECT 10.645 73.525 10.975 74.285 ;
        RECT 11.155 73.695 11.325 74.455 ;
        RECT 11.585 74.600 11.755 75.400 ;
        RECT 12.040 75.355 12.705 75.525 ;
        RECT 12.040 75.100 12.210 75.355 ;
        RECT 13.025 75.255 13.235 76.075 ;
        RECT 13.405 75.275 13.735 75.905 ;
        RECT 11.925 74.770 12.210 75.100 ;
        RECT 12.445 74.805 12.775 75.175 ;
        RECT 12.040 74.625 12.210 74.770 ;
        RECT 13.405 74.675 13.655 75.275 ;
        RECT 13.905 75.255 14.135 76.075 ;
        RECT 14.810 75.335 15.065 75.905 ;
        RECT 15.235 75.675 15.565 76.075 ;
        RECT 15.990 75.540 16.520 75.905 ;
        RECT 15.990 75.505 16.165 75.540 ;
        RECT 15.235 75.335 16.165 75.505 ;
        RECT 16.710 75.395 16.985 75.905 ;
        RECT 13.825 74.835 14.155 75.085 ;
        RECT 11.585 73.695 11.855 74.600 ;
        RECT 12.040 74.455 12.705 74.625 ;
        RECT 12.025 73.525 12.355 74.285 ;
        RECT 12.535 73.695 12.705 74.455 ;
        RECT 13.025 73.525 13.235 74.665 ;
        RECT 13.405 73.695 13.735 74.675 ;
        RECT 14.810 74.665 14.980 75.335 ;
        RECT 15.235 75.165 15.405 75.335 ;
        RECT 15.150 74.835 15.405 75.165 ;
        RECT 15.630 74.835 15.825 75.165 ;
        RECT 13.905 73.525 14.135 74.665 ;
        RECT 14.810 73.695 15.145 74.665 ;
        RECT 15.315 73.525 15.485 74.665 ;
        RECT 15.655 73.865 15.825 74.835 ;
        RECT 15.995 74.205 16.165 75.335 ;
        RECT 16.335 74.545 16.505 75.345 ;
        RECT 16.705 75.225 16.985 75.395 ;
        RECT 16.710 74.745 16.985 75.225 ;
        RECT 17.155 74.545 17.345 75.905 ;
        RECT 17.525 75.540 18.035 76.075 ;
        RECT 18.255 75.265 18.500 75.870 ;
        RECT 18.945 75.305 22.455 76.075 ;
        RECT 17.545 75.095 18.775 75.265 ;
        RECT 16.335 74.375 17.345 74.545 ;
        RECT 17.515 74.530 18.265 74.720 ;
        RECT 15.995 74.035 17.120 74.205 ;
        RECT 17.515 73.865 17.685 74.530 ;
        RECT 18.435 74.285 18.775 75.095 ;
        RECT 18.945 74.785 20.595 75.305 ;
        RECT 23.085 75.275 23.425 75.905 ;
        RECT 23.595 75.275 23.845 76.075 ;
        RECT 24.035 75.425 24.365 75.905 ;
        RECT 24.535 75.615 24.760 76.075 ;
        RECT 24.930 75.425 25.260 75.905 ;
        RECT 20.765 74.615 22.455 75.135 ;
        RECT 15.655 73.695 17.685 73.865 ;
        RECT 17.855 73.525 18.025 74.285 ;
        RECT 18.260 73.875 18.775 74.285 ;
        RECT 18.945 73.525 22.455 74.615 ;
        RECT 23.085 74.665 23.260 75.275 ;
        RECT 24.035 75.255 25.260 75.425 ;
        RECT 25.890 75.295 26.390 75.905 ;
        RECT 23.430 74.915 24.125 75.085 ;
        RECT 23.955 74.665 24.125 74.915 ;
        RECT 24.300 74.885 24.720 75.085 ;
        RECT 24.890 74.885 25.220 75.085 ;
        RECT 25.390 74.885 25.720 75.085 ;
        RECT 25.890 74.665 26.060 75.295 ;
        RECT 26.765 75.275 27.105 75.905 ;
        RECT 27.275 75.275 27.525 76.075 ;
        RECT 27.715 75.425 28.045 75.905 ;
        RECT 28.215 75.615 28.440 76.075 ;
        RECT 28.610 75.425 28.940 75.905 ;
        RECT 26.245 74.835 26.595 75.085 ;
        RECT 26.765 74.665 26.940 75.275 ;
        RECT 27.715 75.255 28.940 75.425 ;
        RECT 29.570 75.295 30.070 75.905 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 31.825 75.530 37.170 76.075 ;
        RECT 27.110 74.915 27.805 75.085 ;
        RECT 27.635 74.665 27.805 74.915 ;
        RECT 27.980 74.885 28.400 75.085 ;
        RECT 28.570 74.885 28.900 75.085 ;
        RECT 29.070 74.885 29.400 75.085 ;
        RECT 29.570 74.665 29.740 75.295 ;
        RECT 29.925 74.835 30.275 75.085 ;
        RECT 33.410 74.700 33.750 75.530 ;
        RECT 37.345 75.305 39.015 76.075 ;
        RECT 23.085 73.695 23.425 74.665 ;
        RECT 23.595 73.525 23.765 74.665 ;
        RECT 23.955 74.495 26.390 74.665 ;
        RECT 24.035 73.525 24.285 74.325 ;
        RECT 24.930 73.695 25.260 74.495 ;
        RECT 25.560 73.525 25.890 74.325 ;
        RECT 26.060 73.695 26.390 74.495 ;
        RECT 26.765 73.695 27.105 74.665 ;
        RECT 27.275 73.525 27.445 74.665 ;
        RECT 27.635 74.495 30.070 74.665 ;
        RECT 27.715 73.525 27.965 74.325 ;
        RECT 28.610 73.695 28.940 74.495 ;
        RECT 29.240 73.525 29.570 74.325 ;
        RECT 29.740 73.695 30.070 74.495 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 35.230 73.960 35.580 75.210 ;
        RECT 37.345 74.785 38.095 75.305 ;
        RECT 39.685 75.255 39.915 76.075 ;
        RECT 40.085 75.275 40.415 75.905 ;
        RECT 38.265 74.615 39.015 75.135 ;
        RECT 39.665 74.835 39.995 75.085 ;
        RECT 40.165 74.675 40.415 75.275 ;
        RECT 40.585 75.255 40.795 76.075 ;
        RECT 41.025 75.530 46.370 76.075 ;
        RECT 46.545 75.530 51.890 76.075 ;
        RECT 42.610 74.700 42.950 75.530 ;
        RECT 31.825 73.525 37.170 73.960 ;
        RECT 37.345 73.525 39.015 74.615 ;
        RECT 39.685 73.525 39.915 74.665 ;
        RECT 40.085 73.695 40.415 74.675 ;
        RECT 40.585 73.525 40.795 74.665 ;
        RECT 44.430 73.960 44.780 75.210 ;
        RECT 48.130 74.700 48.470 75.530 ;
        RECT 53.190 75.295 53.690 75.905 ;
        RECT 49.950 73.960 50.300 75.210 ;
        RECT 52.985 74.835 53.335 75.085 ;
        RECT 53.520 74.665 53.690 75.295 ;
        RECT 54.320 75.425 54.650 75.905 ;
        RECT 54.820 75.615 55.045 76.075 ;
        RECT 55.215 75.425 55.545 75.905 ;
        RECT 54.320 75.255 55.545 75.425 ;
        RECT 55.735 75.275 55.985 76.075 ;
        RECT 56.155 75.275 56.495 75.905 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 57.645 75.595 57.925 76.075 ;
        RECT 58.095 75.425 58.355 75.815 ;
        RECT 58.530 75.595 58.785 76.075 ;
        RECT 58.955 75.425 59.250 75.815 ;
        RECT 59.430 75.595 59.705 76.075 ;
        RECT 59.875 75.575 60.175 75.905 ;
        RECT 53.860 74.885 54.190 75.085 ;
        RECT 54.360 74.885 54.690 75.085 ;
        RECT 54.860 74.885 55.280 75.085 ;
        RECT 55.455 74.915 56.150 75.085 ;
        RECT 55.455 74.665 55.625 74.915 ;
        RECT 56.320 74.665 56.495 75.275 ;
        RECT 57.600 75.255 59.250 75.425 ;
        RECT 57.600 74.745 58.005 75.255 ;
        RECT 58.175 74.915 59.315 75.085 ;
        RECT 53.190 74.495 55.625 74.665 ;
        RECT 41.025 73.525 46.370 73.960 ;
        RECT 46.545 73.525 51.890 73.960 ;
        RECT 53.190 73.695 53.520 74.495 ;
        RECT 53.690 73.525 54.020 74.325 ;
        RECT 54.320 73.695 54.650 74.495 ;
        RECT 55.295 73.525 55.545 74.325 ;
        RECT 55.815 73.525 55.985 74.665 ;
        RECT 56.155 73.695 56.495 74.665 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 57.600 74.575 58.355 74.745 ;
        RECT 57.640 73.525 57.925 74.395 ;
        RECT 58.095 74.325 58.355 74.575 ;
        RECT 59.145 74.665 59.315 74.915 ;
        RECT 59.485 74.835 59.835 75.405 ;
        RECT 60.005 74.665 60.175 75.575 ;
        RECT 60.345 75.305 62.015 76.075 ;
        RECT 60.345 74.785 61.095 75.305 ;
        RECT 62.190 75.235 62.450 76.075 ;
        RECT 62.625 75.330 62.880 75.905 ;
        RECT 63.050 75.695 63.380 76.075 ;
        RECT 63.595 75.525 63.765 75.905 ;
        RECT 64.025 75.565 64.330 76.075 ;
        RECT 63.050 75.355 63.765 75.525 ;
        RECT 59.145 74.495 60.175 74.665 ;
        RECT 61.265 74.615 62.015 75.135 ;
        RECT 58.095 74.155 59.215 74.325 ;
        RECT 58.095 73.695 58.355 74.155 ;
        RECT 58.530 73.525 58.785 73.985 ;
        RECT 58.955 73.695 59.215 74.155 ;
        RECT 59.385 73.525 59.695 74.325 ;
        RECT 59.865 73.695 60.175 74.495 ;
        RECT 60.345 73.525 62.015 74.615 ;
        RECT 62.190 73.525 62.450 74.675 ;
        RECT 62.625 74.600 62.795 75.330 ;
        RECT 63.050 75.165 63.220 75.355 ;
        RECT 62.965 74.835 63.220 75.165 ;
        RECT 63.050 74.625 63.220 74.835 ;
        RECT 63.500 74.805 63.855 75.175 ;
        RECT 64.025 74.835 64.340 75.395 ;
        RECT 64.510 75.085 64.760 75.895 ;
        RECT 64.930 75.550 65.190 76.075 ;
        RECT 65.370 75.085 65.620 75.895 ;
        RECT 65.790 75.515 66.050 76.075 ;
        RECT 66.220 75.425 66.480 75.880 ;
        RECT 66.650 75.595 66.910 76.075 ;
        RECT 67.080 75.425 67.340 75.880 ;
        RECT 67.510 75.595 67.770 76.075 ;
        RECT 67.940 75.425 68.200 75.880 ;
        RECT 68.370 75.595 68.615 76.075 ;
        RECT 68.785 75.425 69.060 75.880 ;
        RECT 69.230 75.595 69.475 76.075 ;
        RECT 69.645 75.425 69.905 75.880 ;
        RECT 70.085 75.595 70.335 76.075 ;
        RECT 70.505 75.425 70.765 75.880 ;
        RECT 70.945 75.595 71.195 76.075 ;
        RECT 71.365 75.425 71.625 75.880 ;
        RECT 71.805 75.595 72.065 76.075 ;
        RECT 72.235 75.425 72.495 75.880 ;
        RECT 72.665 75.595 72.965 76.075 ;
        RECT 73.225 75.530 78.570 76.075 ;
        RECT 66.220 75.255 72.965 75.425 ;
        RECT 64.510 74.835 71.630 75.085 ;
        RECT 62.625 73.695 62.880 74.600 ;
        RECT 63.050 74.455 63.765 74.625 ;
        RECT 63.050 73.525 63.380 74.285 ;
        RECT 63.595 73.695 63.765 74.455 ;
        RECT 64.035 73.525 64.330 74.335 ;
        RECT 64.510 73.695 64.755 74.835 ;
        RECT 64.930 73.525 65.190 74.335 ;
        RECT 65.370 73.700 65.620 74.835 ;
        RECT 71.800 74.665 72.965 75.255 ;
        RECT 74.810 74.700 75.150 75.530 ;
        RECT 79.410 75.295 79.910 75.905 ;
        RECT 66.220 74.440 72.965 74.665 ;
        RECT 66.220 74.425 71.625 74.440 ;
        RECT 65.790 73.530 66.050 74.325 ;
        RECT 66.220 73.700 66.480 74.425 ;
        RECT 66.650 73.530 66.910 74.255 ;
        RECT 67.080 73.700 67.340 74.425 ;
        RECT 67.510 73.530 67.770 74.255 ;
        RECT 67.940 73.700 68.200 74.425 ;
        RECT 68.370 73.530 68.630 74.255 ;
        RECT 68.800 73.700 69.060 74.425 ;
        RECT 69.230 73.530 69.475 74.255 ;
        RECT 69.645 73.700 69.905 74.425 ;
        RECT 70.090 73.530 70.335 74.255 ;
        RECT 70.505 73.700 70.765 74.425 ;
        RECT 70.950 73.530 71.195 74.255 ;
        RECT 71.365 73.700 71.625 74.425 ;
        RECT 71.810 73.530 72.065 74.255 ;
        RECT 72.235 73.700 72.525 74.440 ;
        RECT 65.790 73.525 72.065 73.530 ;
        RECT 72.695 73.525 72.965 74.270 ;
        RECT 76.630 73.960 76.980 75.210 ;
        RECT 79.205 74.835 79.555 75.085 ;
        RECT 79.740 74.665 79.910 75.295 ;
        RECT 80.540 75.425 80.870 75.905 ;
        RECT 81.040 75.615 81.265 76.075 ;
        RECT 81.435 75.425 81.765 75.905 ;
        RECT 80.540 75.255 81.765 75.425 ;
        RECT 81.955 75.275 82.205 76.075 ;
        RECT 82.375 75.275 82.715 75.905 ;
        RECT 82.885 75.350 83.175 76.075 ;
        RECT 83.550 75.295 84.050 75.905 ;
        RECT 80.080 74.885 80.410 75.085 ;
        RECT 80.580 74.885 80.910 75.085 ;
        RECT 81.080 74.885 81.500 75.085 ;
        RECT 81.675 74.915 82.370 75.085 ;
        RECT 81.675 74.665 81.845 74.915 ;
        RECT 82.540 74.665 82.715 75.275 ;
        RECT 83.345 74.835 83.695 75.085 ;
        RECT 79.410 74.495 81.845 74.665 ;
        RECT 73.225 73.525 78.570 73.960 ;
        RECT 79.410 73.695 79.740 74.495 ;
        RECT 79.910 73.525 80.240 74.325 ;
        RECT 80.540 73.695 80.870 74.495 ;
        RECT 81.515 73.525 81.765 74.325 ;
        RECT 82.035 73.525 82.205 74.665 ;
        RECT 82.375 73.695 82.715 74.665 ;
        RECT 82.885 73.525 83.175 74.690 ;
        RECT 83.880 74.665 84.050 75.295 ;
        RECT 84.680 75.425 85.010 75.905 ;
        RECT 85.180 75.615 85.405 76.075 ;
        RECT 85.575 75.425 85.905 75.905 ;
        RECT 84.680 75.255 85.905 75.425 ;
        RECT 86.095 75.275 86.345 76.075 ;
        RECT 86.515 75.275 86.855 75.905 ;
        RECT 87.035 75.575 87.365 76.075 ;
        RECT 87.565 75.505 87.735 75.855 ;
        RECT 87.935 75.675 88.265 76.075 ;
        RECT 88.435 75.505 88.605 75.855 ;
        RECT 88.775 75.675 89.155 76.075 ;
        RECT 86.625 75.225 86.855 75.275 ;
        RECT 84.220 74.885 84.550 75.085 ;
        RECT 84.720 74.885 85.050 75.085 ;
        RECT 85.220 74.885 85.640 75.085 ;
        RECT 85.815 74.915 86.510 75.085 ;
        RECT 85.815 74.665 85.985 74.915 ;
        RECT 86.680 74.665 86.855 75.225 ;
        RECT 87.030 74.835 87.380 75.405 ;
        RECT 87.565 75.335 89.175 75.505 ;
        RECT 89.345 75.400 89.615 75.745 ;
        RECT 89.795 75.575 90.125 76.075 ;
        RECT 90.325 75.505 90.495 75.855 ;
        RECT 90.695 75.675 91.025 76.075 ;
        RECT 91.195 75.505 91.365 75.855 ;
        RECT 91.535 75.675 91.915 76.075 ;
        RECT 89.005 75.165 89.175 75.335 ;
        RECT 87.550 74.715 88.260 75.165 ;
        RECT 88.430 74.835 88.835 75.165 ;
        RECT 89.005 74.835 89.275 75.165 ;
        RECT 83.550 74.495 85.985 74.665 ;
        RECT 83.550 73.695 83.880 74.495 ;
        RECT 84.050 73.525 84.380 74.325 ;
        RECT 84.680 73.695 85.010 74.495 ;
        RECT 85.655 73.525 85.905 74.325 ;
        RECT 86.175 73.525 86.345 74.665 ;
        RECT 86.515 73.695 86.855 74.665 ;
        RECT 87.030 74.375 87.350 74.665 ;
        RECT 87.545 74.545 88.260 74.715 ;
        RECT 89.005 74.665 89.175 74.835 ;
        RECT 89.445 74.665 89.615 75.400 ;
        RECT 89.790 74.835 90.140 75.405 ;
        RECT 90.325 75.335 91.935 75.505 ;
        RECT 92.105 75.400 92.375 75.745 ;
        RECT 91.765 75.165 91.935 75.335 ;
        RECT 88.450 74.495 89.175 74.665 ;
        RECT 88.450 74.375 88.620 74.495 ;
        RECT 87.030 74.205 88.620 74.375 ;
        RECT 87.030 73.745 88.685 74.035 ;
        RECT 88.855 73.525 89.135 74.325 ;
        RECT 89.345 73.695 89.615 74.665 ;
        RECT 89.790 74.375 90.110 74.665 ;
        RECT 90.310 74.545 91.020 75.165 ;
        RECT 91.190 74.835 91.595 75.165 ;
        RECT 91.765 74.835 92.035 75.165 ;
        RECT 91.765 74.665 91.935 74.835 ;
        RECT 92.205 74.665 92.375 75.400 ;
        RECT 92.545 75.325 93.755 76.075 ;
        RECT 92.545 74.785 93.065 75.325 ;
        RECT 93.925 75.275 94.265 75.905 ;
        RECT 94.435 75.275 94.685 76.075 ;
        RECT 94.875 75.425 95.205 75.905 ;
        RECT 95.375 75.615 95.600 76.075 ;
        RECT 95.770 75.425 96.100 75.905 ;
        RECT 91.210 74.495 91.935 74.665 ;
        RECT 91.210 74.375 91.380 74.495 ;
        RECT 89.790 74.205 91.380 74.375 ;
        RECT 89.790 73.745 91.445 74.035 ;
        RECT 91.615 73.525 91.895 74.325 ;
        RECT 92.105 73.695 92.375 74.665 ;
        RECT 93.235 74.615 93.755 75.155 ;
        RECT 92.545 73.525 93.755 74.615 ;
        RECT 93.925 74.665 94.100 75.275 ;
        RECT 94.875 75.255 96.100 75.425 ;
        RECT 96.730 75.295 97.230 75.905 ;
        RECT 94.270 74.915 94.965 75.085 ;
        RECT 94.795 74.665 94.965 74.915 ;
        RECT 95.140 74.885 95.560 75.085 ;
        RECT 95.730 74.885 96.060 75.085 ;
        RECT 96.230 74.885 96.560 75.085 ;
        RECT 96.730 74.665 96.900 75.295 ;
        RECT 97.605 75.275 97.945 75.905 ;
        RECT 98.115 75.275 98.365 76.075 ;
        RECT 98.555 75.425 98.885 75.905 ;
        RECT 99.055 75.615 99.280 76.075 ;
        RECT 99.450 75.425 99.780 75.905 ;
        RECT 97.085 74.835 97.435 75.085 ;
        RECT 97.605 74.665 97.780 75.275 ;
        RECT 98.555 75.255 99.780 75.425 ;
        RECT 100.410 75.295 100.910 75.905 ;
        RECT 101.285 75.400 101.545 75.905 ;
        RECT 101.725 75.695 102.055 76.075 ;
        RECT 102.235 75.525 102.405 75.905 ;
        RECT 102.665 75.530 108.010 76.075 ;
        RECT 97.950 74.915 98.645 75.085 ;
        RECT 98.475 74.665 98.645 74.915 ;
        RECT 98.820 74.885 99.240 75.085 ;
        RECT 99.410 74.885 99.740 75.085 ;
        RECT 99.910 74.885 100.240 75.085 ;
        RECT 100.410 74.665 100.580 75.295 ;
        RECT 100.765 74.835 101.115 75.085 ;
        RECT 93.925 73.695 94.265 74.665 ;
        RECT 94.435 73.525 94.605 74.665 ;
        RECT 94.795 74.495 97.230 74.665 ;
        RECT 94.875 73.525 95.125 74.325 ;
        RECT 95.770 73.695 96.100 74.495 ;
        RECT 96.400 73.525 96.730 74.325 ;
        RECT 96.900 73.695 97.230 74.495 ;
        RECT 97.605 73.695 97.945 74.665 ;
        RECT 98.115 73.525 98.285 74.665 ;
        RECT 98.475 74.495 100.910 74.665 ;
        RECT 98.555 73.525 98.805 74.325 ;
        RECT 99.450 73.695 99.780 74.495 ;
        RECT 100.080 73.525 100.410 74.325 ;
        RECT 100.580 73.695 100.910 74.495 ;
        RECT 101.285 74.600 101.455 75.400 ;
        RECT 101.740 75.355 102.405 75.525 ;
        RECT 101.740 75.100 101.910 75.355 ;
        RECT 101.625 74.770 101.910 75.100 ;
        RECT 102.145 74.805 102.475 75.175 ;
        RECT 101.740 74.625 101.910 74.770 ;
        RECT 104.250 74.700 104.590 75.530 ;
        RECT 108.645 75.350 108.935 76.075 ;
        RECT 109.105 75.305 111.695 76.075 ;
        RECT 112.330 75.335 112.585 75.905 ;
        RECT 112.755 75.675 113.085 76.075 ;
        RECT 113.510 75.540 114.040 75.905 ;
        RECT 113.510 75.505 113.685 75.540 ;
        RECT 112.755 75.335 113.685 75.505 ;
        RECT 101.285 73.695 101.555 74.600 ;
        RECT 101.740 74.455 102.405 74.625 ;
        RECT 101.725 73.525 102.055 74.285 ;
        RECT 102.235 73.695 102.405 74.455 ;
        RECT 106.070 73.960 106.420 75.210 ;
        RECT 109.105 74.785 110.315 75.305 ;
        RECT 102.665 73.525 108.010 73.960 ;
        RECT 108.645 73.525 108.935 74.690 ;
        RECT 110.485 74.615 111.695 75.135 ;
        RECT 109.105 73.525 111.695 74.615 ;
        RECT 112.330 74.665 112.500 75.335 ;
        RECT 112.755 75.165 112.925 75.335 ;
        RECT 112.670 74.835 112.925 75.165 ;
        RECT 113.150 74.835 113.345 75.165 ;
        RECT 112.330 73.695 112.665 74.665 ;
        RECT 112.835 73.525 113.005 74.665 ;
        RECT 113.175 73.865 113.345 74.835 ;
        RECT 113.515 74.205 113.685 75.335 ;
        RECT 113.855 74.545 114.025 75.345 ;
        RECT 114.230 75.055 114.505 75.905 ;
        RECT 114.225 74.885 114.505 75.055 ;
        RECT 114.230 74.745 114.505 74.885 ;
        RECT 114.675 74.545 114.865 75.905 ;
        RECT 115.045 75.540 115.555 76.075 ;
        RECT 115.775 75.265 116.020 75.870 ;
        RECT 116.465 75.530 121.810 76.075 ;
        RECT 115.065 75.095 116.295 75.265 ;
        RECT 113.855 74.375 114.865 74.545 ;
        RECT 115.035 74.530 115.785 74.720 ;
        RECT 113.515 74.035 114.640 74.205 ;
        RECT 115.035 73.865 115.205 74.530 ;
        RECT 115.955 74.285 116.295 75.095 ;
        RECT 118.050 74.700 118.390 75.530 ;
        RECT 122.445 75.325 123.655 76.075 ;
        RECT 113.175 73.695 115.205 73.865 ;
        RECT 115.375 73.525 115.545 74.285 ;
        RECT 115.780 73.875 116.295 74.285 ;
        RECT 119.870 73.960 120.220 75.210 ;
        RECT 122.445 74.615 122.965 75.155 ;
        RECT 123.135 74.785 123.655 75.325 ;
        RECT 116.465 73.525 121.810 73.960 ;
        RECT 122.445 73.525 123.655 74.615 ;
        RECT 5.520 73.355 123.740 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 7.535 72.685 7.705 73.185 ;
        RECT 7.875 72.855 8.205 73.355 ;
        RECT 7.535 72.515 8.200 72.685 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 7.450 71.695 7.800 72.345 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 7.970 71.525 8.200 72.515 ;
        RECT 7.535 71.355 8.200 71.525 ;
        RECT 7.535 71.065 7.705 71.355 ;
        RECT 7.875 70.805 8.205 71.185 ;
        RECT 8.375 71.065 8.600 73.185 ;
        RECT 8.815 72.855 9.145 73.355 ;
        RECT 9.315 72.685 9.485 73.185 ;
        RECT 9.720 72.970 10.550 73.140 ;
        RECT 10.790 72.975 11.170 73.355 ;
        RECT 8.790 72.515 9.485 72.685 ;
        RECT 8.790 71.545 8.960 72.515 ;
        RECT 9.130 71.725 9.540 72.345 ;
        RECT 9.710 72.295 10.210 72.675 ;
        RECT 8.790 71.355 9.485 71.545 ;
        RECT 9.710 71.425 9.930 72.295 ;
        RECT 10.380 72.125 10.550 72.970 ;
        RECT 11.350 72.805 11.520 73.095 ;
        RECT 11.690 72.975 12.020 73.355 ;
        RECT 12.490 72.885 13.120 73.135 ;
        RECT 13.300 72.975 13.720 73.355 ;
        RECT 12.950 72.805 13.120 72.885 ;
        RECT 13.920 72.805 14.160 73.095 ;
        RECT 10.720 72.555 12.090 72.805 ;
        RECT 10.720 72.295 10.970 72.555 ;
        RECT 11.480 72.125 11.730 72.285 ;
        RECT 10.380 71.955 11.730 72.125 ;
        RECT 10.380 71.915 10.800 71.955 ;
        RECT 10.110 71.365 10.460 71.735 ;
        RECT 8.815 70.805 9.145 71.185 ;
        RECT 9.315 71.025 9.485 71.355 ;
        RECT 10.630 71.185 10.800 71.915 ;
        RECT 11.900 71.785 12.090 72.555 ;
        RECT 10.970 71.455 11.380 71.785 ;
        RECT 11.670 71.445 12.090 71.785 ;
        RECT 12.260 72.375 12.780 72.685 ;
        RECT 12.950 72.635 14.160 72.805 ;
        RECT 14.390 72.665 14.720 73.355 ;
        RECT 12.260 71.615 12.430 72.375 ;
        RECT 12.600 71.785 12.780 72.195 ;
        RECT 12.950 72.125 13.120 72.635 ;
        RECT 14.890 72.485 15.060 73.095 ;
        RECT 15.330 72.635 15.660 73.145 ;
        RECT 14.890 72.465 15.210 72.485 ;
        RECT 13.290 72.295 15.210 72.465 ;
        RECT 12.950 71.955 14.850 72.125 ;
        RECT 13.180 71.615 13.510 71.735 ;
        RECT 12.260 71.445 13.510 71.615 ;
        RECT 9.785 70.985 10.800 71.185 ;
        RECT 10.970 70.805 11.380 71.245 ;
        RECT 11.670 71.015 11.920 71.445 ;
        RECT 12.120 70.805 12.440 71.265 ;
        RECT 13.680 71.195 13.850 71.955 ;
        RECT 14.520 71.895 14.850 71.955 ;
        RECT 14.040 71.725 14.370 71.785 ;
        RECT 14.040 71.455 14.700 71.725 ;
        RECT 15.020 71.400 15.210 72.295 ;
        RECT 13.000 71.025 13.850 71.195 ;
        RECT 14.050 70.805 14.710 71.285 ;
        RECT 14.890 71.070 15.210 71.400 ;
        RECT 15.410 72.045 15.660 72.635 ;
        RECT 15.840 72.555 16.125 73.355 ;
        RECT 16.305 73.015 16.560 73.045 ;
        RECT 16.305 72.845 16.645 73.015 ;
        RECT 16.305 72.375 16.560 72.845 ;
        RECT 15.410 71.715 16.210 72.045 ;
        RECT 15.410 71.065 15.660 71.715 ;
        RECT 16.380 71.515 16.560 72.375 ;
        RECT 17.165 72.215 17.375 73.355 ;
        RECT 17.545 72.205 17.875 73.185 ;
        RECT 18.045 72.215 18.275 73.355 ;
        RECT 15.840 70.805 16.125 71.265 ;
        RECT 16.305 70.985 16.560 71.515 ;
        RECT 17.165 70.805 17.375 71.625 ;
        RECT 17.545 71.605 17.795 72.205 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 18.945 72.265 22.455 73.355 ;
        RECT 22.625 72.265 23.835 73.355 ;
        RECT 17.965 71.795 18.295 72.045 ;
        RECT 17.545 70.975 17.875 71.605 ;
        RECT 18.045 70.805 18.275 71.625 ;
        RECT 18.945 71.575 20.595 72.095 ;
        RECT 20.765 71.745 22.455 72.265 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 18.945 70.805 22.455 71.575 ;
        RECT 22.625 71.555 23.145 72.095 ;
        RECT 23.315 71.725 23.835 72.265 ;
        RECT 24.005 72.215 24.345 73.185 ;
        RECT 24.515 72.215 24.685 73.355 ;
        RECT 24.955 72.555 25.205 73.355 ;
        RECT 25.850 72.385 26.180 73.185 ;
        RECT 26.480 72.555 26.810 73.355 ;
        RECT 26.980 72.385 27.310 73.185 ;
        RECT 24.875 72.215 27.310 72.385 ;
        RECT 27.890 72.385 28.220 73.185 ;
        RECT 28.390 72.555 28.720 73.355 ;
        RECT 29.020 72.385 29.350 73.185 ;
        RECT 29.995 72.555 30.245 73.355 ;
        RECT 27.890 72.215 30.325 72.385 ;
        RECT 30.515 72.215 30.685 73.355 ;
        RECT 30.855 72.215 31.195 73.185 ;
        RECT 31.365 72.265 33.035 73.355 ;
        RECT 24.005 71.605 24.180 72.215 ;
        RECT 24.875 71.965 25.045 72.215 ;
        RECT 24.350 71.795 25.045 71.965 ;
        RECT 25.220 71.795 25.640 71.995 ;
        RECT 25.810 71.795 26.140 71.995 ;
        RECT 26.310 71.795 26.640 71.995 ;
        RECT 22.625 70.805 23.835 71.555 ;
        RECT 24.005 70.975 24.345 71.605 ;
        RECT 24.515 70.805 24.765 71.605 ;
        RECT 24.955 71.455 26.180 71.625 ;
        RECT 24.955 70.975 25.285 71.455 ;
        RECT 25.455 70.805 25.680 71.265 ;
        RECT 25.850 70.975 26.180 71.455 ;
        RECT 26.810 71.585 26.980 72.215 ;
        RECT 27.165 71.795 27.515 72.045 ;
        RECT 27.685 71.795 28.035 72.045 ;
        RECT 28.220 71.585 28.390 72.215 ;
        RECT 28.560 71.795 28.890 71.995 ;
        RECT 29.060 71.795 29.390 71.995 ;
        RECT 29.560 71.795 29.980 71.995 ;
        RECT 30.155 71.965 30.325 72.215 ;
        RECT 30.155 71.795 30.850 71.965 ;
        RECT 26.810 70.975 27.310 71.585 ;
        RECT 27.890 70.975 28.390 71.585 ;
        RECT 29.020 71.455 30.245 71.625 ;
        RECT 31.020 71.605 31.195 72.215 ;
        RECT 29.020 70.975 29.350 71.455 ;
        RECT 29.520 70.805 29.745 71.265 ;
        RECT 29.915 70.975 30.245 71.455 ;
        RECT 30.435 70.805 30.685 71.605 ;
        RECT 30.855 70.975 31.195 71.605 ;
        RECT 31.365 71.575 32.115 72.095 ;
        RECT 32.285 71.745 33.035 72.265 ;
        RECT 33.410 72.385 33.740 73.185 ;
        RECT 33.910 72.555 34.240 73.355 ;
        RECT 34.540 72.385 34.870 73.185 ;
        RECT 35.515 72.555 35.765 73.355 ;
        RECT 33.410 72.215 35.845 72.385 ;
        RECT 36.035 72.215 36.205 73.355 ;
        RECT 36.375 72.215 36.715 73.185 ;
        RECT 36.885 72.920 42.230 73.355 ;
        RECT 33.205 71.795 33.555 72.045 ;
        RECT 33.740 71.585 33.910 72.215 ;
        RECT 34.080 71.795 34.410 71.995 ;
        RECT 34.580 71.795 34.910 71.995 ;
        RECT 35.080 71.795 35.500 71.995 ;
        RECT 35.675 71.965 35.845 72.215 ;
        RECT 35.675 71.795 36.370 71.965 ;
        RECT 31.365 70.805 33.035 71.575 ;
        RECT 33.410 70.975 33.910 71.585 ;
        RECT 34.540 71.455 35.765 71.625 ;
        RECT 36.540 71.605 36.715 72.215 ;
        RECT 34.540 70.975 34.870 71.455 ;
        RECT 35.040 70.805 35.265 71.265 ;
        RECT 35.435 70.975 35.765 71.455 ;
        RECT 35.955 70.805 36.205 71.605 ;
        RECT 36.375 70.975 36.715 71.605 ;
        RECT 38.470 71.350 38.810 72.180 ;
        RECT 40.290 71.670 40.640 72.920 ;
        RECT 42.405 72.265 44.075 73.355 ;
        RECT 42.405 71.575 43.155 72.095 ;
        RECT 43.325 71.745 44.075 72.265 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.705 72.265 48.215 73.355 ;
        RECT 44.705 71.575 46.355 72.095 ;
        RECT 46.525 71.745 48.215 72.265 ;
        RECT 48.885 72.215 49.115 73.355 ;
        RECT 49.285 72.205 49.615 73.185 ;
        RECT 49.785 72.215 49.995 73.355 ;
        RECT 50.430 72.385 50.760 73.185 ;
        RECT 50.930 72.555 51.260 73.355 ;
        RECT 51.560 72.385 51.890 73.185 ;
        RECT 52.535 72.555 52.785 73.355 ;
        RECT 50.430 72.215 52.865 72.385 ;
        RECT 53.055 72.215 53.225 73.355 ;
        RECT 53.395 72.215 53.735 73.185 ;
        RECT 54.110 72.385 54.440 73.185 ;
        RECT 54.610 72.555 54.940 73.355 ;
        RECT 55.240 72.385 55.570 73.185 ;
        RECT 56.215 72.555 56.465 73.355 ;
        RECT 54.110 72.215 56.545 72.385 ;
        RECT 56.735 72.215 56.905 73.355 ;
        RECT 57.075 72.215 57.415 73.185 ;
        RECT 48.865 71.795 49.195 72.045 ;
        RECT 36.885 70.805 42.230 71.350 ;
        RECT 42.405 70.805 44.075 71.575 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.705 70.805 48.215 71.575 ;
        RECT 48.885 70.805 49.115 71.625 ;
        RECT 49.365 71.605 49.615 72.205 ;
        RECT 50.225 71.795 50.575 72.045 ;
        RECT 49.285 70.975 49.615 71.605 ;
        RECT 49.785 70.805 49.995 71.625 ;
        RECT 50.760 71.585 50.930 72.215 ;
        RECT 51.100 71.795 51.430 71.995 ;
        RECT 51.600 71.795 51.930 71.995 ;
        RECT 52.100 71.795 52.520 71.995 ;
        RECT 52.695 71.965 52.865 72.215 ;
        RECT 52.695 71.795 53.390 71.965 ;
        RECT 50.430 70.975 50.930 71.585 ;
        RECT 51.560 71.455 52.785 71.625 ;
        RECT 53.560 71.605 53.735 72.215 ;
        RECT 53.905 71.795 54.255 72.045 ;
        RECT 51.560 70.975 51.890 71.455 ;
        RECT 52.060 70.805 52.285 71.265 ;
        RECT 52.455 70.975 52.785 71.455 ;
        RECT 52.975 70.805 53.225 71.605 ;
        RECT 53.395 70.975 53.735 71.605 ;
        RECT 54.440 71.585 54.610 72.215 ;
        RECT 54.780 71.795 55.110 71.995 ;
        RECT 55.280 71.795 55.610 71.995 ;
        RECT 55.780 71.795 56.200 71.995 ;
        RECT 56.375 71.965 56.545 72.215 ;
        RECT 56.375 71.795 57.070 71.965 ;
        RECT 54.110 70.975 54.610 71.585 ;
        RECT 55.240 71.455 56.465 71.625 ;
        RECT 57.240 71.605 57.415 72.215 ;
        RECT 55.240 70.975 55.570 71.455 ;
        RECT 55.740 70.805 55.965 71.265 ;
        RECT 56.135 70.975 56.465 71.455 ;
        RECT 56.655 70.805 56.905 71.605 ;
        RECT 57.075 70.975 57.415 71.605 ;
        RECT 57.585 72.215 57.925 73.185 ;
        RECT 58.095 72.215 58.265 73.355 ;
        RECT 58.535 72.555 58.785 73.355 ;
        RECT 59.430 72.385 59.760 73.185 ;
        RECT 60.060 72.555 60.390 73.355 ;
        RECT 60.560 72.385 60.890 73.185 ;
        RECT 58.455 72.215 60.890 72.385 ;
        RECT 61.265 72.265 62.935 73.355 ;
        RECT 57.585 71.605 57.760 72.215 ;
        RECT 58.455 71.965 58.625 72.215 ;
        RECT 57.930 71.795 58.625 71.965 ;
        RECT 58.800 71.795 59.220 71.995 ;
        RECT 59.390 71.795 59.720 71.995 ;
        RECT 59.890 71.795 60.220 71.995 ;
        RECT 57.585 70.975 57.925 71.605 ;
        RECT 58.095 70.805 58.345 71.605 ;
        RECT 58.535 71.455 59.760 71.625 ;
        RECT 58.535 70.975 58.865 71.455 ;
        RECT 59.035 70.805 59.260 71.265 ;
        RECT 59.430 70.975 59.760 71.455 ;
        RECT 60.390 71.585 60.560 72.215 ;
        RECT 60.745 71.795 61.095 72.045 ;
        RECT 60.390 70.975 60.890 71.585 ;
        RECT 61.265 71.575 62.015 72.095 ;
        RECT 62.185 71.745 62.935 72.265 ;
        RECT 63.105 72.385 63.415 73.185 ;
        RECT 63.585 72.555 63.895 73.355 ;
        RECT 64.065 72.725 64.325 73.185 ;
        RECT 64.495 72.895 64.750 73.355 ;
        RECT 64.925 72.725 65.185 73.185 ;
        RECT 64.065 72.555 65.185 72.725 ;
        RECT 63.105 72.215 64.135 72.385 ;
        RECT 61.265 70.805 62.935 71.575 ;
        RECT 63.105 71.305 63.275 72.215 ;
        RECT 63.445 71.475 63.795 72.045 ;
        RECT 63.965 71.965 64.135 72.215 ;
        RECT 64.925 72.305 65.185 72.555 ;
        RECT 65.355 72.485 65.640 73.355 ;
        RECT 64.925 72.135 65.680 72.305 ;
        RECT 65.865 72.265 67.075 73.355 ;
        RECT 63.965 71.795 65.105 71.965 ;
        RECT 65.275 71.625 65.680 72.135 ;
        RECT 64.030 71.455 65.680 71.625 ;
        RECT 65.865 71.555 66.385 72.095 ;
        RECT 66.555 71.725 67.075 72.265 ;
        RECT 67.335 72.425 67.505 73.185 ;
        RECT 67.720 72.595 68.050 73.355 ;
        RECT 67.335 72.255 68.050 72.425 ;
        RECT 68.220 72.280 68.475 73.185 ;
        RECT 67.245 71.705 67.600 72.075 ;
        RECT 67.880 72.045 68.050 72.255 ;
        RECT 67.880 71.715 68.135 72.045 ;
        RECT 63.105 70.975 63.405 71.305 ;
        RECT 63.575 70.805 63.850 71.285 ;
        RECT 64.030 71.065 64.325 71.455 ;
        RECT 64.495 70.805 64.750 71.285 ;
        RECT 64.925 71.065 65.185 71.455 ;
        RECT 65.355 70.805 65.635 71.285 ;
        RECT 65.865 70.805 67.075 71.555 ;
        RECT 67.880 71.525 68.050 71.715 ;
        RECT 68.305 71.550 68.475 72.280 ;
        RECT 68.650 72.205 68.910 73.355 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 71.390 72.215 71.725 73.185 ;
        RECT 71.895 72.215 72.065 73.355 ;
        RECT 72.235 73.015 74.265 73.185 ;
        RECT 67.335 71.355 68.050 71.525 ;
        RECT 67.335 70.975 67.505 71.355 ;
        RECT 67.720 70.805 68.050 71.185 ;
        RECT 68.220 70.975 68.475 71.550 ;
        RECT 68.650 70.805 68.910 71.645 ;
        RECT 71.390 71.545 71.560 72.215 ;
        RECT 72.235 72.045 72.405 73.015 ;
        RECT 71.730 71.715 71.985 72.045 ;
        RECT 72.210 71.715 72.405 72.045 ;
        RECT 72.575 72.675 73.700 72.845 ;
        RECT 71.815 71.545 71.985 71.715 ;
        RECT 72.575 71.545 72.745 72.675 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 71.390 70.975 71.645 71.545 ;
        RECT 71.815 71.375 72.745 71.545 ;
        RECT 72.915 72.335 73.925 72.505 ;
        RECT 72.915 71.535 73.085 72.335 ;
        RECT 73.290 71.995 73.565 72.135 ;
        RECT 73.285 71.825 73.565 71.995 ;
        RECT 72.570 71.340 72.745 71.375 ;
        RECT 71.815 70.805 72.145 71.205 ;
        RECT 72.570 70.975 73.100 71.340 ;
        RECT 73.290 70.975 73.565 71.825 ;
        RECT 73.735 70.975 73.925 72.335 ;
        RECT 74.095 72.350 74.265 73.015 ;
        RECT 74.435 72.595 74.605 73.355 ;
        RECT 74.840 72.595 75.355 73.005 ;
        RECT 75.525 72.920 80.870 73.355 ;
        RECT 81.045 72.920 86.390 73.355 ;
        RECT 74.095 72.160 74.845 72.350 ;
        RECT 75.015 71.785 75.355 72.595 ;
        RECT 74.125 71.615 75.355 71.785 ;
        RECT 74.105 70.805 74.615 71.340 ;
        RECT 74.835 71.010 75.080 71.615 ;
        RECT 77.110 71.350 77.450 72.180 ;
        RECT 78.930 71.670 79.280 72.920 ;
        RECT 82.630 71.350 82.970 72.180 ;
        RECT 84.450 71.670 84.800 72.920 ;
        RECT 86.565 72.265 88.235 73.355 ;
        RECT 86.565 71.575 87.315 72.095 ;
        RECT 87.485 71.745 88.235 72.265 ;
        RECT 89.070 72.385 89.400 73.185 ;
        RECT 89.570 72.555 89.900 73.355 ;
        RECT 90.200 72.385 90.530 73.185 ;
        RECT 91.175 72.555 91.425 73.355 ;
        RECT 89.070 72.215 91.505 72.385 ;
        RECT 91.695 72.215 91.865 73.355 ;
        RECT 92.035 72.215 92.375 73.185 ;
        RECT 92.545 72.265 95.135 73.355 ;
        RECT 88.865 71.795 89.215 72.045 ;
        RECT 89.400 71.585 89.570 72.215 ;
        RECT 89.740 71.795 90.070 71.995 ;
        RECT 90.240 71.795 90.570 71.995 ;
        RECT 90.740 71.795 91.160 71.995 ;
        RECT 91.335 71.965 91.505 72.215 ;
        RECT 91.335 71.795 92.030 71.965 ;
        RECT 75.525 70.805 80.870 71.350 ;
        RECT 81.045 70.805 86.390 71.350 ;
        RECT 86.565 70.805 88.235 71.575 ;
        RECT 89.070 70.975 89.570 71.585 ;
        RECT 90.200 71.455 91.425 71.625 ;
        RECT 92.200 71.605 92.375 72.215 ;
        RECT 90.200 70.975 90.530 71.455 ;
        RECT 90.700 70.805 90.925 71.265 ;
        RECT 91.095 70.975 91.425 71.455 ;
        RECT 91.615 70.805 91.865 71.605 ;
        RECT 92.035 70.975 92.375 71.605 ;
        RECT 92.545 71.575 93.755 72.095 ;
        RECT 93.925 71.745 95.135 72.265 ;
        RECT 95.765 72.190 96.055 73.355 ;
        RECT 96.225 72.265 98.815 73.355 ;
        RECT 99.535 72.685 99.705 73.185 ;
        RECT 99.875 72.855 100.205 73.355 ;
        RECT 99.535 72.515 100.200 72.685 ;
        RECT 96.225 71.575 97.435 72.095 ;
        RECT 97.605 71.745 98.815 72.265 ;
        RECT 99.450 71.695 99.800 72.345 ;
        RECT 92.545 70.805 95.135 71.575 ;
        RECT 95.765 70.805 96.055 71.530 ;
        RECT 96.225 70.805 98.815 71.575 ;
        RECT 99.970 71.525 100.200 72.515 ;
        RECT 99.535 71.355 100.200 71.525 ;
        RECT 99.535 71.065 99.705 71.355 ;
        RECT 99.875 70.805 100.205 71.185 ;
        RECT 100.375 71.065 100.600 73.185 ;
        RECT 100.815 72.855 101.145 73.355 ;
        RECT 101.315 72.685 101.485 73.185 ;
        RECT 101.720 72.970 102.550 73.140 ;
        RECT 102.790 72.975 103.170 73.355 ;
        RECT 100.790 72.515 101.485 72.685 ;
        RECT 100.790 71.545 100.960 72.515 ;
        RECT 101.130 71.725 101.540 72.345 ;
        RECT 101.710 72.295 102.210 72.675 ;
        RECT 100.790 71.355 101.485 71.545 ;
        RECT 101.710 71.425 101.930 72.295 ;
        RECT 102.380 72.125 102.550 72.970 ;
        RECT 103.350 72.805 103.520 73.095 ;
        RECT 103.690 72.975 104.020 73.355 ;
        RECT 104.490 72.885 105.120 73.135 ;
        RECT 105.300 72.975 105.720 73.355 ;
        RECT 104.950 72.805 105.120 72.885 ;
        RECT 105.920 72.805 106.160 73.095 ;
        RECT 102.720 72.555 104.090 72.805 ;
        RECT 102.720 72.295 102.970 72.555 ;
        RECT 103.480 72.125 103.730 72.285 ;
        RECT 102.380 71.955 103.730 72.125 ;
        RECT 102.380 71.915 102.800 71.955 ;
        RECT 102.110 71.365 102.460 71.735 ;
        RECT 100.815 70.805 101.145 71.185 ;
        RECT 101.315 71.025 101.485 71.355 ;
        RECT 102.630 71.185 102.800 71.915 ;
        RECT 103.900 71.785 104.090 72.555 ;
        RECT 102.970 71.455 103.380 71.785 ;
        RECT 103.670 71.445 104.090 71.785 ;
        RECT 104.260 72.375 104.780 72.685 ;
        RECT 104.950 72.635 106.160 72.805 ;
        RECT 106.390 72.665 106.720 73.355 ;
        RECT 104.260 71.615 104.430 72.375 ;
        RECT 104.600 71.785 104.780 72.195 ;
        RECT 104.950 72.125 105.120 72.635 ;
        RECT 106.890 72.485 107.060 73.095 ;
        RECT 107.330 72.635 107.660 73.145 ;
        RECT 106.890 72.465 107.210 72.485 ;
        RECT 105.290 72.295 107.210 72.465 ;
        RECT 104.950 71.955 106.850 72.125 ;
        RECT 105.180 71.615 105.510 71.735 ;
        RECT 104.260 71.445 105.510 71.615 ;
        RECT 101.785 70.985 102.800 71.185 ;
        RECT 102.970 70.805 103.380 71.245 ;
        RECT 103.670 71.015 103.920 71.445 ;
        RECT 104.120 70.805 104.440 71.265 ;
        RECT 105.680 71.195 105.850 71.955 ;
        RECT 106.520 71.895 106.850 71.955 ;
        RECT 106.040 71.725 106.370 71.785 ;
        RECT 106.040 71.455 106.700 71.725 ;
        RECT 107.020 71.400 107.210 72.295 ;
        RECT 105.000 71.025 105.850 71.195 ;
        RECT 106.050 70.805 106.710 71.285 ;
        RECT 106.890 71.070 107.210 71.400 ;
        RECT 107.410 72.045 107.660 72.635 ;
        RECT 107.840 72.555 108.125 73.355 ;
        RECT 108.305 72.375 108.560 73.045 ;
        RECT 107.410 71.715 108.210 72.045 ;
        RECT 107.410 71.065 107.660 71.715 ;
        RECT 108.380 71.515 108.560 72.375 ;
        RECT 109.165 72.215 109.375 73.355 ;
        RECT 109.545 72.205 109.875 73.185 ;
        RECT 110.045 72.215 110.275 73.355 ;
        RECT 110.485 72.265 112.155 73.355 ;
        RECT 108.305 71.315 108.560 71.515 ;
        RECT 107.840 70.805 108.125 71.265 ;
        RECT 108.305 71.145 108.645 71.315 ;
        RECT 108.305 70.985 108.560 71.145 ;
        RECT 109.165 70.805 109.375 71.625 ;
        RECT 109.545 71.605 109.795 72.205 ;
        RECT 109.965 71.795 110.295 72.045 ;
        RECT 109.545 70.975 109.875 71.605 ;
        RECT 110.045 70.805 110.275 71.625 ;
        RECT 110.485 71.575 111.235 72.095 ;
        RECT 111.405 71.745 112.155 72.265 ;
        RECT 112.785 72.595 113.300 73.005 ;
        RECT 113.535 72.595 113.705 73.355 ;
        RECT 113.875 73.015 115.905 73.185 ;
        RECT 112.785 71.785 113.125 72.595 ;
        RECT 113.875 72.350 114.045 73.015 ;
        RECT 114.440 72.675 115.565 72.845 ;
        RECT 113.295 72.160 114.045 72.350 ;
        RECT 114.215 72.335 115.225 72.505 ;
        RECT 112.785 71.615 114.015 71.785 ;
        RECT 110.485 70.805 112.155 71.575 ;
        RECT 113.060 71.010 113.305 71.615 ;
        RECT 113.525 70.805 114.035 71.340 ;
        RECT 114.215 70.975 114.405 72.335 ;
        RECT 114.575 71.995 114.850 72.135 ;
        RECT 114.575 71.825 114.855 71.995 ;
        RECT 114.575 70.975 114.850 71.825 ;
        RECT 115.055 71.535 115.225 72.335 ;
        RECT 115.395 71.545 115.565 72.675 ;
        RECT 115.735 72.045 115.905 73.015 ;
        RECT 116.075 72.215 116.245 73.355 ;
        RECT 116.415 72.215 116.750 73.185 ;
        RECT 115.735 71.715 115.930 72.045 ;
        RECT 116.155 71.715 116.410 72.045 ;
        RECT 116.155 71.545 116.325 71.715 ;
        RECT 116.580 71.545 116.750 72.215 ;
        RECT 115.395 71.375 116.325 71.545 ;
        RECT 115.395 71.340 115.570 71.375 ;
        RECT 115.040 70.975 115.570 71.340 ;
        RECT 115.995 70.805 116.325 71.205 ;
        RECT 116.495 70.975 116.750 71.545 ;
        RECT 116.925 72.280 117.195 73.185 ;
        RECT 117.365 72.595 117.695 73.355 ;
        RECT 117.875 72.425 118.045 73.185 ;
        RECT 116.925 71.480 117.095 72.280 ;
        RECT 117.380 72.255 118.045 72.425 ;
        RECT 118.305 72.265 120.895 73.355 ;
        RECT 117.380 72.110 117.550 72.255 ;
        RECT 117.265 71.780 117.550 72.110 ;
        RECT 117.380 71.525 117.550 71.780 ;
        RECT 117.785 71.705 118.115 72.075 ;
        RECT 118.305 71.575 119.515 72.095 ;
        RECT 119.685 71.745 120.895 72.265 ;
        RECT 121.525 72.190 121.815 73.355 ;
        RECT 122.445 72.265 123.655 73.355 ;
        RECT 122.445 71.725 122.965 72.265 ;
        RECT 116.925 70.975 117.185 71.480 ;
        RECT 117.380 71.355 118.045 71.525 ;
        RECT 117.365 70.805 117.695 71.185 ;
        RECT 117.875 70.975 118.045 71.355 ;
        RECT 118.305 70.805 120.895 71.575 ;
        RECT 123.135 71.555 123.655 72.095 ;
        RECT 121.525 70.805 121.815 71.530 ;
        RECT 122.445 70.805 123.655 71.555 ;
        RECT 5.520 70.635 123.740 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 6.985 69.885 8.195 70.635 ;
        RECT 8.370 70.085 8.625 70.375 ;
        RECT 8.795 70.255 9.125 70.635 ;
        RECT 8.370 69.915 9.120 70.085 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 6.985 69.345 7.505 69.885 ;
        RECT 7.675 69.175 8.195 69.715 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 6.985 68.085 8.195 69.175 ;
        RECT 8.370 69.095 8.720 69.745 ;
        RECT 8.890 68.925 9.120 69.915 ;
        RECT 8.370 68.755 9.120 68.925 ;
        RECT 8.370 68.255 8.625 68.755 ;
        RECT 8.795 68.085 9.125 68.585 ;
        RECT 9.295 68.255 9.465 70.375 ;
        RECT 9.825 70.275 10.155 70.635 ;
        RECT 10.325 70.245 10.820 70.415 ;
        RECT 11.025 70.245 11.880 70.415 ;
        RECT 9.695 69.055 10.155 70.105 ;
        RECT 9.635 68.270 9.960 69.055 ;
        RECT 10.325 68.885 10.495 70.245 ;
        RECT 10.665 69.335 11.015 69.955 ;
        RECT 11.185 69.735 11.540 69.955 ;
        RECT 11.185 69.145 11.355 69.735 ;
        RECT 11.710 69.535 11.880 70.245 ;
        RECT 12.755 70.175 13.085 70.635 ;
        RECT 13.295 70.275 13.645 70.445 ;
        RECT 12.085 69.705 12.875 69.955 ;
        RECT 13.295 69.885 13.555 70.275 ;
        RECT 13.865 70.185 14.815 70.465 ;
        RECT 14.985 70.195 15.175 70.635 ;
        RECT 15.345 70.255 16.415 70.425 ;
        RECT 13.045 69.535 13.215 69.715 ;
        RECT 10.325 68.715 10.720 68.885 ;
        RECT 10.890 68.755 11.355 69.145 ;
        RECT 11.525 69.365 13.215 69.535 ;
        RECT 10.550 68.585 10.720 68.715 ;
        RECT 11.525 68.585 11.695 69.365 ;
        RECT 13.385 69.195 13.555 69.885 ;
        RECT 12.055 69.025 13.555 69.195 ;
        RECT 13.745 69.225 13.955 70.015 ;
        RECT 14.125 69.395 14.475 70.015 ;
        RECT 14.645 69.405 14.815 70.185 ;
        RECT 15.345 70.025 15.515 70.255 ;
        RECT 14.985 69.855 15.515 70.025 ;
        RECT 14.985 69.575 15.205 69.855 ;
        RECT 15.685 69.685 15.925 70.085 ;
        RECT 14.645 69.235 15.050 69.405 ;
        RECT 15.385 69.315 15.925 69.685 ;
        RECT 16.095 69.900 16.415 70.255 ;
        RECT 16.660 70.175 16.965 70.635 ;
        RECT 17.135 69.925 17.390 70.455 ;
        RECT 16.095 69.725 16.420 69.900 ;
        RECT 16.095 69.425 17.010 69.725 ;
        RECT 16.270 69.395 17.010 69.425 ;
        RECT 13.745 69.065 14.420 69.225 ;
        RECT 14.880 69.145 15.050 69.235 ;
        RECT 13.745 69.055 14.710 69.065 ;
        RECT 13.385 68.885 13.555 69.025 ;
        RECT 10.130 68.085 10.380 68.545 ;
        RECT 10.550 68.255 10.800 68.585 ;
        RECT 11.015 68.255 11.695 68.585 ;
        RECT 11.865 68.685 12.940 68.855 ;
        RECT 13.385 68.715 13.945 68.885 ;
        RECT 14.250 68.765 14.710 69.055 ;
        RECT 14.880 68.975 16.100 69.145 ;
        RECT 11.865 68.345 12.035 68.685 ;
        RECT 12.270 68.085 12.600 68.515 ;
        RECT 12.770 68.345 12.940 68.685 ;
        RECT 13.235 68.085 13.605 68.545 ;
        RECT 13.775 68.255 13.945 68.715 ;
        RECT 14.880 68.595 15.050 68.975 ;
        RECT 16.270 68.805 16.440 69.395 ;
        RECT 17.180 69.275 17.390 69.925 ;
        RECT 17.715 69.835 18.045 70.635 ;
        RECT 18.215 69.985 18.385 70.465 ;
        RECT 18.555 70.155 18.885 70.635 ;
        RECT 19.055 69.985 19.225 70.465 ;
        RECT 19.475 70.155 19.715 70.635 ;
        RECT 19.895 69.985 20.065 70.465 ;
        RECT 14.180 68.255 15.050 68.595 ;
        RECT 15.640 68.635 16.440 68.805 ;
        RECT 15.220 68.085 15.470 68.545 ;
        RECT 15.640 68.345 15.810 68.635 ;
        RECT 15.990 68.085 16.320 68.465 ;
        RECT 16.660 68.085 16.965 69.225 ;
        RECT 17.135 68.395 17.390 69.275 ;
        RECT 18.215 69.815 19.225 69.985 ;
        RECT 19.430 69.815 20.065 69.985 ;
        RECT 20.325 69.865 23.835 70.635 ;
        RECT 18.215 69.275 18.710 69.815 ;
        RECT 19.430 69.645 19.600 69.815 ;
        RECT 19.100 69.475 19.600 69.645 ;
        RECT 17.715 68.085 18.045 69.235 ;
        RECT 18.215 69.105 19.225 69.275 ;
        RECT 18.215 68.255 18.385 69.105 ;
        RECT 18.555 68.085 18.885 68.885 ;
        RECT 19.055 68.255 19.225 69.105 ;
        RECT 19.430 69.235 19.600 69.475 ;
        RECT 19.770 69.405 20.150 69.645 ;
        RECT 20.325 69.345 21.975 69.865 ;
        RECT 24.005 69.835 24.345 70.465 ;
        RECT 24.515 69.835 24.765 70.635 ;
        RECT 24.955 69.985 25.285 70.465 ;
        RECT 25.455 70.175 25.680 70.635 ;
        RECT 25.850 69.985 26.180 70.465 ;
        RECT 19.430 69.065 20.145 69.235 ;
        RECT 22.145 69.175 23.835 69.695 ;
        RECT 19.405 68.085 19.645 68.885 ;
        RECT 19.815 68.255 20.145 69.065 ;
        RECT 20.325 68.085 23.835 69.175 ;
        RECT 24.005 69.225 24.180 69.835 ;
        RECT 24.955 69.815 26.180 69.985 ;
        RECT 26.810 69.855 27.310 70.465 ;
        RECT 27.685 69.865 31.195 70.635 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 31.825 69.865 35.335 70.635 ;
        RECT 35.505 69.885 36.715 70.635 ;
        RECT 36.885 69.960 37.145 70.465 ;
        RECT 37.325 70.255 37.655 70.635 ;
        RECT 37.835 70.085 38.005 70.465 ;
        RECT 24.350 69.475 25.045 69.645 ;
        RECT 24.875 69.225 25.045 69.475 ;
        RECT 25.220 69.445 25.640 69.645 ;
        RECT 25.810 69.445 26.140 69.645 ;
        RECT 26.310 69.445 26.640 69.645 ;
        RECT 26.810 69.225 26.980 69.855 ;
        RECT 27.165 69.395 27.515 69.645 ;
        RECT 27.685 69.345 29.335 69.865 ;
        RECT 24.005 68.255 24.345 69.225 ;
        RECT 24.515 68.085 24.685 69.225 ;
        RECT 24.875 69.055 27.310 69.225 ;
        RECT 29.505 69.175 31.195 69.695 ;
        RECT 31.825 69.345 33.475 69.865 ;
        RECT 24.955 68.085 25.205 68.885 ;
        RECT 25.850 68.255 26.180 69.055 ;
        RECT 26.480 68.085 26.810 68.885 ;
        RECT 26.980 68.255 27.310 69.055 ;
        RECT 27.685 68.085 31.195 69.175 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 33.645 69.175 35.335 69.695 ;
        RECT 35.505 69.345 36.025 69.885 ;
        RECT 36.195 69.175 36.715 69.715 ;
        RECT 31.825 68.085 35.335 69.175 ;
        RECT 35.505 68.085 36.715 69.175 ;
        RECT 36.885 69.160 37.055 69.960 ;
        RECT 37.340 69.915 38.005 70.085 ;
        RECT 37.340 69.660 37.510 69.915 ;
        RECT 38.265 69.865 39.935 70.635 ;
        RECT 37.225 69.330 37.510 69.660 ;
        RECT 37.745 69.365 38.075 69.735 ;
        RECT 38.265 69.345 39.015 69.865 ;
        RECT 40.165 69.815 40.375 70.635 ;
        RECT 40.545 69.835 40.875 70.465 ;
        RECT 37.340 69.185 37.510 69.330 ;
        RECT 36.885 68.255 37.155 69.160 ;
        RECT 37.340 69.015 38.005 69.185 ;
        RECT 39.185 69.175 39.935 69.695 ;
        RECT 40.545 69.235 40.795 69.835 ;
        RECT 41.045 69.815 41.275 70.635 ;
        RECT 41.485 69.865 44.075 70.635 ;
        RECT 44.795 70.085 44.965 70.375 ;
        RECT 45.135 70.255 45.465 70.635 ;
        RECT 44.795 69.915 45.460 70.085 ;
        RECT 40.965 69.395 41.295 69.645 ;
        RECT 41.485 69.345 42.695 69.865 ;
        RECT 37.325 68.085 37.655 68.845 ;
        RECT 37.835 68.255 38.005 69.015 ;
        RECT 38.265 68.085 39.935 69.175 ;
        RECT 40.165 68.085 40.375 69.225 ;
        RECT 40.545 68.255 40.875 69.235 ;
        RECT 41.045 68.085 41.275 69.225 ;
        RECT 42.865 69.175 44.075 69.695 ;
        RECT 41.485 68.085 44.075 69.175 ;
        RECT 44.710 69.095 45.060 69.745 ;
        RECT 45.230 68.925 45.460 69.915 ;
        RECT 44.795 68.755 45.460 68.925 ;
        RECT 44.795 68.255 44.965 68.755 ;
        RECT 45.135 68.085 45.465 68.585 ;
        RECT 45.635 68.255 45.860 70.375 ;
        RECT 46.075 70.255 46.405 70.635 ;
        RECT 46.575 70.085 46.745 70.415 ;
        RECT 47.045 70.255 48.060 70.455 ;
        RECT 46.050 69.895 46.745 70.085 ;
        RECT 46.050 68.925 46.220 69.895 ;
        RECT 46.390 69.095 46.800 69.715 ;
        RECT 46.970 69.145 47.190 70.015 ;
        RECT 47.370 69.705 47.720 70.075 ;
        RECT 47.890 69.525 48.060 70.255 ;
        RECT 48.230 70.195 48.640 70.635 ;
        RECT 48.930 69.995 49.180 70.425 ;
        RECT 49.380 70.175 49.700 70.635 ;
        RECT 50.260 70.245 51.110 70.415 ;
        RECT 48.230 69.655 48.640 69.985 ;
        RECT 48.930 69.655 49.350 69.995 ;
        RECT 47.640 69.485 48.060 69.525 ;
        RECT 47.640 69.315 48.990 69.485 ;
        RECT 46.050 68.755 46.745 68.925 ;
        RECT 46.970 68.765 47.470 69.145 ;
        RECT 46.075 68.085 46.405 68.585 ;
        RECT 46.575 68.255 46.745 68.755 ;
        RECT 47.640 68.470 47.810 69.315 ;
        RECT 48.740 69.155 48.990 69.315 ;
        RECT 47.980 68.885 48.230 69.145 ;
        RECT 49.160 68.885 49.350 69.655 ;
        RECT 47.980 68.635 49.350 68.885 ;
        RECT 49.520 69.825 50.770 69.995 ;
        RECT 49.520 69.065 49.690 69.825 ;
        RECT 50.440 69.705 50.770 69.825 ;
        RECT 49.860 69.245 50.040 69.655 ;
        RECT 50.940 69.485 51.110 70.245 ;
        RECT 51.310 70.155 51.970 70.635 ;
        RECT 52.150 70.040 52.470 70.370 ;
        RECT 51.300 69.715 51.960 69.985 ;
        RECT 51.300 69.655 51.630 69.715 ;
        RECT 51.780 69.485 52.110 69.545 ;
        RECT 50.210 69.315 52.110 69.485 ;
        RECT 49.520 68.755 50.040 69.065 ;
        RECT 50.210 68.805 50.380 69.315 ;
        RECT 52.280 69.145 52.470 70.040 ;
        RECT 50.550 68.975 52.470 69.145 ;
        RECT 52.150 68.955 52.470 68.975 ;
        RECT 52.670 69.725 52.920 70.375 ;
        RECT 53.100 70.175 53.385 70.635 ;
        RECT 53.565 69.925 53.820 70.455 ;
        RECT 52.670 69.395 53.470 69.725 ;
        RECT 53.640 69.615 53.820 69.925 ;
        RECT 54.365 69.865 56.955 70.635 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 57.585 69.865 60.175 70.635 ;
        RECT 60.805 69.875 61.515 70.465 ;
        RECT 62.025 70.105 62.355 70.465 ;
        RECT 62.555 70.275 62.885 70.635 ;
        RECT 63.055 70.105 63.385 70.465 ;
        RECT 62.025 69.895 63.385 70.105 ;
        RECT 53.640 69.445 53.905 69.615 ;
        RECT 50.210 68.635 51.420 68.805 ;
        RECT 46.980 68.300 47.810 68.470 ;
        RECT 48.050 68.085 48.430 68.465 ;
        RECT 48.610 68.345 48.780 68.635 ;
        RECT 50.210 68.555 50.380 68.635 ;
        RECT 48.950 68.085 49.280 68.465 ;
        RECT 49.750 68.305 50.380 68.555 ;
        RECT 50.560 68.085 50.980 68.465 ;
        RECT 51.180 68.345 51.420 68.635 ;
        RECT 51.650 68.085 51.980 68.775 ;
        RECT 52.150 68.345 52.320 68.955 ;
        RECT 52.670 68.805 52.920 69.395 ;
        RECT 53.640 69.065 53.820 69.445 ;
        RECT 54.365 69.345 55.575 69.865 ;
        RECT 55.745 69.175 56.955 69.695 ;
        RECT 57.585 69.345 58.795 69.865 ;
        RECT 52.590 68.295 52.920 68.805 ;
        RECT 53.100 68.085 53.385 68.885 ;
        RECT 53.565 68.395 53.820 69.065 ;
        RECT 54.365 68.085 56.955 69.175 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 58.965 69.175 60.175 69.695 ;
        RECT 57.585 68.085 60.175 69.175 ;
        RECT 60.805 68.905 61.010 69.875 ;
        RECT 64.030 69.795 64.290 70.635 ;
        RECT 64.465 69.890 64.720 70.465 ;
        RECT 64.890 70.255 65.220 70.635 ;
        RECT 65.435 70.085 65.605 70.465 ;
        RECT 64.890 69.915 65.605 70.085 ;
        RECT 65.955 70.085 66.125 70.465 ;
        RECT 66.340 70.255 66.670 70.635 ;
        RECT 65.955 69.915 66.670 70.085 ;
        RECT 61.180 69.105 61.510 69.645 ;
        RECT 61.685 69.395 62.180 69.725 ;
        RECT 62.500 69.395 62.875 69.725 ;
        RECT 63.085 69.395 63.395 69.725 ;
        RECT 61.685 69.105 62.010 69.395 ;
        RECT 62.205 68.905 62.535 69.125 ;
        RECT 60.805 68.675 62.535 68.905 ;
        RECT 60.805 68.255 61.505 68.675 ;
        RECT 61.705 68.085 62.035 68.445 ;
        RECT 62.205 68.275 62.535 68.675 ;
        RECT 62.705 68.470 62.875 69.395 ;
        RECT 63.055 68.085 63.385 69.145 ;
        RECT 64.030 68.085 64.290 69.235 ;
        RECT 64.465 69.160 64.635 69.890 ;
        RECT 64.890 69.725 65.060 69.915 ;
        RECT 64.805 69.395 65.060 69.725 ;
        RECT 64.890 69.185 65.060 69.395 ;
        RECT 65.340 69.365 65.695 69.735 ;
        RECT 65.865 69.365 66.220 69.735 ;
        RECT 66.500 69.725 66.670 69.915 ;
        RECT 66.840 69.890 67.095 70.465 ;
        RECT 66.500 69.395 66.755 69.725 ;
        RECT 66.500 69.185 66.670 69.395 ;
        RECT 64.465 68.255 64.720 69.160 ;
        RECT 64.890 69.015 65.605 69.185 ;
        RECT 64.890 68.085 65.220 68.845 ;
        RECT 65.435 68.255 65.605 69.015 ;
        RECT 65.955 69.015 66.670 69.185 ;
        RECT 66.925 69.160 67.095 69.890 ;
        RECT 67.270 69.795 67.530 70.635 ;
        RECT 67.795 70.085 67.965 70.465 ;
        RECT 68.180 70.255 68.510 70.635 ;
        RECT 67.795 69.915 68.510 70.085 ;
        RECT 67.705 69.365 68.060 69.735 ;
        RECT 68.340 69.725 68.510 69.915 ;
        RECT 68.680 69.890 68.935 70.465 ;
        RECT 68.340 69.395 68.595 69.725 ;
        RECT 65.955 68.255 66.125 69.015 ;
        RECT 66.340 68.085 66.670 68.845 ;
        RECT 66.840 68.255 67.095 69.160 ;
        RECT 67.270 68.085 67.530 69.235 ;
        RECT 68.340 69.185 68.510 69.395 ;
        RECT 67.795 69.015 68.510 69.185 ;
        RECT 68.765 69.160 68.935 69.890 ;
        RECT 69.110 69.795 69.370 70.635 ;
        RECT 69.635 70.085 69.805 70.465 ;
        RECT 70.020 70.255 70.350 70.635 ;
        RECT 69.635 69.915 70.350 70.085 ;
        RECT 69.545 69.365 69.900 69.735 ;
        RECT 70.180 69.725 70.350 69.915 ;
        RECT 70.520 69.890 70.775 70.465 ;
        RECT 70.180 69.395 70.435 69.725 ;
        RECT 67.795 68.255 67.965 69.015 ;
        RECT 68.180 68.085 68.510 68.845 ;
        RECT 68.680 68.255 68.935 69.160 ;
        RECT 69.110 68.085 69.370 69.235 ;
        RECT 70.180 69.185 70.350 69.395 ;
        RECT 69.635 69.015 70.350 69.185 ;
        RECT 70.605 69.160 70.775 69.890 ;
        RECT 70.950 69.795 71.210 70.635 ;
        RECT 71.475 70.085 71.645 70.465 ;
        RECT 71.825 70.255 72.155 70.635 ;
        RECT 71.475 69.915 72.140 70.085 ;
        RECT 72.335 69.960 72.595 70.465 ;
        RECT 71.405 69.365 71.735 69.735 ;
        RECT 71.970 69.660 72.140 69.915 ;
        RECT 71.970 69.330 72.255 69.660 ;
        RECT 69.635 68.255 69.805 69.015 ;
        RECT 70.020 68.085 70.350 68.845 ;
        RECT 70.520 68.255 70.775 69.160 ;
        RECT 70.950 68.085 71.210 69.235 ;
        RECT 71.970 69.185 72.140 69.330 ;
        RECT 71.475 69.015 72.140 69.185 ;
        RECT 72.425 69.160 72.595 69.960 ;
        RECT 72.765 69.865 76.275 70.635 ;
        RECT 76.450 69.895 76.705 70.465 ;
        RECT 76.875 70.235 77.205 70.635 ;
        RECT 77.630 70.100 78.160 70.465 ;
        RECT 77.630 70.065 77.805 70.100 ;
        RECT 76.875 69.895 77.805 70.065 ;
        RECT 72.765 69.345 74.415 69.865 ;
        RECT 74.585 69.175 76.275 69.695 ;
        RECT 71.475 68.255 71.645 69.015 ;
        RECT 71.825 68.085 72.155 68.845 ;
        RECT 72.325 68.255 72.595 69.160 ;
        RECT 72.765 68.085 76.275 69.175 ;
        RECT 76.450 69.225 76.620 69.895 ;
        RECT 76.875 69.725 77.045 69.895 ;
        RECT 76.790 69.395 77.045 69.725 ;
        RECT 77.270 69.395 77.465 69.725 ;
        RECT 76.450 68.255 76.785 69.225 ;
        RECT 76.955 68.085 77.125 69.225 ;
        RECT 77.295 68.425 77.465 69.395 ;
        RECT 77.635 68.765 77.805 69.895 ;
        RECT 77.975 69.105 78.145 69.905 ;
        RECT 78.350 69.615 78.625 70.465 ;
        RECT 78.345 69.445 78.625 69.615 ;
        RECT 78.350 69.305 78.625 69.445 ;
        RECT 78.795 69.105 78.985 70.465 ;
        RECT 79.165 70.100 79.675 70.635 ;
        RECT 79.895 69.825 80.140 70.430 ;
        RECT 79.185 69.655 80.415 69.825 ;
        RECT 80.645 69.815 80.855 70.635 ;
        RECT 81.025 69.835 81.355 70.465 ;
        RECT 77.975 68.935 78.985 69.105 ;
        RECT 79.155 69.090 79.905 69.280 ;
        RECT 77.635 68.595 78.760 68.765 ;
        RECT 79.155 68.425 79.325 69.090 ;
        RECT 80.075 68.845 80.415 69.655 ;
        RECT 81.025 69.235 81.275 69.835 ;
        RECT 81.525 69.815 81.755 70.635 ;
        RECT 82.885 69.910 83.175 70.635 ;
        RECT 83.345 70.090 88.690 70.635 ;
        RECT 81.445 69.395 81.775 69.645 ;
        RECT 84.930 69.260 85.270 70.090 ;
        RECT 88.865 69.865 90.535 70.635 ;
        RECT 77.295 68.255 79.325 68.425 ;
        RECT 79.495 68.085 79.665 68.845 ;
        RECT 79.900 68.435 80.415 68.845 ;
        RECT 80.645 68.085 80.855 69.225 ;
        RECT 81.025 68.255 81.355 69.235 ;
        RECT 81.525 68.085 81.755 69.225 ;
        RECT 82.885 68.085 83.175 69.250 ;
        RECT 86.750 68.520 87.100 69.770 ;
        RECT 88.865 69.345 89.615 69.865 ;
        RECT 90.705 69.835 91.045 70.465 ;
        RECT 91.215 69.835 91.465 70.635 ;
        RECT 91.655 69.985 91.985 70.465 ;
        RECT 92.155 70.175 92.380 70.635 ;
        RECT 92.550 69.985 92.880 70.465 ;
        RECT 89.785 69.175 90.535 69.695 ;
        RECT 83.345 68.085 88.690 68.520 ;
        RECT 88.865 68.085 90.535 69.175 ;
        RECT 90.705 69.225 90.880 69.835 ;
        RECT 91.655 69.815 92.880 69.985 ;
        RECT 93.510 69.855 94.010 70.465 ;
        RECT 91.050 69.475 91.745 69.645 ;
        RECT 91.575 69.225 91.745 69.475 ;
        RECT 91.920 69.445 92.340 69.645 ;
        RECT 92.510 69.445 92.840 69.645 ;
        RECT 93.010 69.445 93.340 69.645 ;
        RECT 93.510 69.225 93.680 69.855 ;
        RECT 94.385 69.835 94.725 70.465 ;
        RECT 94.895 69.835 95.145 70.635 ;
        RECT 95.335 69.985 95.665 70.465 ;
        RECT 95.835 70.175 96.060 70.635 ;
        RECT 96.230 69.985 96.560 70.465 ;
        RECT 93.865 69.395 94.215 69.645 ;
        RECT 94.385 69.225 94.560 69.835 ;
        RECT 95.335 69.815 96.560 69.985 ;
        RECT 97.190 69.855 97.690 70.465 ;
        RECT 98.270 69.855 98.770 70.465 ;
        RECT 94.730 69.475 95.425 69.645 ;
        RECT 95.255 69.225 95.425 69.475 ;
        RECT 95.600 69.445 96.020 69.645 ;
        RECT 96.190 69.445 96.520 69.645 ;
        RECT 96.690 69.445 97.020 69.645 ;
        RECT 97.190 69.225 97.360 69.855 ;
        RECT 97.545 69.395 97.895 69.645 ;
        RECT 98.065 69.395 98.415 69.645 ;
        RECT 98.600 69.225 98.770 69.855 ;
        RECT 99.400 69.985 99.730 70.465 ;
        RECT 99.900 70.175 100.125 70.635 ;
        RECT 100.295 69.985 100.625 70.465 ;
        RECT 99.400 69.815 100.625 69.985 ;
        RECT 100.815 69.835 101.065 70.635 ;
        RECT 101.235 69.835 101.575 70.465 ;
        RECT 98.940 69.445 99.270 69.645 ;
        RECT 99.440 69.445 99.770 69.645 ;
        RECT 99.940 69.445 100.360 69.645 ;
        RECT 100.535 69.475 101.230 69.645 ;
        RECT 100.535 69.225 100.705 69.475 ;
        RECT 101.400 69.275 101.575 69.835 ;
        RECT 101.345 69.225 101.575 69.275 ;
        RECT 90.705 68.255 91.045 69.225 ;
        RECT 91.215 68.085 91.385 69.225 ;
        RECT 91.575 69.055 94.010 69.225 ;
        RECT 91.655 68.085 91.905 68.885 ;
        RECT 92.550 68.255 92.880 69.055 ;
        RECT 93.180 68.085 93.510 68.885 ;
        RECT 93.680 68.255 94.010 69.055 ;
        RECT 94.385 68.255 94.725 69.225 ;
        RECT 94.895 68.085 95.065 69.225 ;
        RECT 95.255 69.055 97.690 69.225 ;
        RECT 95.335 68.085 95.585 68.885 ;
        RECT 96.230 68.255 96.560 69.055 ;
        RECT 96.860 68.085 97.190 68.885 ;
        RECT 97.360 68.255 97.690 69.055 ;
        RECT 98.270 69.055 100.705 69.225 ;
        RECT 98.270 68.255 98.600 69.055 ;
        RECT 98.770 68.085 99.100 68.885 ;
        RECT 99.400 68.255 99.730 69.055 ;
        RECT 100.375 68.085 100.625 68.885 ;
        RECT 100.895 68.085 101.065 69.225 ;
        RECT 101.235 68.255 101.575 69.225 ;
        RECT 101.750 69.895 102.005 70.465 ;
        RECT 102.175 70.235 102.505 70.635 ;
        RECT 102.930 70.100 103.460 70.465 ;
        RECT 103.650 70.295 103.925 70.465 ;
        RECT 103.645 70.125 103.925 70.295 ;
        RECT 102.930 70.065 103.105 70.100 ;
        RECT 102.175 69.895 103.105 70.065 ;
        RECT 101.750 69.225 101.920 69.895 ;
        RECT 102.175 69.725 102.345 69.895 ;
        RECT 102.090 69.395 102.345 69.725 ;
        RECT 102.570 69.395 102.765 69.725 ;
        RECT 101.750 68.255 102.085 69.225 ;
        RECT 102.255 68.085 102.425 69.225 ;
        RECT 102.595 68.425 102.765 69.395 ;
        RECT 102.935 68.765 103.105 69.895 ;
        RECT 103.275 69.105 103.445 69.905 ;
        RECT 103.650 69.305 103.925 70.125 ;
        RECT 104.095 69.105 104.285 70.465 ;
        RECT 104.465 70.100 104.975 70.635 ;
        RECT 105.195 69.825 105.440 70.430 ;
        RECT 105.885 69.865 108.475 70.635 ;
        RECT 108.645 69.910 108.935 70.635 ;
        RECT 109.105 69.865 110.775 70.635 ;
        RECT 111.495 70.085 111.665 70.375 ;
        RECT 111.835 70.255 112.165 70.635 ;
        RECT 111.495 69.915 112.160 70.085 ;
        RECT 104.485 69.655 105.715 69.825 ;
        RECT 103.275 68.935 104.285 69.105 ;
        RECT 104.455 69.090 105.205 69.280 ;
        RECT 102.935 68.595 104.060 68.765 ;
        RECT 104.455 68.425 104.625 69.090 ;
        RECT 105.375 68.845 105.715 69.655 ;
        RECT 105.885 69.345 107.095 69.865 ;
        RECT 107.265 69.175 108.475 69.695 ;
        RECT 109.105 69.345 109.855 69.865 ;
        RECT 102.595 68.255 104.625 68.425 ;
        RECT 104.795 68.085 104.965 68.845 ;
        RECT 105.200 68.435 105.715 68.845 ;
        RECT 105.885 68.085 108.475 69.175 ;
        RECT 108.645 68.085 108.935 69.250 ;
        RECT 110.025 69.175 110.775 69.695 ;
        RECT 109.105 68.085 110.775 69.175 ;
        RECT 111.410 69.095 111.760 69.745 ;
        RECT 111.930 68.925 112.160 69.915 ;
        RECT 111.495 68.755 112.160 68.925 ;
        RECT 111.495 68.255 111.665 68.755 ;
        RECT 111.835 68.085 112.165 68.585 ;
        RECT 112.335 68.255 112.560 70.375 ;
        RECT 112.775 70.255 113.105 70.635 ;
        RECT 113.275 70.085 113.445 70.415 ;
        RECT 113.745 70.255 114.760 70.455 ;
        RECT 112.750 69.895 113.445 70.085 ;
        RECT 112.750 68.925 112.920 69.895 ;
        RECT 113.090 69.095 113.500 69.715 ;
        RECT 113.670 69.145 113.890 70.015 ;
        RECT 114.070 69.705 114.420 70.075 ;
        RECT 114.590 69.525 114.760 70.255 ;
        RECT 114.930 70.195 115.340 70.635 ;
        RECT 115.630 69.995 115.880 70.425 ;
        RECT 116.080 70.175 116.400 70.635 ;
        RECT 116.960 70.245 117.810 70.415 ;
        RECT 114.930 69.655 115.340 69.985 ;
        RECT 115.630 69.655 116.050 69.995 ;
        RECT 114.340 69.485 114.760 69.525 ;
        RECT 114.340 69.315 115.690 69.485 ;
        RECT 112.750 68.755 113.445 68.925 ;
        RECT 113.670 68.765 114.170 69.145 ;
        RECT 112.775 68.085 113.105 68.585 ;
        RECT 113.275 68.255 113.445 68.755 ;
        RECT 114.340 68.470 114.510 69.315 ;
        RECT 115.440 69.155 115.690 69.315 ;
        RECT 114.680 68.885 114.930 69.145 ;
        RECT 115.860 68.885 116.050 69.655 ;
        RECT 114.680 68.635 116.050 68.885 ;
        RECT 116.220 69.825 117.470 69.995 ;
        RECT 116.220 69.065 116.390 69.825 ;
        RECT 117.140 69.705 117.470 69.825 ;
        RECT 116.560 69.245 116.740 69.655 ;
        RECT 117.640 69.485 117.810 70.245 ;
        RECT 118.010 70.155 118.670 70.635 ;
        RECT 118.850 70.040 119.170 70.370 ;
        RECT 118.000 69.715 118.660 69.985 ;
        RECT 118.000 69.655 118.330 69.715 ;
        RECT 118.480 69.485 118.810 69.545 ;
        RECT 116.910 69.315 118.810 69.485 ;
        RECT 116.220 68.755 116.740 69.065 ;
        RECT 116.910 68.805 117.080 69.315 ;
        RECT 118.980 69.145 119.170 70.040 ;
        RECT 117.250 68.975 119.170 69.145 ;
        RECT 118.850 68.955 119.170 68.975 ;
        RECT 119.370 69.725 119.620 70.375 ;
        RECT 119.800 70.175 120.085 70.635 ;
        RECT 120.265 70.295 120.520 70.455 ;
        RECT 120.265 70.125 120.605 70.295 ;
        RECT 120.265 69.925 120.520 70.125 ;
        RECT 119.370 69.395 120.170 69.725 ;
        RECT 116.910 68.635 118.120 68.805 ;
        RECT 113.680 68.300 114.510 68.470 ;
        RECT 114.750 68.085 115.130 68.465 ;
        RECT 115.310 68.345 115.480 68.635 ;
        RECT 116.910 68.555 117.080 68.635 ;
        RECT 115.650 68.085 115.980 68.465 ;
        RECT 116.450 68.305 117.080 68.555 ;
        RECT 117.260 68.085 117.680 68.465 ;
        RECT 117.880 68.345 118.120 68.635 ;
        RECT 118.350 68.085 118.680 68.775 ;
        RECT 118.850 68.345 119.020 68.955 ;
        RECT 119.370 68.805 119.620 69.395 ;
        RECT 120.340 69.065 120.520 69.925 ;
        RECT 121.065 69.885 122.275 70.635 ;
        RECT 122.445 69.885 123.655 70.635 ;
        RECT 121.065 69.345 121.585 69.885 ;
        RECT 121.755 69.175 122.275 69.715 ;
        RECT 119.290 68.295 119.620 68.805 ;
        RECT 119.800 68.085 120.085 68.885 ;
        RECT 120.265 68.395 120.520 69.065 ;
        RECT 121.065 68.085 122.275 69.175 ;
        RECT 122.445 69.175 122.965 69.715 ;
        RECT 123.135 69.345 123.655 69.885 ;
        RECT 122.445 68.085 123.655 69.175 ;
        RECT 5.520 67.915 123.740 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 6.985 67.480 12.330 67.915 ;
        RECT 12.505 67.480 17.850 67.915 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 8.570 65.910 8.910 66.740 ;
        RECT 10.390 66.230 10.740 67.480 ;
        RECT 14.090 65.910 14.430 66.740 ;
        RECT 15.910 66.230 16.260 67.480 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.945 67.480 24.290 67.915 ;
        RECT 6.985 65.365 12.330 65.910 ;
        RECT 12.505 65.365 17.850 65.910 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 20.530 65.910 20.870 66.740 ;
        RECT 22.350 66.230 22.700 67.480 ;
        RECT 24.465 66.825 27.975 67.915 ;
        RECT 24.465 66.135 26.115 66.655 ;
        RECT 26.285 66.305 27.975 66.825 ;
        RECT 28.145 66.840 28.415 67.745 ;
        RECT 28.585 67.155 28.915 67.915 ;
        RECT 29.095 66.985 29.265 67.745 ;
        RECT 18.945 65.365 24.290 65.910 ;
        RECT 24.465 65.365 27.975 66.135 ;
        RECT 28.145 66.040 28.315 66.840 ;
        RECT 28.600 66.815 29.265 66.985 ;
        RECT 28.600 66.670 28.770 66.815 ;
        RECT 28.485 66.340 28.770 66.670 ;
        RECT 29.530 66.775 29.865 67.745 ;
        RECT 30.035 66.775 30.205 67.915 ;
        RECT 30.375 67.575 32.405 67.745 ;
        RECT 28.600 66.085 28.770 66.340 ;
        RECT 29.005 66.265 29.335 66.635 ;
        RECT 29.530 66.105 29.700 66.775 ;
        RECT 30.375 66.605 30.545 67.575 ;
        RECT 29.870 66.275 30.125 66.605 ;
        RECT 30.350 66.275 30.545 66.605 ;
        RECT 30.715 67.235 31.840 67.405 ;
        RECT 29.955 66.105 30.125 66.275 ;
        RECT 30.715 66.105 30.885 67.235 ;
        RECT 28.145 65.535 28.405 66.040 ;
        RECT 28.600 65.915 29.265 66.085 ;
        RECT 28.585 65.365 28.915 65.745 ;
        RECT 29.095 65.535 29.265 65.915 ;
        RECT 29.530 65.535 29.785 66.105 ;
        RECT 29.955 65.935 30.885 66.105 ;
        RECT 31.055 66.895 32.065 67.065 ;
        RECT 31.055 66.095 31.225 66.895 ;
        RECT 31.430 66.555 31.705 66.695 ;
        RECT 31.425 66.385 31.705 66.555 ;
        RECT 30.710 65.900 30.885 65.935 ;
        RECT 29.955 65.365 30.285 65.765 ;
        RECT 30.710 65.535 31.240 65.900 ;
        RECT 31.430 65.535 31.705 66.385 ;
        RECT 31.875 65.535 32.065 66.895 ;
        RECT 32.235 66.910 32.405 67.575 ;
        RECT 32.575 67.155 32.745 67.915 ;
        RECT 32.980 67.155 33.495 67.565 ;
        RECT 32.235 66.720 32.985 66.910 ;
        RECT 33.155 66.345 33.495 67.155 ;
        RECT 34.675 67.245 34.845 67.745 ;
        RECT 35.015 67.415 35.345 67.915 ;
        RECT 34.675 67.075 35.340 67.245 ;
        RECT 32.265 66.175 33.495 66.345 ;
        RECT 34.590 66.255 34.940 66.905 ;
        RECT 32.245 65.365 32.755 65.900 ;
        RECT 32.975 65.570 33.220 66.175 ;
        RECT 35.110 66.085 35.340 67.075 ;
        RECT 34.675 65.915 35.340 66.085 ;
        RECT 34.675 65.625 34.845 65.915 ;
        RECT 35.015 65.365 35.345 65.745 ;
        RECT 35.515 65.625 35.740 67.745 ;
        RECT 35.955 67.415 36.285 67.915 ;
        RECT 36.455 67.245 36.625 67.745 ;
        RECT 36.860 67.530 37.690 67.700 ;
        RECT 37.930 67.535 38.310 67.915 ;
        RECT 35.930 67.075 36.625 67.245 ;
        RECT 35.930 66.105 36.100 67.075 ;
        RECT 36.270 66.285 36.680 66.905 ;
        RECT 36.850 66.855 37.350 67.235 ;
        RECT 35.930 65.915 36.625 66.105 ;
        RECT 36.850 65.985 37.070 66.855 ;
        RECT 37.520 66.685 37.690 67.530 ;
        RECT 38.490 67.365 38.660 67.655 ;
        RECT 38.830 67.535 39.160 67.915 ;
        RECT 39.630 67.445 40.260 67.695 ;
        RECT 40.440 67.535 40.860 67.915 ;
        RECT 40.090 67.365 40.260 67.445 ;
        RECT 41.060 67.365 41.300 67.655 ;
        RECT 37.860 67.115 39.230 67.365 ;
        RECT 37.860 66.855 38.110 67.115 ;
        RECT 38.620 66.685 38.870 66.845 ;
        RECT 37.520 66.515 38.870 66.685 ;
        RECT 37.520 66.475 37.940 66.515 ;
        RECT 37.250 65.925 37.600 66.295 ;
        RECT 35.955 65.365 36.285 65.745 ;
        RECT 36.455 65.585 36.625 65.915 ;
        RECT 37.770 65.745 37.940 66.475 ;
        RECT 39.040 66.345 39.230 67.115 ;
        RECT 38.110 66.015 38.520 66.345 ;
        RECT 38.810 66.005 39.230 66.345 ;
        RECT 39.400 66.935 39.920 67.245 ;
        RECT 40.090 67.195 41.300 67.365 ;
        RECT 41.530 67.225 41.860 67.915 ;
        RECT 39.400 66.175 39.570 66.935 ;
        RECT 39.740 66.345 39.920 66.755 ;
        RECT 40.090 66.685 40.260 67.195 ;
        RECT 42.030 67.045 42.200 67.655 ;
        RECT 42.470 67.195 42.800 67.705 ;
        RECT 42.030 67.025 42.350 67.045 ;
        RECT 40.430 66.855 42.350 67.025 ;
        RECT 40.090 66.515 41.990 66.685 ;
        RECT 40.320 66.175 40.650 66.295 ;
        RECT 39.400 66.005 40.650 66.175 ;
        RECT 36.925 65.545 37.940 65.745 ;
        RECT 38.110 65.365 38.520 65.805 ;
        RECT 38.810 65.575 39.060 66.005 ;
        RECT 39.260 65.365 39.580 65.825 ;
        RECT 40.820 65.755 40.990 66.515 ;
        RECT 41.660 66.455 41.990 66.515 ;
        RECT 41.180 66.285 41.510 66.345 ;
        RECT 41.180 66.015 41.840 66.285 ;
        RECT 42.160 65.960 42.350 66.855 ;
        RECT 40.140 65.585 40.990 65.755 ;
        RECT 41.190 65.365 41.850 65.845 ;
        RECT 42.030 65.630 42.350 65.960 ;
        RECT 42.550 66.605 42.800 67.195 ;
        RECT 42.980 67.115 43.265 67.915 ;
        RECT 43.445 66.935 43.700 67.605 ;
        RECT 42.550 66.275 43.350 66.605 ;
        RECT 42.550 65.625 42.800 66.275 ;
        RECT 43.520 66.215 43.700 66.935 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.705 66.825 47.295 67.915 ;
        RECT 43.520 66.075 43.785 66.215 ;
        RECT 44.705 66.135 45.915 66.655 ;
        RECT 46.085 66.305 47.295 66.825 ;
        RECT 47.465 66.840 47.735 67.745 ;
        RECT 47.905 67.155 48.235 67.915 ;
        RECT 48.415 66.985 48.585 67.745 ;
        RECT 43.445 66.045 43.785 66.075 ;
        RECT 42.980 65.365 43.265 65.825 ;
        RECT 43.445 65.545 43.700 66.045 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 44.705 65.365 47.295 66.135 ;
        RECT 47.465 66.040 47.635 66.840 ;
        RECT 47.920 66.815 48.585 66.985 ;
        RECT 47.920 66.670 48.090 66.815 ;
        RECT 47.805 66.340 48.090 66.670 ;
        RECT 48.850 66.775 49.185 67.745 ;
        RECT 49.355 66.775 49.525 67.915 ;
        RECT 49.695 67.575 51.725 67.745 ;
        RECT 47.920 66.085 48.090 66.340 ;
        RECT 48.325 66.265 48.655 66.635 ;
        RECT 48.850 66.105 49.020 66.775 ;
        RECT 49.695 66.605 49.865 67.575 ;
        RECT 49.190 66.275 49.445 66.605 ;
        RECT 49.670 66.275 49.865 66.605 ;
        RECT 50.035 67.235 51.160 67.405 ;
        RECT 49.275 66.105 49.445 66.275 ;
        RECT 50.035 66.105 50.205 67.235 ;
        RECT 47.465 65.535 47.725 66.040 ;
        RECT 47.920 65.915 48.585 66.085 ;
        RECT 47.905 65.365 48.235 65.745 ;
        RECT 48.415 65.535 48.585 65.915 ;
        RECT 48.850 65.535 49.105 66.105 ;
        RECT 49.275 65.935 50.205 66.105 ;
        RECT 50.375 66.895 51.385 67.065 ;
        RECT 50.375 66.095 50.545 66.895 ;
        RECT 50.750 66.555 51.025 66.695 ;
        RECT 50.745 66.385 51.025 66.555 ;
        RECT 50.030 65.900 50.205 65.935 ;
        RECT 49.275 65.365 49.605 65.765 ;
        RECT 50.030 65.535 50.560 65.900 ;
        RECT 50.750 65.535 51.025 66.385 ;
        RECT 51.195 65.535 51.385 66.895 ;
        RECT 51.555 66.910 51.725 67.575 ;
        RECT 51.895 67.155 52.065 67.915 ;
        RECT 52.300 67.155 52.815 67.565 ;
        RECT 52.985 67.480 58.330 67.915 ;
        RECT 51.555 66.720 52.305 66.910 ;
        RECT 52.475 66.345 52.815 67.155 ;
        RECT 51.585 66.175 52.815 66.345 ;
        RECT 51.565 65.365 52.075 65.900 ;
        RECT 52.295 65.570 52.540 66.175 ;
        RECT 54.570 65.910 54.910 66.740 ;
        RECT 56.390 66.230 56.740 67.480 ;
        RECT 58.505 66.825 62.015 67.915 ;
        RECT 58.505 66.135 60.155 66.655 ;
        RECT 60.325 66.305 62.015 66.825 ;
        RECT 62.650 66.765 62.910 67.915 ;
        RECT 63.085 66.840 63.340 67.745 ;
        RECT 63.510 67.155 63.840 67.915 ;
        RECT 64.055 66.985 64.225 67.745 ;
        RECT 52.985 65.365 58.330 65.910 ;
        RECT 58.505 65.365 62.015 66.135 ;
        RECT 62.650 65.365 62.910 66.205 ;
        RECT 63.085 66.110 63.255 66.840 ;
        RECT 63.510 66.815 64.225 66.985 ;
        RECT 63.510 66.605 63.680 66.815 ;
        RECT 64.490 66.765 64.750 67.915 ;
        RECT 64.925 66.840 65.180 67.745 ;
        RECT 65.350 67.155 65.680 67.915 ;
        RECT 65.895 66.985 66.065 67.745 ;
        RECT 63.425 66.275 63.680 66.605 ;
        RECT 63.085 65.535 63.340 66.110 ;
        RECT 63.510 66.085 63.680 66.275 ;
        RECT 63.960 66.265 64.315 66.635 ;
        RECT 63.510 65.915 64.225 66.085 ;
        RECT 63.510 65.365 63.840 65.745 ;
        RECT 64.055 65.535 64.225 65.915 ;
        RECT 64.490 65.365 64.750 66.205 ;
        RECT 64.925 66.110 65.095 66.840 ;
        RECT 65.350 66.815 66.065 66.985 ;
        RECT 66.325 66.825 67.535 67.915 ;
        RECT 65.350 66.605 65.520 66.815 ;
        RECT 65.265 66.275 65.520 66.605 ;
        RECT 64.925 65.535 65.180 66.110 ;
        RECT 65.350 66.085 65.520 66.275 ;
        RECT 65.800 66.265 66.155 66.635 ;
        RECT 66.325 66.115 66.845 66.655 ;
        RECT 67.015 66.285 67.535 66.825 ;
        RECT 67.710 66.765 67.970 67.915 ;
        RECT 68.145 66.840 68.400 67.745 ;
        RECT 68.570 67.155 68.900 67.915 ;
        RECT 69.115 66.985 69.285 67.745 ;
        RECT 65.350 65.915 66.065 66.085 ;
        RECT 65.350 65.365 65.680 65.745 ;
        RECT 65.895 65.535 66.065 65.915 ;
        RECT 66.325 65.365 67.535 66.115 ;
        RECT 67.710 65.365 67.970 66.205 ;
        RECT 68.145 66.110 68.315 66.840 ;
        RECT 68.570 66.815 69.285 66.985 ;
        RECT 68.570 66.605 68.740 66.815 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 70.465 66.825 72.135 67.915 ;
        RECT 68.485 66.275 68.740 66.605 ;
        RECT 68.145 65.535 68.400 66.110 ;
        RECT 68.570 66.085 68.740 66.275 ;
        RECT 69.020 66.265 69.375 66.635 ;
        RECT 70.465 66.135 71.215 66.655 ;
        RECT 71.385 66.305 72.135 66.825 ;
        RECT 72.395 66.985 72.565 67.745 ;
        RECT 72.745 67.155 73.075 67.915 ;
        RECT 72.395 66.815 73.060 66.985 ;
        RECT 73.245 66.840 73.515 67.745 ;
        RECT 73.775 67.245 73.945 67.745 ;
        RECT 74.115 67.415 74.445 67.915 ;
        RECT 73.775 67.075 74.440 67.245 ;
        RECT 72.890 66.670 73.060 66.815 ;
        RECT 72.325 66.265 72.655 66.635 ;
        RECT 72.890 66.340 73.175 66.670 ;
        RECT 68.570 65.915 69.285 66.085 ;
        RECT 68.570 65.365 68.900 65.745 ;
        RECT 69.115 65.535 69.285 65.915 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 70.465 65.365 72.135 66.135 ;
        RECT 72.890 66.085 73.060 66.340 ;
        RECT 72.395 65.915 73.060 66.085 ;
        RECT 73.345 66.040 73.515 66.840 ;
        RECT 73.690 66.255 74.040 66.905 ;
        RECT 74.210 66.085 74.440 67.075 ;
        RECT 72.395 65.535 72.565 65.915 ;
        RECT 72.745 65.365 73.075 65.745 ;
        RECT 73.255 65.535 73.515 66.040 ;
        RECT 73.775 65.915 74.440 66.085 ;
        RECT 73.775 65.625 73.945 65.915 ;
        RECT 74.115 65.365 74.445 65.745 ;
        RECT 74.615 65.625 74.840 67.745 ;
        RECT 75.055 67.415 75.385 67.915 ;
        RECT 75.555 67.245 75.725 67.745 ;
        RECT 75.960 67.530 76.790 67.700 ;
        RECT 77.030 67.535 77.410 67.915 ;
        RECT 75.030 67.075 75.725 67.245 ;
        RECT 75.030 66.105 75.200 67.075 ;
        RECT 75.370 66.285 75.780 66.905 ;
        RECT 75.950 66.855 76.450 67.235 ;
        RECT 75.030 65.915 75.725 66.105 ;
        RECT 75.950 65.985 76.170 66.855 ;
        RECT 76.620 66.685 76.790 67.530 ;
        RECT 77.590 67.365 77.760 67.655 ;
        RECT 77.930 67.535 78.260 67.915 ;
        RECT 78.730 67.445 79.360 67.695 ;
        RECT 79.540 67.535 79.960 67.915 ;
        RECT 79.190 67.365 79.360 67.445 ;
        RECT 80.160 67.365 80.400 67.655 ;
        RECT 76.960 67.115 78.330 67.365 ;
        RECT 76.960 66.855 77.210 67.115 ;
        RECT 77.720 66.685 77.970 66.845 ;
        RECT 76.620 66.515 77.970 66.685 ;
        RECT 76.620 66.475 77.040 66.515 ;
        RECT 76.350 65.925 76.700 66.295 ;
        RECT 75.055 65.365 75.385 65.745 ;
        RECT 75.555 65.585 75.725 65.915 ;
        RECT 76.870 65.745 77.040 66.475 ;
        RECT 78.140 66.345 78.330 67.115 ;
        RECT 77.210 66.015 77.620 66.345 ;
        RECT 77.910 66.005 78.330 66.345 ;
        RECT 78.500 66.935 79.020 67.245 ;
        RECT 79.190 67.195 80.400 67.365 ;
        RECT 80.630 67.225 80.960 67.915 ;
        RECT 78.500 66.175 78.670 66.935 ;
        RECT 78.840 66.345 79.020 66.755 ;
        RECT 79.190 66.685 79.360 67.195 ;
        RECT 81.130 67.045 81.300 67.655 ;
        RECT 81.570 67.195 81.900 67.705 ;
        RECT 81.130 67.025 81.450 67.045 ;
        RECT 79.530 66.855 81.450 67.025 ;
        RECT 79.190 66.515 81.090 66.685 ;
        RECT 79.420 66.175 79.750 66.295 ;
        RECT 78.500 66.005 79.750 66.175 ;
        RECT 76.025 65.545 77.040 65.745 ;
        RECT 77.210 65.365 77.620 65.805 ;
        RECT 77.910 65.575 78.160 66.005 ;
        RECT 78.360 65.365 78.680 65.825 ;
        RECT 79.920 65.755 80.090 66.515 ;
        RECT 80.760 66.455 81.090 66.515 ;
        RECT 80.280 66.285 80.610 66.345 ;
        RECT 80.280 66.015 80.940 66.285 ;
        RECT 81.260 65.960 81.450 66.855 ;
        RECT 79.240 65.585 80.090 65.755 ;
        RECT 80.290 65.365 80.950 65.845 ;
        RECT 81.130 65.630 81.450 65.960 ;
        RECT 81.650 66.605 81.900 67.195 ;
        RECT 82.080 67.115 82.365 67.915 ;
        RECT 82.545 67.575 82.800 67.605 ;
        RECT 82.545 67.405 82.885 67.575 ;
        RECT 82.545 66.935 82.800 67.405 ;
        RECT 81.650 66.275 82.450 66.605 ;
        RECT 81.650 65.625 81.900 66.275 ;
        RECT 82.620 66.075 82.800 66.935 ;
        RECT 83.355 66.935 83.685 67.745 ;
        RECT 83.855 67.115 84.095 67.915 ;
        RECT 83.355 66.765 84.070 66.935 ;
        RECT 83.350 66.355 83.730 66.595 ;
        RECT 83.900 66.525 84.070 66.765 ;
        RECT 84.275 66.895 84.445 67.745 ;
        RECT 84.615 67.115 84.945 67.915 ;
        RECT 85.115 66.895 85.285 67.745 ;
        RECT 84.275 66.725 85.285 66.895 ;
        RECT 85.455 66.765 85.785 67.915 ;
        RECT 86.105 66.825 89.615 67.915 ;
        RECT 83.900 66.355 84.400 66.525 ;
        RECT 83.900 66.185 84.070 66.355 ;
        RECT 84.790 66.185 85.285 66.725 ;
        RECT 82.080 65.365 82.365 65.825 ;
        RECT 82.545 65.545 82.800 66.075 ;
        RECT 83.435 66.015 84.070 66.185 ;
        RECT 84.275 66.015 85.285 66.185 ;
        RECT 83.435 65.535 83.605 66.015 ;
        RECT 83.785 65.365 84.025 65.845 ;
        RECT 84.275 65.535 84.445 66.015 ;
        RECT 84.615 65.365 84.945 65.845 ;
        RECT 85.115 65.535 85.285 66.015 ;
        RECT 85.455 65.365 85.785 66.165 ;
        RECT 86.105 66.135 87.755 66.655 ;
        RECT 87.925 66.305 89.615 66.825 ;
        RECT 90.250 66.775 90.585 67.745 ;
        RECT 90.755 66.775 90.925 67.915 ;
        RECT 91.095 67.575 93.125 67.745 ;
        RECT 86.105 65.365 89.615 66.135 ;
        RECT 90.250 66.105 90.420 66.775 ;
        RECT 91.095 66.605 91.265 67.575 ;
        RECT 90.590 66.275 90.845 66.605 ;
        RECT 91.070 66.275 91.265 66.605 ;
        RECT 91.435 67.235 92.560 67.405 ;
        RECT 90.675 66.105 90.845 66.275 ;
        RECT 91.435 66.105 91.605 67.235 ;
        RECT 90.250 65.535 90.505 66.105 ;
        RECT 90.675 65.935 91.605 66.105 ;
        RECT 91.775 66.895 92.785 67.065 ;
        RECT 91.775 66.095 91.945 66.895 ;
        RECT 92.150 66.555 92.425 66.695 ;
        RECT 92.145 66.385 92.425 66.555 ;
        RECT 91.430 65.900 91.605 65.935 ;
        RECT 90.675 65.365 91.005 65.765 ;
        RECT 91.430 65.535 91.960 65.900 ;
        RECT 92.150 65.535 92.425 66.385 ;
        RECT 92.595 65.535 92.785 66.895 ;
        RECT 92.955 66.910 93.125 67.575 ;
        RECT 93.295 67.155 93.465 67.915 ;
        RECT 93.700 67.155 94.215 67.565 ;
        RECT 92.955 66.720 93.705 66.910 ;
        RECT 93.875 66.345 94.215 67.155 ;
        RECT 94.385 66.825 95.595 67.915 ;
        RECT 92.985 66.175 94.215 66.345 ;
        RECT 92.965 65.365 93.475 65.900 ;
        RECT 93.695 65.570 93.940 66.175 ;
        RECT 94.385 66.115 94.905 66.655 ;
        RECT 95.075 66.285 95.595 66.825 ;
        RECT 95.765 66.750 96.055 67.915 ;
        RECT 96.225 67.480 101.570 67.915 ;
        RECT 101.745 67.480 107.090 67.915 ;
        RECT 107.265 67.480 112.610 67.915 ;
        RECT 94.385 65.365 95.595 66.115 ;
        RECT 95.765 65.365 96.055 66.090 ;
        RECT 97.810 65.910 98.150 66.740 ;
        RECT 99.630 66.230 99.980 67.480 ;
        RECT 103.330 65.910 103.670 66.740 ;
        RECT 105.150 66.230 105.500 67.480 ;
        RECT 108.850 65.910 109.190 66.740 ;
        RECT 110.670 66.230 111.020 67.480 ;
        RECT 112.785 67.155 113.300 67.565 ;
        RECT 113.535 67.155 113.705 67.915 ;
        RECT 113.875 67.575 115.905 67.745 ;
        RECT 112.785 66.345 113.125 67.155 ;
        RECT 113.875 66.910 114.045 67.575 ;
        RECT 114.440 67.235 115.565 67.405 ;
        RECT 113.295 66.720 114.045 66.910 ;
        RECT 114.215 66.895 115.225 67.065 ;
        RECT 112.785 66.175 114.015 66.345 ;
        RECT 96.225 65.365 101.570 65.910 ;
        RECT 101.745 65.365 107.090 65.910 ;
        RECT 107.265 65.365 112.610 65.910 ;
        RECT 113.060 65.570 113.305 66.175 ;
        RECT 113.525 65.365 114.035 65.900 ;
        RECT 114.215 65.535 114.405 66.895 ;
        RECT 114.575 65.875 114.850 66.695 ;
        RECT 115.055 66.095 115.225 66.895 ;
        RECT 115.395 66.105 115.565 67.235 ;
        RECT 115.735 66.605 115.905 67.575 ;
        RECT 116.075 66.775 116.245 67.915 ;
        RECT 116.415 66.775 116.750 67.745 ;
        RECT 116.985 66.775 117.195 67.915 ;
        RECT 115.735 66.275 115.930 66.605 ;
        RECT 116.155 66.275 116.410 66.605 ;
        RECT 116.155 66.105 116.325 66.275 ;
        RECT 116.580 66.105 116.750 66.775 ;
        RECT 117.365 66.765 117.695 67.745 ;
        RECT 117.865 66.775 118.095 67.915 ;
        RECT 118.305 66.825 120.895 67.915 ;
        RECT 115.395 65.935 116.325 66.105 ;
        RECT 115.395 65.900 115.570 65.935 ;
        RECT 114.575 65.705 114.855 65.875 ;
        RECT 114.575 65.535 114.850 65.705 ;
        RECT 115.040 65.535 115.570 65.900 ;
        RECT 115.995 65.365 116.325 65.765 ;
        RECT 116.495 65.535 116.750 66.105 ;
        RECT 116.985 65.365 117.195 66.185 ;
        RECT 117.365 66.165 117.615 66.765 ;
        RECT 117.785 66.355 118.115 66.605 ;
        RECT 117.365 65.535 117.695 66.165 ;
        RECT 117.865 65.365 118.095 66.185 ;
        RECT 118.305 66.135 119.515 66.655 ;
        RECT 119.685 66.305 120.895 66.825 ;
        RECT 121.525 66.750 121.815 67.915 ;
        RECT 122.445 66.825 123.655 67.915 ;
        RECT 122.445 66.285 122.965 66.825 ;
        RECT 118.305 65.365 120.895 66.135 ;
        RECT 123.135 66.115 123.655 66.655 ;
        RECT 121.525 65.365 121.815 66.090 ;
        RECT 122.445 65.365 123.655 66.115 ;
        RECT 5.520 65.195 123.740 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.985 64.425 10.495 65.195 ;
        RECT 10.665 64.445 11.875 65.195 ;
        RECT 12.045 64.520 12.305 65.025 ;
        RECT 12.485 64.815 12.815 65.195 ;
        RECT 12.995 64.645 13.165 65.025 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 6.985 63.905 8.635 64.425 ;
        RECT 8.805 63.735 10.495 64.255 ;
        RECT 10.665 63.905 11.185 64.445 ;
        RECT 11.355 63.735 11.875 64.275 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 6.985 62.645 10.495 63.735 ;
        RECT 10.665 62.645 11.875 63.735 ;
        RECT 12.045 63.720 12.215 64.520 ;
        RECT 12.500 64.475 13.165 64.645 ;
        RECT 13.515 64.545 13.685 65.025 ;
        RECT 13.865 64.715 14.105 65.195 ;
        RECT 14.355 64.545 14.525 65.025 ;
        RECT 14.695 64.715 15.025 65.195 ;
        RECT 15.195 64.545 15.365 65.025 ;
        RECT 12.500 64.220 12.670 64.475 ;
        RECT 13.515 64.375 14.150 64.545 ;
        RECT 14.355 64.375 15.365 64.545 ;
        RECT 15.535 64.395 15.865 65.195 ;
        RECT 17.110 64.455 17.365 65.025 ;
        RECT 17.535 64.795 17.865 65.195 ;
        RECT 18.290 64.660 18.820 65.025 ;
        RECT 18.290 64.625 18.465 64.660 ;
        RECT 17.535 64.455 18.465 64.625 ;
        RECT 12.385 63.890 12.670 64.220 ;
        RECT 12.905 63.925 13.235 64.295 ;
        RECT 13.980 64.205 14.150 64.375 ;
        RECT 14.865 64.345 15.365 64.375 ;
        RECT 13.430 63.965 13.810 64.205 ;
        RECT 13.980 64.035 14.480 64.205 ;
        RECT 12.500 63.745 12.670 63.890 ;
        RECT 13.980 63.795 14.150 64.035 ;
        RECT 14.870 63.835 15.365 64.345 ;
        RECT 12.045 62.815 12.315 63.720 ;
        RECT 12.500 63.575 13.165 63.745 ;
        RECT 12.485 62.645 12.815 63.405 ;
        RECT 12.995 62.815 13.165 63.575 ;
        RECT 13.435 63.625 14.150 63.795 ;
        RECT 14.355 63.665 15.365 63.835 ;
        RECT 13.435 62.815 13.765 63.625 ;
        RECT 13.935 62.645 14.175 63.445 ;
        RECT 14.355 62.815 14.525 63.665 ;
        RECT 14.695 62.645 15.025 63.445 ;
        RECT 15.195 62.815 15.365 63.665 ;
        RECT 15.535 62.645 15.865 63.795 ;
        RECT 17.110 63.785 17.280 64.455 ;
        RECT 17.535 64.285 17.705 64.455 ;
        RECT 17.450 63.955 17.705 64.285 ;
        RECT 17.930 63.955 18.125 64.285 ;
        RECT 17.110 62.815 17.445 63.785 ;
        RECT 17.615 62.645 17.785 63.785 ;
        RECT 17.955 62.985 18.125 63.955 ;
        RECT 18.295 63.325 18.465 64.455 ;
        RECT 18.635 63.665 18.805 64.465 ;
        RECT 19.010 64.175 19.285 65.025 ;
        RECT 19.005 64.005 19.285 64.175 ;
        RECT 19.010 63.865 19.285 64.005 ;
        RECT 19.455 63.665 19.645 65.025 ;
        RECT 19.825 64.660 20.335 65.195 ;
        RECT 20.555 64.385 20.800 64.990 ;
        RECT 21.250 64.455 21.505 65.025 ;
        RECT 21.675 64.795 22.005 65.195 ;
        RECT 22.430 64.660 22.960 65.025 ;
        RECT 23.150 64.855 23.425 65.025 ;
        RECT 23.145 64.685 23.425 64.855 ;
        RECT 22.430 64.625 22.605 64.660 ;
        RECT 21.675 64.455 22.605 64.625 ;
        RECT 19.845 64.215 21.075 64.385 ;
        RECT 18.635 63.495 19.645 63.665 ;
        RECT 19.815 63.650 20.565 63.840 ;
        RECT 18.295 63.155 19.420 63.325 ;
        RECT 19.815 62.985 19.985 63.650 ;
        RECT 20.735 63.405 21.075 64.215 ;
        RECT 17.955 62.815 19.985 62.985 ;
        RECT 20.155 62.645 20.325 63.405 ;
        RECT 20.560 62.995 21.075 63.405 ;
        RECT 21.250 63.785 21.420 64.455 ;
        RECT 21.675 64.285 21.845 64.455 ;
        RECT 21.590 63.955 21.845 64.285 ;
        RECT 22.070 63.955 22.265 64.285 ;
        RECT 21.250 62.815 21.585 63.785 ;
        RECT 21.755 62.645 21.925 63.785 ;
        RECT 22.095 62.985 22.265 63.955 ;
        RECT 22.435 63.325 22.605 64.455 ;
        RECT 22.775 63.665 22.945 64.465 ;
        RECT 23.150 63.865 23.425 64.685 ;
        RECT 23.595 63.665 23.785 65.025 ;
        RECT 23.965 64.660 24.475 65.195 ;
        RECT 24.695 64.385 24.940 64.990 ;
        RECT 25.850 64.455 26.105 65.025 ;
        RECT 26.275 64.795 26.605 65.195 ;
        RECT 27.030 64.660 27.560 65.025 ;
        RECT 27.750 64.855 28.025 65.025 ;
        RECT 27.745 64.685 28.025 64.855 ;
        RECT 27.030 64.625 27.205 64.660 ;
        RECT 26.275 64.455 27.205 64.625 ;
        RECT 23.985 64.215 25.215 64.385 ;
        RECT 22.775 63.495 23.785 63.665 ;
        RECT 23.955 63.650 24.705 63.840 ;
        RECT 22.435 63.155 23.560 63.325 ;
        RECT 23.955 62.985 24.125 63.650 ;
        RECT 24.875 63.405 25.215 64.215 ;
        RECT 22.095 62.815 24.125 62.985 ;
        RECT 24.295 62.645 24.465 63.405 ;
        RECT 24.700 62.995 25.215 63.405 ;
        RECT 25.850 63.785 26.020 64.455 ;
        RECT 26.275 64.285 26.445 64.455 ;
        RECT 26.190 63.955 26.445 64.285 ;
        RECT 26.670 63.955 26.865 64.285 ;
        RECT 25.850 62.815 26.185 63.785 ;
        RECT 26.355 62.645 26.525 63.785 ;
        RECT 26.695 62.985 26.865 63.955 ;
        RECT 27.035 63.325 27.205 64.455 ;
        RECT 27.375 63.665 27.545 64.465 ;
        RECT 27.750 63.865 28.025 64.685 ;
        RECT 28.195 63.665 28.385 65.025 ;
        RECT 28.565 64.660 29.075 65.195 ;
        RECT 29.295 64.385 29.540 64.990 ;
        RECT 29.985 64.445 31.195 65.195 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 28.585 64.215 29.815 64.385 ;
        RECT 27.375 63.495 28.385 63.665 ;
        RECT 28.555 63.650 29.305 63.840 ;
        RECT 27.035 63.155 28.160 63.325 ;
        RECT 28.555 62.985 28.725 63.650 ;
        RECT 29.475 63.405 29.815 64.215 ;
        RECT 29.985 63.905 30.505 64.445 ;
        RECT 31.865 64.375 32.095 65.195 ;
        RECT 32.265 64.395 32.595 65.025 ;
        RECT 30.675 63.735 31.195 64.275 ;
        RECT 31.845 63.955 32.175 64.205 ;
        RECT 26.695 62.815 28.725 62.985 ;
        RECT 28.895 62.645 29.065 63.405 ;
        RECT 29.300 62.995 29.815 63.405 ;
        RECT 29.985 62.645 31.195 63.735 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 32.345 63.795 32.595 64.395 ;
        RECT 32.765 64.375 32.975 65.195 ;
        RECT 33.205 64.425 36.715 65.195 ;
        RECT 36.890 64.455 37.145 65.025 ;
        RECT 37.315 64.795 37.645 65.195 ;
        RECT 38.070 64.660 38.600 65.025 ;
        RECT 38.070 64.625 38.245 64.660 ;
        RECT 37.315 64.455 38.245 64.625 ;
        RECT 38.790 64.515 39.065 65.025 ;
        RECT 33.205 63.905 34.855 64.425 ;
        RECT 31.865 62.645 32.095 63.785 ;
        RECT 32.265 62.815 32.595 63.795 ;
        RECT 32.765 62.645 32.975 63.785 ;
        RECT 35.025 63.735 36.715 64.255 ;
        RECT 33.205 62.645 36.715 63.735 ;
        RECT 36.890 63.785 37.060 64.455 ;
        RECT 37.315 64.285 37.485 64.455 ;
        RECT 37.230 63.955 37.485 64.285 ;
        RECT 37.710 63.955 37.905 64.285 ;
        RECT 36.890 62.815 37.225 63.785 ;
        RECT 37.395 62.645 37.565 63.785 ;
        RECT 37.735 62.985 37.905 63.955 ;
        RECT 38.075 63.325 38.245 64.455 ;
        RECT 38.415 63.665 38.585 64.465 ;
        RECT 38.785 64.345 39.065 64.515 ;
        RECT 38.790 63.865 39.065 64.345 ;
        RECT 39.235 63.665 39.425 65.025 ;
        RECT 39.605 64.660 40.115 65.195 ;
        RECT 40.335 64.385 40.580 64.990 ;
        RECT 41.025 64.650 46.370 65.195 ;
        RECT 39.625 64.215 40.855 64.385 ;
        RECT 38.415 63.495 39.425 63.665 ;
        RECT 39.595 63.650 40.345 63.840 ;
        RECT 38.075 63.155 39.200 63.325 ;
        RECT 39.595 62.985 39.765 63.650 ;
        RECT 40.515 63.405 40.855 64.215 ;
        RECT 42.610 63.820 42.950 64.650 ;
        RECT 46.545 64.425 50.055 65.195 ;
        RECT 50.225 64.520 50.485 65.025 ;
        RECT 50.665 64.815 50.995 65.195 ;
        RECT 51.175 64.645 51.345 65.025 ;
        RECT 37.735 62.815 39.765 62.985 ;
        RECT 39.935 62.645 40.105 63.405 ;
        RECT 40.340 62.995 40.855 63.405 ;
        RECT 44.430 63.080 44.780 64.330 ;
        RECT 46.545 63.905 48.195 64.425 ;
        RECT 48.365 63.735 50.055 64.255 ;
        RECT 41.025 62.645 46.370 63.080 ;
        RECT 46.545 62.645 50.055 63.735 ;
        RECT 50.225 63.720 50.395 64.520 ;
        RECT 50.680 64.475 51.345 64.645 ;
        RECT 50.680 64.220 50.850 64.475 ;
        RECT 51.610 64.455 51.865 65.025 ;
        RECT 52.035 64.795 52.365 65.195 ;
        RECT 52.790 64.660 53.320 65.025 ;
        RECT 53.510 64.855 53.785 65.025 ;
        RECT 53.505 64.685 53.785 64.855 ;
        RECT 52.790 64.625 52.965 64.660 ;
        RECT 52.035 64.455 52.965 64.625 ;
        RECT 50.565 63.890 50.850 64.220 ;
        RECT 51.085 63.925 51.415 64.295 ;
        RECT 50.680 63.745 50.850 63.890 ;
        RECT 51.610 63.785 51.780 64.455 ;
        RECT 52.035 64.285 52.205 64.455 ;
        RECT 51.950 63.955 52.205 64.285 ;
        RECT 52.430 63.955 52.625 64.285 ;
        RECT 50.225 62.815 50.495 63.720 ;
        RECT 50.680 63.575 51.345 63.745 ;
        RECT 50.665 62.645 50.995 63.405 ;
        RECT 51.175 62.815 51.345 63.575 ;
        RECT 51.610 62.815 51.945 63.785 ;
        RECT 52.115 62.645 52.285 63.785 ;
        RECT 52.455 62.985 52.625 63.955 ;
        RECT 52.795 63.325 52.965 64.455 ;
        RECT 53.135 63.665 53.305 64.465 ;
        RECT 53.510 63.865 53.785 64.685 ;
        RECT 53.955 63.665 54.145 65.025 ;
        RECT 54.325 64.660 54.835 65.195 ;
        RECT 55.055 64.385 55.300 64.990 ;
        RECT 55.745 64.445 56.955 65.195 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 57.585 64.650 62.930 65.195 ;
        RECT 54.345 64.215 55.575 64.385 ;
        RECT 53.135 63.495 54.145 63.665 ;
        RECT 54.315 63.650 55.065 63.840 ;
        RECT 52.795 63.155 53.920 63.325 ;
        RECT 54.315 62.985 54.485 63.650 ;
        RECT 55.235 63.405 55.575 64.215 ;
        RECT 55.745 63.905 56.265 64.445 ;
        RECT 56.435 63.735 56.955 64.275 ;
        RECT 59.170 63.820 59.510 64.650 ;
        RECT 63.105 64.425 65.695 65.195 ;
        RECT 65.955 64.645 66.125 65.025 ;
        RECT 66.340 64.815 66.670 65.195 ;
        RECT 65.955 64.475 66.670 64.645 ;
        RECT 52.455 62.815 54.485 62.985 ;
        RECT 54.655 62.645 54.825 63.405 ;
        RECT 55.060 62.995 55.575 63.405 ;
        RECT 55.745 62.645 56.955 63.735 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 60.990 63.080 61.340 64.330 ;
        RECT 63.105 63.905 64.315 64.425 ;
        RECT 64.485 63.735 65.695 64.255 ;
        RECT 65.865 63.925 66.220 64.295 ;
        RECT 66.500 64.285 66.670 64.475 ;
        RECT 66.840 64.450 67.095 65.025 ;
        RECT 66.500 63.955 66.755 64.285 ;
        RECT 66.500 63.745 66.670 63.955 ;
        RECT 57.585 62.645 62.930 63.080 ;
        RECT 63.105 62.645 65.695 63.735 ;
        RECT 65.955 63.575 66.670 63.745 ;
        RECT 66.925 63.720 67.095 64.450 ;
        RECT 67.270 64.355 67.530 65.195 ;
        RECT 67.795 64.645 67.965 65.025 ;
        RECT 68.180 64.815 68.510 65.195 ;
        RECT 67.795 64.475 68.510 64.645 ;
        RECT 67.705 63.925 68.060 64.295 ;
        RECT 68.340 64.285 68.510 64.475 ;
        RECT 68.680 64.450 68.935 65.025 ;
        RECT 68.340 63.955 68.595 64.285 ;
        RECT 65.955 62.815 66.125 63.575 ;
        RECT 66.340 62.645 66.670 63.405 ;
        RECT 66.840 62.815 67.095 63.720 ;
        RECT 67.270 62.645 67.530 63.795 ;
        RECT 68.340 63.745 68.510 63.955 ;
        RECT 67.795 63.575 68.510 63.745 ;
        RECT 68.765 63.720 68.935 64.450 ;
        RECT 69.110 64.355 69.370 65.195 ;
        RECT 70.470 64.645 70.725 64.935 ;
        RECT 70.895 64.815 71.225 65.195 ;
        RECT 70.470 64.475 71.220 64.645 ;
        RECT 67.795 62.815 67.965 63.575 ;
        RECT 68.180 62.645 68.510 63.405 ;
        RECT 68.680 62.815 68.935 63.720 ;
        RECT 69.110 62.645 69.370 63.795 ;
        RECT 70.470 63.655 70.820 64.305 ;
        RECT 70.990 63.485 71.220 64.475 ;
        RECT 70.470 63.315 71.220 63.485 ;
        RECT 70.470 62.815 70.725 63.315 ;
        RECT 70.895 62.645 71.225 63.145 ;
        RECT 71.395 62.815 71.565 64.935 ;
        RECT 71.925 64.835 72.255 65.195 ;
        RECT 72.425 64.805 72.920 64.975 ;
        RECT 73.125 64.805 73.980 64.975 ;
        RECT 71.795 63.615 72.255 64.665 ;
        RECT 71.735 62.830 72.060 63.615 ;
        RECT 72.425 63.445 72.595 64.805 ;
        RECT 72.765 63.895 73.115 64.515 ;
        RECT 73.285 64.295 73.640 64.515 ;
        RECT 73.285 63.705 73.455 64.295 ;
        RECT 73.810 64.095 73.980 64.805 ;
        RECT 74.855 64.735 75.185 65.195 ;
        RECT 75.395 64.835 75.745 65.005 ;
        RECT 74.185 64.265 74.975 64.515 ;
        RECT 75.395 64.445 75.655 64.835 ;
        RECT 75.965 64.745 76.915 65.025 ;
        RECT 77.085 64.755 77.275 65.195 ;
        RECT 77.445 64.815 78.515 64.985 ;
        RECT 75.145 64.095 75.315 64.275 ;
        RECT 72.425 63.275 72.820 63.445 ;
        RECT 72.990 63.315 73.455 63.705 ;
        RECT 73.625 63.925 75.315 64.095 ;
        RECT 72.650 63.145 72.820 63.275 ;
        RECT 73.625 63.145 73.795 63.925 ;
        RECT 75.485 63.755 75.655 64.445 ;
        RECT 74.155 63.585 75.655 63.755 ;
        RECT 75.845 63.785 76.055 64.575 ;
        RECT 76.225 63.955 76.575 64.575 ;
        RECT 76.745 63.965 76.915 64.745 ;
        RECT 77.445 64.585 77.615 64.815 ;
        RECT 77.085 64.415 77.615 64.585 ;
        RECT 77.085 64.135 77.305 64.415 ;
        RECT 77.785 64.245 78.025 64.645 ;
        RECT 76.745 63.795 77.150 63.965 ;
        RECT 77.485 63.875 78.025 64.245 ;
        RECT 78.195 64.460 78.515 64.815 ;
        RECT 78.760 64.735 79.065 65.195 ;
        RECT 79.235 64.485 79.490 65.015 ;
        RECT 78.195 64.285 78.520 64.460 ;
        RECT 78.195 63.985 79.110 64.285 ;
        RECT 78.370 63.955 79.110 63.985 ;
        RECT 75.845 63.625 76.520 63.785 ;
        RECT 76.980 63.705 77.150 63.795 ;
        RECT 75.845 63.615 76.810 63.625 ;
        RECT 75.485 63.445 75.655 63.585 ;
        RECT 72.230 62.645 72.480 63.105 ;
        RECT 72.650 62.815 72.900 63.145 ;
        RECT 73.115 62.815 73.795 63.145 ;
        RECT 73.965 63.245 75.040 63.415 ;
        RECT 75.485 63.275 76.045 63.445 ;
        RECT 76.350 63.325 76.810 63.615 ;
        RECT 76.980 63.535 78.200 63.705 ;
        RECT 73.965 62.905 74.135 63.245 ;
        RECT 74.370 62.645 74.700 63.075 ;
        RECT 74.870 62.905 75.040 63.245 ;
        RECT 75.335 62.645 75.705 63.105 ;
        RECT 75.875 62.815 76.045 63.275 ;
        RECT 76.980 63.155 77.150 63.535 ;
        RECT 78.370 63.365 78.540 63.955 ;
        RECT 79.280 63.835 79.490 64.485 ;
        RECT 79.725 64.375 79.935 65.195 ;
        RECT 80.105 64.395 80.435 65.025 ;
        RECT 76.280 62.815 77.150 63.155 ;
        RECT 77.740 63.195 78.540 63.365 ;
        RECT 77.320 62.645 77.570 63.105 ;
        RECT 77.740 62.905 77.910 63.195 ;
        RECT 78.090 62.645 78.420 63.025 ;
        RECT 78.760 62.645 79.065 63.785 ;
        RECT 79.235 62.955 79.490 63.835 ;
        RECT 80.105 63.795 80.355 64.395 ;
        RECT 80.605 64.375 80.835 65.195 ;
        RECT 81.045 64.425 82.715 65.195 ;
        RECT 82.885 64.470 83.175 65.195 ;
        RECT 83.345 64.425 86.855 65.195 ;
        RECT 87.025 64.520 87.285 65.025 ;
        RECT 87.465 64.815 87.795 65.195 ;
        RECT 87.975 64.645 88.145 65.025 ;
        RECT 80.525 63.955 80.855 64.205 ;
        RECT 81.045 63.905 81.795 64.425 ;
        RECT 79.725 62.645 79.935 63.785 ;
        RECT 80.105 62.815 80.435 63.795 ;
        RECT 80.605 62.645 80.835 63.785 ;
        RECT 81.965 63.735 82.715 64.255 ;
        RECT 83.345 63.905 84.995 64.425 ;
        RECT 81.045 62.645 82.715 63.735 ;
        RECT 82.885 62.645 83.175 63.810 ;
        RECT 85.165 63.735 86.855 64.255 ;
        RECT 83.345 62.645 86.855 63.735 ;
        RECT 87.025 63.720 87.195 64.520 ;
        RECT 87.480 64.475 88.145 64.645 ;
        RECT 88.405 64.695 88.705 65.025 ;
        RECT 88.875 64.715 89.150 65.195 ;
        RECT 87.480 64.220 87.650 64.475 ;
        RECT 87.365 63.890 87.650 64.220 ;
        RECT 87.885 63.925 88.215 64.295 ;
        RECT 87.480 63.745 87.650 63.890 ;
        RECT 88.405 63.785 88.575 64.695 ;
        RECT 89.330 64.545 89.625 64.935 ;
        RECT 89.795 64.715 90.050 65.195 ;
        RECT 90.225 64.545 90.485 64.935 ;
        RECT 90.655 64.715 90.935 65.195 ;
        RECT 88.745 63.955 89.095 64.525 ;
        RECT 89.330 64.375 90.980 64.545 ;
        RECT 92.360 64.385 92.605 64.990 ;
        RECT 92.825 64.660 93.335 65.195 ;
        RECT 89.265 64.035 90.405 64.205 ;
        RECT 89.265 63.785 89.435 64.035 ;
        RECT 90.575 63.865 90.980 64.375 ;
        RECT 87.025 62.815 87.295 63.720 ;
        RECT 87.480 63.575 88.145 63.745 ;
        RECT 87.465 62.645 87.795 63.405 ;
        RECT 87.975 62.815 88.145 63.575 ;
        RECT 88.405 63.615 89.435 63.785 ;
        RECT 90.225 63.695 90.980 63.865 ;
        RECT 92.085 64.215 93.315 64.385 ;
        RECT 88.405 62.815 88.715 63.615 ;
        RECT 90.225 63.445 90.485 63.695 ;
        RECT 88.885 62.645 89.195 63.445 ;
        RECT 89.365 63.275 90.485 63.445 ;
        RECT 89.365 62.815 89.625 63.275 ;
        RECT 89.795 62.645 90.050 63.105 ;
        RECT 90.225 62.815 90.485 63.275 ;
        RECT 90.655 62.645 90.940 63.515 ;
        RECT 92.085 63.405 92.425 64.215 ;
        RECT 92.595 63.650 93.345 63.840 ;
        RECT 92.085 62.995 92.600 63.405 ;
        RECT 92.835 62.645 93.005 63.405 ;
        RECT 93.175 62.985 93.345 63.650 ;
        RECT 93.515 63.665 93.705 65.025 ;
        RECT 93.875 64.855 94.150 65.025 ;
        RECT 93.875 64.685 94.155 64.855 ;
        RECT 93.875 63.865 94.150 64.685 ;
        RECT 94.340 64.660 94.870 65.025 ;
        RECT 95.295 64.795 95.625 65.195 ;
        RECT 94.695 64.625 94.870 64.660 ;
        RECT 94.355 63.665 94.525 64.465 ;
        RECT 93.515 63.495 94.525 63.665 ;
        RECT 94.695 64.455 95.625 64.625 ;
        RECT 95.795 64.455 96.050 65.025 ;
        RECT 96.315 64.645 96.485 65.025 ;
        RECT 96.665 64.815 96.995 65.195 ;
        RECT 96.315 64.475 96.980 64.645 ;
        RECT 97.175 64.520 97.435 65.025 ;
        RECT 94.695 63.325 94.865 64.455 ;
        RECT 95.455 64.285 95.625 64.455 ;
        RECT 93.740 63.155 94.865 63.325 ;
        RECT 95.035 63.955 95.230 64.285 ;
        RECT 95.455 63.955 95.710 64.285 ;
        RECT 95.035 62.985 95.205 63.955 ;
        RECT 95.880 63.785 96.050 64.455 ;
        RECT 96.245 63.925 96.575 64.295 ;
        RECT 96.810 64.220 96.980 64.475 ;
        RECT 93.175 62.815 95.205 62.985 ;
        RECT 95.375 62.645 95.545 63.785 ;
        RECT 95.715 62.815 96.050 63.785 ;
        RECT 96.810 63.890 97.095 64.220 ;
        RECT 96.810 63.745 96.980 63.890 ;
        RECT 96.315 63.575 96.980 63.745 ;
        RECT 97.265 63.720 97.435 64.520 ;
        RECT 97.605 64.425 100.195 65.195 ;
        RECT 100.370 64.455 100.625 65.025 ;
        RECT 100.795 64.795 101.125 65.195 ;
        RECT 101.550 64.660 102.080 65.025 ;
        RECT 101.550 64.625 101.725 64.660 ;
        RECT 100.795 64.455 101.725 64.625 ;
        RECT 102.270 64.515 102.545 65.025 ;
        RECT 97.605 63.905 98.815 64.425 ;
        RECT 98.985 63.735 100.195 64.255 ;
        RECT 96.315 62.815 96.485 63.575 ;
        RECT 96.665 62.645 96.995 63.405 ;
        RECT 97.165 62.815 97.435 63.720 ;
        RECT 97.605 62.645 100.195 63.735 ;
        RECT 100.370 63.785 100.540 64.455 ;
        RECT 100.795 64.285 100.965 64.455 ;
        RECT 100.710 63.955 100.965 64.285 ;
        RECT 101.190 63.955 101.385 64.285 ;
        RECT 100.370 62.815 100.705 63.785 ;
        RECT 100.875 62.645 101.045 63.785 ;
        RECT 101.215 62.985 101.385 63.955 ;
        RECT 101.555 63.325 101.725 64.455 ;
        RECT 101.895 63.665 102.065 64.465 ;
        RECT 102.265 64.345 102.545 64.515 ;
        RECT 102.270 63.865 102.545 64.345 ;
        RECT 102.715 63.665 102.905 65.025 ;
        RECT 103.085 64.660 103.595 65.195 ;
        RECT 103.815 64.385 104.060 64.990 ;
        RECT 104.505 64.425 108.015 65.195 ;
        RECT 108.645 64.470 108.935 65.195 ;
        RECT 109.105 64.425 111.695 65.195 ;
        RECT 111.870 64.645 112.125 64.935 ;
        RECT 112.295 64.815 112.625 65.195 ;
        RECT 111.870 64.475 112.620 64.645 ;
        RECT 103.105 64.215 104.335 64.385 ;
        RECT 101.895 63.495 102.905 63.665 ;
        RECT 103.075 63.650 103.825 63.840 ;
        RECT 101.555 63.155 102.680 63.325 ;
        RECT 103.075 62.985 103.245 63.650 ;
        RECT 103.995 63.405 104.335 64.215 ;
        RECT 104.505 63.905 106.155 64.425 ;
        RECT 106.325 63.735 108.015 64.255 ;
        RECT 109.105 63.905 110.315 64.425 ;
        RECT 101.215 62.815 103.245 62.985 ;
        RECT 103.415 62.645 103.585 63.405 ;
        RECT 103.820 62.995 104.335 63.405 ;
        RECT 104.505 62.645 108.015 63.735 ;
        RECT 108.645 62.645 108.935 63.810 ;
        RECT 110.485 63.735 111.695 64.255 ;
        RECT 109.105 62.645 111.695 63.735 ;
        RECT 111.870 63.655 112.220 64.305 ;
        RECT 112.390 63.485 112.620 64.475 ;
        RECT 111.870 63.315 112.620 63.485 ;
        RECT 111.870 62.815 112.125 63.315 ;
        RECT 112.295 62.645 112.625 63.145 ;
        RECT 112.795 62.815 112.965 64.935 ;
        RECT 113.325 64.835 113.655 65.195 ;
        RECT 113.825 64.805 114.320 64.975 ;
        RECT 114.525 64.805 115.380 64.975 ;
        RECT 113.195 63.615 113.655 64.665 ;
        RECT 113.135 62.830 113.460 63.615 ;
        RECT 113.825 63.445 113.995 64.805 ;
        RECT 114.165 63.895 114.515 64.515 ;
        RECT 114.685 64.295 115.040 64.515 ;
        RECT 114.685 63.705 114.855 64.295 ;
        RECT 115.210 64.095 115.380 64.805 ;
        RECT 116.255 64.735 116.585 65.195 ;
        RECT 116.795 64.835 117.145 65.005 ;
        RECT 115.585 64.265 116.375 64.515 ;
        RECT 116.795 64.445 117.055 64.835 ;
        RECT 117.365 64.745 118.315 65.025 ;
        RECT 118.485 64.755 118.675 65.195 ;
        RECT 118.845 64.815 119.915 64.985 ;
        RECT 116.545 64.095 116.715 64.275 ;
        RECT 113.825 63.275 114.220 63.445 ;
        RECT 114.390 63.315 114.855 63.705 ;
        RECT 115.025 63.925 116.715 64.095 ;
        RECT 114.050 63.145 114.220 63.275 ;
        RECT 115.025 63.145 115.195 63.925 ;
        RECT 116.885 63.755 117.055 64.445 ;
        RECT 115.555 63.585 117.055 63.755 ;
        RECT 117.245 63.785 117.455 64.575 ;
        RECT 117.625 63.955 117.975 64.575 ;
        RECT 118.145 63.965 118.315 64.745 ;
        RECT 118.845 64.585 119.015 64.815 ;
        RECT 118.485 64.415 119.015 64.585 ;
        RECT 118.485 64.135 118.705 64.415 ;
        RECT 119.185 64.245 119.425 64.645 ;
        RECT 118.145 63.795 118.550 63.965 ;
        RECT 118.885 63.875 119.425 64.245 ;
        RECT 119.595 64.460 119.915 64.815 ;
        RECT 120.160 64.735 120.465 65.195 ;
        RECT 120.635 64.485 120.890 65.015 ;
        RECT 119.595 64.285 119.920 64.460 ;
        RECT 119.595 63.985 120.510 64.285 ;
        RECT 119.770 63.955 120.510 63.985 ;
        RECT 117.245 63.625 117.920 63.785 ;
        RECT 118.380 63.705 118.550 63.795 ;
        RECT 117.245 63.615 118.210 63.625 ;
        RECT 116.885 63.445 117.055 63.585 ;
        RECT 113.630 62.645 113.880 63.105 ;
        RECT 114.050 62.815 114.300 63.145 ;
        RECT 114.515 62.815 115.195 63.145 ;
        RECT 115.365 63.245 116.440 63.415 ;
        RECT 116.885 63.275 117.445 63.445 ;
        RECT 117.750 63.325 118.210 63.615 ;
        RECT 118.380 63.535 119.600 63.705 ;
        RECT 115.365 62.905 115.535 63.245 ;
        RECT 115.770 62.645 116.100 63.075 ;
        RECT 116.270 62.905 116.440 63.245 ;
        RECT 116.735 62.645 117.105 63.105 ;
        RECT 117.275 62.815 117.445 63.275 ;
        RECT 118.380 63.155 118.550 63.535 ;
        RECT 119.770 63.365 119.940 63.955 ;
        RECT 120.680 63.835 120.890 64.485 ;
        RECT 121.065 64.445 122.275 65.195 ;
        RECT 122.445 64.445 123.655 65.195 ;
        RECT 121.065 63.905 121.585 64.445 ;
        RECT 117.680 62.815 118.550 63.155 ;
        RECT 119.140 63.195 119.940 63.365 ;
        RECT 118.720 62.645 118.970 63.105 ;
        RECT 119.140 62.905 119.310 63.195 ;
        RECT 119.490 62.645 119.820 63.025 ;
        RECT 120.160 62.645 120.465 63.785 ;
        RECT 120.635 62.955 120.890 63.835 ;
        RECT 121.755 63.735 122.275 64.275 ;
        RECT 121.065 62.645 122.275 63.735 ;
        RECT 122.445 63.735 122.965 64.275 ;
        RECT 123.135 63.905 123.655 64.445 ;
        RECT 122.445 62.645 123.655 63.735 ;
        RECT 5.520 62.475 123.740 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 7.910 61.805 8.165 62.305 ;
        RECT 8.335 61.975 8.665 62.475 ;
        RECT 7.910 61.635 8.660 61.805 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 7.910 60.815 8.260 61.465 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 8.430 60.645 8.660 61.635 ;
        RECT 7.910 60.475 8.660 60.645 ;
        RECT 7.910 60.185 8.165 60.475 ;
        RECT 8.335 59.925 8.665 60.305 ;
        RECT 8.835 60.185 9.005 62.305 ;
        RECT 9.175 61.505 9.500 62.290 ;
        RECT 9.670 62.015 9.920 62.475 ;
        RECT 10.090 61.975 10.340 62.305 ;
        RECT 10.555 61.975 11.235 62.305 ;
        RECT 10.090 61.845 10.260 61.975 ;
        RECT 9.865 61.675 10.260 61.845 ;
        RECT 9.235 60.455 9.695 61.505 ;
        RECT 9.865 60.315 10.035 61.675 ;
        RECT 10.430 61.415 10.895 61.805 ;
        RECT 10.205 60.605 10.555 61.225 ;
        RECT 10.725 60.825 10.895 61.415 ;
        RECT 11.065 61.195 11.235 61.975 ;
        RECT 11.405 61.875 11.575 62.215 ;
        RECT 11.810 62.045 12.140 62.475 ;
        RECT 12.310 61.875 12.480 62.215 ;
        RECT 12.775 62.015 13.145 62.475 ;
        RECT 11.405 61.705 12.480 61.875 ;
        RECT 13.315 61.845 13.485 62.305 ;
        RECT 13.720 61.965 14.590 62.305 ;
        RECT 14.760 62.015 15.010 62.475 ;
        RECT 12.925 61.675 13.485 61.845 ;
        RECT 12.925 61.535 13.095 61.675 ;
        RECT 11.595 61.365 13.095 61.535 ;
        RECT 13.790 61.505 14.250 61.795 ;
        RECT 11.065 61.025 12.755 61.195 ;
        RECT 10.725 60.605 11.080 60.825 ;
        RECT 11.250 60.315 11.420 61.025 ;
        RECT 11.625 60.605 12.415 60.855 ;
        RECT 12.585 60.845 12.755 61.025 ;
        RECT 12.925 60.675 13.095 61.365 ;
        RECT 9.365 59.925 9.695 60.285 ;
        RECT 9.865 60.145 10.360 60.315 ;
        RECT 10.565 60.145 11.420 60.315 ;
        RECT 12.295 59.925 12.625 60.385 ;
        RECT 12.835 60.285 13.095 60.675 ;
        RECT 13.285 61.495 14.250 61.505 ;
        RECT 14.420 61.585 14.590 61.965 ;
        RECT 15.180 61.925 15.350 62.215 ;
        RECT 15.530 62.095 15.860 62.475 ;
        RECT 15.180 61.755 15.980 61.925 ;
        RECT 13.285 61.335 13.960 61.495 ;
        RECT 14.420 61.415 15.640 61.585 ;
        RECT 13.285 60.545 13.495 61.335 ;
        RECT 14.420 61.325 14.590 61.415 ;
        RECT 13.665 60.545 14.015 61.165 ;
        RECT 14.185 61.155 14.590 61.325 ;
        RECT 14.185 60.375 14.355 61.155 ;
        RECT 14.525 60.705 14.745 60.985 ;
        RECT 14.925 60.875 15.465 61.245 ;
        RECT 15.810 61.165 15.980 61.755 ;
        RECT 16.200 61.335 16.505 62.475 ;
        RECT 16.675 61.285 16.930 62.165 ;
        RECT 15.810 61.135 16.550 61.165 ;
        RECT 14.525 60.535 15.055 60.705 ;
        RECT 12.835 60.115 13.185 60.285 ;
        RECT 13.405 60.095 14.355 60.375 ;
        RECT 14.525 59.925 14.715 60.365 ;
        RECT 14.885 60.305 15.055 60.535 ;
        RECT 15.225 60.475 15.465 60.875 ;
        RECT 15.635 60.835 16.550 61.135 ;
        RECT 15.635 60.660 15.960 60.835 ;
        RECT 15.635 60.305 15.955 60.660 ;
        RECT 16.720 60.635 16.930 61.285 ;
        RECT 14.885 60.135 15.955 60.305 ;
        RECT 16.200 59.925 16.505 60.385 ;
        RECT 16.675 60.105 16.930 60.635 ;
        RECT 17.105 61.400 17.375 62.305 ;
        RECT 17.545 61.715 17.875 62.475 ;
        RECT 18.055 61.545 18.225 62.305 ;
        RECT 17.105 60.600 17.275 61.400 ;
        RECT 17.560 61.375 18.225 61.545 ;
        RECT 17.560 61.230 17.730 61.375 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 19.870 61.335 20.205 62.305 ;
        RECT 20.375 61.335 20.545 62.475 ;
        RECT 20.715 62.135 22.745 62.305 ;
        RECT 17.445 60.900 17.730 61.230 ;
        RECT 17.560 60.645 17.730 60.900 ;
        RECT 17.965 60.825 18.295 61.195 ;
        RECT 19.870 60.665 20.040 61.335 ;
        RECT 20.715 61.165 20.885 62.135 ;
        RECT 20.210 60.835 20.465 61.165 ;
        RECT 20.690 60.835 20.885 61.165 ;
        RECT 21.055 61.795 22.180 61.965 ;
        RECT 20.295 60.665 20.465 60.835 ;
        RECT 21.055 60.665 21.225 61.795 ;
        RECT 17.105 60.095 17.365 60.600 ;
        RECT 17.560 60.475 18.225 60.645 ;
        RECT 17.545 59.925 17.875 60.305 ;
        RECT 18.055 60.095 18.225 60.475 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 19.870 60.095 20.125 60.665 ;
        RECT 20.295 60.495 21.225 60.665 ;
        RECT 21.395 61.455 22.405 61.625 ;
        RECT 21.395 60.655 21.565 61.455 ;
        RECT 21.770 60.775 22.045 61.255 ;
        RECT 21.765 60.605 22.045 60.775 ;
        RECT 21.050 60.460 21.225 60.495 ;
        RECT 20.295 59.925 20.625 60.325 ;
        RECT 21.050 60.095 21.580 60.460 ;
        RECT 21.770 60.095 22.045 60.605 ;
        RECT 22.215 60.095 22.405 61.455 ;
        RECT 22.575 61.470 22.745 62.135 ;
        RECT 22.915 61.715 23.085 62.475 ;
        RECT 23.320 61.715 23.835 62.125 ;
        RECT 22.575 61.280 23.325 61.470 ;
        RECT 23.495 60.905 23.835 61.715 ;
        RECT 24.005 61.385 26.595 62.475 ;
        RECT 27.315 61.805 27.485 62.305 ;
        RECT 27.655 61.975 27.985 62.475 ;
        RECT 27.315 61.635 27.980 61.805 ;
        RECT 22.605 60.735 23.835 60.905 ;
        RECT 22.585 59.925 23.095 60.460 ;
        RECT 23.315 60.130 23.560 60.735 ;
        RECT 24.005 60.695 25.215 61.215 ;
        RECT 25.385 60.865 26.595 61.385 ;
        RECT 27.230 60.815 27.580 61.465 ;
        RECT 24.005 59.925 26.595 60.695 ;
        RECT 27.750 60.645 27.980 61.635 ;
        RECT 27.315 60.475 27.980 60.645 ;
        RECT 27.315 60.185 27.485 60.475 ;
        RECT 27.655 59.925 27.985 60.305 ;
        RECT 28.155 60.185 28.380 62.305 ;
        RECT 28.595 61.975 28.925 62.475 ;
        RECT 29.095 61.805 29.265 62.305 ;
        RECT 29.500 62.090 30.330 62.260 ;
        RECT 30.570 62.095 30.950 62.475 ;
        RECT 28.570 61.635 29.265 61.805 ;
        RECT 28.570 60.665 28.740 61.635 ;
        RECT 28.910 60.845 29.320 61.465 ;
        RECT 29.490 61.415 29.990 61.795 ;
        RECT 28.570 60.475 29.265 60.665 ;
        RECT 29.490 60.545 29.710 61.415 ;
        RECT 30.160 61.245 30.330 62.090 ;
        RECT 31.130 61.925 31.300 62.215 ;
        RECT 31.470 62.095 31.800 62.475 ;
        RECT 32.270 62.005 32.900 62.255 ;
        RECT 33.080 62.095 33.500 62.475 ;
        RECT 32.730 61.925 32.900 62.005 ;
        RECT 33.700 61.925 33.940 62.215 ;
        RECT 30.500 61.675 31.870 61.925 ;
        RECT 30.500 61.415 30.750 61.675 ;
        RECT 31.260 61.245 31.510 61.405 ;
        RECT 30.160 61.075 31.510 61.245 ;
        RECT 30.160 61.035 30.580 61.075 ;
        RECT 29.890 60.485 30.240 60.855 ;
        RECT 28.595 59.925 28.925 60.305 ;
        RECT 29.095 60.145 29.265 60.475 ;
        RECT 30.410 60.305 30.580 61.035 ;
        RECT 31.680 60.905 31.870 61.675 ;
        RECT 30.750 60.575 31.160 60.905 ;
        RECT 31.450 60.565 31.870 60.905 ;
        RECT 32.040 61.495 32.560 61.805 ;
        RECT 32.730 61.755 33.940 61.925 ;
        RECT 34.170 61.785 34.500 62.475 ;
        RECT 32.040 60.735 32.210 61.495 ;
        RECT 32.380 60.905 32.560 61.315 ;
        RECT 32.730 61.245 32.900 61.755 ;
        RECT 34.670 61.605 34.840 62.215 ;
        RECT 35.110 61.755 35.440 62.265 ;
        RECT 34.670 61.585 34.990 61.605 ;
        RECT 33.070 61.415 34.990 61.585 ;
        RECT 32.730 61.075 34.630 61.245 ;
        RECT 32.960 60.735 33.290 60.855 ;
        RECT 32.040 60.565 33.290 60.735 ;
        RECT 29.565 60.105 30.580 60.305 ;
        RECT 30.750 59.925 31.160 60.365 ;
        RECT 31.450 60.135 31.700 60.565 ;
        RECT 31.900 59.925 32.220 60.385 ;
        RECT 33.460 60.315 33.630 61.075 ;
        RECT 34.300 61.015 34.630 61.075 ;
        RECT 33.820 60.845 34.150 60.905 ;
        RECT 33.820 60.575 34.480 60.845 ;
        RECT 34.800 60.520 34.990 61.415 ;
        RECT 32.780 60.145 33.630 60.315 ;
        RECT 33.830 59.925 34.490 60.405 ;
        RECT 34.670 60.190 34.990 60.520 ;
        RECT 35.190 61.165 35.440 61.755 ;
        RECT 35.620 61.675 35.905 62.475 ;
        RECT 36.085 62.135 36.340 62.165 ;
        RECT 36.085 61.965 36.425 62.135 ;
        RECT 36.885 62.040 42.230 62.475 ;
        RECT 36.085 61.495 36.340 61.965 ;
        RECT 35.190 60.835 35.990 61.165 ;
        RECT 35.190 60.185 35.440 60.835 ;
        RECT 36.160 60.635 36.340 61.495 ;
        RECT 35.620 59.925 35.905 60.385 ;
        RECT 36.085 60.105 36.340 60.635 ;
        RECT 38.470 60.470 38.810 61.300 ;
        RECT 40.290 60.790 40.640 62.040 ;
        RECT 42.405 61.385 44.075 62.475 ;
        RECT 42.405 60.695 43.155 61.215 ;
        RECT 43.325 60.865 44.075 61.385 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 44.705 61.385 45.915 62.475 ;
        RECT 36.885 59.925 42.230 60.470 ;
        RECT 42.405 59.925 44.075 60.695 ;
        RECT 44.705 60.675 45.225 61.215 ;
        RECT 45.395 60.845 45.915 61.385 ;
        RECT 46.125 61.335 46.355 62.475 ;
        RECT 46.525 61.325 46.855 62.305 ;
        RECT 47.025 61.335 47.235 62.475 ;
        RECT 47.505 61.335 47.735 62.475 ;
        RECT 47.905 61.325 48.235 62.305 ;
        RECT 48.405 61.335 48.615 62.475 ;
        RECT 48.935 61.805 49.105 62.305 ;
        RECT 49.275 61.975 49.605 62.475 ;
        RECT 48.935 61.635 49.600 61.805 ;
        RECT 46.105 60.915 46.435 61.165 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 44.705 59.925 45.915 60.675 ;
        RECT 46.125 59.925 46.355 60.745 ;
        RECT 46.605 60.725 46.855 61.325 ;
        RECT 47.485 60.915 47.815 61.165 ;
        RECT 46.525 60.095 46.855 60.725 ;
        RECT 47.025 59.925 47.235 60.745 ;
        RECT 47.505 59.925 47.735 60.745 ;
        RECT 47.985 60.725 48.235 61.325 ;
        RECT 48.850 60.815 49.200 61.465 ;
        RECT 47.905 60.095 48.235 60.725 ;
        RECT 48.405 59.925 48.615 60.745 ;
        RECT 49.370 60.645 49.600 61.635 ;
        RECT 48.935 60.475 49.600 60.645 ;
        RECT 48.935 60.185 49.105 60.475 ;
        RECT 49.275 59.925 49.605 60.305 ;
        RECT 49.775 60.185 50.000 62.305 ;
        RECT 50.215 61.975 50.545 62.475 ;
        RECT 50.715 61.805 50.885 62.305 ;
        RECT 51.120 62.090 51.950 62.260 ;
        RECT 52.190 62.095 52.570 62.475 ;
        RECT 50.190 61.635 50.885 61.805 ;
        RECT 50.190 60.665 50.360 61.635 ;
        RECT 50.530 60.845 50.940 61.465 ;
        RECT 51.110 61.415 51.610 61.795 ;
        RECT 50.190 60.475 50.885 60.665 ;
        RECT 51.110 60.545 51.330 61.415 ;
        RECT 51.780 61.245 51.950 62.090 ;
        RECT 52.750 61.925 52.920 62.215 ;
        RECT 53.090 62.095 53.420 62.475 ;
        RECT 53.890 62.005 54.520 62.255 ;
        RECT 54.700 62.095 55.120 62.475 ;
        RECT 54.350 61.925 54.520 62.005 ;
        RECT 55.320 61.925 55.560 62.215 ;
        RECT 52.120 61.675 53.490 61.925 ;
        RECT 52.120 61.415 52.370 61.675 ;
        RECT 52.880 61.245 53.130 61.405 ;
        RECT 51.780 61.075 53.130 61.245 ;
        RECT 51.780 61.035 52.200 61.075 ;
        RECT 51.510 60.485 51.860 60.855 ;
        RECT 50.215 59.925 50.545 60.305 ;
        RECT 50.715 60.145 50.885 60.475 ;
        RECT 52.030 60.305 52.200 61.035 ;
        RECT 53.300 60.905 53.490 61.675 ;
        RECT 52.370 60.575 52.780 60.905 ;
        RECT 53.070 60.565 53.490 60.905 ;
        RECT 53.660 61.495 54.180 61.805 ;
        RECT 54.350 61.755 55.560 61.925 ;
        RECT 55.790 61.785 56.120 62.475 ;
        RECT 53.660 60.735 53.830 61.495 ;
        RECT 54.000 60.905 54.180 61.315 ;
        RECT 54.350 61.245 54.520 61.755 ;
        RECT 56.290 61.605 56.460 62.215 ;
        RECT 56.730 61.755 57.060 62.265 ;
        RECT 56.290 61.585 56.610 61.605 ;
        RECT 54.690 61.415 56.610 61.585 ;
        RECT 54.350 61.075 56.250 61.245 ;
        RECT 54.580 60.735 54.910 60.855 ;
        RECT 53.660 60.565 54.910 60.735 ;
        RECT 51.185 60.105 52.200 60.305 ;
        RECT 52.370 59.925 52.780 60.365 ;
        RECT 53.070 60.135 53.320 60.565 ;
        RECT 53.520 59.925 53.840 60.385 ;
        RECT 55.080 60.315 55.250 61.075 ;
        RECT 55.920 61.015 56.250 61.075 ;
        RECT 55.440 60.845 55.770 60.905 ;
        RECT 55.440 60.575 56.100 60.845 ;
        RECT 56.420 60.520 56.610 61.415 ;
        RECT 54.400 60.145 55.250 60.315 ;
        RECT 55.450 59.925 56.110 60.405 ;
        RECT 56.290 60.190 56.610 60.520 ;
        RECT 56.810 61.165 57.060 61.755 ;
        RECT 57.240 61.675 57.525 62.475 ;
        RECT 57.705 61.495 57.960 62.165 ;
        RECT 59.480 61.605 59.765 62.475 ;
        RECT 59.935 61.845 60.195 62.305 ;
        RECT 60.370 62.015 60.625 62.475 ;
        RECT 60.795 61.845 61.055 62.305 ;
        RECT 59.935 61.675 61.055 61.845 ;
        RECT 61.225 61.675 61.535 62.475 ;
        RECT 56.810 60.835 57.610 61.165 ;
        RECT 56.810 60.185 57.060 60.835 ;
        RECT 57.780 60.635 57.960 61.495 ;
        RECT 59.935 61.425 60.195 61.675 ;
        RECT 61.705 61.505 62.015 62.305 ;
        RECT 57.705 60.435 57.960 60.635 ;
        RECT 59.440 61.255 60.195 61.425 ;
        RECT 60.985 61.335 62.015 61.505 ;
        RECT 59.440 60.745 59.845 61.255 ;
        RECT 60.985 61.085 61.155 61.335 ;
        RECT 60.015 60.915 61.155 61.085 ;
        RECT 59.440 60.575 61.090 60.745 ;
        RECT 61.325 60.595 61.675 61.165 ;
        RECT 57.240 59.925 57.525 60.385 ;
        RECT 57.705 60.265 58.045 60.435 ;
        RECT 57.705 60.105 57.960 60.265 ;
        RECT 59.485 59.925 59.765 60.405 ;
        RECT 59.935 60.185 60.195 60.575 ;
        RECT 60.370 59.925 60.625 60.405 ;
        RECT 60.795 60.185 61.090 60.575 ;
        RECT 61.845 60.425 62.015 61.335 ;
        RECT 61.270 59.925 61.545 60.405 ;
        RECT 61.715 60.095 62.015 60.425 ;
        RECT 62.645 61.885 63.345 62.305 ;
        RECT 63.545 62.115 63.875 62.475 ;
        RECT 64.045 61.885 64.375 62.285 ;
        RECT 62.645 61.655 64.375 61.885 ;
        RECT 62.645 60.685 62.850 61.655 ;
        RECT 63.020 60.915 63.350 61.455 ;
        RECT 63.525 61.165 63.850 61.455 ;
        RECT 64.045 61.435 64.375 61.655 ;
        RECT 64.545 61.165 64.715 62.090 ;
        RECT 64.895 61.415 65.225 62.475 ;
        RECT 65.495 61.545 65.665 62.305 ;
        RECT 65.880 61.715 66.210 62.475 ;
        RECT 65.495 61.375 66.210 61.545 ;
        RECT 66.380 61.400 66.635 62.305 ;
        RECT 63.525 60.835 64.020 61.165 ;
        RECT 64.340 60.835 64.715 61.165 ;
        RECT 64.925 60.835 65.235 61.165 ;
        RECT 65.405 60.825 65.760 61.195 ;
        RECT 66.040 61.165 66.210 61.375 ;
        RECT 66.040 60.835 66.295 61.165 ;
        RECT 62.645 60.095 63.355 60.685 ;
        RECT 63.865 60.455 65.225 60.665 ;
        RECT 66.040 60.645 66.210 60.835 ;
        RECT 66.465 60.670 66.635 61.400 ;
        RECT 66.810 61.325 67.070 62.475 ;
        RECT 67.245 61.385 69.835 62.475 ;
        RECT 63.865 60.095 64.195 60.455 ;
        RECT 64.395 59.925 64.725 60.285 ;
        RECT 64.895 60.095 65.225 60.455 ;
        RECT 65.495 60.475 66.210 60.645 ;
        RECT 65.495 60.095 65.665 60.475 ;
        RECT 65.880 59.925 66.210 60.305 ;
        RECT 66.380 60.095 66.635 60.670 ;
        RECT 66.810 59.925 67.070 60.765 ;
        RECT 67.245 60.695 68.455 61.215 ;
        RECT 68.625 60.865 69.835 61.385 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.475 61.495 70.805 62.305 ;
        RECT 70.975 61.675 71.215 62.475 ;
        RECT 70.475 61.325 71.190 61.495 ;
        RECT 70.470 60.915 70.850 61.155 ;
        RECT 71.020 61.085 71.190 61.325 ;
        RECT 71.395 61.455 71.565 62.305 ;
        RECT 71.735 61.675 72.065 62.475 ;
        RECT 72.235 61.455 72.405 62.305 ;
        RECT 71.395 61.285 72.405 61.455 ;
        RECT 72.575 61.325 72.905 62.475 ;
        RECT 73.225 62.040 78.570 62.475 ;
        RECT 78.745 62.040 84.090 62.475 ;
        RECT 71.020 60.915 71.520 61.085 ;
        RECT 71.020 60.745 71.190 60.915 ;
        RECT 71.910 60.775 72.405 61.285 ;
        RECT 71.905 60.745 72.405 60.775 ;
        RECT 67.245 59.925 69.835 60.695 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 70.555 60.575 71.190 60.745 ;
        RECT 71.395 60.575 72.405 60.745 ;
        RECT 70.555 60.095 70.725 60.575 ;
        RECT 70.905 59.925 71.145 60.405 ;
        RECT 71.395 60.095 71.565 60.575 ;
        RECT 71.735 59.925 72.065 60.405 ;
        RECT 72.235 60.095 72.405 60.575 ;
        RECT 72.575 59.925 72.905 60.725 ;
        RECT 74.810 60.470 75.150 61.300 ;
        RECT 76.630 60.790 76.980 62.040 ;
        RECT 80.330 60.470 80.670 61.300 ;
        RECT 82.150 60.790 82.500 62.040 ;
        RECT 85.190 61.805 85.445 62.305 ;
        RECT 85.615 61.975 85.945 62.475 ;
        RECT 85.190 61.635 85.940 61.805 ;
        RECT 85.190 60.815 85.540 61.465 ;
        RECT 85.710 60.645 85.940 61.635 ;
        RECT 85.190 60.475 85.940 60.645 ;
        RECT 73.225 59.925 78.570 60.470 ;
        RECT 78.745 59.925 84.090 60.470 ;
        RECT 85.190 60.185 85.445 60.475 ;
        RECT 85.615 59.925 85.945 60.305 ;
        RECT 86.115 60.185 86.285 62.305 ;
        RECT 86.455 61.505 86.780 62.290 ;
        RECT 86.950 62.015 87.200 62.475 ;
        RECT 87.370 61.975 87.620 62.305 ;
        RECT 87.835 61.975 88.515 62.305 ;
        RECT 87.370 61.845 87.540 61.975 ;
        RECT 87.145 61.675 87.540 61.845 ;
        RECT 86.515 60.455 86.975 61.505 ;
        RECT 87.145 60.315 87.315 61.675 ;
        RECT 87.710 61.415 88.175 61.805 ;
        RECT 87.485 60.605 87.835 61.225 ;
        RECT 88.005 60.825 88.175 61.415 ;
        RECT 88.345 61.195 88.515 61.975 ;
        RECT 88.685 61.875 88.855 62.215 ;
        RECT 89.090 62.045 89.420 62.475 ;
        RECT 89.590 61.875 89.760 62.215 ;
        RECT 90.055 62.015 90.425 62.475 ;
        RECT 88.685 61.705 89.760 61.875 ;
        RECT 90.595 61.845 90.765 62.305 ;
        RECT 91.000 61.965 91.870 62.305 ;
        RECT 92.040 62.015 92.290 62.475 ;
        RECT 90.205 61.675 90.765 61.845 ;
        RECT 90.205 61.535 90.375 61.675 ;
        RECT 88.875 61.365 90.375 61.535 ;
        RECT 91.070 61.505 91.530 61.795 ;
        RECT 88.345 61.025 90.035 61.195 ;
        RECT 88.005 60.605 88.360 60.825 ;
        RECT 88.530 60.315 88.700 61.025 ;
        RECT 88.905 60.605 89.695 60.855 ;
        RECT 89.865 60.845 90.035 61.025 ;
        RECT 90.205 60.675 90.375 61.365 ;
        RECT 86.645 59.925 86.975 60.285 ;
        RECT 87.145 60.145 87.640 60.315 ;
        RECT 87.845 60.145 88.700 60.315 ;
        RECT 89.575 59.925 89.905 60.385 ;
        RECT 90.115 60.285 90.375 60.675 ;
        RECT 90.565 61.495 91.530 61.505 ;
        RECT 91.700 61.585 91.870 61.965 ;
        RECT 92.460 61.925 92.630 62.215 ;
        RECT 92.810 62.095 93.140 62.475 ;
        RECT 92.460 61.755 93.260 61.925 ;
        RECT 90.565 61.335 91.240 61.495 ;
        RECT 91.700 61.415 92.920 61.585 ;
        RECT 90.565 60.545 90.775 61.335 ;
        RECT 91.700 61.325 91.870 61.415 ;
        RECT 90.945 60.545 91.295 61.165 ;
        RECT 91.465 61.155 91.870 61.325 ;
        RECT 91.465 60.375 91.635 61.155 ;
        RECT 91.805 60.705 92.025 60.985 ;
        RECT 92.205 60.875 92.745 61.245 ;
        RECT 93.090 61.165 93.260 61.755 ;
        RECT 93.480 61.335 93.785 62.475 ;
        RECT 93.955 61.285 94.210 62.165 ;
        RECT 94.385 61.385 95.595 62.475 ;
        RECT 93.090 61.135 93.830 61.165 ;
        RECT 91.805 60.535 92.335 60.705 ;
        RECT 90.115 60.115 90.465 60.285 ;
        RECT 90.685 60.095 91.635 60.375 ;
        RECT 91.805 59.925 91.995 60.365 ;
        RECT 92.165 60.305 92.335 60.535 ;
        RECT 92.505 60.475 92.745 60.875 ;
        RECT 92.915 60.835 93.830 61.135 ;
        RECT 92.915 60.660 93.240 60.835 ;
        RECT 92.915 60.305 93.235 60.660 ;
        RECT 94.000 60.635 94.210 61.285 ;
        RECT 92.165 60.135 93.235 60.305 ;
        RECT 93.480 59.925 93.785 60.385 ;
        RECT 93.955 60.105 94.210 60.635 ;
        RECT 94.385 60.675 94.905 61.215 ;
        RECT 95.075 60.845 95.595 61.385 ;
        RECT 95.765 61.310 96.055 62.475 ;
        RECT 96.230 61.805 96.485 62.305 ;
        RECT 96.655 61.975 96.985 62.475 ;
        RECT 96.230 61.635 96.980 61.805 ;
        RECT 96.230 60.815 96.580 61.465 ;
        RECT 94.385 59.925 95.595 60.675 ;
        RECT 95.765 59.925 96.055 60.650 ;
        RECT 96.750 60.645 96.980 61.635 ;
        RECT 96.230 60.475 96.980 60.645 ;
        RECT 96.230 60.185 96.485 60.475 ;
        RECT 96.655 59.925 96.985 60.305 ;
        RECT 97.155 60.185 97.325 62.305 ;
        RECT 97.495 61.505 97.820 62.290 ;
        RECT 97.990 62.015 98.240 62.475 ;
        RECT 98.410 61.975 98.660 62.305 ;
        RECT 98.875 61.975 99.555 62.305 ;
        RECT 98.410 61.845 98.580 61.975 ;
        RECT 98.185 61.675 98.580 61.845 ;
        RECT 97.555 60.455 98.015 61.505 ;
        RECT 98.185 60.315 98.355 61.675 ;
        RECT 98.750 61.415 99.215 61.805 ;
        RECT 98.525 60.605 98.875 61.225 ;
        RECT 99.045 60.825 99.215 61.415 ;
        RECT 99.385 61.195 99.555 61.975 ;
        RECT 99.725 61.875 99.895 62.215 ;
        RECT 100.130 62.045 100.460 62.475 ;
        RECT 100.630 61.875 100.800 62.215 ;
        RECT 101.095 62.015 101.465 62.475 ;
        RECT 99.725 61.705 100.800 61.875 ;
        RECT 101.635 61.845 101.805 62.305 ;
        RECT 102.040 61.965 102.910 62.305 ;
        RECT 103.080 62.015 103.330 62.475 ;
        RECT 101.245 61.675 101.805 61.845 ;
        RECT 101.245 61.535 101.415 61.675 ;
        RECT 99.915 61.365 101.415 61.535 ;
        RECT 102.110 61.505 102.570 61.795 ;
        RECT 99.385 61.025 101.075 61.195 ;
        RECT 99.045 60.605 99.400 60.825 ;
        RECT 99.570 60.315 99.740 61.025 ;
        RECT 99.945 60.605 100.735 60.855 ;
        RECT 100.905 60.845 101.075 61.025 ;
        RECT 101.245 60.675 101.415 61.365 ;
        RECT 97.685 59.925 98.015 60.285 ;
        RECT 98.185 60.145 98.680 60.315 ;
        RECT 98.885 60.145 99.740 60.315 ;
        RECT 100.615 59.925 100.945 60.385 ;
        RECT 101.155 60.285 101.415 60.675 ;
        RECT 101.605 61.495 102.570 61.505 ;
        RECT 102.740 61.585 102.910 61.965 ;
        RECT 103.500 61.925 103.670 62.215 ;
        RECT 103.850 62.095 104.180 62.475 ;
        RECT 103.500 61.755 104.300 61.925 ;
        RECT 101.605 61.335 102.280 61.495 ;
        RECT 102.740 61.415 103.960 61.585 ;
        RECT 101.605 60.545 101.815 61.335 ;
        RECT 102.740 61.325 102.910 61.415 ;
        RECT 101.985 60.545 102.335 61.165 ;
        RECT 102.505 61.155 102.910 61.325 ;
        RECT 102.505 60.375 102.675 61.155 ;
        RECT 102.845 60.705 103.065 60.985 ;
        RECT 103.245 60.875 103.785 61.245 ;
        RECT 104.130 61.165 104.300 61.755 ;
        RECT 104.520 61.335 104.825 62.475 ;
        RECT 104.995 61.285 105.250 62.165 ;
        RECT 105.430 61.805 105.685 62.305 ;
        RECT 105.855 61.975 106.185 62.475 ;
        RECT 105.430 61.635 106.180 61.805 ;
        RECT 104.130 61.135 104.870 61.165 ;
        RECT 102.845 60.535 103.375 60.705 ;
        RECT 101.155 60.115 101.505 60.285 ;
        RECT 101.725 60.095 102.675 60.375 ;
        RECT 102.845 59.925 103.035 60.365 ;
        RECT 103.205 60.305 103.375 60.535 ;
        RECT 103.545 60.475 103.785 60.875 ;
        RECT 103.955 60.835 104.870 61.135 ;
        RECT 103.955 60.660 104.280 60.835 ;
        RECT 103.955 60.305 104.275 60.660 ;
        RECT 105.040 60.635 105.250 61.285 ;
        RECT 105.430 60.815 105.780 61.465 ;
        RECT 105.950 60.645 106.180 61.635 ;
        RECT 103.205 60.135 104.275 60.305 ;
        RECT 104.520 59.925 104.825 60.385 ;
        RECT 104.995 60.105 105.250 60.635 ;
        RECT 105.430 60.475 106.180 60.645 ;
        RECT 105.430 60.185 105.685 60.475 ;
        RECT 105.855 59.925 106.185 60.305 ;
        RECT 106.355 60.185 106.525 62.305 ;
        RECT 106.695 61.505 107.020 62.290 ;
        RECT 107.190 62.015 107.440 62.475 ;
        RECT 107.610 61.975 107.860 62.305 ;
        RECT 108.075 61.975 108.755 62.305 ;
        RECT 107.610 61.845 107.780 61.975 ;
        RECT 107.385 61.675 107.780 61.845 ;
        RECT 106.755 60.455 107.215 61.505 ;
        RECT 107.385 60.315 107.555 61.675 ;
        RECT 107.950 61.415 108.415 61.805 ;
        RECT 107.725 60.605 108.075 61.225 ;
        RECT 108.245 60.825 108.415 61.415 ;
        RECT 108.585 61.195 108.755 61.975 ;
        RECT 108.925 61.875 109.095 62.215 ;
        RECT 109.330 62.045 109.660 62.475 ;
        RECT 109.830 61.875 110.000 62.215 ;
        RECT 110.295 62.015 110.665 62.475 ;
        RECT 108.925 61.705 110.000 61.875 ;
        RECT 110.835 61.845 111.005 62.305 ;
        RECT 111.240 61.965 112.110 62.305 ;
        RECT 112.280 62.015 112.530 62.475 ;
        RECT 110.445 61.675 111.005 61.845 ;
        RECT 110.445 61.535 110.615 61.675 ;
        RECT 109.115 61.365 110.615 61.535 ;
        RECT 111.310 61.505 111.770 61.795 ;
        RECT 108.585 61.025 110.275 61.195 ;
        RECT 108.245 60.605 108.600 60.825 ;
        RECT 108.770 60.315 108.940 61.025 ;
        RECT 109.145 60.605 109.935 60.855 ;
        RECT 110.105 60.845 110.275 61.025 ;
        RECT 110.445 60.675 110.615 61.365 ;
        RECT 106.885 59.925 107.215 60.285 ;
        RECT 107.385 60.145 107.880 60.315 ;
        RECT 108.085 60.145 108.940 60.315 ;
        RECT 109.815 59.925 110.145 60.385 ;
        RECT 110.355 60.285 110.615 60.675 ;
        RECT 110.805 61.495 111.770 61.505 ;
        RECT 111.940 61.585 112.110 61.965 ;
        RECT 112.700 61.925 112.870 62.215 ;
        RECT 113.050 62.095 113.380 62.475 ;
        RECT 112.700 61.755 113.500 61.925 ;
        RECT 110.805 61.335 111.480 61.495 ;
        RECT 111.940 61.415 113.160 61.585 ;
        RECT 110.805 60.545 111.015 61.335 ;
        RECT 111.940 61.325 112.110 61.415 ;
        RECT 111.185 60.545 111.535 61.165 ;
        RECT 111.705 61.155 112.110 61.325 ;
        RECT 111.705 60.375 111.875 61.155 ;
        RECT 112.045 60.705 112.265 60.985 ;
        RECT 112.445 60.875 112.985 61.245 ;
        RECT 113.330 61.165 113.500 61.755 ;
        RECT 113.720 61.335 114.025 62.475 ;
        RECT 114.195 61.285 114.450 62.165 ;
        RECT 113.330 61.135 114.070 61.165 ;
        RECT 112.045 60.535 112.575 60.705 ;
        RECT 110.355 60.115 110.705 60.285 ;
        RECT 110.925 60.095 111.875 60.375 ;
        RECT 112.045 59.925 112.235 60.365 ;
        RECT 112.405 60.305 112.575 60.535 ;
        RECT 112.745 60.475 112.985 60.875 ;
        RECT 113.155 60.835 114.070 61.135 ;
        RECT 113.155 60.660 113.480 60.835 ;
        RECT 113.155 60.305 113.475 60.660 ;
        RECT 114.240 60.635 114.450 61.285 ;
        RECT 112.405 60.135 113.475 60.305 ;
        RECT 113.720 59.925 114.025 60.385 ;
        RECT 114.195 60.105 114.450 60.635 ;
        RECT 114.630 61.335 114.965 62.305 ;
        RECT 115.135 61.335 115.305 62.475 ;
        RECT 115.475 62.135 117.505 62.305 ;
        RECT 114.630 60.665 114.800 61.335 ;
        RECT 115.475 61.165 115.645 62.135 ;
        RECT 114.970 60.835 115.225 61.165 ;
        RECT 115.450 60.835 115.645 61.165 ;
        RECT 115.815 61.795 116.940 61.965 ;
        RECT 115.055 60.665 115.225 60.835 ;
        RECT 115.815 60.665 115.985 61.795 ;
        RECT 114.630 60.095 114.885 60.665 ;
        RECT 115.055 60.495 115.985 60.665 ;
        RECT 116.155 61.455 117.165 61.625 ;
        RECT 116.155 60.655 116.325 61.455 ;
        RECT 116.530 61.115 116.805 61.255 ;
        RECT 116.525 60.945 116.805 61.115 ;
        RECT 115.810 60.460 115.985 60.495 ;
        RECT 115.055 59.925 115.385 60.325 ;
        RECT 115.810 60.095 116.340 60.460 ;
        RECT 116.530 60.095 116.805 60.945 ;
        RECT 116.975 60.095 117.165 61.455 ;
        RECT 117.335 61.470 117.505 62.135 ;
        RECT 117.675 61.715 117.845 62.475 ;
        RECT 118.080 61.715 118.595 62.125 ;
        RECT 117.335 61.280 118.085 61.470 ;
        RECT 118.255 60.905 118.595 61.715 ;
        RECT 117.365 60.735 118.595 60.905 ;
        RECT 118.765 61.400 119.035 62.305 ;
        RECT 119.205 61.715 119.535 62.475 ;
        RECT 119.715 61.545 119.885 62.305 ;
        RECT 117.345 59.925 117.855 60.460 ;
        RECT 118.075 60.130 118.320 60.735 ;
        RECT 118.765 60.600 118.935 61.400 ;
        RECT 119.220 61.375 119.885 61.545 ;
        RECT 120.145 61.385 121.355 62.475 ;
        RECT 119.220 61.230 119.390 61.375 ;
        RECT 119.105 60.900 119.390 61.230 ;
        RECT 119.220 60.645 119.390 60.900 ;
        RECT 119.625 60.825 119.955 61.195 ;
        RECT 120.145 60.675 120.665 61.215 ;
        RECT 120.835 60.845 121.355 61.385 ;
        RECT 121.525 61.310 121.815 62.475 ;
        RECT 122.445 61.385 123.655 62.475 ;
        RECT 122.445 60.845 122.965 61.385 ;
        RECT 123.135 60.675 123.655 61.215 ;
        RECT 118.765 60.095 119.025 60.600 ;
        RECT 119.220 60.475 119.885 60.645 ;
        RECT 119.205 59.925 119.535 60.305 ;
        RECT 119.715 60.095 119.885 60.475 ;
        RECT 120.145 59.925 121.355 60.675 ;
        RECT 121.525 59.925 121.815 60.650 ;
        RECT 122.445 59.925 123.655 60.675 ;
        RECT 5.520 59.755 123.740 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.985 58.985 9.575 59.755 ;
        RECT 10.205 59.080 10.465 59.585 ;
        RECT 10.645 59.375 10.975 59.755 ;
        RECT 11.155 59.205 11.325 59.585 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 6.985 58.465 8.195 58.985 ;
        RECT 8.365 58.295 9.575 58.815 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 6.985 57.205 9.575 58.295 ;
        RECT 10.205 58.280 10.375 59.080 ;
        RECT 10.660 59.035 11.325 59.205 ;
        RECT 10.660 58.780 10.830 59.035 ;
        RECT 11.645 58.935 11.855 59.755 ;
        RECT 12.025 58.955 12.355 59.585 ;
        RECT 10.545 58.450 10.830 58.780 ;
        RECT 11.065 58.485 11.395 58.855 ;
        RECT 10.660 58.305 10.830 58.450 ;
        RECT 12.025 58.355 12.275 58.955 ;
        RECT 12.525 58.935 12.755 59.755 ;
        RECT 12.970 59.205 13.225 59.495 ;
        RECT 13.395 59.375 13.725 59.755 ;
        RECT 12.970 59.035 13.720 59.205 ;
        RECT 12.445 58.515 12.775 58.765 ;
        RECT 10.205 57.375 10.475 58.280 ;
        RECT 10.660 58.135 11.325 58.305 ;
        RECT 10.645 57.205 10.975 57.965 ;
        RECT 11.155 57.375 11.325 58.135 ;
        RECT 11.645 57.205 11.855 58.345 ;
        RECT 12.025 57.375 12.355 58.355 ;
        RECT 12.525 57.205 12.755 58.345 ;
        RECT 12.970 58.215 13.320 58.865 ;
        RECT 13.490 58.045 13.720 59.035 ;
        RECT 12.970 57.875 13.720 58.045 ;
        RECT 12.970 57.375 13.225 57.875 ;
        RECT 13.395 57.205 13.725 57.705 ;
        RECT 13.895 57.375 14.065 59.495 ;
        RECT 14.425 59.395 14.755 59.755 ;
        RECT 14.925 59.365 15.420 59.535 ;
        RECT 15.625 59.365 16.480 59.535 ;
        RECT 14.295 58.175 14.755 59.225 ;
        RECT 14.235 57.390 14.560 58.175 ;
        RECT 14.925 58.005 15.095 59.365 ;
        RECT 15.265 58.455 15.615 59.075 ;
        RECT 15.785 58.855 16.140 59.075 ;
        RECT 15.785 58.265 15.955 58.855 ;
        RECT 16.310 58.655 16.480 59.365 ;
        RECT 17.355 59.295 17.685 59.755 ;
        RECT 17.895 59.395 18.245 59.565 ;
        RECT 16.685 58.825 17.475 59.075 ;
        RECT 17.895 59.005 18.155 59.395 ;
        RECT 18.465 59.305 19.415 59.585 ;
        RECT 19.585 59.315 19.775 59.755 ;
        RECT 19.945 59.375 21.015 59.545 ;
        RECT 17.645 58.655 17.815 58.835 ;
        RECT 14.925 57.835 15.320 58.005 ;
        RECT 15.490 57.875 15.955 58.265 ;
        RECT 16.125 58.485 17.815 58.655 ;
        RECT 15.150 57.705 15.320 57.835 ;
        RECT 16.125 57.705 16.295 58.485 ;
        RECT 17.985 58.315 18.155 59.005 ;
        RECT 16.655 58.145 18.155 58.315 ;
        RECT 18.345 58.345 18.555 59.135 ;
        RECT 18.725 58.515 19.075 59.135 ;
        RECT 19.245 58.525 19.415 59.305 ;
        RECT 19.945 59.145 20.115 59.375 ;
        RECT 19.585 58.975 20.115 59.145 ;
        RECT 19.585 58.695 19.805 58.975 ;
        RECT 20.285 58.805 20.525 59.205 ;
        RECT 19.245 58.355 19.650 58.525 ;
        RECT 19.985 58.435 20.525 58.805 ;
        RECT 20.695 59.020 21.015 59.375 ;
        RECT 21.260 59.295 21.565 59.755 ;
        RECT 21.735 59.045 21.990 59.575 ;
        RECT 20.695 58.845 21.020 59.020 ;
        RECT 20.695 58.545 21.610 58.845 ;
        RECT 20.870 58.515 21.610 58.545 ;
        RECT 18.345 58.185 19.020 58.345 ;
        RECT 19.480 58.265 19.650 58.355 ;
        RECT 18.345 58.175 19.310 58.185 ;
        RECT 17.985 58.005 18.155 58.145 ;
        RECT 14.730 57.205 14.980 57.665 ;
        RECT 15.150 57.375 15.400 57.705 ;
        RECT 15.615 57.375 16.295 57.705 ;
        RECT 16.465 57.805 17.540 57.975 ;
        RECT 17.985 57.835 18.545 58.005 ;
        RECT 18.850 57.885 19.310 58.175 ;
        RECT 19.480 58.095 20.700 58.265 ;
        RECT 16.465 57.465 16.635 57.805 ;
        RECT 16.870 57.205 17.200 57.635 ;
        RECT 17.370 57.465 17.540 57.805 ;
        RECT 17.835 57.205 18.205 57.665 ;
        RECT 18.375 57.375 18.545 57.835 ;
        RECT 19.480 57.715 19.650 58.095 ;
        RECT 20.870 57.925 21.040 58.515 ;
        RECT 21.780 58.395 21.990 59.045 ;
        RECT 22.170 59.205 22.425 59.495 ;
        RECT 22.595 59.375 22.925 59.755 ;
        RECT 22.170 59.035 22.920 59.205 ;
        RECT 18.780 57.375 19.650 57.715 ;
        RECT 20.240 57.755 21.040 57.925 ;
        RECT 19.820 57.205 20.070 57.665 ;
        RECT 20.240 57.465 20.410 57.755 ;
        RECT 20.590 57.205 20.920 57.585 ;
        RECT 21.260 57.205 21.565 58.345 ;
        RECT 21.735 57.515 21.990 58.395 ;
        RECT 22.170 58.215 22.520 58.865 ;
        RECT 22.690 58.045 22.920 59.035 ;
        RECT 22.170 57.875 22.920 58.045 ;
        RECT 22.170 57.375 22.425 57.875 ;
        RECT 22.595 57.205 22.925 57.705 ;
        RECT 23.095 57.375 23.265 59.495 ;
        RECT 23.625 59.395 23.955 59.755 ;
        RECT 24.125 59.365 24.620 59.535 ;
        RECT 24.825 59.365 25.680 59.535 ;
        RECT 23.495 58.175 23.955 59.225 ;
        RECT 23.435 57.390 23.760 58.175 ;
        RECT 24.125 58.005 24.295 59.365 ;
        RECT 24.465 58.455 24.815 59.075 ;
        RECT 24.985 58.855 25.340 59.075 ;
        RECT 24.985 58.265 25.155 58.855 ;
        RECT 25.510 58.655 25.680 59.365 ;
        RECT 26.555 59.295 26.885 59.755 ;
        RECT 27.095 59.395 27.445 59.565 ;
        RECT 25.885 58.825 26.675 59.075 ;
        RECT 27.095 59.005 27.355 59.395 ;
        RECT 27.665 59.305 28.615 59.585 ;
        RECT 28.785 59.315 28.975 59.755 ;
        RECT 29.145 59.375 30.215 59.545 ;
        RECT 26.845 58.655 27.015 58.835 ;
        RECT 24.125 57.835 24.520 58.005 ;
        RECT 24.690 57.875 25.155 58.265 ;
        RECT 25.325 58.485 27.015 58.655 ;
        RECT 24.350 57.705 24.520 57.835 ;
        RECT 25.325 57.705 25.495 58.485 ;
        RECT 27.185 58.315 27.355 59.005 ;
        RECT 25.855 58.145 27.355 58.315 ;
        RECT 27.545 58.345 27.755 59.135 ;
        RECT 27.925 58.515 28.275 59.135 ;
        RECT 28.445 58.525 28.615 59.305 ;
        RECT 29.145 59.145 29.315 59.375 ;
        RECT 28.785 58.975 29.315 59.145 ;
        RECT 28.785 58.695 29.005 58.975 ;
        RECT 29.485 58.805 29.725 59.205 ;
        RECT 28.445 58.355 28.850 58.525 ;
        RECT 29.185 58.435 29.725 58.805 ;
        RECT 29.895 59.020 30.215 59.375 ;
        RECT 30.460 59.295 30.765 59.755 ;
        RECT 30.935 59.045 31.190 59.575 ;
        RECT 29.895 58.845 30.220 59.020 ;
        RECT 29.895 58.545 30.810 58.845 ;
        RECT 30.070 58.515 30.810 58.545 ;
        RECT 27.545 58.185 28.220 58.345 ;
        RECT 28.680 58.265 28.850 58.355 ;
        RECT 27.545 58.175 28.510 58.185 ;
        RECT 27.185 58.005 27.355 58.145 ;
        RECT 23.930 57.205 24.180 57.665 ;
        RECT 24.350 57.375 24.600 57.705 ;
        RECT 24.815 57.375 25.495 57.705 ;
        RECT 25.665 57.805 26.740 57.975 ;
        RECT 27.185 57.835 27.745 58.005 ;
        RECT 28.050 57.885 28.510 58.175 ;
        RECT 28.680 58.095 29.900 58.265 ;
        RECT 25.665 57.465 25.835 57.805 ;
        RECT 26.070 57.205 26.400 57.635 ;
        RECT 26.570 57.465 26.740 57.805 ;
        RECT 27.035 57.205 27.405 57.665 ;
        RECT 27.575 57.375 27.745 57.835 ;
        RECT 28.680 57.715 28.850 58.095 ;
        RECT 30.070 57.925 30.240 58.515 ;
        RECT 30.980 58.395 31.190 59.045 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.825 58.985 35.335 59.755 ;
        RECT 36.425 59.080 36.685 59.585 ;
        RECT 36.865 59.375 37.195 59.755 ;
        RECT 37.375 59.205 37.545 59.585 ;
        RECT 31.825 58.465 33.475 58.985 ;
        RECT 27.980 57.375 28.850 57.715 ;
        RECT 29.440 57.755 30.240 57.925 ;
        RECT 29.020 57.205 29.270 57.665 ;
        RECT 29.440 57.465 29.610 57.755 ;
        RECT 29.790 57.205 30.120 57.585 ;
        RECT 30.460 57.205 30.765 58.345 ;
        RECT 30.935 57.515 31.190 58.395 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 33.645 58.295 35.335 58.815 ;
        RECT 31.825 57.205 35.335 58.295 ;
        RECT 36.425 58.280 36.595 59.080 ;
        RECT 36.880 59.035 37.545 59.205 ;
        RECT 36.880 58.780 37.050 59.035 ;
        RECT 37.810 59.015 38.065 59.585 ;
        RECT 38.235 59.355 38.565 59.755 ;
        RECT 38.990 59.220 39.520 59.585 ;
        RECT 38.990 59.185 39.165 59.220 ;
        RECT 38.235 59.015 39.165 59.185 ;
        RECT 36.765 58.450 37.050 58.780 ;
        RECT 37.285 58.485 37.615 58.855 ;
        RECT 36.880 58.305 37.050 58.450 ;
        RECT 37.810 58.345 37.980 59.015 ;
        RECT 38.235 58.845 38.405 59.015 ;
        RECT 38.150 58.515 38.405 58.845 ;
        RECT 38.630 58.515 38.825 58.845 ;
        RECT 36.425 57.375 36.695 58.280 ;
        RECT 36.880 58.135 37.545 58.305 ;
        RECT 36.865 57.205 37.195 57.965 ;
        RECT 37.375 57.375 37.545 58.135 ;
        RECT 37.810 57.375 38.145 58.345 ;
        RECT 38.315 57.205 38.485 58.345 ;
        RECT 38.655 57.545 38.825 58.515 ;
        RECT 38.995 57.885 39.165 59.015 ;
        RECT 39.335 58.225 39.505 59.025 ;
        RECT 39.710 58.735 39.985 59.585 ;
        RECT 39.705 58.565 39.985 58.735 ;
        RECT 39.710 58.425 39.985 58.565 ;
        RECT 40.155 58.225 40.345 59.585 ;
        RECT 40.525 59.220 41.035 59.755 ;
        RECT 41.255 58.945 41.500 59.550 ;
        RECT 42.955 59.205 43.125 59.495 ;
        RECT 43.295 59.375 43.625 59.755 ;
        RECT 42.955 59.035 43.620 59.205 ;
        RECT 40.545 58.775 41.775 58.945 ;
        RECT 39.335 58.055 40.345 58.225 ;
        RECT 40.515 58.210 41.265 58.400 ;
        RECT 38.995 57.715 40.120 57.885 ;
        RECT 40.515 57.545 40.685 58.210 ;
        RECT 41.435 57.965 41.775 58.775 ;
        RECT 42.870 58.215 43.220 58.865 ;
        RECT 43.390 58.045 43.620 59.035 ;
        RECT 38.655 57.375 40.685 57.545 ;
        RECT 40.855 57.205 41.025 57.965 ;
        RECT 41.260 57.555 41.775 57.965 ;
        RECT 42.955 57.875 43.620 58.045 ;
        RECT 42.955 57.375 43.125 57.875 ;
        RECT 43.295 57.205 43.625 57.705 ;
        RECT 43.795 57.375 44.020 59.495 ;
        RECT 44.235 59.375 44.565 59.755 ;
        RECT 44.735 59.205 44.905 59.535 ;
        RECT 45.205 59.375 46.220 59.575 ;
        RECT 44.210 59.015 44.905 59.205 ;
        RECT 44.210 58.045 44.380 59.015 ;
        RECT 44.550 58.215 44.960 58.835 ;
        RECT 45.130 58.265 45.350 59.135 ;
        RECT 45.530 58.825 45.880 59.195 ;
        RECT 46.050 58.645 46.220 59.375 ;
        RECT 46.390 59.315 46.800 59.755 ;
        RECT 47.090 59.115 47.340 59.545 ;
        RECT 47.540 59.295 47.860 59.755 ;
        RECT 48.420 59.365 49.270 59.535 ;
        RECT 46.390 58.775 46.800 59.105 ;
        RECT 47.090 58.775 47.510 59.115 ;
        RECT 45.800 58.605 46.220 58.645 ;
        RECT 45.800 58.435 47.150 58.605 ;
        RECT 44.210 57.875 44.905 58.045 ;
        RECT 45.130 57.885 45.630 58.265 ;
        RECT 44.235 57.205 44.565 57.705 ;
        RECT 44.735 57.375 44.905 57.875 ;
        RECT 45.800 57.590 45.970 58.435 ;
        RECT 46.900 58.275 47.150 58.435 ;
        RECT 46.140 58.005 46.390 58.265 ;
        RECT 47.320 58.005 47.510 58.775 ;
        RECT 46.140 57.755 47.510 58.005 ;
        RECT 47.680 58.945 48.930 59.115 ;
        RECT 47.680 58.185 47.850 58.945 ;
        RECT 48.600 58.825 48.930 58.945 ;
        RECT 48.020 58.365 48.200 58.775 ;
        RECT 49.100 58.605 49.270 59.365 ;
        RECT 49.470 59.275 50.130 59.755 ;
        RECT 50.310 59.160 50.630 59.490 ;
        RECT 49.460 58.835 50.120 59.105 ;
        RECT 49.460 58.775 49.790 58.835 ;
        RECT 49.940 58.605 50.270 58.665 ;
        RECT 48.370 58.435 50.270 58.605 ;
        RECT 47.680 57.875 48.200 58.185 ;
        RECT 48.370 57.925 48.540 58.435 ;
        RECT 50.440 58.265 50.630 59.160 ;
        RECT 48.710 58.095 50.630 58.265 ;
        RECT 50.310 58.075 50.630 58.095 ;
        RECT 50.830 58.845 51.080 59.495 ;
        RECT 51.260 59.295 51.545 59.755 ;
        RECT 51.725 59.075 51.980 59.575 ;
        RECT 51.725 59.045 52.065 59.075 ;
        RECT 51.800 58.905 52.065 59.045 ;
        RECT 52.530 59.015 52.785 59.585 ;
        RECT 52.955 59.355 53.285 59.755 ;
        RECT 53.710 59.220 54.240 59.585 ;
        RECT 54.430 59.415 54.705 59.585 ;
        RECT 54.425 59.245 54.705 59.415 ;
        RECT 53.710 59.185 53.885 59.220 ;
        RECT 52.955 59.015 53.885 59.185 ;
        RECT 50.830 58.515 51.630 58.845 ;
        RECT 48.370 57.755 49.580 57.925 ;
        RECT 45.140 57.420 45.970 57.590 ;
        RECT 46.210 57.205 46.590 57.585 ;
        RECT 46.770 57.465 46.940 57.755 ;
        RECT 48.370 57.675 48.540 57.755 ;
        RECT 47.110 57.205 47.440 57.585 ;
        RECT 47.910 57.425 48.540 57.675 ;
        RECT 48.720 57.205 49.140 57.585 ;
        RECT 49.340 57.465 49.580 57.755 ;
        RECT 49.810 57.205 50.140 57.895 ;
        RECT 50.310 57.465 50.480 58.075 ;
        RECT 50.830 57.925 51.080 58.515 ;
        RECT 51.800 58.185 51.980 58.905 ;
        RECT 50.750 57.415 51.080 57.925 ;
        RECT 51.260 57.205 51.545 58.005 ;
        RECT 51.725 57.515 51.980 58.185 ;
        RECT 52.530 58.345 52.700 59.015 ;
        RECT 52.955 58.845 53.125 59.015 ;
        RECT 52.870 58.515 53.125 58.845 ;
        RECT 53.350 58.515 53.545 58.845 ;
        RECT 52.530 57.375 52.865 58.345 ;
        RECT 53.035 57.205 53.205 58.345 ;
        RECT 53.375 57.545 53.545 58.515 ;
        RECT 53.715 57.885 53.885 59.015 ;
        RECT 54.055 58.225 54.225 59.025 ;
        RECT 54.430 58.425 54.705 59.245 ;
        RECT 54.875 58.225 55.065 59.585 ;
        RECT 55.245 59.220 55.755 59.755 ;
        RECT 55.975 58.945 56.220 59.550 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 57.585 59.210 62.930 59.755 ;
        RECT 63.105 59.210 68.450 59.755 ;
        RECT 68.625 59.210 73.970 59.755 ;
        RECT 55.265 58.775 56.495 58.945 ;
        RECT 54.055 58.055 55.065 58.225 ;
        RECT 55.235 58.210 55.985 58.400 ;
        RECT 53.715 57.715 54.840 57.885 ;
        RECT 55.235 57.545 55.405 58.210 ;
        RECT 56.155 57.965 56.495 58.775 ;
        RECT 59.170 58.380 59.510 59.210 ;
        RECT 53.375 57.375 55.405 57.545 ;
        RECT 55.575 57.205 55.745 57.965 ;
        RECT 55.980 57.555 56.495 57.965 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 60.990 57.640 61.340 58.890 ;
        RECT 64.690 58.380 65.030 59.210 ;
        RECT 66.510 57.640 66.860 58.890 ;
        RECT 70.210 58.380 70.550 59.210 ;
        RECT 74.145 59.005 75.355 59.755 ;
        RECT 75.615 59.105 75.785 59.585 ;
        RECT 75.965 59.275 76.205 59.755 ;
        RECT 76.455 59.105 76.625 59.585 ;
        RECT 76.795 59.275 77.125 59.755 ;
        RECT 77.295 59.105 77.465 59.585 ;
        RECT 72.030 57.640 72.380 58.890 ;
        RECT 74.145 58.465 74.665 59.005 ;
        RECT 75.615 58.935 76.250 59.105 ;
        RECT 76.455 58.935 77.465 59.105 ;
        RECT 77.635 58.955 77.965 59.755 ;
        RECT 78.285 58.985 81.795 59.755 ;
        RECT 82.885 59.030 83.175 59.755 ;
        RECT 83.435 59.105 83.605 59.585 ;
        RECT 83.785 59.275 84.025 59.755 ;
        RECT 84.275 59.105 84.445 59.585 ;
        RECT 84.615 59.275 84.945 59.755 ;
        RECT 85.115 59.105 85.285 59.585 ;
        RECT 74.835 58.295 75.355 58.835 ;
        RECT 76.080 58.765 76.250 58.935 ;
        RECT 76.965 58.905 77.465 58.935 ;
        RECT 75.530 58.525 75.910 58.765 ;
        RECT 76.080 58.595 76.580 58.765 ;
        RECT 76.080 58.355 76.250 58.595 ;
        RECT 76.970 58.395 77.465 58.905 ;
        RECT 78.285 58.465 79.935 58.985 ;
        RECT 83.435 58.935 84.070 59.105 ;
        RECT 84.275 58.935 85.285 59.105 ;
        RECT 85.455 58.955 85.785 59.755 ;
        RECT 86.105 58.985 89.615 59.755 ;
        RECT 57.585 57.205 62.930 57.640 ;
        RECT 63.105 57.205 68.450 57.640 ;
        RECT 68.625 57.205 73.970 57.640 ;
        RECT 74.145 57.205 75.355 58.295 ;
        RECT 75.535 58.185 76.250 58.355 ;
        RECT 76.455 58.225 77.465 58.395 ;
        RECT 75.535 57.375 75.865 58.185 ;
        RECT 76.035 57.205 76.275 58.005 ;
        RECT 76.455 57.375 76.625 58.225 ;
        RECT 76.795 57.205 77.125 58.005 ;
        RECT 77.295 57.375 77.465 58.225 ;
        RECT 77.635 57.205 77.965 58.355 ;
        RECT 80.105 58.295 81.795 58.815 ;
        RECT 83.900 58.765 84.070 58.935 ;
        RECT 83.350 58.525 83.730 58.765 ;
        RECT 83.900 58.595 84.400 58.765 ;
        RECT 84.790 58.735 85.285 58.935 ;
        RECT 78.285 57.205 81.795 58.295 ;
        RECT 82.885 57.205 83.175 58.370 ;
        RECT 83.900 58.355 84.070 58.595 ;
        RECT 84.785 58.565 85.285 58.735 ;
        RECT 84.790 58.395 85.285 58.565 ;
        RECT 86.105 58.465 87.755 58.985 ;
        RECT 89.825 58.935 90.055 59.755 ;
        RECT 90.225 58.955 90.555 59.585 ;
        RECT 83.355 58.185 84.070 58.355 ;
        RECT 84.275 58.225 85.285 58.395 ;
        RECT 83.355 57.375 83.685 58.185 ;
        RECT 83.855 57.205 84.095 58.005 ;
        RECT 84.275 57.375 84.445 58.225 ;
        RECT 84.615 57.205 84.945 58.005 ;
        RECT 85.115 57.375 85.285 58.225 ;
        RECT 85.455 57.205 85.785 58.355 ;
        RECT 87.925 58.295 89.615 58.815 ;
        RECT 89.805 58.515 90.135 58.765 ;
        RECT 90.305 58.355 90.555 58.955 ;
        RECT 90.725 58.935 90.935 59.755 ;
        RECT 91.165 59.210 96.510 59.755 ;
        RECT 92.750 58.380 93.090 59.210 ;
        RECT 96.685 58.985 99.275 59.755 ;
        RECT 99.535 59.205 99.705 59.585 ;
        RECT 99.885 59.375 100.215 59.755 ;
        RECT 99.535 59.035 100.200 59.205 ;
        RECT 100.395 59.080 100.655 59.585 ;
        RECT 86.105 57.205 89.615 58.295 ;
        RECT 89.825 57.205 90.055 58.345 ;
        RECT 90.225 57.375 90.555 58.355 ;
        RECT 90.725 57.205 90.935 58.345 ;
        RECT 94.570 57.640 94.920 58.890 ;
        RECT 96.685 58.465 97.895 58.985 ;
        RECT 98.065 58.295 99.275 58.815 ;
        RECT 99.465 58.485 99.795 58.855 ;
        RECT 100.030 58.780 100.200 59.035 ;
        RECT 100.030 58.450 100.315 58.780 ;
        RECT 100.030 58.305 100.200 58.450 ;
        RECT 91.165 57.205 96.510 57.640 ;
        RECT 96.685 57.205 99.275 58.295 ;
        RECT 99.535 58.135 100.200 58.305 ;
        RECT 100.485 58.280 100.655 59.080 ;
        RECT 100.865 58.935 101.095 59.755 ;
        RECT 101.265 58.955 101.595 59.585 ;
        RECT 100.845 58.515 101.175 58.765 ;
        RECT 101.345 58.355 101.595 58.955 ;
        RECT 101.765 58.935 101.975 59.755 ;
        RECT 102.205 58.985 105.715 59.755 ;
        RECT 102.205 58.465 103.855 58.985 ;
        RECT 105.925 58.935 106.155 59.755 ;
        RECT 106.325 58.955 106.655 59.585 ;
        RECT 99.535 57.375 99.705 58.135 ;
        RECT 99.885 57.205 100.215 57.965 ;
        RECT 100.385 57.375 100.655 58.280 ;
        RECT 100.865 57.205 101.095 58.345 ;
        RECT 101.265 57.375 101.595 58.355 ;
        RECT 101.765 57.205 101.975 58.345 ;
        RECT 104.025 58.295 105.715 58.815 ;
        RECT 105.905 58.515 106.235 58.765 ;
        RECT 106.405 58.355 106.655 58.955 ;
        RECT 106.825 58.935 107.035 59.755 ;
        RECT 107.355 59.205 107.525 59.585 ;
        RECT 107.705 59.375 108.035 59.755 ;
        RECT 107.355 59.035 108.020 59.205 ;
        RECT 108.215 59.080 108.475 59.585 ;
        RECT 107.285 58.485 107.615 58.855 ;
        RECT 107.850 58.780 108.020 59.035 ;
        RECT 102.205 57.205 105.715 58.295 ;
        RECT 105.925 57.205 106.155 58.345 ;
        RECT 106.325 57.375 106.655 58.355 ;
        RECT 107.850 58.450 108.135 58.780 ;
        RECT 106.825 57.205 107.035 58.345 ;
        RECT 107.850 58.305 108.020 58.450 ;
        RECT 107.355 58.135 108.020 58.305 ;
        RECT 108.305 58.280 108.475 59.080 ;
        RECT 108.645 59.030 108.935 59.755 ;
        RECT 109.110 59.205 109.365 59.495 ;
        RECT 109.535 59.375 109.865 59.755 ;
        RECT 109.110 59.035 109.860 59.205 ;
        RECT 107.355 57.375 107.525 58.135 ;
        RECT 107.705 57.205 108.035 57.965 ;
        RECT 108.205 57.375 108.475 58.280 ;
        RECT 108.645 57.205 108.935 58.370 ;
        RECT 109.110 58.215 109.460 58.865 ;
        RECT 109.630 58.045 109.860 59.035 ;
        RECT 109.110 57.875 109.860 58.045 ;
        RECT 109.110 57.375 109.365 57.875 ;
        RECT 109.535 57.205 109.865 57.705 ;
        RECT 110.035 57.375 110.205 59.495 ;
        RECT 110.565 59.395 110.895 59.755 ;
        RECT 111.065 59.365 111.560 59.535 ;
        RECT 111.765 59.365 112.620 59.535 ;
        RECT 110.435 58.175 110.895 59.225 ;
        RECT 110.375 57.390 110.700 58.175 ;
        RECT 111.065 58.005 111.235 59.365 ;
        RECT 111.405 58.455 111.755 59.075 ;
        RECT 111.925 58.855 112.280 59.075 ;
        RECT 111.925 58.265 112.095 58.855 ;
        RECT 112.450 58.655 112.620 59.365 ;
        RECT 113.495 59.295 113.825 59.755 ;
        RECT 114.035 59.395 114.385 59.565 ;
        RECT 112.825 58.825 113.615 59.075 ;
        RECT 114.035 59.005 114.295 59.395 ;
        RECT 114.605 59.305 115.555 59.585 ;
        RECT 115.725 59.315 115.915 59.755 ;
        RECT 116.085 59.375 117.155 59.545 ;
        RECT 113.785 58.655 113.955 58.835 ;
        RECT 111.065 57.835 111.460 58.005 ;
        RECT 111.630 57.875 112.095 58.265 ;
        RECT 112.265 58.485 113.955 58.655 ;
        RECT 111.290 57.705 111.460 57.835 ;
        RECT 112.265 57.705 112.435 58.485 ;
        RECT 114.125 58.315 114.295 59.005 ;
        RECT 112.795 58.145 114.295 58.315 ;
        RECT 114.485 58.345 114.695 59.135 ;
        RECT 114.865 58.515 115.215 59.135 ;
        RECT 115.385 58.525 115.555 59.305 ;
        RECT 116.085 59.145 116.255 59.375 ;
        RECT 115.725 58.975 116.255 59.145 ;
        RECT 115.725 58.695 115.945 58.975 ;
        RECT 116.425 58.805 116.665 59.205 ;
        RECT 115.385 58.355 115.790 58.525 ;
        RECT 116.125 58.435 116.665 58.805 ;
        RECT 116.835 59.020 117.155 59.375 ;
        RECT 117.400 59.295 117.705 59.755 ;
        RECT 117.875 59.045 118.130 59.575 ;
        RECT 116.835 58.845 117.160 59.020 ;
        RECT 116.835 58.545 117.750 58.845 ;
        RECT 117.010 58.515 117.750 58.545 ;
        RECT 114.485 58.185 115.160 58.345 ;
        RECT 115.620 58.265 115.790 58.355 ;
        RECT 114.485 58.175 115.450 58.185 ;
        RECT 114.125 58.005 114.295 58.145 ;
        RECT 110.870 57.205 111.120 57.665 ;
        RECT 111.290 57.375 111.540 57.705 ;
        RECT 111.755 57.375 112.435 57.705 ;
        RECT 112.605 57.805 113.680 57.975 ;
        RECT 114.125 57.835 114.685 58.005 ;
        RECT 114.990 57.885 115.450 58.175 ;
        RECT 115.620 58.095 116.840 58.265 ;
        RECT 112.605 57.465 112.775 57.805 ;
        RECT 113.010 57.205 113.340 57.635 ;
        RECT 113.510 57.465 113.680 57.805 ;
        RECT 113.975 57.205 114.345 57.665 ;
        RECT 114.515 57.375 114.685 57.835 ;
        RECT 115.620 57.715 115.790 58.095 ;
        RECT 117.010 57.925 117.180 58.515 ;
        RECT 117.920 58.395 118.130 59.045 ;
        RECT 118.345 58.935 118.575 59.755 ;
        RECT 118.745 58.955 119.075 59.585 ;
        RECT 118.325 58.515 118.655 58.765 ;
        RECT 114.920 57.375 115.790 57.715 ;
        RECT 116.380 57.755 117.180 57.925 ;
        RECT 115.960 57.205 116.210 57.665 ;
        RECT 116.380 57.465 116.550 57.755 ;
        RECT 116.730 57.205 117.060 57.585 ;
        RECT 117.400 57.205 117.705 58.345 ;
        RECT 117.875 57.515 118.130 58.395 ;
        RECT 118.825 58.355 119.075 58.955 ;
        RECT 119.245 58.935 119.455 59.755 ;
        RECT 119.685 58.985 122.275 59.755 ;
        RECT 122.445 59.005 123.655 59.755 ;
        RECT 119.685 58.465 120.895 58.985 ;
        RECT 118.345 57.205 118.575 58.345 ;
        RECT 118.745 57.375 119.075 58.355 ;
        RECT 119.245 57.205 119.455 58.345 ;
        RECT 121.065 58.295 122.275 58.815 ;
        RECT 119.685 57.205 122.275 58.295 ;
        RECT 122.445 58.295 122.965 58.835 ;
        RECT 123.135 58.465 123.655 59.005 ;
        RECT 122.445 57.205 123.655 58.295 ;
        RECT 5.520 57.035 123.740 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 6.985 55.945 8.655 57.035 ;
        RECT 9.290 56.365 9.545 56.865 ;
        RECT 9.715 56.535 10.045 57.035 ;
        RECT 9.290 56.195 10.040 56.365 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 6.985 55.255 7.735 55.775 ;
        RECT 7.905 55.425 8.655 55.945 ;
        RECT 9.290 55.375 9.640 56.025 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 6.985 54.485 8.655 55.255 ;
        RECT 9.810 55.205 10.040 56.195 ;
        RECT 9.290 55.035 10.040 55.205 ;
        RECT 9.290 54.745 9.545 55.035 ;
        RECT 9.715 54.485 10.045 54.865 ;
        RECT 10.215 54.745 10.385 56.865 ;
        RECT 10.555 56.065 10.880 56.850 ;
        RECT 11.050 56.575 11.300 57.035 ;
        RECT 11.470 56.535 11.720 56.865 ;
        RECT 11.935 56.535 12.615 56.865 ;
        RECT 11.470 56.405 11.640 56.535 ;
        RECT 11.245 56.235 11.640 56.405 ;
        RECT 10.615 55.015 11.075 56.065 ;
        RECT 11.245 54.875 11.415 56.235 ;
        RECT 11.810 55.975 12.275 56.365 ;
        RECT 11.585 55.165 11.935 55.785 ;
        RECT 12.105 55.385 12.275 55.975 ;
        RECT 12.445 55.755 12.615 56.535 ;
        RECT 12.785 56.435 12.955 56.775 ;
        RECT 13.190 56.605 13.520 57.035 ;
        RECT 13.690 56.435 13.860 56.775 ;
        RECT 14.155 56.575 14.525 57.035 ;
        RECT 12.785 56.265 13.860 56.435 ;
        RECT 14.695 56.405 14.865 56.865 ;
        RECT 15.100 56.525 15.970 56.865 ;
        RECT 16.140 56.575 16.390 57.035 ;
        RECT 14.305 56.235 14.865 56.405 ;
        RECT 14.305 56.095 14.475 56.235 ;
        RECT 12.975 55.925 14.475 56.095 ;
        RECT 15.170 56.065 15.630 56.355 ;
        RECT 12.445 55.585 14.135 55.755 ;
        RECT 12.105 55.165 12.460 55.385 ;
        RECT 12.630 54.875 12.800 55.585 ;
        RECT 13.005 55.165 13.795 55.415 ;
        RECT 13.965 55.405 14.135 55.585 ;
        RECT 14.305 55.235 14.475 55.925 ;
        RECT 10.745 54.485 11.075 54.845 ;
        RECT 11.245 54.705 11.740 54.875 ;
        RECT 11.945 54.705 12.800 54.875 ;
        RECT 13.675 54.485 14.005 54.945 ;
        RECT 14.215 54.845 14.475 55.235 ;
        RECT 14.665 56.055 15.630 56.065 ;
        RECT 15.800 56.145 15.970 56.525 ;
        RECT 16.560 56.485 16.730 56.775 ;
        RECT 16.910 56.655 17.240 57.035 ;
        RECT 16.560 56.315 17.360 56.485 ;
        RECT 14.665 55.895 15.340 56.055 ;
        RECT 15.800 55.975 17.020 56.145 ;
        RECT 14.665 55.105 14.875 55.895 ;
        RECT 15.800 55.885 15.970 55.975 ;
        RECT 15.045 55.105 15.395 55.725 ;
        RECT 15.565 55.715 15.970 55.885 ;
        RECT 15.565 54.935 15.735 55.715 ;
        RECT 15.905 55.265 16.125 55.545 ;
        RECT 16.305 55.435 16.845 55.805 ;
        RECT 17.190 55.725 17.360 56.315 ;
        RECT 17.580 55.895 17.885 57.035 ;
        RECT 18.055 55.845 18.310 56.725 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 19.005 55.895 19.215 57.035 ;
        RECT 19.385 55.885 19.715 56.865 ;
        RECT 19.885 55.895 20.115 57.035 ;
        RECT 20.875 56.105 21.045 56.865 ;
        RECT 21.225 56.275 21.555 57.035 ;
        RECT 20.875 55.935 21.540 56.105 ;
        RECT 21.725 55.960 21.995 56.865 ;
        RECT 22.165 56.065 22.425 57.035 ;
        RECT 17.190 55.695 17.930 55.725 ;
        RECT 15.905 55.095 16.435 55.265 ;
        RECT 14.215 54.675 14.565 54.845 ;
        RECT 14.785 54.655 15.735 54.935 ;
        RECT 15.905 54.485 16.095 54.925 ;
        RECT 16.265 54.865 16.435 55.095 ;
        RECT 16.605 55.035 16.845 55.435 ;
        RECT 17.015 55.395 17.930 55.695 ;
        RECT 17.015 55.220 17.340 55.395 ;
        RECT 17.015 54.865 17.335 55.220 ;
        RECT 18.100 55.195 18.310 55.845 ;
        RECT 16.265 54.695 17.335 54.865 ;
        RECT 17.580 54.485 17.885 54.945 ;
        RECT 18.055 54.665 18.310 55.195 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 19.005 54.485 19.215 55.305 ;
        RECT 19.385 55.285 19.635 55.885 ;
        RECT 21.370 55.790 21.540 55.935 ;
        RECT 19.805 55.475 20.135 55.725 ;
        RECT 20.805 55.385 21.135 55.755 ;
        RECT 21.370 55.460 21.655 55.790 ;
        RECT 19.385 54.655 19.715 55.285 ;
        RECT 19.885 54.485 20.115 55.305 ;
        RECT 21.370 55.205 21.540 55.460 ;
        RECT 20.875 55.035 21.540 55.205 ;
        RECT 21.825 55.160 21.995 55.960 ;
        RECT 20.875 54.655 21.045 55.035 ;
        RECT 21.225 54.485 21.555 54.865 ;
        RECT 21.735 54.655 21.995 55.160 ;
        RECT 22.165 54.775 22.405 55.725 ;
        RECT 22.595 55.690 22.925 56.865 ;
        RECT 23.095 56.065 23.375 57.035 ;
        RECT 23.635 56.290 23.905 57.035 ;
        RECT 24.535 57.030 30.810 57.035 ;
        RECT 24.075 56.120 24.365 56.860 ;
        RECT 24.535 56.305 24.790 57.030 ;
        RECT 24.975 56.135 25.235 56.860 ;
        RECT 25.405 56.305 25.650 57.030 ;
        RECT 25.835 56.135 26.095 56.860 ;
        RECT 26.265 56.305 26.510 57.030 ;
        RECT 26.695 56.135 26.955 56.860 ;
        RECT 27.125 56.305 27.370 57.030 ;
        RECT 27.540 56.135 27.800 56.860 ;
        RECT 27.970 56.305 28.230 57.030 ;
        RECT 28.400 56.135 28.660 56.860 ;
        RECT 28.830 56.305 29.090 57.030 ;
        RECT 29.260 56.135 29.520 56.860 ;
        RECT 29.690 56.305 29.950 57.030 ;
        RECT 30.120 56.135 30.380 56.860 ;
        RECT 30.550 56.235 30.810 57.030 ;
        RECT 24.975 56.120 30.380 56.135 ;
        RECT 23.635 55.895 30.380 56.120 ;
        RECT 22.595 55.160 23.375 55.690 ;
        RECT 23.635 55.675 24.800 55.895 ;
        RECT 30.980 55.725 31.230 56.860 ;
        RECT 31.410 56.225 31.670 57.035 ;
        RECT 31.845 55.725 32.090 56.865 ;
        RECT 32.270 56.225 32.565 57.035 ;
        RECT 33.670 56.365 33.925 56.865 ;
        RECT 34.095 56.535 34.425 57.035 ;
        RECT 33.670 56.195 34.420 56.365 ;
        RECT 23.605 55.505 24.800 55.675 ;
        RECT 23.635 55.305 24.800 55.505 ;
        RECT 24.970 55.475 32.090 55.725 ;
        RECT 22.595 54.655 22.920 55.160 ;
        RECT 23.635 55.135 30.380 55.305 ;
        RECT 23.090 54.485 23.375 54.990 ;
        RECT 23.635 54.485 23.935 54.965 ;
        RECT 24.105 54.680 24.365 55.135 ;
        RECT 24.535 54.485 24.795 54.965 ;
        RECT 24.975 54.680 25.235 55.135 ;
        RECT 25.405 54.485 25.655 54.965 ;
        RECT 25.835 54.680 26.095 55.135 ;
        RECT 26.265 54.485 26.515 54.965 ;
        RECT 26.695 54.680 26.955 55.135 ;
        RECT 27.125 54.485 27.370 54.965 ;
        RECT 27.540 54.680 27.815 55.135 ;
        RECT 27.985 54.485 28.230 54.965 ;
        RECT 28.400 54.680 28.660 55.135 ;
        RECT 28.830 54.485 29.090 54.965 ;
        RECT 29.260 54.680 29.520 55.135 ;
        RECT 29.690 54.485 29.950 54.965 ;
        RECT 30.120 54.680 30.380 55.135 ;
        RECT 30.550 54.485 30.810 55.045 ;
        RECT 30.980 54.665 31.230 55.475 ;
        RECT 31.410 54.485 31.670 55.010 ;
        RECT 31.840 54.665 32.090 55.475 ;
        RECT 32.260 55.165 32.575 55.725 ;
        RECT 33.670 55.375 34.020 56.025 ;
        RECT 34.190 55.205 34.420 56.195 ;
        RECT 33.670 55.035 34.420 55.205 ;
        RECT 32.270 54.485 32.575 54.995 ;
        RECT 33.670 54.745 33.925 55.035 ;
        RECT 34.095 54.485 34.425 54.865 ;
        RECT 34.595 54.745 34.765 56.865 ;
        RECT 34.935 56.065 35.260 56.850 ;
        RECT 35.430 56.575 35.680 57.035 ;
        RECT 35.850 56.535 36.100 56.865 ;
        RECT 36.315 56.535 36.995 56.865 ;
        RECT 35.850 56.405 36.020 56.535 ;
        RECT 35.625 56.235 36.020 56.405 ;
        RECT 34.995 55.015 35.455 56.065 ;
        RECT 35.625 54.875 35.795 56.235 ;
        RECT 36.190 55.975 36.655 56.365 ;
        RECT 35.965 55.165 36.315 55.785 ;
        RECT 36.485 55.385 36.655 55.975 ;
        RECT 36.825 55.755 36.995 56.535 ;
        RECT 37.165 56.435 37.335 56.775 ;
        RECT 37.570 56.605 37.900 57.035 ;
        RECT 38.070 56.435 38.240 56.775 ;
        RECT 38.535 56.575 38.905 57.035 ;
        RECT 37.165 56.265 38.240 56.435 ;
        RECT 39.075 56.405 39.245 56.865 ;
        RECT 39.480 56.525 40.350 56.865 ;
        RECT 40.520 56.575 40.770 57.035 ;
        RECT 38.685 56.235 39.245 56.405 ;
        RECT 38.685 56.095 38.855 56.235 ;
        RECT 37.355 55.925 38.855 56.095 ;
        RECT 39.550 56.065 40.010 56.355 ;
        RECT 36.825 55.585 38.515 55.755 ;
        RECT 36.485 55.165 36.840 55.385 ;
        RECT 37.010 54.875 37.180 55.585 ;
        RECT 37.385 55.165 38.175 55.415 ;
        RECT 38.345 55.405 38.515 55.585 ;
        RECT 38.685 55.235 38.855 55.925 ;
        RECT 35.125 54.485 35.455 54.845 ;
        RECT 35.625 54.705 36.120 54.875 ;
        RECT 36.325 54.705 37.180 54.875 ;
        RECT 38.055 54.485 38.385 54.945 ;
        RECT 38.595 54.845 38.855 55.235 ;
        RECT 39.045 56.055 40.010 56.065 ;
        RECT 40.180 56.145 40.350 56.525 ;
        RECT 40.940 56.485 41.110 56.775 ;
        RECT 41.290 56.655 41.620 57.035 ;
        RECT 40.940 56.315 41.740 56.485 ;
        RECT 39.045 55.895 39.720 56.055 ;
        RECT 40.180 55.975 41.400 56.145 ;
        RECT 39.045 55.105 39.255 55.895 ;
        RECT 40.180 55.885 40.350 55.975 ;
        RECT 39.425 55.105 39.775 55.725 ;
        RECT 39.945 55.715 40.350 55.885 ;
        RECT 39.945 54.935 40.115 55.715 ;
        RECT 40.285 55.265 40.505 55.545 ;
        RECT 40.685 55.435 41.225 55.805 ;
        RECT 41.570 55.725 41.740 56.315 ;
        RECT 41.960 55.895 42.265 57.035 ;
        RECT 42.435 55.845 42.690 56.725 ;
        RECT 42.925 55.895 43.135 57.035 ;
        RECT 41.570 55.695 42.310 55.725 ;
        RECT 40.285 55.095 40.815 55.265 ;
        RECT 38.595 54.675 38.945 54.845 ;
        RECT 39.165 54.655 40.115 54.935 ;
        RECT 40.285 54.485 40.475 54.925 ;
        RECT 40.645 54.865 40.815 55.095 ;
        RECT 40.985 55.035 41.225 55.435 ;
        RECT 41.395 55.395 42.310 55.695 ;
        RECT 41.395 55.220 41.720 55.395 ;
        RECT 41.395 54.865 41.715 55.220 ;
        RECT 42.480 55.195 42.690 55.845 ;
        RECT 43.305 55.885 43.635 56.865 ;
        RECT 43.805 55.895 44.035 57.035 ;
        RECT 40.645 54.695 41.715 54.865 ;
        RECT 41.960 54.485 42.265 54.945 ;
        RECT 42.435 54.665 42.690 55.195 ;
        RECT 42.925 54.485 43.135 55.305 ;
        RECT 43.305 55.285 43.555 55.885 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 44.705 55.945 46.375 57.035 ;
        RECT 43.725 55.475 44.055 55.725 ;
        RECT 43.305 54.655 43.635 55.285 ;
        RECT 43.805 54.485 44.035 55.305 ;
        RECT 44.705 55.255 45.455 55.775 ;
        RECT 45.625 55.425 46.375 55.945 ;
        RECT 46.545 55.960 46.815 56.865 ;
        RECT 46.985 56.275 47.315 57.035 ;
        RECT 47.495 56.105 47.665 56.865 ;
        RECT 47.925 56.600 53.270 57.035 ;
        RECT 53.445 56.600 58.790 57.035 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 44.705 54.485 46.375 55.255 ;
        RECT 46.545 55.160 46.715 55.960 ;
        RECT 47.000 55.935 47.665 56.105 ;
        RECT 47.000 55.790 47.170 55.935 ;
        RECT 46.885 55.460 47.170 55.790 ;
        RECT 47.000 55.205 47.170 55.460 ;
        RECT 47.405 55.385 47.735 55.755 ;
        RECT 46.545 54.655 46.805 55.160 ;
        RECT 47.000 55.035 47.665 55.205 ;
        RECT 46.985 54.485 47.315 54.865 ;
        RECT 47.495 54.655 47.665 55.035 ;
        RECT 49.510 55.030 49.850 55.860 ;
        RECT 51.330 55.350 51.680 56.600 ;
        RECT 55.030 55.030 55.370 55.860 ;
        RECT 56.850 55.350 57.200 56.600 ;
        RECT 58.965 55.945 62.475 57.035 ;
        RECT 63.815 56.585 64.145 57.035 ;
        RECT 58.965 55.255 60.615 55.775 ;
        RECT 60.785 55.425 62.475 55.945 ;
        RECT 63.105 56.195 65.715 56.405 ;
        RECT 47.925 54.485 53.270 55.030 ;
        RECT 53.445 54.485 58.790 55.030 ;
        RECT 58.965 54.485 62.475 55.255 ;
        RECT 63.105 55.225 63.275 56.195 ;
        RECT 63.445 55.395 63.795 56.015 ;
        RECT 63.965 55.395 64.285 56.015 ;
        RECT 64.455 55.395 64.785 56.015 ;
        RECT 64.955 55.395 65.255 56.015 ;
        RECT 65.495 55.395 65.715 56.195 ;
        RECT 65.895 55.225 66.155 56.850 ;
        RECT 66.330 55.885 66.590 57.035 ;
        RECT 66.765 55.960 67.020 56.865 ;
        RECT 67.190 56.275 67.520 57.035 ;
        RECT 67.735 56.105 67.905 56.865 ;
        RECT 63.105 55.055 63.580 55.225 ;
        RECT 63.410 54.805 63.580 55.055 ;
        RECT 63.815 54.485 64.145 55.225 ;
        RECT 64.315 55.055 66.155 55.225 ;
        RECT 64.315 54.710 64.515 55.055 ;
        RECT 64.685 54.485 65.015 54.885 ;
        RECT 65.185 54.700 65.385 55.055 ;
        RECT 65.555 54.485 65.885 54.880 ;
        RECT 66.330 54.485 66.590 55.325 ;
        RECT 66.765 55.230 66.935 55.960 ;
        RECT 67.190 55.935 67.905 56.105 ;
        RECT 67.190 55.725 67.360 55.935 ;
        RECT 68.205 55.895 68.435 57.035 ;
        RECT 68.605 55.885 68.935 56.865 ;
        RECT 69.105 55.895 69.315 57.035 ;
        RECT 67.105 55.395 67.360 55.725 ;
        RECT 66.765 54.655 67.020 55.230 ;
        RECT 67.190 55.205 67.360 55.395 ;
        RECT 67.640 55.385 67.995 55.755 ;
        RECT 68.185 55.475 68.515 55.725 ;
        RECT 67.190 55.035 67.905 55.205 ;
        RECT 67.190 54.485 67.520 54.865 ;
        RECT 67.735 54.655 67.905 55.035 ;
        RECT 68.205 54.485 68.435 55.305 ;
        RECT 68.685 55.285 68.935 55.885 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 70.555 56.105 70.725 56.865 ;
        RECT 70.940 56.275 71.270 57.035 ;
        RECT 70.555 55.935 71.270 56.105 ;
        RECT 71.440 55.960 71.695 56.865 ;
        RECT 70.465 55.385 70.820 55.755 ;
        RECT 71.100 55.725 71.270 55.935 ;
        RECT 71.100 55.395 71.355 55.725 ;
        RECT 68.605 54.655 68.935 55.285 ;
        RECT 69.105 54.485 69.315 55.305 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 71.100 55.205 71.270 55.395 ;
        RECT 71.525 55.230 71.695 55.960 ;
        RECT 71.870 55.885 72.130 57.035 ;
        RECT 72.305 56.600 77.650 57.035 ;
        RECT 70.555 55.035 71.270 55.205 ;
        RECT 70.555 54.655 70.725 55.035 ;
        RECT 70.940 54.485 71.270 54.865 ;
        RECT 71.440 54.655 71.695 55.230 ;
        RECT 71.870 54.485 72.130 55.325 ;
        RECT 73.890 55.030 74.230 55.860 ;
        RECT 75.710 55.350 76.060 56.600 ;
        RECT 77.825 55.960 78.095 56.865 ;
        RECT 78.265 56.275 78.595 57.035 ;
        RECT 78.775 56.105 78.945 56.865 ;
        RECT 77.825 55.160 77.995 55.960 ;
        RECT 78.280 55.935 78.945 56.105 ;
        RECT 78.280 55.790 78.450 55.935 ;
        RECT 79.265 55.895 79.475 57.035 ;
        RECT 78.165 55.460 78.450 55.790 ;
        RECT 79.645 55.885 79.975 56.865 ;
        RECT 80.145 55.895 80.375 57.035 ;
        RECT 80.595 56.015 80.925 56.865 ;
        RECT 81.095 56.185 81.265 57.035 ;
        RECT 81.435 56.015 81.765 56.865 ;
        RECT 81.935 56.185 82.105 57.035 ;
        RECT 82.275 56.015 82.605 56.865 ;
        RECT 82.775 56.235 82.945 57.035 ;
        RECT 83.115 56.015 83.445 56.865 ;
        RECT 83.615 56.235 83.785 57.035 ;
        RECT 83.955 56.015 84.285 56.865 ;
        RECT 84.455 56.235 84.625 57.035 ;
        RECT 84.795 56.015 85.125 56.865 ;
        RECT 85.295 56.235 85.465 57.035 ;
        RECT 85.635 56.015 85.965 56.865 ;
        RECT 86.135 56.235 86.305 57.035 ;
        RECT 86.475 56.015 86.805 56.865 ;
        RECT 86.975 56.235 87.145 57.035 ;
        RECT 87.315 56.015 87.645 56.865 ;
        RECT 87.815 56.235 87.985 57.035 ;
        RECT 88.155 56.015 88.485 56.865 ;
        RECT 88.655 56.235 88.825 57.035 ;
        RECT 88.995 56.015 89.325 56.865 ;
        RECT 89.495 56.235 89.665 57.035 ;
        RECT 89.835 56.015 90.165 56.865 ;
        RECT 90.335 56.235 90.505 57.035 ;
        RECT 90.675 56.015 91.005 56.865 ;
        RECT 91.175 56.235 91.345 57.035 ;
        RECT 91.830 56.065 92.160 56.865 ;
        RECT 92.330 56.235 92.660 57.035 ;
        RECT 92.960 56.065 93.290 56.865 ;
        RECT 93.935 56.235 94.185 57.035 ;
        RECT 78.280 55.205 78.450 55.460 ;
        RECT 78.685 55.385 79.015 55.755 ;
        RECT 72.305 54.485 77.650 55.030 ;
        RECT 77.825 54.655 78.085 55.160 ;
        RECT 78.280 55.035 78.945 55.205 ;
        RECT 78.265 54.485 78.595 54.865 ;
        RECT 78.775 54.655 78.945 55.035 ;
        RECT 79.265 54.485 79.475 55.305 ;
        RECT 79.645 55.285 79.895 55.885 ;
        RECT 80.595 55.845 82.105 56.015 ;
        RECT 82.275 55.845 84.625 56.015 ;
        RECT 84.795 55.845 91.455 56.015 ;
        RECT 91.830 55.895 94.265 56.065 ;
        RECT 94.455 55.895 94.625 57.035 ;
        RECT 94.795 55.895 95.135 56.865 ;
        RECT 80.065 55.475 80.395 55.725 ;
        RECT 81.935 55.675 82.105 55.845 ;
        RECT 84.450 55.675 84.625 55.845 ;
        RECT 80.590 55.475 81.765 55.675 ;
        RECT 81.935 55.475 84.245 55.675 ;
        RECT 84.450 55.475 91.010 55.675 ;
        RECT 81.935 55.305 82.105 55.475 ;
        RECT 84.450 55.305 84.625 55.475 ;
        RECT 91.180 55.305 91.455 55.845 ;
        RECT 91.625 55.475 91.975 55.725 ;
        RECT 79.645 54.655 79.975 55.285 ;
        RECT 80.145 54.485 80.375 55.305 ;
        RECT 80.595 55.135 82.105 55.305 ;
        RECT 82.275 55.135 84.625 55.305 ;
        RECT 84.795 55.135 91.455 55.305 ;
        RECT 92.160 55.265 92.330 55.895 ;
        RECT 92.500 55.475 92.830 55.675 ;
        RECT 93.000 55.475 93.330 55.675 ;
        RECT 93.500 55.475 93.920 55.675 ;
        RECT 94.095 55.645 94.265 55.895 ;
        RECT 94.095 55.475 94.790 55.645 ;
        RECT 80.595 54.660 80.925 55.135 ;
        RECT 81.095 54.485 81.265 54.965 ;
        RECT 81.435 54.660 81.765 55.135 ;
        RECT 81.935 54.485 82.105 54.965 ;
        RECT 82.275 54.660 82.605 55.135 ;
        RECT 82.775 54.485 82.945 54.965 ;
        RECT 83.115 54.660 83.445 55.135 ;
        RECT 83.615 54.485 83.785 54.965 ;
        RECT 83.955 54.660 84.285 55.135 ;
        RECT 84.455 54.485 84.625 54.965 ;
        RECT 84.795 54.660 85.125 55.135 ;
        RECT 84.795 54.655 85.045 54.660 ;
        RECT 85.295 54.485 85.465 54.965 ;
        RECT 85.635 54.660 85.965 55.135 ;
        RECT 85.715 54.655 85.885 54.660 ;
        RECT 86.135 54.485 86.305 54.965 ;
        RECT 86.475 54.660 86.805 55.135 ;
        RECT 86.555 54.655 86.725 54.660 ;
        RECT 86.975 54.485 87.145 54.965 ;
        RECT 87.315 54.660 87.645 55.135 ;
        RECT 87.815 54.485 87.985 54.965 ;
        RECT 88.155 54.660 88.485 55.135 ;
        RECT 88.655 54.485 88.825 54.965 ;
        RECT 88.995 54.660 89.325 55.135 ;
        RECT 89.495 54.485 89.665 54.965 ;
        RECT 89.835 54.660 90.165 55.135 ;
        RECT 90.335 54.485 90.505 54.965 ;
        RECT 90.675 54.660 91.005 55.135 ;
        RECT 91.175 54.485 91.345 54.965 ;
        RECT 91.830 54.655 92.330 55.265 ;
        RECT 92.960 55.135 94.185 55.305 ;
        RECT 94.960 55.285 95.135 55.895 ;
        RECT 95.765 55.870 96.055 57.035 ;
        RECT 96.225 55.945 98.815 57.035 ;
        RECT 99.445 56.065 99.705 57.035 ;
        RECT 92.960 54.655 93.290 55.135 ;
        RECT 93.460 54.485 93.685 54.945 ;
        RECT 93.855 54.655 94.185 55.135 ;
        RECT 94.375 54.485 94.625 55.285 ;
        RECT 94.795 54.655 95.135 55.285 ;
        RECT 96.225 55.255 97.435 55.775 ;
        RECT 97.605 55.425 98.815 55.945 ;
        RECT 95.765 54.485 96.055 55.210 ;
        RECT 96.225 54.485 98.815 55.255 ;
        RECT 99.445 54.775 99.685 55.725 ;
        RECT 99.875 55.690 100.205 56.865 ;
        RECT 100.375 56.065 100.655 57.035 ;
        RECT 100.835 56.225 101.130 57.035 ;
        RECT 101.310 55.725 101.555 56.865 ;
        RECT 101.730 56.225 101.990 57.035 ;
        RECT 102.590 57.030 108.865 57.035 ;
        RECT 102.170 55.725 102.420 56.860 ;
        RECT 102.590 56.235 102.850 57.030 ;
        RECT 103.020 56.135 103.280 56.860 ;
        RECT 103.450 56.305 103.710 57.030 ;
        RECT 103.880 56.135 104.140 56.860 ;
        RECT 104.310 56.305 104.570 57.030 ;
        RECT 104.740 56.135 105.000 56.860 ;
        RECT 105.170 56.305 105.430 57.030 ;
        RECT 105.600 56.135 105.860 56.860 ;
        RECT 106.030 56.305 106.275 57.030 ;
        RECT 106.445 56.135 106.705 56.860 ;
        RECT 106.890 56.305 107.135 57.030 ;
        RECT 107.305 56.135 107.565 56.860 ;
        RECT 107.750 56.305 107.995 57.030 ;
        RECT 108.165 56.135 108.425 56.860 ;
        RECT 108.610 56.305 108.865 57.030 ;
        RECT 103.020 56.120 108.425 56.135 ;
        RECT 109.035 56.120 109.325 56.860 ;
        RECT 109.495 56.290 109.765 57.035 ;
        RECT 103.020 55.895 109.765 56.120 ;
        RECT 110.025 55.945 112.615 57.035 ;
        RECT 99.875 55.160 100.655 55.690 ;
        RECT 100.825 55.165 101.140 55.725 ;
        RECT 101.310 55.475 108.430 55.725 ;
        RECT 99.875 54.655 100.200 55.160 ;
        RECT 100.370 54.485 100.655 54.990 ;
        RECT 100.825 54.485 101.130 54.995 ;
        RECT 101.310 54.665 101.560 55.475 ;
        RECT 101.730 54.485 101.990 55.010 ;
        RECT 102.170 54.665 102.420 55.475 ;
        RECT 108.600 55.305 109.765 55.895 ;
        RECT 103.020 55.135 109.765 55.305 ;
        RECT 110.025 55.255 111.235 55.775 ;
        RECT 111.405 55.425 112.615 55.945 ;
        RECT 113.285 55.895 113.515 57.035 ;
        RECT 113.685 55.885 114.015 56.865 ;
        RECT 114.185 55.895 114.395 57.035 ;
        RECT 114.625 56.600 119.970 57.035 ;
        RECT 113.265 55.475 113.595 55.725 ;
        RECT 102.590 54.485 102.850 55.045 ;
        RECT 103.020 54.680 103.280 55.135 ;
        RECT 103.450 54.485 103.710 54.965 ;
        RECT 103.880 54.680 104.140 55.135 ;
        RECT 104.310 54.485 104.570 54.965 ;
        RECT 104.740 54.680 105.000 55.135 ;
        RECT 105.170 54.485 105.415 54.965 ;
        RECT 105.585 54.680 105.860 55.135 ;
        RECT 106.030 54.485 106.275 54.965 ;
        RECT 106.445 54.680 106.705 55.135 ;
        RECT 106.885 54.485 107.135 54.965 ;
        RECT 107.305 54.680 107.565 55.135 ;
        RECT 107.745 54.485 107.995 54.965 ;
        RECT 108.165 54.680 108.425 55.135 ;
        RECT 108.605 54.485 108.865 54.965 ;
        RECT 109.035 54.680 109.295 55.135 ;
        RECT 109.465 54.485 109.765 54.965 ;
        RECT 110.025 54.485 112.615 55.255 ;
        RECT 113.285 54.485 113.515 55.305 ;
        RECT 113.765 55.285 114.015 55.885 ;
        RECT 113.685 54.655 114.015 55.285 ;
        RECT 114.185 54.485 114.395 55.305 ;
        RECT 116.210 55.030 116.550 55.860 ;
        RECT 118.030 55.350 118.380 56.600 ;
        RECT 120.145 55.945 121.355 57.035 ;
        RECT 120.145 55.235 120.665 55.775 ;
        RECT 120.835 55.405 121.355 55.945 ;
        RECT 121.525 55.870 121.815 57.035 ;
        RECT 122.445 55.945 123.655 57.035 ;
        RECT 122.445 55.405 122.965 55.945 ;
        RECT 123.135 55.235 123.655 55.775 ;
        RECT 114.625 54.485 119.970 55.030 ;
        RECT 120.145 54.485 121.355 55.235 ;
        RECT 121.525 54.485 121.815 55.210 ;
        RECT 122.445 54.485 123.655 55.235 ;
        RECT 5.520 54.315 123.740 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.985 53.545 9.575 54.315 ;
        RECT 10.205 53.815 10.465 54.145 ;
        RECT 10.675 53.835 10.950 54.315 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 6.985 53.025 8.195 53.545 ;
        RECT 8.365 52.855 9.575 53.375 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 6.985 51.765 9.575 52.855 ;
        RECT 10.205 52.905 10.375 53.815 ;
        RECT 11.160 53.745 11.365 54.145 ;
        RECT 11.535 53.915 11.870 54.315 ;
        RECT 10.545 53.075 10.905 53.655 ;
        RECT 11.160 53.575 11.845 53.745 ;
        RECT 11.085 52.905 11.335 53.405 ;
        RECT 10.205 52.735 11.335 52.905 ;
        RECT 10.205 51.965 10.475 52.735 ;
        RECT 11.505 52.545 11.845 53.575 ;
        RECT 12.045 53.545 13.715 54.315 ;
        RECT 12.045 53.025 12.795 53.545 ;
        RECT 14.405 53.495 14.615 54.315 ;
        RECT 14.785 53.515 15.115 54.145 ;
        RECT 12.965 52.855 13.715 53.375 ;
        RECT 14.785 52.915 15.035 53.515 ;
        RECT 15.285 53.495 15.515 54.315 ;
        RECT 15.725 53.770 21.070 54.315 ;
        RECT 21.245 53.770 26.590 54.315 ;
        RECT 15.205 53.075 15.535 53.325 ;
        RECT 17.310 52.940 17.650 53.770 ;
        RECT 10.645 51.765 10.975 52.545 ;
        RECT 11.180 52.370 11.845 52.545 ;
        RECT 11.180 51.965 11.365 52.370 ;
        RECT 11.535 51.765 11.870 52.190 ;
        RECT 12.045 51.765 13.715 52.855 ;
        RECT 14.405 51.765 14.615 52.905 ;
        RECT 14.785 51.935 15.115 52.915 ;
        RECT 15.285 51.765 15.515 52.905 ;
        RECT 19.130 52.200 19.480 53.450 ;
        RECT 22.830 52.940 23.170 53.770 ;
        RECT 26.765 53.545 29.355 54.315 ;
        RECT 24.650 52.200 25.000 53.450 ;
        RECT 26.765 53.025 27.975 53.545 ;
        RECT 29.585 53.495 29.795 54.315 ;
        RECT 29.965 53.515 30.295 54.145 ;
        RECT 28.145 52.855 29.355 53.375 ;
        RECT 29.965 52.915 30.215 53.515 ;
        RECT 30.465 53.495 30.695 54.315 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 31.825 53.770 37.170 54.315 ;
        RECT 30.385 53.075 30.715 53.325 ;
        RECT 33.410 52.940 33.750 53.770 ;
        RECT 15.725 51.765 21.070 52.200 ;
        RECT 21.245 51.765 26.590 52.200 ;
        RECT 26.765 51.765 29.355 52.855 ;
        RECT 29.585 51.765 29.795 52.905 ;
        RECT 29.965 51.935 30.295 52.915 ;
        RECT 30.465 51.765 30.695 52.905 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 35.230 52.200 35.580 53.450 ;
        RECT 37.805 53.075 38.045 54.025 ;
        RECT 38.235 53.640 38.560 54.145 ;
        RECT 38.730 53.810 39.015 54.315 ;
        RECT 39.275 53.835 39.575 54.315 ;
        RECT 39.745 53.665 40.005 54.120 ;
        RECT 40.175 53.835 40.435 54.315 ;
        RECT 40.615 53.665 40.875 54.120 ;
        RECT 41.045 53.835 41.295 54.315 ;
        RECT 41.475 53.665 41.735 54.120 ;
        RECT 41.905 53.835 42.155 54.315 ;
        RECT 42.335 53.665 42.595 54.120 ;
        RECT 42.765 53.835 43.010 54.315 ;
        RECT 43.180 53.665 43.455 54.120 ;
        RECT 43.625 53.835 43.870 54.315 ;
        RECT 44.040 53.665 44.300 54.120 ;
        RECT 44.470 53.835 44.730 54.315 ;
        RECT 44.900 53.665 45.160 54.120 ;
        RECT 45.330 53.835 45.590 54.315 ;
        RECT 45.760 53.665 46.020 54.120 ;
        RECT 46.190 53.755 46.450 54.315 ;
        RECT 38.235 53.110 39.015 53.640 ;
        RECT 39.275 53.635 46.020 53.665 ;
        RECT 39.245 53.495 46.020 53.635 ;
        RECT 39.245 53.465 40.440 53.495 ;
        RECT 31.825 51.765 37.170 52.200 ;
        RECT 37.805 51.765 38.065 52.735 ;
        RECT 38.235 51.935 38.565 53.110 ;
        RECT 39.275 52.905 40.440 53.465 ;
        RECT 46.620 53.325 46.870 54.135 ;
        RECT 47.050 53.790 47.310 54.315 ;
        RECT 47.480 53.325 47.730 54.135 ;
        RECT 47.910 53.805 48.215 54.315 ;
        RECT 40.610 53.075 47.730 53.325 ;
        RECT 47.900 53.075 48.215 53.635 ;
        RECT 49.050 53.535 49.550 54.145 ;
        RECT 48.845 53.075 49.195 53.325 ;
        RECT 38.735 51.765 39.015 52.735 ;
        RECT 39.275 52.680 46.020 52.905 ;
        RECT 39.275 51.765 39.545 52.510 ;
        RECT 39.715 51.940 40.005 52.680 ;
        RECT 40.615 52.665 46.020 52.680 ;
        RECT 40.175 51.770 40.430 52.495 ;
        RECT 40.615 51.940 40.875 52.665 ;
        RECT 41.045 51.770 41.290 52.495 ;
        RECT 41.475 51.940 41.735 52.665 ;
        RECT 41.905 51.770 42.150 52.495 ;
        RECT 42.335 51.940 42.595 52.665 ;
        RECT 42.765 51.770 43.010 52.495 ;
        RECT 43.180 51.940 43.440 52.665 ;
        RECT 43.610 51.770 43.870 52.495 ;
        RECT 44.040 51.940 44.300 52.665 ;
        RECT 44.470 51.770 44.730 52.495 ;
        RECT 44.900 51.940 45.160 52.665 ;
        RECT 45.330 51.770 45.590 52.495 ;
        RECT 45.760 51.940 46.020 52.665 ;
        RECT 46.190 51.770 46.450 52.565 ;
        RECT 46.620 51.940 46.870 53.075 ;
        RECT 40.175 51.765 46.450 51.770 ;
        RECT 47.050 51.765 47.310 52.575 ;
        RECT 47.485 51.935 47.730 53.075 ;
        RECT 49.380 52.905 49.550 53.535 ;
        RECT 50.180 53.665 50.510 54.145 ;
        RECT 50.680 53.855 50.905 54.315 ;
        RECT 51.075 53.665 51.405 54.145 ;
        RECT 50.180 53.495 51.405 53.665 ;
        RECT 51.595 53.515 51.845 54.315 ;
        RECT 52.015 53.515 52.355 54.145 ;
        RECT 49.720 53.125 50.050 53.325 ;
        RECT 50.220 53.125 50.550 53.325 ;
        RECT 50.720 53.125 51.140 53.325 ;
        RECT 51.315 53.155 52.010 53.325 ;
        RECT 51.315 52.905 51.485 53.155 ;
        RECT 52.180 52.905 52.355 53.515 ;
        RECT 52.525 53.545 56.035 54.315 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 57.585 53.545 61.095 54.315 ;
        RECT 61.265 53.815 61.525 54.145 ;
        RECT 61.835 53.935 62.165 54.315 ;
        RECT 62.345 53.975 63.825 54.145 ;
        RECT 52.525 53.025 54.175 53.545 ;
        RECT 49.050 52.735 51.485 52.905 ;
        RECT 47.910 51.765 48.205 52.575 ;
        RECT 49.050 51.935 49.380 52.735 ;
        RECT 49.550 51.765 49.880 52.565 ;
        RECT 50.180 51.935 50.510 52.735 ;
        RECT 51.155 51.765 51.405 52.565 ;
        RECT 51.675 51.765 51.845 52.905 ;
        RECT 52.015 51.935 52.355 52.905 ;
        RECT 54.345 52.855 56.035 53.375 ;
        RECT 57.585 53.025 59.235 53.545 ;
        RECT 52.525 51.765 56.035 52.855 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 59.405 52.855 61.095 53.375 ;
        RECT 57.585 51.765 61.095 52.855 ;
        RECT 61.265 53.115 61.435 53.815 ;
        RECT 62.345 53.645 62.745 53.975 ;
        RECT 61.785 53.455 61.995 53.635 ;
        RECT 61.785 53.285 62.405 53.455 ;
        RECT 62.575 53.165 62.745 53.645 ;
        RECT 62.935 53.475 63.485 53.805 ;
        RECT 61.265 52.945 62.395 53.115 ;
        RECT 62.575 52.995 63.145 53.165 ;
        RECT 61.265 52.265 61.435 52.945 ;
        RECT 62.225 52.825 62.395 52.945 ;
        RECT 61.605 52.445 61.955 52.775 ;
        RECT 62.225 52.655 62.805 52.825 ;
        RECT 62.975 52.485 63.145 52.995 ;
        RECT 62.405 52.315 63.145 52.485 ;
        RECT 63.315 52.485 63.485 53.475 ;
        RECT 63.655 53.075 63.825 53.975 ;
        RECT 64.075 53.405 64.260 53.985 ;
        RECT 64.530 53.405 64.725 53.980 ;
        RECT 64.935 53.935 65.265 54.315 ;
        RECT 64.075 53.075 64.305 53.405 ;
        RECT 64.530 53.075 64.785 53.405 ;
        RECT 64.075 52.765 64.260 53.075 ;
        RECT 64.530 52.765 64.725 53.075 ;
        RECT 65.095 52.485 65.265 53.405 ;
        RECT 63.315 52.315 65.265 52.485 ;
        RECT 61.265 51.935 61.525 52.265 ;
        RECT 61.835 51.765 62.165 52.145 ;
        RECT 62.405 51.935 62.595 52.315 ;
        RECT 62.845 51.765 63.175 52.145 ;
        RECT 63.385 51.935 63.555 52.315 ;
        RECT 63.750 51.765 64.080 52.145 ;
        RECT 64.340 51.935 64.510 52.315 ;
        RECT 64.935 51.765 65.265 52.145 ;
        RECT 65.435 51.935 65.695 54.145 ;
        RECT 65.875 53.955 67.945 54.145 ;
        RECT 68.175 53.955 68.505 54.315 ;
        RECT 69.035 53.955 69.365 54.315 ;
        RECT 69.895 53.955 70.225 54.315 ;
        RECT 66.825 53.935 67.945 53.955 ;
        RECT 65.865 52.430 66.155 53.405 ;
        RECT 66.325 52.860 66.655 53.730 ;
        RECT 66.825 53.510 67.015 53.935 ;
        RECT 69.535 53.765 69.725 53.885 ;
        RECT 67.185 53.555 69.725 53.765 ;
        RECT 70.555 53.765 70.725 54.145 ;
        RECT 70.940 53.935 71.270 54.315 ;
        RECT 69.895 53.325 70.235 53.635 ;
        RECT 70.555 53.595 71.270 53.765 ;
        RECT 66.825 53.035 67.685 53.325 ;
        RECT 68.145 53.045 69.115 53.325 ;
        RECT 69.285 53.155 70.235 53.325 ;
        RECT 69.340 53.105 70.235 53.155 ;
        RECT 70.465 53.045 70.820 53.415 ;
        RECT 71.100 53.405 71.270 53.595 ;
        RECT 71.440 53.570 71.695 54.145 ;
        RECT 71.100 53.075 71.355 53.405 ;
        RECT 66.325 52.690 68.935 52.860 ;
        RECT 65.895 51.765 66.155 52.225 ;
        RECT 66.325 51.935 66.585 52.690 ;
        RECT 66.755 51.765 67.085 52.485 ;
        RECT 67.255 51.935 67.445 52.690 ;
        RECT 67.615 51.765 67.945 52.485 ;
        RECT 68.175 52.105 68.435 52.300 ;
        RECT 68.605 52.275 68.935 52.690 ;
        RECT 69.105 52.705 70.225 52.875 ;
        RECT 71.100 52.865 71.270 53.075 ;
        RECT 69.105 52.105 69.295 52.705 ;
        RECT 68.175 51.935 69.295 52.105 ;
        RECT 69.465 51.765 69.795 52.535 ;
        RECT 69.965 51.935 70.225 52.705 ;
        RECT 70.555 52.695 71.270 52.865 ;
        RECT 71.525 52.840 71.695 53.570 ;
        RECT 71.870 53.475 72.130 54.315 ;
        RECT 72.305 53.565 73.515 54.315 ;
        RECT 73.690 53.765 73.945 54.055 ;
        RECT 74.115 53.935 74.445 54.315 ;
        RECT 73.690 53.595 74.440 53.765 ;
        RECT 72.305 53.025 72.825 53.565 ;
        RECT 70.555 51.935 70.725 52.695 ;
        RECT 70.940 51.765 71.270 52.525 ;
        RECT 71.440 51.935 71.695 52.840 ;
        RECT 71.870 51.765 72.130 52.915 ;
        RECT 72.995 52.855 73.515 53.395 ;
        RECT 72.305 51.765 73.515 52.855 ;
        RECT 73.690 52.775 74.040 53.425 ;
        RECT 74.210 52.605 74.440 53.595 ;
        RECT 73.690 52.435 74.440 52.605 ;
        RECT 73.690 51.935 73.945 52.435 ;
        RECT 74.115 51.765 74.445 52.265 ;
        RECT 74.615 51.935 74.785 54.055 ;
        RECT 75.145 53.955 75.475 54.315 ;
        RECT 75.645 53.925 76.140 54.095 ;
        RECT 76.345 53.925 77.200 54.095 ;
        RECT 75.015 52.735 75.475 53.785 ;
        RECT 74.955 51.950 75.280 52.735 ;
        RECT 75.645 52.565 75.815 53.925 ;
        RECT 75.985 53.015 76.335 53.635 ;
        RECT 76.505 53.415 76.860 53.635 ;
        RECT 76.505 52.825 76.675 53.415 ;
        RECT 77.030 53.215 77.200 53.925 ;
        RECT 78.075 53.855 78.405 54.315 ;
        RECT 78.615 53.955 78.965 54.125 ;
        RECT 77.405 53.385 78.195 53.635 ;
        RECT 78.615 53.565 78.875 53.955 ;
        RECT 79.185 53.865 80.135 54.145 ;
        RECT 80.305 53.875 80.495 54.315 ;
        RECT 80.665 53.935 81.735 54.105 ;
        RECT 78.365 53.215 78.535 53.395 ;
        RECT 75.645 52.395 76.040 52.565 ;
        RECT 76.210 52.435 76.675 52.825 ;
        RECT 76.845 53.045 78.535 53.215 ;
        RECT 75.870 52.265 76.040 52.395 ;
        RECT 76.845 52.265 77.015 53.045 ;
        RECT 78.705 52.875 78.875 53.565 ;
        RECT 77.375 52.705 78.875 52.875 ;
        RECT 79.065 52.905 79.275 53.695 ;
        RECT 79.445 53.075 79.795 53.695 ;
        RECT 79.965 53.085 80.135 53.865 ;
        RECT 80.665 53.705 80.835 53.935 ;
        RECT 80.305 53.535 80.835 53.705 ;
        RECT 80.305 53.255 80.525 53.535 ;
        RECT 81.005 53.365 81.245 53.765 ;
        RECT 79.965 52.915 80.370 53.085 ;
        RECT 80.705 52.995 81.245 53.365 ;
        RECT 81.415 53.580 81.735 53.935 ;
        RECT 81.980 53.855 82.285 54.315 ;
        RECT 82.455 53.605 82.710 54.135 ;
        RECT 81.415 53.405 81.740 53.580 ;
        RECT 81.415 53.105 82.330 53.405 ;
        RECT 81.590 53.075 82.330 53.105 ;
        RECT 79.065 52.745 79.740 52.905 ;
        RECT 80.200 52.825 80.370 52.915 ;
        RECT 79.065 52.735 80.030 52.745 ;
        RECT 78.705 52.565 78.875 52.705 ;
        RECT 75.450 51.765 75.700 52.225 ;
        RECT 75.870 51.935 76.120 52.265 ;
        RECT 76.335 51.935 77.015 52.265 ;
        RECT 77.185 52.365 78.260 52.535 ;
        RECT 78.705 52.395 79.265 52.565 ;
        RECT 79.570 52.445 80.030 52.735 ;
        RECT 80.200 52.655 81.420 52.825 ;
        RECT 77.185 52.025 77.355 52.365 ;
        RECT 77.590 51.765 77.920 52.195 ;
        RECT 78.090 52.025 78.260 52.365 ;
        RECT 78.555 51.765 78.925 52.225 ;
        RECT 79.095 51.935 79.265 52.395 ;
        RECT 80.200 52.275 80.370 52.655 ;
        RECT 81.590 52.485 81.760 53.075 ;
        RECT 82.500 52.955 82.710 53.605 ;
        RECT 82.885 53.590 83.175 54.315 ;
        RECT 83.435 53.835 83.735 54.315 ;
        RECT 83.905 53.665 84.165 54.120 ;
        RECT 84.335 53.835 84.595 54.315 ;
        RECT 84.775 53.665 85.035 54.120 ;
        RECT 85.205 53.835 85.455 54.315 ;
        RECT 85.635 53.665 85.895 54.120 ;
        RECT 86.065 53.835 86.315 54.315 ;
        RECT 86.495 53.665 86.755 54.120 ;
        RECT 86.925 53.835 87.170 54.315 ;
        RECT 87.340 53.665 87.615 54.120 ;
        RECT 87.785 53.835 88.030 54.315 ;
        RECT 88.200 53.665 88.460 54.120 ;
        RECT 88.630 53.835 88.890 54.315 ;
        RECT 89.060 53.665 89.320 54.120 ;
        RECT 89.490 53.835 89.750 54.315 ;
        RECT 89.920 53.665 90.180 54.120 ;
        RECT 90.350 53.755 90.610 54.315 ;
        RECT 83.435 53.635 90.180 53.665 ;
        RECT 83.405 53.495 90.180 53.635 ;
        RECT 83.405 53.465 84.600 53.495 ;
        RECT 79.500 51.935 80.370 52.275 ;
        RECT 80.960 52.315 81.760 52.485 ;
        RECT 80.540 51.765 80.790 52.225 ;
        RECT 80.960 52.025 81.130 52.315 ;
        RECT 81.310 51.765 81.640 52.145 ;
        RECT 81.980 51.765 82.285 52.905 ;
        RECT 82.455 52.075 82.710 52.955 ;
        RECT 82.885 51.765 83.175 52.930 ;
        RECT 83.435 52.905 84.600 53.465 ;
        RECT 90.780 53.325 91.030 54.135 ;
        RECT 91.210 53.790 91.470 54.315 ;
        RECT 91.640 53.325 91.890 54.135 ;
        RECT 92.070 53.805 92.375 54.315 ;
        RECT 92.545 53.770 97.890 54.315 ;
        RECT 84.770 53.075 91.890 53.325 ;
        RECT 92.060 53.075 92.375 53.635 ;
        RECT 83.435 52.680 90.180 52.905 ;
        RECT 83.435 51.765 83.705 52.510 ;
        RECT 83.875 51.940 84.165 52.680 ;
        RECT 84.775 52.665 90.180 52.680 ;
        RECT 84.335 51.770 84.590 52.495 ;
        RECT 84.775 51.940 85.035 52.665 ;
        RECT 85.205 51.770 85.450 52.495 ;
        RECT 85.635 51.940 85.895 52.665 ;
        RECT 86.065 51.770 86.310 52.495 ;
        RECT 86.495 51.940 86.755 52.665 ;
        RECT 86.925 51.770 87.170 52.495 ;
        RECT 87.340 51.940 87.600 52.665 ;
        RECT 87.770 51.770 88.030 52.495 ;
        RECT 88.200 51.940 88.460 52.665 ;
        RECT 88.630 51.770 88.890 52.495 ;
        RECT 89.060 51.940 89.320 52.665 ;
        RECT 89.490 51.770 89.750 52.495 ;
        RECT 89.920 51.940 90.180 52.665 ;
        RECT 90.350 51.770 90.610 52.565 ;
        RECT 90.780 51.940 91.030 53.075 ;
        RECT 84.335 51.765 90.610 51.770 ;
        RECT 91.210 51.765 91.470 52.575 ;
        RECT 91.645 51.935 91.890 53.075 ;
        RECT 94.130 52.940 94.470 53.770 ;
        RECT 98.985 53.515 99.325 54.145 ;
        RECT 99.495 53.515 99.745 54.315 ;
        RECT 99.935 53.665 100.265 54.145 ;
        RECT 100.435 53.855 100.660 54.315 ;
        RECT 100.830 53.665 101.160 54.145 ;
        RECT 92.070 51.765 92.365 52.575 ;
        RECT 95.950 52.200 96.300 53.450 ;
        RECT 98.985 52.905 99.160 53.515 ;
        RECT 99.935 53.495 101.160 53.665 ;
        RECT 101.790 53.535 102.290 54.145 ;
        RECT 102.665 53.770 108.010 54.315 ;
        RECT 99.330 53.155 100.025 53.325 ;
        RECT 99.855 52.905 100.025 53.155 ;
        RECT 100.200 53.125 100.620 53.325 ;
        RECT 100.790 53.125 101.120 53.325 ;
        RECT 101.290 53.125 101.620 53.325 ;
        RECT 101.790 52.905 101.960 53.535 ;
        RECT 102.145 53.075 102.495 53.325 ;
        RECT 104.250 52.940 104.590 53.770 ;
        RECT 108.645 53.590 108.935 54.315 ;
        RECT 109.105 53.770 114.450 54.315 ;
        RECT 114.625 53.770 119.970 54.315 ;
        RECT 92.545 51.765 97.890 52.200 ;
        RECT 98.985 51.935 99.325 52.905 ;
        RECT 99.495 51.765 99.665 52.905 ;
        RECT 99.855 52.735 102.290 52.905 ;
        RECT 99.935 51.765 100.185 52.565 ;
        RECT 100.830 51.935 101.160 52.735 ;
        RECT 101.460 51.765 101.790 52.565 ;
        RECT 101.960 51.935 102.290 52.735 ;
        RECT 106.070 52.200 106.420 53.450 ;
        RECT 110.690 52.940 111.030 53.770 ;
        RECT 102.665 51.765 108.010 52.200 ;
        RECT 108.645 51.765 108.935 52.930 ;
        RECT 112.510 52.200 112.860 53.450 ;
        RECT 116.210 52.940 116.550 53.770 ;
        RECT 120.145 53.545 121.815 54.315 ;
        RECT 122.445 53.565 123.655 54.315 ;
        RECT 118.030 52.200 118.380 53.450 ;
        RECT 120.145 53.025 120.895 53.545 ;
        RECT 121.065 52.855 121.815 53.375 ;
        RECT 109.105 51.765 114.450 52.200 ;
        RECT 114.625 51.765 119.970 52.200 ;
        RECT 120.145 51.765 121.815 52.855 ;
        RECT 122.445 52.855 122.965 53.395 ;
        RECT 123.135 53.025 123.655 53.565 ;
        RECT 122.445 51.765 123.655 52.855 ;
        RECT 5.520 51.595 123.740 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 6.985 51.160 12.330 51.595 ;
        RECT 12.505 51.160 17.850 51.595 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 8.570 49.590 8.910 50.420 ;
        RECT 10.390 49.910 10.740 51.160 ;
        RECT 14.090 49.590 14.430 50.420 ;
        RECT 15.910 49.910 16.260 51.160 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 18.945 50.505 22.455 51.595 ;
        RECT 18.945 49.815 20.595 50.335 ;
        RECT 20.765 49.985 22.455 50.505 ;
        RECT 23.085 50.455 23.425 51.425 ;
        RECT 23.595 50.455 23.765 51.595 ;
        RECT 24.035 50.795 24.285 51.595 ;
        RECT 24.930 50.625 25.260 51.425 ;
        RECT 25.560 50.795 25.890 51.595 ;
        RECT 26.060 50.625 26.390 51.425 ;
        RECT 23.955 50.455 26.390 50.625 ;
        RECT 26.765 50.455 27.105 51.425 ;
        RECT 27.275 50.455 27.445 51.595 ;
        RECT 27.715 50.795 27.965 51.595 ;
        RECT 28.610 50.625 28.940 51.425 ;
        RECT 29.240 50.795 29.570 51.595 ;
        RECT 29.740 50.625 30.070 51.425 ;
        RECT 30.445 51.160 35.790 51.595 ;
        RECT 35.965 51.160 41.310 51.595 ;
        RECT 27.635 50.455 30.070 50.625 ;
        RECT 23.085 49.845 23.260 50.455 ;
        RECT 23.955 50.205 24.125 50.455 ;
        RECT 23.430 50.035 24.125 50.205 ;
        RECT 24.300 50.035 24.720 50.235 ;
        RECT 24.890 50.035 25.220 50.235 ;
        RECT 25.390 50.035 25.720 50.235 ;
        RECT 6.985 49.045 12.330 49.590 ;
        RECT 12.505 49.045 17.850 49.590 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 18.945 49.045 22.455 49.815 ;
        RECT 23.085 49.215 23.425 49.845 ;
        RECT 23.595 49.045 23.845 49.845 ;
        RECT 24.035 49.695 25.260 49.865 ;
        RECT 24.035 49.215 24.365 49.695 ;
        RECT 24.535 49.045 24.760 49.505 ;
        RECT 24.930 49.215 25.260 49.695 ;
        RECT 25.890 49.825 26.060 50.455 ;
        RECT 26.245 50.035 26.595 50.285 ;
        RECT 26.765 49.845 26.940 50.455 ;
        RECT 27.635 50.205 27.805 50.455 ;
        RECT 27.110 50.035 27.805 50.205 ;
        RECT 27.980 50.035 28.400 50.235 ;
        RECT 28.570 50.035 28.900 50.235 ;
        RECT 29.070 50.035 29.400 50.235 ;
        RECT 25.890 49.215 26.390 49.825 ;
        RECT 26.765 49.215 27.105 49.845 ;
        RECT 27.275 49.045 27.525 49.845 ;
        RECT 27.715 49.695 28.940 49.865 ;
        RECT 27.715 49.215 28.045 49.695 ;
        RECT 28.215 49.045 28.440 49.505 ;
        RECT 28.610 49.215 28.940 49.695 ;
        RECT 29.570 49.825 29.740 50.455 ;
        RECT 29.925 50.035 30.275 50.285 ;
        RECT 29.570 49.215 30.070 49.825 ;
        RECT 32.030 49.590 32.370 50.420 ;
        RECT 33.850 49.910 34.200 51.160 ;
        RECT 37.550 49.590 37.890 50.420 ;
        RECT 39.370 49.910 39.720 51.160 ;
        RECT 41.485 50.505 44.075 51.595 ;
        RECT 41.485 49.815 42.695 50.335 ;
        RECT 42.865 49.985 44.075 50.505 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 45.315 50.445 45.645 51.595 ;
        RECT 45.815 50.575 45.985 51.425 ;
        RECT 46.155 50.795 46.485 51.595 ;
        RECT 46.655 50.575 46.825 51.425 ;
        RECT 47.005 50.795 47.245 51.595 ;
        RECT 47.415 50.615 47.745 51.425 ;
        RECT 45.815 50.405 46.825 50.575 ;
        RECT 47.030 50.445 47.745 50.615 ;
        RECT 47.925 50.505 49.595 51.595 ;
        RECT 45.815 49.895 46.310 50.405 ;
        RECT 47.030 50.205 47.200 50.445 ;
        RECT 46.700 50.035 47.200 50.205 ;
        RECT 47.370 50.035 47.750 50.275 ;
        RECT 45.815 49.865 46.315 49.895 ;
        RECT 47.030 49.865 47.200 50.035 ;
        RECT 30.445 49.045 35.790 49.590 ;
        RECT 35.965 49.045 41.310 49.590 ;
        RECT 41.485 49.045 44.075 49.815 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 45.315 49.045 45.645 49.845 ;
        RECT 45.815 49.695 46.825 49.865 ;
        RECT 47.030 49.695 47.665 49.865 ;
        RECT 45.815 49.215 45.985 49.695 ;
        RECT 46.155 49.045 46.485 49.525 ;
        RECT 46.655 49.215 46.825 49.695 ;
        RECT 47.075 49.045 47.315 49.525 ;
        RECT 47.495 49.215 47.665 49.695 ;
        RECT 47.925 49.815 48.675 50.335 ;
        RECT 48.845 49.985 49.595 50.505 ;
        RECT 49.970 50.625 50.300 51.425 ;
        RECT 50.470 50.795 50.800 51.595 ;
        RECT 51.100 50.625 51.430 51.425 ;
        RECT 52.075 50.795 52.325 51.595 ;
        RECT 49.970 50.455 52.405 50.625 ;
        RECT 52.595 50.455 52.765 51.595 ;
        RECT 52.935 50.455 53.275 51.425 ;
        RECT 53.650 50.625 53.980 51.425 ;
        RECT 54.150 50.795 54.480 51.595 ;
        RECT 54.780 50.625 55.110 51.425 ;
        RECT 55.755 50.795 56.005 51.595 ;
        RECT 53.650 50.455 56.085 50.625 ;
        RECT 56.275 50.455 56.445 51.595 ;
        RECT 56.615 50.455 56.955 51.425 ;
        RECT 57.125 51.160 62.470 51.595 ;
        RECT 49.765 50.035 50.115 50.285 ;
        RECT 50.300 49.825 50.470 50.455 ;
        RECT 50.640 50.035 50.970 50.235 ;
        RECT 51.140 50.035 51.470 50.235 ;
        RECT 51.640 50.035 52.060 50.235 ;
        RECT 52.235 50.205 52.405 50.455 ;
        RECT 53.045 50.405 53.275 50.455 ;
        RECT 52.235 50.035 52.930 50.205 ;
        RECT 47.925 49.045 49.595 49.815 ;
        RECT 49.970 49.215 50.470 49.825 ;
        RECT 51.100 49.695 52.325 49.865 ;
        RECT 53.100 49.845 53.275 50.405 ;
        RECT 53.445 50.035 53.795 50.285 ;
        RECT 51.100 49.215 51.430 49.695 ;
        RECT 51.600 49.045 51.825 49.505 ;
        RECT 51.995 49.215 52.325 49.695 ;
        RECT 52.515 49.045 52.765 49.845 ;
        RECT 52.935 49.215 53.275 49.845 ;
        RECT 53.980 49.825 54.150 50.455 ;
        RECT 54.320 50.035 54.650 50.235 ;
        RECT 54.820 50.035 55.150 50.235 ;
        RECT 55.320 50.035 55.740 50.235 ;
        RECT 55.915 50.205 56.085 50.455 ;
        RECT 55.915 50.035 56.610 50.205 ;
        RECT 53.650 49.215 54.150 49.825 ;
        RECT 54.780 49.695 56.005 49.865 ;
        RECT 56.780 49.845 56.955 50.455 ;
        RECT 54.780 49.215 55.110 49.695 ;
        RECT 55.280 49.045 55.505 49.505 ;
        RECT 55.675 49.215 56.005 49.695 ;
        RECT 56.195 49.045 56.445 49.845 ;
        RECT 56.615 49.215 56.955 49.845 ;
        RECT 58.710 49.590 59.050 50.420 ;
        RECT 60.530 49.910 60.880 51.160 ;
        RECT 62.645 50.505 64.315 51.595 ;
        RECT 65.655 51.145 65.985 51.595 ;
        RECT 62.645 49.815 63.395 50.335 ;
        RECT 63.565 49.985 64.315 50.505 ;
        RECT 64.945 50.755 67.555 50.965 ;
        RECT 57.125 49.045 62.470 49.590 ;
        RECT 62.645 49.045 64.315 49.815 ;
        RECT 64.945 49.785 65.115 50.755 ;
        RECT 65.285 49.955 65.635 50.575 ;
        RECT 65.805 49.955 66.125 50.575 ;
        RECT 66.295 49.955 66.625 50.575 ;
        RECT 66.795 49.955 67.095 50.575 ;
        RECT 67.335 49.955 67.555 50.755 ;
        RECT 67.735 49.785 67.995 51.410 ;
        RECT 68.170 50.445 68.430 51.595 ;
        RECT 68.605 50.520 68.860 51.425 ;
        RECT 69.030 50.835 69.360 51.595 ;
        RECT 69.575 50.665 69.745 51.425 ;
        RECT 64.945 49.615 65.420 49.785 ;
        RECT 65.250 49.365 65.420 49.615 ;
        RECT 65.655 49.045 65.985 49.785 ;
        RECT 66.155 49.615 67.995 49.785 ;
        RECT 66.155 49.270 66.355 49.615 ;
        RECT 66.525 49.045 66.855 49.445 ;
        RECT 67.025 49.260 67.225 49.615 ;
        RECT 67.395 49.045 67.725 49.440 ;
        RECT 68.170 49.045 68.430 49.885 ;
        RECT 68.605 49.790 68.775 50.520 ;
        RECT 69.030 50.495 69.745 50.665 ;
        RECT 69.030 50.285 69.200 50.495 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 68.945 49.955 69.200 50.285 ;
        RECT 68.605 49.215 68.860 49.790 ;
        RECT 69.030 49.765 69.200 49.955 ;
        RECT 69.480 49.945 69.835 50.315 ;
        RECT 70.465 49.785 70.725 51.410 ;
        RECT 72.475 51.145 72.805 51.595 ;
        RECT 70.905 50.755 73.515 50.965 ;
        RECT 70.905 49.955 71.125 50.755 ;
        RECT 71.365 49.955 71.665 50.575 ;
        RECT 71.835 49.955 72.165 50.575 ;
        RECT 72.335 49.955 72.655 50.575 ;
        RECT 72.825 49.955 73.175 50.575 ;
        RECT 73.345 49.785 73.515 50.755 ;
        RECT 73.775 50.665 73.945 51.425 ;
        RECT 74.160 50.835 74.490 51.595 ;
        RECT 73.775 50.495 74.490 50.665 ;
        RECT 74.660 50.520 74.915 51.425 ;
        RECT 73.685 49.945 74.040 50.315 ;
        RECT 74.320 50.285 74.490 50.495 ;
        RECT 74.320 49.955 74.575 50.285 ;
        RECT 69.030 49.595 69.745 49.765 ;
        RECT 69.030 49.045 69.360 49.425 ;
        RECT 69.575 49.215 69.745 49.595 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 70.465 49.615 72.305 49.785 ;
        RECT 70.735 49.045 71.065 49.440 ;
        RECT 71.235 49.260 71.435 49.615 ;
        RECT 71.605 49.045 71.935 49.445 ;
        RECT 72.105 49.270 72.305 49.615 ;
        RECT 72.475 49.045 72.805 49.785 ;
        RECT 73.040 49.615 73.515 49.785 ;
        RECT 74.320 49.765 74.490 49.955 ;
        RECT 74.745 49.790 74.915 50.520 ;
        RECT 75.090 50.445 75.350 51.595 ;
        RECT 75.525 50.505 76.735 51.595 ;
        RECT 73.040 49.365 73.210 49.615 ;
        RECT 73.775 49.595 74.490 49.765 ;
        RECT 73.775 49.215 73.945 49.595 ;
        RECT 74.160 49.045 74.490 49.425 ;
        RECT 74.660 49.215 74.915 49.790 ;
        RECT 75.090 49.045 75.350 49.885 ;
        RECT 75.525 49.795 76.045 50.335 ;
        RECT 76.215 49.965 76.735 50.505 ;
        RECT 76.905 50.625 77.215 51.425 ;
        RECT 77.385 50.795 77.695 51.595 ;
        RECT 77.865 50.965 78.125 51.425 ;
        RECT 78.295 51.135 78.550 51.595 ;
        RECT 78.725 50.965 78.985 51.425 ;
        RECT 77.865 50.795 78.985 50.965 ;
        RECT 76.905 50.455 77.935 50.625 ;
        RECT 75.525 49.045 76.735 49.795 ;
        RECT 76.905 49.545 77.075 50.455 ;
        RECT 77.245 49.715 77.595 50.285 ;
        RECT 77.765 50.205 77.935 50.455 ;
        RECT 78.725 50.545 78.985 50.795 ;
        RECT 79.155 50.725 79.440 51.595 ;
        RECT 78.725 50.375 79.480 50.545 ;
        RECT 77.765 50.035 78.905 50.205 ;
        RECT 79.075 49.865 79.480 50.375 ;
        RECT 77.830 49.695 79.480 49.865 ;
        RECT 79.670 50.455 80.005 51.425 ;
        RECT 80.175 50.455 80.345 51.595 ;
        RECT 80.515 51.255 82.545 51.425 ;
        RECT 79.670 49.785 79.840 50.455 ;
        RECT 80.515 50.285 80.685 51.255 ;
        RECT 80.010 49.955 80.265 50.285 ;
        RECT 80.490 49.955 80.685 50.285 ;
        RECT 80.855 50.915 81.980 51.085 ;
        RECT 80.095 49.785 80.265 49.955 ;
        RECT 80.855 49.785 81.025 50.915 ;
        RECT 76.905 49.215 77.205 49.545 ;
        RECT 77.375 49.045 77.650 49.525 ;
        RECT 77.830 49.305 78.125 49.695 ;
        RECT 78.295 49.045 78.550 49.525 ;
        RECT 78.725 49.305 78.985 49.695 ;
        RECT 79.155 49.045 79.435 49.525 ;
        RECT 79.670 49.215 79.925 49.785 ;
        RECT 80.095 49.615 81.025 49.785 ;
        RECT 81.195 50.575 82.205 50.745 ;
        RECT 81.195 49.775 81.365 50.575 ;
        RECT 81.570 50.235 81.845 50.375 ;
        RECT 81.565 50.065 81.845 50.235 ;
        RECT 80.850 49.580 81.025 49.615 ;
        RECT 80.095 49.045 80.425 49.445 ;
        RECT 80.850 49.215 81.380 49.580 ;
        RECT 81.570 49.215 81.845 50.065 ;
        RECT 82.015 49.215 82.205 50.575 ;
        RECT 82.375 50.590 82.545 51.255 ;
        RECT 82.715 50.835 82.885 51.595 ;
        RECT 83.120 50.835 83.635 51.245 ;
        RECT 82.375 50.400 83.125 50.590 ;
        RECT 83.295 50.025 83.635 50.835 ;
        RECT 84.010 50.625 84.340 51.425 ;
        RECT 84.510 50.795 84.840 51.595 ;
        RECT 85.140 50.625 85.470 51.425 ;
        RECT 86.115 50.795 86.365 51.595 ;
        RECT 84.010 50.455 86.445 50.625 ;
        RECT 86.635 50.455 86.805 51.595 ;
        RECT 86.975 50.455 87.315 51.425 ;
        RECT 83.805 50.035 84.155 50.285 ;
        RECT 82.405 49.855 83.635 50.025 ;
        RECT 82.385 49.045 82.895 49.580 ;
        RECT 83.115 49.250 83.360 49.855 ;
        RECT 84.340 49.825 84.510 50.455 ;
        RECT 84.680 50.035 85.010 50.235 ;
        RECT 85.180 50.035 85.510 50.235 ;
        RECT 85.680 50.035 86.100 50.235 ;
        RECT 86.275 50.205 86.445 50.455 ;
        RECT 86.275 50.035 86.970 50.205 ;
        RECT 84.010 49.215 84.510 49.825 ;
        RECT 85.140 49.695 86.365 49.865 ;
        RECT 87.140 49.845 87.315 50.455 ;
        RECT 85.140 49.215 85.470 49.695 ;
        RECT 85.640 49.045 85.865 49.505 ;
        RECT 86.035 49.215 86.365 49.695 ;
        RECT 86.555 49.045 86.805 49.845 ;
        RECT 86.975 49.215 87.315 49.845 ;
        RECT 87.485 50.455 87.825 51.425 ;
        RECT 87.995 50.455 88.165 51.595 ;
        RECT 88.435 50.795 88.685 51.595 ;
        RECT 89.330 50.625 89.660 51.425 ;
        RECT 89.960 50.795 90.290 51.595 ;
        RECT 90.460 50.625 90.790 51.425 ;
        RECT 88.355 50.455 90.790 50.625 ;
        RECT 91.165 50.455 91.505 51.425 ;
        RECT 91.675 50.455 91.845 51.595 ;
        RECT 92.115 50.795 92.365 51.595 ;
        RECT 93.010 50.625 93.340 51.425 ;
        RECT 93.640 50.795 93.970 51.595 ;
        RECT 94.140 50.625 94.470 51.425 ;
        RECT 92.035 50.455 94.470 50.625 ;
        RECT 87.485 50.405 87.715 50.455 ;
        RECT 87.485 49.845 87.660 50.405 ;
        RECT 88.355 50.205 88.525 50.455 ;
        RECT 87.830 50.035 88.525 50.205 ;
        RECT 88.700 50.035 89.120 50.235 ;
        RECT 89.290 50.035 89.620 50.235 ;
        RECT 89.790 50.035 90.120 50.235 ;
        RECT 87.485 49.215 87.825 49.845 ;
        RECT 87.995 49.045 88.245 49.845 ;
        RECT 88.435 49.695 89.660 49.865 ;
        RECT 88.435 49.215 88.765 49.695 ;
        RECT 88.935 49.045 89.160 49.505 ;
        RECT 89.330 49.215 89.660 49.695 ;
        RECT 90.290 49.825 90.460 50.455 ;
        RECT 90.645 50.035 90.995 50.285 ;
        RECT 91.165 49.845 91.340 50.455 ;
        RECT 92.035 50.205 92.205 50.455 ;
        RECT 91.510 50.035 92.205 50.205 ;
        RECT 92.380 50.035 92.800 50.235 ;
        RECT 92.970 50.035 93.300 50.235 ;
        RECT 93.470 50.035 93.800 50.235 ;
        RECT 90.290 49.215 90.790 49.825 ;
        RECT 91.165 49.215 91.505 49.845 ;
        RECT 91.675 49.045 91.925 49.845 ;
        RECT 92.115 49.695 93.340 49.865 ;
        RECT 92.115 49.215 92.445 49.695 ;
        RECT 92.615 49.045 92.840 49.505 ;
        RECT 93.010 49.215 93.340 49.695 ;
        RECT 93.970 49.825 94.140 50.455 ;
        RECT 95.765 50.430 96.055 51.595 ;
        RECT 96.430 50.625 96.760 51.425 ;
        RECT 96.930 50.795 97.260 51.595 ;
        RECT 97.560 50.625 97.890 51.425 ;
        RECT 98.535 50.795 98.785 51.595 ;
        RECT 96.430 50.455 98.865 50.625 ;
        RECT 99.055 50.455 99.225 51.595 ;
        RECT 99.395 50.455 99.735 51.425 ;
        RECT 94.325 50.035 94.675 50.285 ;
        RECT 96.225 50.035 96.575 50.285 ;
        RECT 96.760 49.825 96.930 50.455 ;
        RECT 97.100 50.035 97.430 50.235 ;
        RECT 97.600 50.035 97.930 50.235 ;
        RECT 98.100 50.035 98.520 50.235 ;
        RECT 98.695 50.205 98.865 50.455 ;
        RECT 98.695 50.035 99.390 50.205 ;
        RECT 93.970 49.215 94.470 49.825 ;
        RECT 95.765 49.045 96.055 49.770 ;
        RECT 96.430 49.215 96.930 49.825 ;
        RECT 97.560 49.695 98.785 49.865 ;
        RECT 99.560 49.845 99.735 50.455 ;
        RECT 97.560 49.215 97.890 49.695 ;
        RECT 98.060 49.045 98.285 49.505 ;
        RECT 98.455 49.215 98.785 49.695 ;
        RECT 98.975 49.045 99.225 49.845 ;
        RECT 99.395 49.215 99.735 49.845 ;
        RECT 99.905 50.455 100.245 51.425 ;
        RECT 100.415 50.455 100.585 51.595 ;
        RECT 100.855 50.795 101.105 51.595 ;
        RECT 101.750 50.625 102.080 51.425 ;
        RECT 102.380 50.795 102.710 51.595 ;
        RECT 102.880 50.625 103.210 51.425 ;
        RECT 100.775 50.455 103.210 50.625 ;
        RECT 103.585 50.455 103.925 51.425 ;
        RECT 104.095 50.455 104.265 51.595 ;
        RECT 104.535 50.795 104.785 51.595 ;
        RECT 105.430 50.625 105.760 51.425 ;
        RECT 106.060 50.795 106.390 51.595 ;
        RECT 106.560 50.625 106.890 51.425 ;
        RECT 107.265 51.160 112.610 51.595 ;
        RECT 112.785 51.160 118.130 51.595 ;
        RECT 104.455 50.455 106.890 50.625 ;
        RECT 99.905 49.845 100.080 50.455 ;
        RECT 100.775 50.205 100.945 50.455 ;
        RECT 100.250 50.035 100.945 50.205 ;
        RECT 101.120 50.035 101.540 50.235 ;
        RECT 101.710 50.035 102.040 50.235 ;
        RECT 102.210 50.035 102.540 50.235 ;
        RECT 99.905 49.215 100.245 49.845 ;
        RECT 100.415 49.045 100.665 49.845 ;
        RECT 100.855 49.695 102.080 49.865 ;
        RECT 100.855 49.215 101.185 49.695 ;
        RECT 101.355 49.045 101.580 49.505 ;
        RECT 101.750 49.215 102.080 49.695 ;
        RECT 102.710 49.825 102.880 50.455 ;
        RECT 103.065 50.035 103.415 50.285 ;
        RECT 103.585 49.845 103.760 50.455 ;
        RECT 104.455 50.205 104.625 50.455 ;
        RECT 103.930 50.035 104.625 50.205 ;
        RECT 104.800 50.035 105.220 50.235 ;
        RECT 105.390 50.035 105.720 50.235 ;
        RECT 105.890 50.035 106.220 50.235 ;
        RECT 102.710 49.215 103.210 49.825 ;
        RECT 103.585 49.215 103.925 49.845 ;
        RECT 104.095 49.045 104.345 49.845 ;
        RECT 104.535 49.695 105.760 49.865 ;
        RECT 104.535 49.215 104.865 49.695 ;
        RECT 105.035 49.045 105.260 49.505 ;
        RECT 105.430 49.215 105.760 49.695 ;
        RECT 106.390 49.825 106.560 50.455 ;
        RECT 106.745 50.035 107.095 50.285 ;
        RECT 106.390 49.215 106.890 49.825 ;
        RECT 108.850 49.590 109.190 50.420 ;
        RECT 110.670 49.910 111.020 51.160 ;
        RECT 114.370 49.590 114.710 50.420 ;
        RECT 116.190 49.910 116.540 51.160 ;
        RECT 118.305 50.505 120.895 51.595 ;
        RECT 118.305 49.815 119.515 50.335 ;
        RECT 119.685 49.985 120.895 50.505 ;
        RECT 121.525 50.430 121.815 51.595 ;
        RECT 122.445 50.505 123.655 51.595 ;
        RECT 122.445 49.965 122.965 50.505 ;
        RECT 107.265 49.045 112.610 49.590 ;
        RECT 112.785 49.045 118.130 49.590 ;
        RECT 118.305 49.045 120.895 49.815 ;
        RECT 123.135 49.795 123.655 50.335 ;
        RECT 121.525 49.045 121.815 49.770 ;
        RECT 122.445 49.045 123.655 49.795 ;
        RECT 5.520 48.875 123.740 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.985 48.105 10.495 48.875 ;
        RECT 10.665 48.125 11.875 48.875 ;
        RECT 12.045 48.200 12.305 48.705 ;
        RECT 12.485 48.495 12.815 48.875 ;
        RECT 12.995 48.325 13.165 48.705 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 6.985 47.585 8.635 48.105 ;
        RECT 8.805 47.415 10.495 47.935 ;
        RECT 10.665 47.585 11.185 48.125 ;
        RECT 11.355 47.415 11.875 47.955 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 6.985 46.325 10.495 47.415 ;
        RECT 10.665 46.325 11.875 47.415 ;
        RECT 12.045 47.400 12.215 48.200 ;
        RECT 12.500 48.155 13.165 48.325 ;
        RECT 13.425 48.200 13.685 48.705 ;
        RECT 13.865 48.495 14.195 48.875 ;
        RECT 14.375 48.325 14.545 48.705 ;
        RECT 12.500 47.900 12.670 48.155 ;
        RECT 12.385 47.570 12.670 47.900 ;
        RECT 12.905 47.605 13.235 47.975 ;
        RECT 12.500 47.425 12.670 47.570 ;
        RECT 12.045 46.495 12.315 47.400 ;
        RECT 12.500 47.255 13.165 47.425 ;
        RECT 12.485 46.325 12.815 47.085 ;
        RECT 12.995 46.495 13.165 47.255 ;
        RECT 13.425 47.400 13.595 48.200 ;
        RECT 13.880 48.155 14.545 48.325 ;
        RECT 13.880 47.900 14.050 48.155 ;
        RECT 14.865 48.055 15.075 48.875 ;
        RECT 15.245 48.075 15.575 48.705 ;
        RECT 13.765 47.570 14.050 47.900 ;
        RECT 14.285 47.605 14.615 47.975 ;
        RECT 13.880 47.425 14.050 47.570 ;
        RECT 15.245 47.475 15.495 48.075 ;
        RECT 15.745 48.055 15.975 48.875 ;
        RECT 16.650 48.135 16.905 48.705 ;
        RECT 17.075 48.475 17.405 48.875 ;
        RECT 17.830 48.340 18.360 48.705 ;
        RECT 17.830 48.305 18.005 48.340 ;
        RECT 17.075 48.135 18.005 48.305 ;
        RECT 15.665 47.635 15.995 47.885 ;
        RECT 13.425 46.495 13.695 47.400 ;
        RECT 13.880 47.255 14.545 47.425 ;
        RECT 13.865 46.325 14.195 47.085 ;
        RECT 14.375 46.495 14.545 47.255 ;
        RECT 14.865 46.325 15.075 47.465 ;
        RECT 15.245 46.495 15.575 47.475 ;
        RECT 16.650 47.465 16.820 48.135 ;
        RECT 17.075 47.965 17.245 48.135 ;
        RECT 16.990 47.635 17.245 47.965 ;
        RECT 17.470 47.635 17.665 47.965 ;
        RECT 15.745 46.325 15.975 47.465 ;
        RECT 16.650 46.495 16.985 47.465 ;
        RECT 17.155 46.325 17.325 47.465 ;
        RECT 17.495 46.665 17.665 47.635 ;
        RECT 17.835 47.005 18.005 48.135 ;
        RECT 18.175 47.345 18.345 48.145 ;
        RECT 18.550 47.855 18.825 48.705 ;
        RECT 18.545 47.685 18.825 47.855 ;
        RECT 18.550 47.545 18.825 47.685 ;
        RECT 18.995 47.345 19.185 48.705 ;
        RECT 19.365 48.340 19.875 48.875 ;
        RECT 20.095 48.065 20.340 48.670 ;
        RECT 20.785 48.105 22.455 48.875 ;
        RECT 19.385 47.895 20.615 48.065 ;
        RECT 18.175 47.175 19.185 47.345 ;
        RECT 19.355 47.330 20.105 47.520 ;
        RECT 17.835 46.835 18.960 47.005 ;
        RECT 19.355 46.665 19.525 47.330 ;
        RECT 20.275 47.085 20.615 47.895 ;
        RECT 20.785 47.585 21.535 48.105 ;
        RECT 23.085 48.075 23.425 48.705 ;
        RECT 23.595 48.075 23.845 48.875 ;
        RECT 24.035 48.225 24.365 48.705 ;
        RECT 24.535 48.415 24.760 48.875 ;
        RECT 24.930 48.225 25.260 48.705 ;
        RECT 23.085 48.025 23.315 48.075 ;
        RECT 24.035 48.055 25.260 48.225 ;
        RECT 25.890 48.095 26.390 48.705 ;
        RECT 26.970 48.095 27.470 48.705 ;
        RECT 21.705 47.415 22.455 47.935 ;
        RECT 17.495 46.495 19.525 46.665 ;
        RECT 19.695 46.325 19.865 47.085 ;
        RECT 20.100 46.675 20.615 47.085 ;
        RECT 20.785 46.325 22.455 47.415 ;
        RECT 23.085 47.465 23.260 48.025 ;
        RECT 23.430 47.715 24.125 47.885 ;
        RECT 23.955 47.465 24.125 47.715 ;
        RECT 24.300 47.685 24.720 47.885 ;
        RECT 24.890 47.685 25.220 47.885 ;
        RECT 25.390 47.685 25.720 47.885 ;
        RECT 25.890 47.465 26.060 48.095 ;
        RECT 26.245 47.635 26.595 47.885 ;
        RECT 26.765 47.635 27.115 47.885 ;
        RECT 27.300 47.465 27.470 48.095 ;
        RECT 28.100 48.225 28.430 48.705 ;
        RECT 28.600 48.415 28.825 48.875 ;
        RECT 28.995 48.225 29.325 48.705 ;
        RECT 28.100 48.055 29.325 48.225 ;
        RECT 29.515 48.075 29.765 48.875 ;
        RECT 29.935 48.075 30.275 48.705 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 32.030 48.095 32.530 48.705 ;
        RECT 30.045 48.025 30.275 48.075 ;
        RECT 27.640 47.685 27.970 47.885 ;
        RECT 28.140 47.685 28.470 47.885 ;
        RECT 28.640 47.685 29.060 47.885 ;
        RECT 29.235 47.715 29.930 47.885 ;
        RECT 29.235 47.465 29.405 47.715 ;
        RECT 30.100 47.465 30.275 48.025 ;
        RECT 31.825 47.635 32.175 47.885 ;
        RECT 23.085 46.495 23.425 47.465 ;
        RECT 23.595 46.325 23.765 47.465 ;
        RECT 23.955 47.295 26.390 47.465 ;
        RECT 24.035 46.325 24.285 47.125 ;
        RECT 24.930 46.495 25.260 47.295 ;
        RECT 25.560 46.325 25.890 47.125 ;
        RECT 26.060 46.495 26.390 47.295 ;
        RECT 26.970 47.295 29.405 47.465 ;
        RECT 26.970 46.495 27.300 47.295 ;
        RECT 27.470 46.325 27.800 47.125 ;
        RECT 28.100 46.495 28.430 47.295 ;
        RECT 29.075 46.325 29.325 47.125 ;
        RECT 29.595 46.325 29.765 47.465 ;
        RECT 29.935 46.495 30.275 47.465 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 32.360 47.465 32.530 48.095 ;
        RECT 33.160 48.225 33.490 48.705 ;
        RECT 33.660 48.415 33.885 48.875 ;
        RECT 34.055 48.225 34.385 48.705 ;
        RECT 33.160 48.055 34.385 48.225 ;
        RECT 34.575 48.075 34.825 48.875 ;
        RECT 34.995 48.075 35.335 48.705 ;
        RECT 35.105 48.025 35.335 48.075 ;
        RECT 32.700 47.685 33.030 47.885 ;
        RECT 33.200 47.685 33.530 47.885 ;
        RECT 33.700 47.685 34.120 47.885 ;
        RECT 34.295 47.715 34.990 47.885 ;
        RECT 34.295 47.465 34.465 47.715 ;
        RECT 35.160 47.465 35.335 48.025 ;
        RECT 35.505 48.125 36.715 48.875 ;
        RECT 36.885 48.200 37.145 48.705 ;
        RECT 37.325 48.495 37.655 48.875 ;
        RECT 37.835 48.325 38.005 48.705 ;
        RECT 38.265 48.330 43.610 48.875 ;
        RECT 35.505 47.585 36.025 48.125 ;
        RECT 32.030 47.295 34.465 47.465 ;
        RECT 32.030 46.495 32.360 47.295 ;
        RECT 32.530 46.325 32.860 47.125 ;
        RECT 33.160 46.495 33.490 47.295 ;
        RECT 34.135 46.325 34.385 47.125 ;
        RECT 34.655 46.325 34.825 47.465 ;
        RECT 34.995 46.495 35.335 47.465 ;
        RECT 36.195 47.415 36.715 47.955 ;
        RECT 35.505 46.325 36.715 47.415 ;
        RECT 36.885 47.400 37.055 48.200 ;
        RECT 37.340 48.155 38.005 48.325 ;
        RECT 37.340 47.900 37.510 48.155 ;
        RECT 37.225 47.570 37.510 47.900 ;
        RECT 37.745 47.605 38.075 47.975 ;
        RECT 37.340 47.425 37.510 47.570 ;
        RECT 39.850 47.500 40.190 48.330 ;
        RECT 43.785 48.105 46.375 48.875 ;
        RECT 46.605 48.395 46.885 48.875 ;
        RECT 47.055 48.225 47.315 48.615 ;
        RECT 47.490 48.395 47.745 48.875 ;
        RECT 47.915 48.225 48.210 48.615 ;
        RECT 48.390 48.395 48.665 48.875 ;
        RECT 48.835 48.375 49.135 48.705 ;
        RECT 36.885 46.495 37.155 47.400 ;
        RECT 37.340 47.255 38.005 47.425 ;
        RECT 37.325 46.325 37.655 47.085 ;
        RECT 37.835 46.495 38.005 47.255 ;
        RECT 41.670 46.760 42.020 48.010 ;
        RECT 43.785 47.585 44.995 48.105 ;
        RECT 46.560 48.055 48.210 48.225 ;
        RECT 45.165 47.415 46.375 47.935 ;
        RECT 38.265 46.325 43.610 46.760 ;
        RECT 43.785 46.325 46.375 47.415 ;
        RECT 46.560 47.545 46.965 48.055 ;
        RECT 47.135 47.715 48.275 47.885 ;
        RECT 46.560 47.375 47.315 47.545 ;
        RECT 46.600 46.325 46.885 47.195 ;
        RECT 47.055 47.125 47.315 47.375 ;
        RECT 48.105 47.465 48.275 47.715 ;
        RECT 48.445 47.635 48.795 48.205 ;
        RECT 48.965 47.465 49.135 48.375 ;
        RECT 49.510 48.095 50.010 48.705 ;
        RECT 49.305 47.635 49.655 47.885 ;
        RECT 49.840 47.465 50.010 48.095 ;
        RECT 50.640 48.225 50.970 48.705 ;
        RECT 51.140 48.415 51.365 48.875 ;
        RECT 51.535 48.225 51.865 48.705 ;
        RECT 50.640 48.055 51.865 48.225 ;
        RECT 52.055 48.075 52.305 48.875 ;
        RECT 52.475 48.075 52.815 48.705 ;
        RECT 52.585 48.025 52.815 48.075 ;
        RECT 50.180 47.685 50.510 47.885 ;
        RECT 50.680 47.685 51.010 47.885 ;
        RECT 51.180 47.685 51.600 47.885 ;
        RECT 51.775 47.715 52.470 47.885 ;
        RECT 51.775 47.465 51.945 47.715 ;
        RECT 52.640 47.465 52.815 48.025 ;
        RECT 52.985 48.105 56.495 48.875 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 52.985 47.585 54.635 48.105 ;
        RECT 57.625 48.055 57.855 48.875 ;
        RECT 58.025 48.075 58.355 48.705 ;
        RECT 48.105 47.295 49.135 47.465 ;
        RECT 47.055 46.955 48.175 47.125 ;
        RECT 47.055 46.495 47.315 46.955 ;
        RECT 47.490 46.325 47.745 46.785 ;
        RECT 47.915 46.495 48.175 46.955 ;
        RECT 48.345 46.325 48.655 47.125 ;
        RECT 48.825 46.495 49.135 47.295 ;
        RECT 49.510 47.295 51.945 47.465 ;
        RECT 49.510 46.495 49.840 47.295 ;
        RECT 50.010 46.325 50.340 47.125 ;
        RECT 50.640 46.495 50.970 47.295 ;
        RECT 51.615 46.325 51.865 47.125 ;
        RECT 52.135 46.325 52.305 47.465 ;
        RECT 52.475 46.495 52.815 47.465 ;
        RECT 54.805 47.415 56.495 47.935 ;
        RECT 57.605 47.635 57.935 47.885 ;
        RECT 52.985 46.325 56.495 47.415 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 58.105 47.475 58.355 48.075 ;
        RECT 58.525 48.055 58.735 48.875 ;
        RECT 58.965 48.330 64.310 48.875 ;
        RECT 60.550 47.500 60.890 48.330 ;
        RECT 65.710 48.305 65.880 48.555 ;
        RECT 65.405 48.135 65.880 48.305 ;
        RECT 66.115 48.135 66.445 48.875 ;
        RECT 66.615 48.305 66.815 48.650 ;
        RECT 66.985 48.475 67.315 48.875 ;
        RECT 67.485 48.305 67.685 48.660 ;
        RECT 67.855 48.480 68.185 48.875 ;
        RECT 68.625 48.330 73.970 48.875 ;
        RECT 74.145 48.330 79.490 48.875 ;
        RECT 66.615 48.135 68.455 48.305 ;
        RECT 57.625 46.325 57.855 47.465 ;
        RECT 58.025 46.495 58.355 47.475 ;
        RECT 58.525 46.325 58.735 47.465 ;
        RECT 62.370 46.760 62.720 48.010 ;
        RECT 65.405 47.165 65.575 48.135 ;
        RECT 65.745 47.345 66.095 47.965 ;
        RECT 66.265 47.345 66.585 47.965 ;
        RECT 66.755 47.345 67.085 47.965 ;
        RECT 67.255 47.345 67.555 47.965 ;
        RECT 67.795 47.165 68.015 47.965 ;
        RECT 65.405 46.955 68.015 47.165 ;
        RECT 58.965 46.325 64.310 46.760 ;
        RECT 66.115 46.325 66.445 46.775 ;
        RECT 68.195 46.510 68.455 48.135 ;
        RECT 70.210 47.500 70.550 48.330 ;
        RECT 72.030 46.760 72.380 48.010 ;
        RECT 75.730 47.500 76.070 48.330 ;
        RECT 79.665 48.105 82.255 48.875 ;
        RECT 82.885 48.150 83.175 48.875 ;
        RECT 83.350 48.135 83.605 48.705 ;
        RECT 83.775 48.475 84.105 48.875 ;
        RECT 84.530 48.340 85.060 48.705 ;
        RECT 84.530 48.305 84.705 48.340 ;
        RECT 83.775 48.135 84.705 48.305 ;
        RECT 85.250 48.195 85.525 48.705 ;
        RECT 77.550 46.760 77.900 48.010 ;
        RECT 79.665 47.585 80.875 48.105 ;
        RECT 81.045 47.415 82.255 47.935 ;
        RECT 68.625 46.325 73.970 46.760 ;
        RECT 74.145 46.325 79.490 46.760 ;
        RECT 79.665 46.325 82.255 47.415 ;
        RECT 82.885 46.325 83.175 47.490 ;
        RECT 83.350 47.465 83.520 48.135 ;
        RECT 83.775 47.965 83.945 48.135 ;
        RECT 83.690 47.635 83.945 47.965 ;
        RECT 84.170 47.635 84.365 47.965 ;
        RECT 83.350 46.495 83.685 47.465 ;
        RECT 83.855 46.325 84.025 47.465 ;
        RECT 84.195 46.665 84.365 47.635 ;
        RECT 84.535 47.005 84.705 48.135 ;
        RECT 84.875 47.345 85.045 48.145 ;
        RECT 85.245 48.025 85.525 48.195 ;
        RECT 85.250 47.545 85.525 48.025 ;
        RECT 85.695 47.345 85.885 48.705 ;
        RECT 86.065 48.340 86.575 48.875 ;
        RECT 86.795 48.065 87.040 48.670 ;
        RECT 87.690 48.095 88.190 48.705 ;
        RECT 86.085 47.895 87.315 48.065 ;
        RECT 84.875 47.175 85.885 47.345 ;
        RECT 86.055 47.330 86.805 47.520 ;
        RECT 84.535 46.835 85.660 47.005 ;
        RECT 86.055 46.665 86.225 47.330 ;
        RECT 86.975 47.085 87.315 47.895 ;
        RECT 87.485 47.635 87.835 47.885 ;
        RECT 88.020 47.465 88.190 48.095 ;
        RECT 88.820 48.225 89.150 48.705 ;
        RECT 89.320 48.415 89.545 48.875 ;
        RECT 89.715 48.225 90.045 48.705 ;
        RECT 88.820 48.055 90.045 48.225 ;
        RECT 90.235 48.075 90.485 48.875 ;
        RECT 90.655 48.075 90.995 48.705 ;
        RECT 91.370 48.095 91.870 48.705 ;
        RECT 90.765 48.025 90.995 48.075 ;
        RECT 88.360 47.685 88.690 47.885 ;
        RECT 88.860 47.685 89.190 47.885 ;
        RECT 89.360 47.685 89.780 47.885 ;
        RECT 89.955 47.715 90.650 47.885 ;
        RECT 89.955 47.465 90.125 47.715 ;
        RECT 90.820 47.465 90.995 48.025 ;
        RECT 91.165 47.635 91.515 47.885 ;
        RECT 91.700 47.465 91.870 48.095 ;
        RECT 92.500 48.225 92.830 48.705 ;
        RECT 93.000 48.415 93.225 48.875 ;
        RECT 93.395 48.225 93.725 48.705 ;
        RECT 92.500 48.055 93.725 48.225 ;
        RECT 93.915 48.075 94.165 48.875 ;
        RECT 94.335 48.075 94.675 48.705 ;
        RECT 94.445 48.025 94.675 48.075 ;
        RECT 92.040 47.685 92.370 47.885 ;
        RECT 92.540 47.685 92.870 47.885 ;
        RECT 93.040 47.685 93.460 47.885 ;
        RECT 93.635 47.715 94.330 47.885 ;
        RECT 93.635 47.465 93.805 47.715 ;
        RECT 94.500 47.465 94.675 48.025 ;
        RECT 94.845 48.105 98.355 48.875 ;
        RECT 94.845 47.585 96.495 48.105 ;
        RECT 99.720 48.065 99.965 48.670 ;
        RECT 100.185 48.340 100.695 48.875 ;
        RECT 84.195 46.495 86.225 46.665 ;
        RECT 86.395 46.325 86.565 47.085 ;
        RECT 86.800 46.675 87.315 47.085 ;
        RECT 87.690 47.295 90.125 47.465 ;
        RECT 87.690 46.495 88.020 47.295 ;
        RECT 88.190 46.325 88.520 47.125 ;
        RECT 88.820 46.495 89.150 47.295 ;
        RECT 89.795 46.325 90.045 47.125 ;
        RECT 90.315 46.325 90.485 47.465 ;
        RECT 90.655 46.495 90.995 47.465 ;
        RECT 91.370 47.295 93.805 47.465 ;
        RECT 91.370 46.495 91.700 47.295 ;
        RECT 91.870 46.325 92.200 47.125 ;
        RECT 92.500 46.495 92.830 47.295 ;
        RECT 93.475 46.325 93.725 47.125 ;
        RECT 93.995 46.325 94.165 47.465 ;
        RECT 94.335 46.495 94.675 47.465 ;
        RECT 96.665 47.415 98.355 47.935 ;
        RECT 94.845 46.325 98.355 47.415 ;
        RECT 99.445 47.895 100.675 48.065 ;
        RECT 99.445 47.085 99.785 47.895 ;
        RECT 99.955 47.330 100.705 47.520 ;
        RECT 99.445 46.675 99.960 47.085 ;
        RECT 100.195 46.325 100.365 47.085 ;
        RECT 100.535 46.665 100.705 47.330 ;
        RECT 100.875 47.345 101.065 48.705 ;
        RECT 101.235 47.855 101.510 48.705 ;
        RECT 101.700 48.340 102.230 48.705 ;
        RECT 102.655 48.475 102.985 48.875 ;
        RECT 102.055 48.305 102.230 48.340 ;
        RECT 101.235 47.685 101.515 47.855 ;
        RECT 101.235 47.545 101.510 47.685 ;
        RECT 101.715 47.345 101.885 48.145 ;
        RECT 100.875 47.175 101.885 47.345 ;
        RECT 102.055 48.135 102.985 48.305 ;
        RECT 103.155 48.135 103.410 48.705 ;
        RECT 102.055 47.005 102.225 48.135 ;
        RECT 102.815 47.965 102.985 48.135 ;
        RECT 101.100 46.835 102.225 47.005 ;
        RECT 102.395 47.635 102.590 47.965 ;
        RECT 102.815 47.635 103.070 47.965 ;
        RECT 102.395 46.665 102.565 47.635 ;
        RECT 103.240 47.465 103.410 48.135 ;
        RECT 100.535 46.495 102.565 46.665 ;
        RECT 102.735 46.325 102.905 47.465 ;
        RECT 103.075 46.495 103.410 47.465 ;
        RECT 103.585 48.200 103.845 48.705 ;
        RECT 104.025 48.495 104.355 48.875 ;
        RECT 104.535 48.325 104.705 48.705 ;
        RECT 103.585 47.400 103.755 48.200 ;
        RECT 104.040 48.155 104.705 48.325 ;
        RECT 105.975 48.325 106.145 48.705 ;
        RECT 106.325 48.495 106.655 48.875 ;
        RECT 105.975 48.155 106.640 48.325 ;
        RECT 106.835 48.200 107.095 48.705 ;
        RECT 104.040 47.900 104.210 48.155 ;
        RECT 103.925 47.570 104.210 47.900 ;
        RECT 104.445 47.605 104.775 47.975 ;
        RECT 105.905 47.605 106.235 47.975 ;
        RECT 106.470 47.900 106.640 48.155 ;
        RECT 104.040 47.425 104.210 47.570 ;
        RECT 106.470 47.570 106.755 47.900 ;
        RECT 106.470 47.425 106.640 47.570 ;
        RECT 103.585 46.495 103.855 47.400 ;
        RECT 104.040 47.255 104.705 47.425 ;
        RECT 104.025 46.325 104.355 47.085 ;
        RECT 104.535 46.495 104.705 47.255 ;
        RECT 105.975 47.255 106.640 47.425 ;
        RECT 106.925 47.400 107.095 48.200 ;
        RECT 107.265 48.125 108.475 48.875 ;
        RECT 108.645 48.150 108.935 48.875 ;
        RECT 107.265 47.585 107.785 48.125 ;
        RECT 109.165 48.055 109.375 48.875 ;
        RECT 109.545 48.075 109.875 48.705 ;
        RECT 107.955 47.415 108.475 47.955 ;
        RECT 105.975 46.495 106.145 47.255 ;
        RECT 106.325 46.325 106.655 47.085 ;
        RECT 106.825 46.495 107.095 47.400 ;
        RECT 107.265 46.325 108.475 47.415 ;
        RECT 108.645 46.325 108.935 47.490 ;
        RECT 109.545 47.475 109.795 48.075 ;
        RECT 110.045 48.055 110.275 48.875 ;
        RECT 110.485 48.330 115.830 48.875 ;
        RECT 116.005 48.330 121.350 48.875 ;
        RECT 109.965 47.635 110.295 47.885 ;
        RECT 112.070 47.500 112.410 48.330 ;
        RECT 109.165 46.325 109.375 47.465 ;
        RECT 109.545 46.495 109.875 47.475 ;
        RECT 110.045 46.325 110.275 47.465 ;
        RECT 113.890 46.760 114.240 48.010 ;
        RECT 117.590 47.500 117.930 48.330 ;
        RECT 122.445 48.125 123.655 48.875 ;
        RECT 119.410 46.760 119.760 48.010 ;
        RECT 122.445 47.415 122.965 47.955 ;
        RECT 123.135 47.585 123.655 48.125 ;
        RECT 110.485 46.325 115.830 46.760 ;
        RECT 116.005 46.325 121.350 46.760 ;
        RECT 122.445 46.325 123.655 47.415 ;
        RECT 5.520 46.155 123.740 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 6.985 45.065 8.655 46.155 ;
        RECT 9.290 45.485 9.545 45.985 ;
        RECT 9.715 45.655 10.045 46.155 ;
        RECT 9.290 45.315 10.040 45.485 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 6.985 44.375 7.735 44.895 ;
        RECT 7.905 44.545 8.655 45.065 ;
        RECT 9.290 44.495 9.640 45.145 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 6.985 43.605 8.655 44.375 ;
        RECT 9.810 44.325 10.040 45.315 ;
        RECT 9.290 44.155 10.040 44.325 ;
        RECT 9.290 43.865 9.545 44.155 ;
        RECT 9.715 43.605 10.045 43.985 ;
        RECT 10.215 43.865 10.385 45.985 ;
        RECT 10.555 45.185 10.880 45.970 ;
        RECT 11.050 45.695 11.300 46.155 ;
        RECT 11.470 45.655 11.720 45.985 ;
        RECT 11.935 45.655 12.615 45.985 ;
        RECT 11.470 45.525 11.640 45.655 ;
        RECT 11.245 45.355 11.640 45.525 ;
        RECT 10.615 44.135 11.075 45.185 ;
        RECT 11.245 43.995 11.415 45.355 ;
        RECT 11.810 45.095 12.275 45.485 ;
        RECT 11.585 44.285 11.935 44.905 ;
        RECT 12.105 44.505 12.275 45.095 ;
        RECT 12.445 44.875 12.615 45.655 ;
        RECT 12.785 45.555 12.955 45.895 ;
        RECT 13.190 45.725 13.520 46.155 ;
        RECT 13.690 45.555 13.860 45.895 ;
        RECT 14.155 45.695 14.525 46.155 ;
        RECT 12.785 45.385 13.860 45.555 ;
        RECT 14.695 45.525 14.865 45.985 ;
        RECT 15.100 45.645 15.970 45.985 ;
        RECT 16.140 45.695 16.390 46.155 ;
        RECT 14.305 45.355 14.865 45.525 ;
        RECT 14.305 45.215 14.475 45.355 ;
        RECT 12.975 45.045 14.475 45.215 ;
        RECT 15.170 45.185 15.630 45.475 ;
        RECT 12.445 44.705 14.135 44.875 ;
        RECT 12.105 44.285 12.460 44.505 ;
        RECT 12.630 43.995 12.800 44.705 ;
        RECT 13.005 44.285 13.795 44.535 ;
        RECT 13.965 44.525 14.135 44.705 ;
        RECT 14.305 44.355 14.475 45.045 ;
        RECT 10.745 43.605 11.075 43.965 ;
        RECT 11.245 43.825 11.740 43.995 ;
        RECT 11.945 43.825 12.800 43.995 ;
        RECT 13.675 43.605 14.005 44.065 ;
        RECT 14.215 43.965 14.475 44.355 ;
        RECT 14.665 45.175 15.630 45.185 ;
        RECT 15.800 45.265 15.970 45.645 ;
        RECT 16.560 45.605 16.730 45.895 ;
        RECT 16.910 45.775 17.240 46.155 ;
        RECT 16.560 45.435 17.360 45.605 ;
        RECT 14.665 45.015 15.340 45.175 ;
        RECT 15.800 45.095 17.020 45.265 ;
        RECT 14.665 44.225 14.875 45.015 ;
        RECT 15.800 45.005 15.970 45.095 ;
        RECT 15.045 44.225 15.395 44.845 ;
        RECT 15.565 44.835 15.970 45.005 ;
        RECT 15.565 44.055 15.735 44.835 ;
        RECT 15.905 44.385 16.125 44.665 ;
        RECT 16.305 44.555 16.845 44.925 ;
        RECT 17.190 44.845 17.360 45.435 ;
        RECT 17.580 45.015 17.885 46.155 ;
        RECT 18.055 44.965 18.310 45.845 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 18.950 45.015 19.285 45.985 ;
        RECT 19.455 45.015 19.625 46.155 ;
        RECT 19.795 45.815 21.825 45.985 ;
        RECT 17.190 44.815 17.930 44.845 ;
        RECT 15.905 44.215 16.435 44.385 ;
        RECT 14.215 43.795 14.565 43.965 ;
        RECT 14.785 43.775 15.735 44.055 ;
        RECT 15.905 43.605 16.095 44.045 ;
        RECT 16.265 43.985 16.435 44.215 ;
        RECT 16.605 44.155 16.845 44.555 ;
        RECT 17.015 44.515 17.930 44.815 ;
        RECT 17.015 44.340 17.340 44.515 ;
        RECT 17.015 43.985 17.335 44.340 ;
        RECT 18.100 44.315 18.310 44.965 ;
        RECT 18.950 44.345 19.120 45.015 ;
        RECT 19.795 44.845 19.965 45.815 ;
        RECT 19.290 44.515 19.545 44.845 ;
        RECT 19.770 44.515 19.965 44.845 ;
        RECT 20.135 45.475 21.260 45.645 ;
        RECT 19.375 44.345 19.545 44.515 ;
        RECT 20.135 44.345 20.305 45.475 ;
        RECT 16.265 43.815 17.335 43.985 ;
        RECT 17.580 43.605 17.885 44.065 ;
        RECT 18.055 43.785 18.310 44.315 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 18.950 43.775 19.205 44.345 ;
        RECT 19.375 44.175 20.305 44.345 ;
        RECT 20.475 45.135 21.485 45.305 ;
        RECT 20.475 44.335 20.645 45.135 ;
        RECT 20.130 44.140 20.305 44.175 ;
        RECT 19.375 43.605 19.705 44.005 ;
        RECT 20.130 43.775 20.660 44.140 ;
        RECT 20.850 44.115 21.125 44.935 ;
        RECT 20.845 43.945 21.125 44.115 ;
        RECT 20.850 43.775 21.125 43.945 ;
        RECT 21.295 43.775 21.485 45.135 ;
        RECT 21.655 45.150 21.825 45.815 ;
        RECT 21.995 45.395 22.165 46.155 ;
        RECT 22.400 45.395 22.915 45.805 ;
        RECT 21.655 44.960 22.405 45.150 ;
        RECT 22.575 44.585 22.915 45.395 ;
        RECT 23.085 45.065 25.675 46.155 ;
        RECT 21.685 44.415 22.915 44.585 ;
        RECT 21.665 43.605 22.175 44.140 ;
        RECT 22.395 43.810 22.640 44.415 ;
        RECT 23.085 44.375 24.295 44.895 ;
        RECT 24.465 44.545 25.675 45.065 ;
        RECT 26.050 45.185 26.380 45.985 ;
        RECT 26.550 45.355 26.880 46.155 ;
        RECT 27.180 45.185 27.510 45.985 ;
        RECT 28.155 45.355 28.405 46.155 ;
        RECT 26.050 45.015 28.485 45.185 ;
        RECT 28.675 45.015 28.845 46.155 ;
        RECT 29.015 45.015 29.355 45.985 ;
        RECT 29.525 45.720 34.870 46.155 ;
        RECT 25.845 44.595 26.195 44.845 ;
        RECT 26.380 44.385 26.550 45.015 ;
        RECT 26.720 44.595 27.050 44.795 ;
        RECT 27.220 44.595 27.550 44.795 ;
        RECT 27.720 44.595 28.140 44.795 ;
        RECT 28.315 44.765 28.485 45.015 ;
        RECT 28.315 44.595 29.010 44.765 ;
        RECT 23.085 43.605 25.675 44.375 ;
        RECT 26.050 43.775 26.550 44.385 ;
        RECT 27.180 44.255 28.405 44.425 ;
        RECT 29.180 44.405 29.355 45.015 ;
        RECT 27.180 43.775 27.510 44.255 ;
        RECT 27.680 43.605 27.905 44.065 ;
        RECT 28.075 43.775 28.405 44.255 ;
        RECT 28.595 43.605 28.845 44.405 ;
        RECT 29.015 43.775 29.355 44.405 ;
        RECT 31.110 44.150 31.450 44.980 ;
        RECT 32.930 44.470 33.280 45.720 ;
        RECT 35.050 45.485 35.305 45.985 ;
        RECT 35.475 45.655 35.805 46.155 ;
        RECT 35.050 45.315 35.800 45.485 ;
        RECT 35.050 44.495 35.400 45.145 ;
        RECT 35.570 44.325 35.800 45.315 ;
        RECT 35.050 44.155 35.800 44.325 ;
        RECT 29.525 43.605 34.870 44.150 ;
        RECT 35.050 43.865 35.305 44.155 ;
        RECT 35.475 43.605 35.805 43.985 ;
        RECT 35.975 43.865 36.145 45.985 ;
        RECT 36.315 45.185 36.640 45.970 ;
        RECT 36.810 45.695 37.060 46.155 ;
        RECT 37.230 45.655 37.480 45.985 ;
        RECT 37.695 45.655 38.375 45.985 ;
        RECT 37.230 45.525 37.400 45.655 ;
        RECT 37.005 45.355 37.400 45.525 ;
        RECT 36.375 44.135 36.835 45.185 ;
        RECT 37.005 43.995 37.175 45.355 ;
        RECT 37.570 45.095 38.035 45.485 ;
        RECT 37.345 44.285 37.695 44.905 ;
        RECT 37.865 44.505 38.035 45.095 ;
        RECT 38.205 44.875 38.375 45.655 ;
        RECT 38.545 45.555 38.715 45.895 ;
        RECT 38.950 45.725 39.280 46.155 ;
        RECT 39.450 45.555 39.620 45.895 ;
        RECT 39.915 45.695 40.285 46.155 ;
        RECT 38.545 45.385 39.620 45.555 ;
        RECT 40.455 45.525 40.625 45.985 ;
        RECT 40.860 45.645 41.730 45.985 ;
        RECT 41.900 45.695 42.150 46.155 ;
        RECT 40.065 45.355 40.625 45.525 ;
        RECT 40.065 45.215 40.235 45.355 ;
        RECT 38.735 45.045 40.235 45.215 ;
        RECT 40.930 45.185 41.390 45.475 ;
        RECT 38.205 44.705 39.895 44.875 ;
        RECT 37.865 44.285 38.220 44.505 ;
        RECT 38.390 43.995 38.560 44.705 ;
        RECT 38.765 44.285 39.555 44.535 ;
        RECT 39.725 44.525 39.895 44.705 ;
        RECT 40.065 44.355 40.235 45.045 ;
        RECT 36.505 43.605 36.835 43.965 ;
        RECT 37.005 43.825 37.500 43.995 ;
        RECT 37.705 43.825 38.560 43.995 ;
        RECT 39.435 43.605 39.765 44.065 ;
        RECT 39.975 43.965 40.235 44.355 ;
        RECT 40.425 45.175 41.390 45.185 ;
        RECT 41.560 45.265 41.730 45.645 ;
        RECT 42.320 45.605 42.490 45.895 ;
        RECT 42.670 45.775 43.000 46.155 ;
        RECT 42.320 45.435 43.120 45.605 ;
        RECT 40.425 45.015 41.100 45.175 ;
        RECT 41.560 45.095 42.780 45.265 ;
        RECT 40.425 44.225 40.635 45.015 ;
        RECT 41.560 45.005 41.730 45.095 ;
        RECT 40.805 44.225 41.155 44.845 ;
        RECT 41.325 44.835 41.730 45.005 ;
        RECT 41.325 44.055 41.495 44.835 ;
        RECT 41.665 44.385 41.885 44.665 ;
        RECT 42.065 44.555 42.605 44.925 ;
        RECT 42.950 44.845 43.120 45.435 ;
        RECT 43.340 45.015 43.645 46.155 ;
        RECT 43.815 44.965 44.070 45.845 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 44.765 45.015 44.975 46.155 ;
        RECT 45.145 45.005 45.475 45.985 ;
        RECT 45.645 45.015 45.875 46.155 ;
        RECT 46.085 45.065 47.295 46.155 ;
        RECT 42.950 44.815 43.690 44.845 ;
        RECT 41.665 44.215 42.195 44.385 ;
        RECT 39.975 43.795 40.325 43.965 ;
        RECT 40.545 43.775 41.495 44.055 ;
        RECT 41.665 43.605 41.855 44.045 ;
        RECT 42.025 43.985 42.195 44.215 ;
        RECT 42.365 44.155 42.605 44.555 ;
        RECT 42.775 44.515 43.690 44.815 ;
        RECT 42.775 44.340 43.100 44.515 ;
        RECT 42.775 43.985 43.095 44.340 ;
        RECT 43.860 44.315 44.070 44.965 ;
        RECT 42.025 43.815 43.095 43.985 ;
        RECT 43.340 43.605 43.645 44.065 ;
        RECT 43.815 43.785 44.070 44.315 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 44.765 43.605 44.975 44.425 ;
        RECT 45.145 44.405 45.395 45.005 ;
        RECT 45.565 44.595 45.895 44.845 ;
        RECT 45.145 43.775 45.475 44.405 ;
        RECT 45.645 43.605 45.875 44.425 ;
        RECT 46.085 44.355 46.605 44.895 ;
        RECT 46.775 44.525 47.295 45.065 ;
        RECT 47.615 45.005 47.945 46.155 ;
        RECT 48.115 45.135 48.285 45.985 ;
        RECT 48.455 45.355 48.785 46.155 ;
        RECT 48.955 45.135 49.125 45.985 ;
        RECT 49.305 45.355 49.545 46.155 ;
        RECT 49.715 45.175 50.045 45.985 ;
        RECT 48.115 44.965 49.125 45.135 ;
        RECT 49.330 45.005 50.045 45.175 ;
        RECT 50.225 45.065 52.815 46.155 ;
        RECT 52.990 45.485 53.245 45.985 ;
        RECT 53.415 45.655 53.745 46.155 ;
        RECT 52.990 45.315 53.740 45.485 ;
        RECT 48.115 44.455 48.610 44.965 ;
        RECT 49.330 44.765 49.500 45.005 ;
        RECT 49.000 44.595 49.500 44.765 ;
        RECT 49.670 44.595 50.050 44.835 ;
        RECT 48.115 44.425 48.615 44.455 ;
        RECT 49.330 44.425 49.500 44.595 ;
        RECT 46.085 43.605 47.295 44.355 ;
        RECT 47.615 43.605 47.945 44.405 ;
        RECT 48.115 44.255 49.125 44.425 ;
        RECT 49.330 44.255 49.965 44.425 ;
        RECT 48.115 43.775 48.285 44.255 ;
        RECT 48.455 43.605 48.785 44.085 ;
        RECT 48.955 43.775 49.125 44.255 ;
        RECT 49.375 43.605 49.615 44.085 ;
        RECT 49.795 43.775 49.965 44.255 ;
        RECT 50.225 44.375 51.435 44.895 ;
        RECT 51.605 44.545 52.815 45.065 ;
        RECT 52.990 44.495 53.340 45.145 ;
        RECT 50.225 43.605 52.815 44.375 ;
        RECT 53.510 44.325 53.740 45.315 ;
        RECT 52.990 44.155 53.740 44.325 ;
        RECT 52.990 43.865 53.245 44.155 ;
        RECT 53.415 43.605 53.745 43.985 ;
        RECT 53.915 43.865 54.085 45.985 ;
        RECT 54.255 45.185 54.580 45.970 ;
        RECT 54.750 45.695 55.000 46.155 ;
        RECT 55.170 45.655 55.420 45.985 ;
        RECT 55.635 45.655 56.315 45.985 ;
        RECT 55.170 45.525 55.340 45.655 ;
        RECT 54.945 45.355 55.340 45.525 ;
        RECT 54.315 44.135 54.775 45.185 ;
        RECT 54.945 43.995 55.115 45.355 ;
        RECT 55.510 45.095 55.975 45.485 ;
        RECT 55.285 44.285 55.635 44.905 ;
        RECT 55.805 44.505 55.975 45.095 ;
        RECT 56.145 44.875 56.315 45.655 ;
        RECT 56.485 45.555 56.655 45.895 ;
        RECT 56.890 45.725 57.220 46.155 ;
        RECT 57.390 45.555 57.560 45.895 ;
        RECT 57.855 45.695 58.225 46.155 ;
        RECT 56.485 45.385 57.560 45.555 ;
        RECT 58.395 45.525 58.565 45.985 ;
        RECT 58.800 45.645 59.670 45.985 ;
        RECT 59.840 45.695 60.090 46.155 ;
        RECT 58.005 45.355 58.565 45.525 ;
        RECT 58.005 45.215 58.175 45.355 ;
        RECT 56.675 45.045 58.175 45.215 ;
        RECT 58.870 45.185 59.330 45.475 ;
        RECT 56.145 44.705 57.835 44.875 ;
        RECT 55.805 44.285 56.160 44.505 ;
        RECT 56.330 43.995 56.500 44.705 ;
        RECT 56.705 44.285 57.495 44.535 ;
        RECT 57.665 44.525 57.835 44.705 ;
        RECT 58.005 44.355 58.175 45.045 ;
        RECT 54.445 43.605 54.775 43.965 ;
        RECT 54.945 43.825 55.440 43.995 ;
        RECT 55.645 43.825 56.500 43.995 ;
        RECT 57.375 43.605 57.705 44.065 ;
        RECT 57.915 43.965 58.175 44.355 ;
        RECT 58.365 45.175 59.330 45.185 ;
        RECT 59.500 45.265 59.670 45.645 ;
        RECT 60.260 45.605 60.430 45.895 ;
        RECT 60.610 45.775 60.940 46.155 ;
        RECT 60.260 45.435 61.060 45.605 ;
        RECT 58.365 45.015 59.040 45.175 ;
        RECT 59.500 45.095 60.720 45.265 ;
        RECT 58.365 44.225 58.575 45.015 ;
        RECT 59.500 45.005 59.670 45.095 ;
        RECT 58.745 44.225 59.095 44.845 ;
        RECT 59.265 44.835 59.670 45.005 ;
        RECT 59.265 44.055 59.435 44.835 ;
        RECT 59.605 44.385 59.825 44.665 ;
        RECT 60.005 44.555 60.545 44.925 ;
        RECT 60.890 44.845 61.060 45.435 ;
        RECT 61.280 45.015 61.585 46.155 ;
        RECT 61.755 44.965 62.010 45.845 ;
        RECT 60.890 44.815 61.630 44.845 ;
        RECT 59.605 44.215 60.135 44.385 ;
        RECT 57.915 43.795 58.265 43.965 ;
        RECT 58.485 43.775 59.435 44.055 ;
        RECT 59.605 43.605 59.795 44.045 ;
        RECT 59.965 43.985 60.135 44.215 ;
        RECT 60.305 44.155 60.545 44.555 ;
        RECT 60.715 44.515 61.630 44.815 ;
        RECT 60.715 44.340 61.040 44.515 ;
        RECT 60.715 43.985 61.035 44.340 ;
        RECT 61.800 44.315 62.010 44.965 ;
        RECT 59.965 43.815 61.035 43.985 ;
        RECT 61.280 43.605 61.585 44.065 ;
        RECT 61.755 43.785 62.010 44.315 ;
        RECT 62.185 45.655 62.445 45.985 ;
        RECT 62.755 45.775 63.085 46.155 ;
        RECT 62.185 44.975 62.355 45.655 ;
        RECT 63.325 45.605 63.515 45.985 ;
        RECT 63.765 45.775 64.095 46.155 ;
        RECT 64.305 45.605 64.475 45.985 ;
        RECT 64.670 45.775 65.000 46.155 ;
        RECT 65.260 45.605 65.430 45.985 ;
        RECT 65.855 45.775 66.185 46.155 ;
        RECT 62.525 45.145 62.875 45.475 ;
        RECT 63.325 45.435 64.065 45.605 ;
        RECT 63.145 45.095 63.725 45.265 ;
        RECT 63.145 44.975 63.315 45.095 ;
        RECT 62.185 44.805 63.315 44.975 ;
        RECT 63.895 44.925 64.065 45.435 ;
        RECT 62.185 44.105 62.355 44.805 ;
        RECT 63.495 44.755 64.065 44.925 ;
        RECT 64.235 45.435 66.185 45.605 ;
        RECT 62.705 44.465 63.325 44.635 ;
        RECT 62.705 44.285 62.915 44.465 ;
        RECT 63.495 44.275 63.665 44.755 ;
        RECT 64.235 44.445 64.405 45.435 ;
        RECT 64.995 44.845 65.180 45.155 ;
        RECT 65.450 44.845 65.645 45.155 ;
        RECT 62.185 43.775 62.445 44.105 ;
        RECT 62.755 43.605 63.085 43.985 ;
        RECT 63.265 43.945 63.665 44.275 ;
        RECT 63.855 44.115 64.405 44.445 ;
        RECT 64.575 43.945 64.745 44.845 ;
        RECT 63.265 43.775 64.745 43.945 ;
        RECT 64.995 44.515 65.225 44.845 ;
        RECT 65.450 44.515 65.705 44.845 ;
        RECT 66.015 44.515 66.185 45.435 ;
        RECT 64.995 43.935 65.180 44.515 ;
        RECT 65.450 43.940 65.645 44.515 ;
        RECT 65.855 43.605 66.185 43.985 ;
        RECT 66.355 43.775 66.615 45.985 ;
        RECT 66.875 45.225 67.045 45.985 ;
        RECT 67.260 45.395 67.590 46.155 ;
        RECT 66.875 45.055 67.590 45.225 ;
        RECT 67.760 45.080 68.015 45.985 ;
        RECT 66.785 44.505 67.140 44.875 ;
        RECT 67.420 44.845 67.590 45.055 ;
        RECT 67.420 44.515 67.675 44.845 ;
        RECT 67.420 44.325 67.590 44.515 ;
        RECT 67.845 44.350 68.015 45.080 ;
        RECT 68.190 45.005 68.450 46.155 ;
        RECT 68.625 45.065 69.835 46.155 ;
        RECT 66.875 44.155 67.590 44.325 ;
        RECT 66.875 43.775 67.045 44.155 ;
        RECT 67.260 43.605 67.590 43.985 ;
        RECT 67.760 43.775 68.015 44.350 ;
        RECT 68.190 43.605 68.450 44.445 ;
        RECT 68.625 44.355 69.145 44.895 ;
        RECT 69.315 44.525 69.835 45.065 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.465 45.720 75.810 46.155 ;
        RECT 68.625 43.605 69.835 44.355 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 72.050 44.150 72.390 44.980 ;
        RECT 73.870 44.470 74.220 45.720 ;
        RECT 75.985 45.065 78.575 46.155 ;
        RECT 75.985 44.375 77.195 44.895 ;
        RECT 77.365 44.545 78.575 45.065 ;
        RECT 78.745 45.080 79.015 45.985 ;
        RECT 79.185 45.395 79.515 46.155 ;
        RECT 79.695 45.225 79.865 45.985 ;
        RECT 70.465 43.605 75.810 44.150 ;
        RECT 75.985 43.605 78.575 44.375 ;
        RECT 78.745 44.280 78.915 45.080 ;
        RECT 79.200 45.055 79.865 45.225 ;
        RECT 79.200 44.910 79.370 45.055 ;
        RECT 80.645 45.015 80.855 46.155 ;
        RECT 79.085 44.580 79.370 44.910 ;
        RECT 81.025 45.005 81.355 45.985 ;
        RECT 81.525 45.015 81.755 46.155 ;
        RECT 81.965 45.720 87.310 46.155 ;
        RECT 79.200 44.325 79.370 44.580 ;
        RECT 79.605 44.505 79.935 44.875 ;
        RECT 78.745 43.775 79.005 44.280 ;
        RECT 79.200 44.155 79.865 44.325 ;
        RECT 79.185 43.605 79.515 43.985 ;
        RECT 79.695 43.775 79.865 44.155 ;
        RECT 80.645 43.605 80.855 44.425 ;
        RECT 81.025 44.405 81.275 45.005 ;
        RECT 81.445 44.595 81.775 44.845 ;
        RECT 81.025 43.775 81.355 44.405 ;
        RECT 81.525 43.605 81.755 44.425 ;
        RECT 83.550 44.150 83.890 44.980 ;
        RECT 85.370 44.470 85.720 45.720 ;
        RECT 87.485 45.065 89.155 46.155 ;
        RECT 87.485 44.375 88.235 44.895 ;
        RECT 88.405 44.545 89.155 45.065 ;
        RECT 89.415 45.225 89.585 45.985 ;
        RECT 89.765 45.395 90.095 46.155 ;
        RECT 89.415 45.055 90.080 45.225 ;
        RECT 90.265 45.080 90.535 45.985 ;
        RECT 89.910 44.910 90.080 45.055 ;
        RECT 89.345 44.505 89.675 44.875 ;
        RECT 89.910 44.580 90.195 44.910 ;
        RECT 81.965 43.605 87.310 44.150 ;
        RECT 87.485 43.605 89.155 44.375 ;
        RECT 89.910 44.325 90.080 44.580 ;
        RECT 89.415 44.155 90.080 44.325 ;
        RECT 90.365 44.280 90.535 45.080 ;
        RECT 89.415 43.775 89.585 44.155 ;
        RECT 89.765 43.605 90.095 43.985 ;
        RECT 90.275 43.775 90.535 44.280 ;
        RECT 90.710 45.015 91.045 45.985 ;
        RECT 91.215 45.015 91.385 46.155 ;
        RECT 91.555 45.815 93.585 45.985 ;
        RECT 90.710 44.345 90.880 45.015 ;
        RECT 91.555 44.845 91.725 45.815 ;
        RECT 91.050 44.515 91.305 44.845 ;
        RECT 91.530 44.515 91.725 44.845 ;
        RECT 91.895 45.475 93.020 45.645 ;
        RECT 91.135 44.345 91.305 44.515 ;
        RECT 91.895 44.345 92.065 45.475 ;
        RECT 90.710 43.775 90.965 44.345 ;
        RECT 91.135 44.175 92.065 44.345 ;
        RECT 92.235 45.135 93.245 45.305 ;
        RECT 92.235 44.335 92.405 45.135 ;
        RECT 92.610 44.795 92.885 44.935 ;
        RECT 92.605 44.625 92.885 44.795 ;
        RECT 91.890 44.140 92.065 44.175 ;
        RECT 91.135 43.605 91.465 44.005 ;
        RECT 91.890 43.775 92.420 44.140 ;
        RECT 92.610 43.775 92.885 44.625 ;
        RECT 93.055 43.775 93.245 45.135 ;
        RECT 93.415 45.150 93.585 45.815 ;
        RECT 93.755 45.395 93.925 46.155 ;
        RECT 94.160 45.395 94.675 45.805 ;
        RECT 93.415 44.960 94.165 45.150 ;
        RECT 94.335 44.585 94.675 45.395 ;
        RECT 95.765 44.990 96.055 46.155 ;
        RECT 96.225 45.720 101.570 46.155 ;
        RECT 93.445 44.415 94.675 44.585 ;
        RECT 93.425 43.605 93.935 44.140 ;
        RECT 94.155 43.810 94.400 44.415 ;
        RECT 95.765 43.605 96.055 44.330 ;
        RECT 97.810 44.150 98.150 44.980 ;
        RECT 99.630 44.470 99.980 45.720 ;
        RECT 102.210 45.485 102.465 45.985 ;
        RECT 102.635 45.655 102.965 46.155 ;
        RECT 102.210 45.315 102.960 45.485 ;
        RECT 102.210 44.495 102.560 45.145 ;
        RECT 102.730 44.325 102.960 45.315 ;
        RECT 102.210 44.155 102.960 44.325 ;
        RECT 96.225 43.605 101.570 44.150 ;
        RECT 102.210 43.865 102.465 44.155 ;
        RECT 102.635 43.605 102.965 43.985 ;
        RECT 103.135 43.865 103.305 45.985 ;
        RECT 103.475 45.185 103.800 45.970 ;
        RECT 103.970 45.695 104.220 46.155 ;
        RECT 104.390 45.655 104.640 45.985 ;
        RECT 104.855 45.655 105.535 45.985 ;
        RECT 104.390 45.525 104.560 45.655 ;
        RECT 104.165 45.355 104.560 45.525 ;
        RECT 103.535 44.135 103.995 45.185 ;
        RECT 104.165 43.995 104.335 45.355 ;
        RECT 104.730 45.095 105.195 45.485 ;
        RECT 104.505 44.285 104.855 44.905 ;
        RECT 105.025 44.505 105.195 45.095 ;
        RECT 105.365 44.875 105.535 45.655 ;
        RECT 105.705 45.555 105.875 45.895 ;
        RECT 106.110 45.725 106.440 46.155 ;
        RECT 106.610 45.555 106.780 45.895 ;
        RECT 107.075 45.695 107.445 46.155 ;
        RECT 105.705 45.385 106.780 45.555 ;
        RECT 107.615 45.525 107.785 45.985 ;
        RECT 108.020 45.645 108.890 45.985 ;
        RECT 109.060 45.695 109.310 46.155 ;
        RECT 107.225 45.355 107.785 45.525 ;
        RECT 107.225 45.215 107.395 45.355 ;
        RECT 105.895 45.045 107.395 45.215 ;
        RECT 108.090 45.185 108.550 45.475 ;
        RECT 105.365 44.705 107.055 44.875 ;
        RECT 105.025 44.285 105.380 44.505 ;
        RECT 105.550 43.995 105.720 44.705 ;
        RECT 105.925 44.285 106.715 44.535 ;
        RECT 106.885 44.525 107.055 44.705 ;
        RECT 107.225 44.355 107.395 45.045 ;
        RECT 103.665 43.605 103.995 43.965 ;
        RECT 104.165 43.825 104.660 43.995 ;
        RECT 104.865 43.825 105.720 43.995 ;
        RECT 106.595 43.605 106.925 44.065 ;
        RECT 107.135 43.965 107.395 44.355 ;
        RECT 107.585 45.175 108.550 45.185 ;
        RECT 108.720 45.265 108.890 45.645 ;
        RECT 109.480 45.605 109.650 45.895 ;
        RECT 109.830 45.775 110.160 46.155 ;
        RECT 109.480 45.435 110.280 45.605 ;
        RECT 107.585 45.015 108.260 45.175 ;
        RECT 108.720 45.095 109.940 45.265 ;
        RECT 107.585 44.225 107.795 45.015 ;
        RECT 108.720 45.005 108.890 45.095 ;
        RECT 107.965 44.225 108.315 44.845 ;
        RECT 108.485 44.835 108.890 45.005 ;
        RECT 108.485 44.055 108.655 44.835 ;
        RECT 108.825 44.385 109.045 44.665 ;
        RECT 109.225 44.555 109.765 44.925 ;
        RECT 110.110 44.845 110.280 45.435 ;
        RECT 110.500 45.015 110.805 46.155 ;
        RECT 110.975 44.965 111.230 45.845 ;
        RECT 111.405 45.720 116.750 46.155 ;
        RECT 110.110 44.815 110.850 44.845 ;
        RECT 108.825 44.215 109.355 44.385 ;
        RECT 107.135 43.795 107.485 43.965 ;
        RECT 107.705 43.775 108.655 44.055 ;
        RECT 108.825 43.605 109.015 44.045 ;
        RECT 109.185 43.985 109.355 44.215 ;
        RECT 109.525 44.155 109.765 44.555 ;
        RECT 109.935 44.515 110.850 44.815 ;
        RECT 109.935 44.340 110.260 44.515 ;
        RECT 109.935 43.985 110.255 44.340 ;
        RECT 111.020 44.315 111.230 44.965 ;
        RECT 109.185 43.815 110.255 43.985 ;
        RECT 110.500 43.605 110.805 44.065 ;
        RECT 110.975 43.785 111.230 44.315 ;
        RECT 112.990 44.150 113.330 44.980 ;
        RECT 114.810 44.470 115.160 45.720 ;
        RECT 116.925 45.065 120.435 46.155 ;
        RECT 116.925 44.375 118.575 44.895 ;
        RECT 118.745 44.545 120.435 45.065 ;
        RECT 121.525 44.990 121.815 46.155 ;
        RECT 122.445 45.065 123.655 46.155 ;
        RECT 122.445 44.525 122.965 45.065 ;
        RECT 111.405 43.605 116.750 44.150 ;
        RECT 116.925 43.605 120.435 44.375 ;
        RECT 123.135 44.355 123.655 44.895 ;
        RECT 121.525 43.605 121.815 44.330 ;
        RECT 122.445 43.605 123.655 44.355 ;
        RECT 5.520 43.435 123.740 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.985 42.665 8.655 43.435 ;
        RECT 8.830 42.885 9.085 43.175 ;
        RECT 9.255 43.055 9.585 43.435 ;
        RECT 8.830 42.715 9.580 42.885 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 6.985 42.145 7.735 42.665 ;
        RECT 7.905 41.975 8.655 42.495 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 6.985 40.885 8.655 41.975 ;
        RECT 8.830 41.895 9.180 42.545 ;
        RECT 9.350 41.725 9.580 42.715 ;
        RECT 8.830 41.555 9.580 41.725 ;
        RECT 8.830 41.055 9.085 41.555 ;
        RECT 9.255 40.885 9.585 41.385 ;
        RECT 9.755 41.055 9.925 43.175 ;
        RECT 10.285 43.075 10.615 43.435 ;
        RECT 10.785 43.045 11.280 43.215 ;
        RECT 11.485 43.045 12.340 43.215 ;
        RECT 10.155 41.855 10.615 42.905 ;
        RECT 10.095 41.070 10.420 41.855 ;
        RECT 10.785 41.685 10.955 43.045 ;
        RECT 11.125 42.135 11.475 42.755 ;
        RECT 11.645 42.535 12.000 42.755 ;
        RECT 11.645 41.945 11.815 42.535 ;
        RECT 12.170 42.335 12.340 43.045 ;
        RECT 13.215 42.975 13.545 43.435 ;
        RECT 13.755 43.075 14.105 43.245 ;
        RECT 12.545 42.505 13.335 42.755 ;
        RECT 13.755 42.685 14.015 43.075 ;
        RECT 14.325 42.985 15.275 43.265 ;
        RECT 15.445 42.995 15.635 43.435 ;
        RECT 15.805 43.055 16.875 43.225 ;
        RECT 13.505 42.335 13.675 42.515 ;
        RECT 10.785 41.515 11.180 41.685 ;
        RECT 11.350 41.555 11.815 41.945 ;
        RECT 11.985 42.165 13.675 42.335 ;
        RECT 11.010 41.385 11.180 41.515 ;
        RECT 11.985 41.385 12.155 42.165 ;
        RECT 13.845 41.995 14.015 42.685 ;
        RECT 12.515 41.825 14.015 41.995 ;
        RECT 14.205 42.025 14.415 42.815 ;
        RECT 14.585 42.195 14.935 42.815 ;
        RECT 15.105 42.205 15.275 42.985 ;
        RECT 15.805 42.825 15.975 43.055 ;
        RECT 15.445 42.655 15.975 42.825 ;
        RECT 15.445 42.375 15.665 42.655 ;
        RECT 16.145 42.485 16.385 42.885 ;
        RECT 15.105 42.035 15.510 42.205 ;
        RECT 15.845 42.115 16.385 42.485 ;
        RECT 16.555 42.700 16.875 43.055 ;
        RECT 17.120 42.975 17.425 43.435 ;
        RECT 17.595 42.725 17.850 43.255 ;
        RECT 16.555 42.525 16.880 42.700 ;
        RECT 16.555 42.225 17.470 42.525 ;
        RECT 16.730 42.195 17.470 42.225 ;
        RECT 14.205 41.865 14.880 42.025 ;
        RECT 15.340 41.945 15.510 42.035 ;
        RECT 14.205 41.855 15.170 41.865 ;
        RECT 13.845 41.685 14.015 41.825 ;
        RECT 10.590 40.885 10.840 41.345 ;
        RECT 11.010 41.055 11.260 41.385 ;
        RECT 11.475 41.055 12.155 41.385 ;
        RECT 12.325 41.485 13.400 41.655 ;
        RECT 13.845 41.515 14.405 41.685 ;
        RECT 14.710 41.565 15.170 41.855 ;
        RECT 15.340 41.775 16.560 41.945 ;
        RECT 12.325 41.145 12.495 41.485 ;
        RECT 12.730 40.885 13.060 41.315 ;
        RECT 13.230 41.145 13.400 41.485 ;
        RECT 13.695 40.885 14.065 41.345 ;
        RECT 14.235 41.055 14.405 41.515 ;
        RECT 15.340 41.395 15.510 41.775 ;
        RECT 16.730 41.605 16.900 42.195 ;
        RECT 17.640 42.075 17.850 42.725 ;
        RECT 18.085 42.615 18.295 43.435 ;
        RECT 18.465 42.635 18.795 43.265 ;
        RECT 14.640 41.055 15.510 41.395 ;
        RECT 16.100 41.435 16.900 41.605 ;
        RECT 15.680 40.885 15.930 41.345 ;
        RECT 16.100 41.145 16.270 41.435 ;
        RECT 16.450 40.885 16.780 41.265 ;
        RECT 17.120 40.885 17.425 42.025 ;
        RECT 17.595 41.195 17.850 42.075 ;
        RECT 18.465 42.035 18.715 42.635 ;
        RECT 18.965 42.615 19.195 43.435 ;
        RECT 19.405 42.890 24.750 43.435 ;
        RECT 18.885 42.195 19.215 42.445 ;
        RECT 20.990 42.060 21.330 42.890 ;
        RECT 25.015 42.885 25.185 43.265 ;
        RECT 25.365 43.055 25.695 43.435 ;
        RECT 25.015 42.715 25.680 42.885 ;
        RECT 25.875 42.760 26.135 43.265 ;
        RECT 18.085 40.885 18.295 42.025 ;
        RECT 18.465 41.055 18.795 42.035 ;
        RECT 18.965 40.885 19.195 42.025 ;
        RECT 22.810 41.320 23.160 42.570 ;
        RECT 24.945 42.165 25.275 42.535 ;
        RECT 25.510 42.460 25.680 42.715 ;
        RECT 25.510 42.130 25.795 42.460 ;
        RECT 25.510 41.985 25.680 42.130 ;
        RECT 25.015 41.815 25.680 41.985 ;
        RECT 25.965 41.960 26.135 42.760 ;
        RECT 19.405 40.885 24.750 41.320 ;
        RECT 25.015 41.055 25.185 41.815 ;
        RECT 25.365 40.885 25.695 41.645 ;
        RECT 25.865 41.055 26.135 41.960 ;
        RECT 26.310 42.695 26.565 43.265 ;
        RECT 26.735 43.035 27.065 43.435 ;
        RECT 27.490 42.900 28.020 43.265 ;
        RECT 28.210 43.095 28.485 43.265 ;
        RECT 28.205 42.925 28.485 43.095 ;
        RECT 27.490 42.865 27.665 42.900 ;
        RECT 26.735 42.695 27.665 42.865 ;
        RECT 26.310 42.025 26.480 42.695 ;
        RECT 26.735 42.525 26.905 42.695 ;
        RECT 26.650 42.195 26.905 42.525 ;
        RECT 27.130 42.195 27.325 42.525 ;
        RECT 26.310 41.055 26.645 42.025 ;
        RECT 26.815 40.885 26.985 42.025 ;
        RECT 27.155 41.225 27.325 42.195 ;
        RECT 27.495 41.565 27.665 42.695 ;
        RECT 27.835 41.905 28.005 42.705 ;
        RECT 28.210 42.105 28.485 42.925 ;
        RECT 28.655 41.905 28.845 43.265 ;
        RECT 29.025 42.900 29.535 43.435 ;
        RECT 29.755 42.625 30.000 43.230 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.825 42.665 35.335 43.435 ;
        RECT 36.430 42.695 36.685 43.265 ;
        RECT 36.855 43.035 37.185 43.435 ;
        RECT 37.610 42.900 38.140 43.265 ;
        RECT 37.610 42.865 37.785 42.900 ;
        RECT 36.855 42.695 37.785 42.865 ;
        RECT 38.330 42.755 38.605 43.265 ;
        RECT 29.045 42.455 30.275 42.625 ;
        RECT 27.835 41.735 28.845 41.905 ;
        RECT 29.015 41.890 29.765 42.080 ;
        RECT 27.495 41.395 28.620 41.565 ;
        RECT 29.015 41.225 29.185 41.890 ;
        RECT 29.935 41.645 30.275 42.455 ;
        RECT 31.825 42.145 33.475 42.665 ;
        RECT 27.155 41.055 29.185 41.225 ;
        RECT 29.355 40.885 29.525 41.645 ;
        RECT 29.760 41.235 30.275 41.645 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 33.645 41.975 35.335 42.495 ;
        RECT 31.825 40.885 35.335 41.975 ;
        RECT 36.430 42.025 36.600 42.695 ;
        RECT 36.855 42.525 37.025 42.695 ;
        RECT 36.770 42.195 37.025 42.525 ;
        RECT 37.250 42.195 37.445 42.525 ;
        RECT 36.430 41.055 36.765 42.025 ;
        RECT 36.935 40.885 37.105 42.025 ;
        RECT 37.275 41.225 37.445 42.195 ;
        RECT 37.615 41.565 37.785 42.695 ;
        RECT 37.955 41.905 38.125 42.705 ;
        RECT 38.325 42.585 38.605 42.755 ;
        RECT 38.330 42.105 38.605 42.585 ;
        RECT 38.775 41.905 38.965 43.265 ;
        RECT 39.145 42.900 39.655 43.435 ;
        RECT 39.875 42.625 40.120 43.230 ;
        RECT 41.490 42.695 41.745 43.265 ;
        RECT 41.915 43.035 42.245 43.435 ;
        RECT 42.670 42.900 43.200 43.265 ;
        RECT 42.670 42.865 42.845 42.900 ;
        RECT 41.915 42.695 42.845 42.865 ;
        RECT 43.390 42.755 43.665 43.265 ;
        RECT 39.165 42.455 40.395 42.625 ;
        RECT 37.955 41.735 38.965 41.905 ;
        RECT 39.135 41.890 39.885 42.080 ;
        RECT 37.615 41.395 38.740 41.565 ;
        RECT 39.135 41.225 39.305 41.890 ;
        RECT 40.055 41.645 40.395 42.455 ;
        RECT 37.275 41.055 39.305 41.225 ;
        RECT 39.475 40.885 39.645 41.645 ;
        RECT 39.880 41.235 40.395 41.645 ;
        RECT 41.490 42.025 41.660 42.695 ;
        RECT 41.915 42.525 42.085 42.695 ;
        RECT 41.830 42.195 42.085 42.525 ;
        RECT 42.310 42.195 42.505 42.525 ;
        RECT 41.490 41.055 41.825 42.025 ;
        RECT 41.995 40.885 42.165 42.025 ;
        RECT 42.335 41.225 42.505 42.195 ;
        RECT 42.675 41.565 42.845 42.695 ;
        RECT 43.015 41.905 43.185 42.705 ;
        RECT 43.385 42.585 43.665 42.755 ;
        RECT 43.390 42.105 43.665 42.585 ;
        RECT 43.835 41.905 44.025 43.265 ;
        RECT 44.205 42.900 44.715 43.435 ;
        RECT 44.935 42.625 45.180 43.230 ;
        RECT 45.625 42.890 50.970 43.435 ;
        RECT 51.145 42.890 56.490 43.435 ;
        RECT 44.225 42.455 45.455 42.625 ;
        RECT 43.015 41.735 44.025 41.905 ;
        RECT 44.195 41.890 44.945 42.080 ;
        RECT 42.675 41.395 43.800 41.565 ;
        RECT 44.195 41.225 44.365 41.890 ;
        RECT 45.115 41.645 45.455 42.455 ;
        RECT 47.210 42.060 47.550 42.890 ;
        RECT 42.335 41.055 44.365 41.225 ;
        RECT 44.535 40.885 44.705 41.645 ;
        RECT 44.940 41.235 45.455 41.645 ;
        RECT 49.030 41.320 49.380 42.570 ;
        RECT 52.730 42.060 53.070 42.890 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 58.565 42.615 58.775 43.435 ;
        RECT 58.945 42.635 59.275 43.265 ;
        RECT 54.550 41.320 54.900 42.570 ;
        RECT 45.625 40.885 50.970 41.320 ;
        RECT 51.145 40.885 56.490 41.320 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 58.945 42.035 59.195 42.635 ;
        RECT 59.445 42.615 59.675 43.435 ;
        RECT 59.885 42.685 61.095 43.435 ;
        RECT 61.350 42.865 61.525 43.265 ;
        RECT 61.695 43.055 62.025 43.435 ;
        RECT 62.270 42.935 62.500 43.265 ;
        RECT 61.350 42.695 61.980 42.865 ;
        RECT 59.365 42.195 59.695 42.445 ;
        RECT 59.885 42.145 60.405 42.685 ;
        RECT 61.810 42.525 61.980 42.695 ;
        RECT 58.565 40.885 58.775 42.025 ;
        RECT 58.945 41.055 59.275 42.035 ;
        RECT 59.445 40.885 59.675 42.025 ;
        RECT 60.575 41.975 61.095 42.515 ;
        RECT 59.885 40.885 61.095 41.975 ;
        RECT 61.265 41.845 61.630 42.525 ;
        RECT 61.810 42.195 62.160 42.525 ;
        RECT 61.810 41.675 61.980 42.195 ;
        RECT 61.350 41.505 61.980 41.675 ;
        RECT 62.330 41.645 62.500 42.935 ;
        RECT 62.700 41.825 62.980 43.100 ;
        RECT 63.205 43.095 63.475 43.100 ;
        RECT 63.165 42.925 63.475 43.095 ;
        RECT 63.935 43.055 64.265 43.435 ;
        RECT 64.435 43.180 64.770 43.225 ;
        RECT 63.205 41.825 63.475 42.925 ;
        RECT 63.665 41.825 64.005 42.855 ;
        RECT 64.435 42.715 64.775 43.180 ;
        RECT 64.175 42.195 64.435 42.525 ;
        RECT 64.175 41.645 64.345 42.195 ;
        RECT 64.605 42.025 64.775 42.715 ;
        RECT 61.350 41.055 61.525 41.505 ;
        RECT 62.330 41.475 64.345 41.645 ;
        RECT 61.695 40.885 62.025 41.325 ;
        RECT 62.330 41.055 62.500 41.475 ;
        RECT 62.735 40.885 63.405 41.295 ;
        RECT 63.620 41.055 63.790 41.475 ;
        RECT 63.990 40.885 64.320 41.295 ;
        RECT 64.515 41.055 64.775 42.025 ;
        RECT 64.945 42.935 65.205 43.265 ;
        RECT 65.415 42.955 65.690 43.435 ;
        RECT 64.945 42.025 65.115 42.935 ;
        RECT 65.900 42.865 66.105 43.265 ;
        RECT 66.275 43.035 66.610 43.435 ;
        RECT 66.785 42.890 72.130 43.435 ;
        RECT 65.285 42.195 65.645 42.775 ;
        RECT 65.900 42.695 66.585 42.865 ;
        RECT 65.825 42.025 66.075 42.525 ;
        RECT 64.945 41.855 66.075 42.025 ;
        RECT 64.945 41.085 65.215 41.855 ;
        RECT 66.245 41.665 66.585 42.695 ;
        RECT 68.370 42.060 68.710 42.890 ;
        RECT 72.305 42.685 73.515 43.435 ;
        RECT 73.690 42.885 73.945 43.175 ;
        RECT 74.115 43.055 74.445 43.435 ;
        RECT 73.690 42.715 74.440 42.885 ;
        RECT 65.385 40.885 65.715 41.665 ;
        RECT 65.920 41.490 66.585 41.665 ;
        RECT 65.920 41.085 66.105 41.490 ;
        RECT 70.190 41.320 70.540 42.570 ;
        RECT 72.305 42.145 72.825 42.685 ;
        RECT 72.995 41.975 73.515 42.515 ;
        RECT 66.275 40.885 66.610 41.310 ;
        RECT 66.785 40.885 72.130 41.320 ;
        RECT 72.305 40.885 73.515 41.975 ;
        RECT 73.690 41.895 74.040 42.545 ;
        RECT 74.210 41.725 74.440 42.715 ;
        RECT 73.690 41.555 74.440 41.725 ;
        RECT 73.690 41.055 73.945 41.555 ;
        RECT 74.115 40.885 74.445 41.385 ;
        RECT 74.615 41.055 74.785 43.175 ;
        RECT 75.145 43.075 75.475 43.435 ;
        RECT 75.645 43.045 76.140 43.215 ;
        RECT 76.345 43.045 77.200 43.215 ;
        RECT 75.015 41.855 75.475 42.905 ;
        RECT 74.955 41.070 75.280 41.855 ;
        RECT 75.645 41.685 75.815 43.045 ;
        RECT 75.985 42.135 76.335 42.755 ;
        RECT 76.505 42.535 76.860 42.755 ;
        RECT 76.505 41.945 76.675 42.535 ;
        RECT 77.030 42.335 77.200 43.045 ;
        RECT 78.075 42.975 78.405 43.435 ;
        RECT 78.615 43.075 78.965 43.245 ;
        RECT 77.405 42.505 78.195 42.755 ;
        RECT 78.615 42.685 78.875 43.075 ;
        RECT 79.185 42.985 80.135 43.265 ;
        RECT 80.305 42.995 80.495 43.435 ;
        RECT 80.665 43.055 81.735 43.225 ;
        RECT 78.365 42.335 78.535 42.515 ;
        RECT 75.645 41.515 76.040 41.685 ;
        RECT 76.210 41.555 76.675 41.945 ;
        RECT 76.845 42.165 78.535 42.335 ;
        RECT 75.870 41.385 76.040 41.515 ;
        RECT 76.845 41.385 77.015 42.165 ;
        RECT 78.705 41.995 78.875 42.685 ;
        RECT 77.375 41.825 78.875 41.995 ;
        RECT 79.065 42.025 79.275 42.815 ;
        RECT 79.445 42.195 79.795 42.815 ;
        RECT 79.965 42.205 80.135 42.985 ;
        RECT 80.665 42.825 80.835 43.055 ;
        RECT 80.305 42.655 80.835 42.825 ;
        RECT 80.305 42.375 80.525 42.655 ;
        RECT 81.005 42.485 81.245 42.885 ;
        RECT 79.965 42.035 80.370 42.205 ;
        RECT 80.705 42.115 81.245 42.485 ;
        RECT 81.415 42.700 81.735 43.055 ;
        RECT 81.980 42.975 82.285 43.435 ;
        RECT 82.455 42.725 82.710 43.255 ;
        RECT 81.415 42.525 81.740 42.700 ;
        RECT 81.415 42.225 82.330 42.525 ;
        RECT 81.590 42.195 82.330 42.225 ;
        RECT 79.065 41.865 79.740 42.025 ;
        RECT 80.200 41.945 80.370 42.035 ;
        RECT 79.065 41.855 80.030 41.865 ;
        RECT 78.705 41.685 78.875 41.825 ;
        RECT 75.450 40.885 75.700 41.345 ;
        RECT 75.870 41.055 76.120 41.385 ;
        RECT 76.335 41.055 77.015 41.385 ;
        RECT 77.185 41.485 78.260 41.655 ;
        RECT 78.705 41.515 79.265 41.685 ;
        RECT 79.570 41.565 80.030 41.855 ;
        RECT 80.200 41.775 81.420 41.945 ;
        RECT 77.185 41.145 77.355 41.485 ;
        RECT 77.590 40.885 77.920 41.315 ;
        RECT 78.090 41.145 78.260 41.485 ;
        RECT 78.555 40.885 78.925 41.345 ;
        RECT 79.095 41.055 79.265 41.515 ;
        RECT 80.200 41.395 80.370 41.775 ;
        RECT 81.590 41.605 81.760 42.195 ;
        RECT 82.500 42.075 82.710 42.725 ;
        RECT 82.885 42.710 83.175 43.435 ;
        RECT 79.500 41.055 80.370 41.395 ;
        RECT 80.960 41.435 81.760 41.605 ;
        RECT 80.540 40.885 80.790 41.345 ;
        RECT 80.960 41.145 81.130 41.435 ;
        RECT 81.310 40.885 81.640 41.265 ;
        RECT 81.980 40.885 82.285 42.025 ;
        RECT 82.455 41.195 82.710 42.075 ;
        RECT 84.270 42.695 84.525 43.265 ;
        RECT 84.695 43.035 85.025 43.435 ;
        RECT 85.450 42.900 85.980 43.265 ;
        RECT 86.170 43.095 86.445 43.265 ;
        RECT 86.165 42.925 86.445 43.095 ;
        RECT 85.450 42.865 85.625 42.900 ;
        RECT 84.695 42.695 85.625 42.865 ;
        RECT 82.885 40.885 83.175 42.050 ;
        RECT 84.270 42.025 84.440 42.695 ;
        RECT 84.695 42.525 84.865 42.695 ;
        RECT 84.610 42.195 84.865 42.525 ;
        RECT 85.090 42.195 85.285 42.525 ;
        RECT 84.270 41.055 84.605 42.025 ;
        RECT 84.775 40.885 84.945 42.025 ;
        RECT 85.115 41.225 85.285 42.195 ;
        RECT 85.455 41.565 85.625 42.695 ;
        RECT 85.795 41.905 85.965 42.705 ;
        RECT 86.170 42.105 86.445 42.925 ;
        RECT 86.615 41.905 86.805 43.265 ;
        RECT 86.985 42.900 87.495 43.435 ;
        RECT 87.715 42.625 87.960 43.230 ;
        RECT 88.405 42.665 90.075 43.435 ;
        RECT 90.710 42.885 90.965 43.175 ;
        RECT 91.135 43.055 91.465 43.435 ;
        RECT 90.710 42.715 91.460 42.885 ;
        RECT 87.005 42.455 88.235 42.625 ;
        RECT 85.795 41.735 86.805 41.905 ;
        RECT 86.975 41.890 87.725 42.080 ;
        RECT 85.455 41.395 86.580 41.565 ;
        RECT 86.975 41.225 87.145 41.890 ;
        RECT 87.895 41.645 88.235 42.455 ;
        RECT 88.405 42.145 89.155 42.665 ;
        RECT 89.325 41.975 90.075 42.495 ;
        RECT 85.115 41.055 87.145 41.225 ;
        RECT 87.315 40.885 87.485 41.645 ;
        RECT 87.720 41.235 88.235 41.645 ;
        RECT 88.405 40.885 90.075 41.975 ;
        RECT 90.710 41.895 91.060 42.545 ;
        RECT 91.230 41.725 91.460 42.715 ;
        RECT 90.710 41.555 91.460 41.725 ;
        RECT 90.710 41.055 90.965 41.555 ;
        RECT 91.135 40.885 91.465 41.385 ;
        RECT 91.635 41.055 91.805 43.175 ;
        RECT 92.165 43.075 92.495 43.435 ;
        RECT 92.665 43.045 93.160 43.215 ;
        RECT 93.365 43.045 94.220 43.215 ;
        RECT 92.035 41.855 92.495 42.905 ;
        RECT 91.975 41.070 92.300 41.855 ;
        RECT 92.665 41.685 92.835 43.045 ;
        RECT 93.005 42.135 93.355 42.755 ;
        RECT 93.525 42.535 93.880 42.755 ;
        RECT 93.525 41.945 93.695 42.535 ;
        RECT 94.050 42.335 94.220 43.045 ;
        RECT 95.095 42.975 95.425 43.435 ;
        RECT 95.635 43.075 95.985 43.245 ;
        RECT 94.425 42.505 95.215 42.755 ;
        RECT 95.635 42.685 95.895 43.075 ;
        RECT 96.205 42.985 97.155 43.265 ;
        RECT 97.325 42.995 97.515 43.435 ;
        RECT 97.685 43.055 98.755 43.225 ;
        RECT 95.385 42.335 95.555 42.515 ;
        RECT 92.665 41.515 93.060 41.685 ;
        RECT 93.230 41.555 93.695 41.945 ;
        RECT 93.865 42.165 95.555 42.335 ;
        RECT 92.890 41.385 93.060 41.515 ;
        RECT 93.865 41.385 94.035 42.165 ;
        RECT 95.725 41.995 95.895 42.685 ;
        RECT 94.395 41.825 95.895 41.995 ;
        RECT 96.085 42.025 96.295 42.815 ;
        RECT 96.465 42.195 96.815 42.815 ;
        RECT 96.985 42.205 97.155 42.985 ;
        RECT 97.685 42.825 97.855 43.055 ;
        RECT 97.325 42.655 97.855 42.825 ;
        RECT 97.325 42.375 97.545 42.655 ;
        RECT 98.025 42.485 98.265 42.885 ;
        RECT 96.985 42.035 97.390 42.205 ;
        RECT 97.725 42.115 98.265 42.485 ;
        RECT 98.435 42.700 98.755 43.055 ;
        RECT 99.000 42.975 99.305 43.435 ;
        RECT 99.475 42.725 99.730 43.255 ;
        RECT 98.435 42.525 98.760 42.700 ;
        RECT 98.435 42.225 99.350 42.525 ;
        RECT 98.610 42.195 99.350 42.225 ;
        RECT 96.085 41.865 96.760 42.025 ;
        RECT 97.220 41.945 97.390 42.035 ;
        RECT 96.085 41.855 97.050 41.865 ;
        RECT 95.725 41.685 95.895 41.825 ;
        RECT 92.470 40.885 92.720 41.345 ;
        RECT 92.890 41.055 93.140 41.385 ;
        RECT 93.355 41.055 94.035 41.385 ;
        RECT 94.205 41.485 95.280 41.655 ;
        RECT 95.725 41.515 96.285 41.685 ;
        RECT 96.590 41.565 97.050 41.855 ;
        RECT 97.220 41.775 98.440 41.945 ;
        RECT 94.205 41.145 94.375 41.485 ;
        RECT 94.610 40.885 94.940 41.315 ;
        RECT 95.110 41.145 95.280 41.485 ;
        RECT 95.575 40.885 95.945 41.345 ;
        RECT 96.115 41.055 96.285 41.515 ;
        RECT 97.220 41.395 97.390 41.775 ;
        RECT 98.610 41.605 98.780 42.195 ;
        RECT 99.520 42.075 99.730 42.725 ;
        RECT 99.905 42.665 103.415 43.435 ;
        RECT 99.905 42.145 101.555 42.665 ;
        RECT 104.780 42.625 105.025 43.230 ;
        RECT 105.245 42.900 105.755 43.435 ;
        RECT 96.520 41.055 97.390 41.395 ;
        RECT 97.980 41.435 98.780 41.605 ;
        RECT 97.560 40.885 97.810 41.345 ;
        RECT 97.980 41.145 98.150 41.435 ;
        RECT 98.330 40.885 98.660 41.265 ;
        RECT 99.000 40.885 99.305 42.025 ;
        RECT 99.475 41.195 99.730 42.075 ;
        RECT 101.725 41.975 103.415 42.495 ;
        RECT 99.905 40.885 103.415 41.975 ;
        RECT 104.505 42.455 105.735 42.625 ;
        RECT 104.505 41.645 104.845 42.455 ;
        RECT 105.015 41.890 105.765 42.080 ;
        RECT 104.505 41.235 105.020 41.645 ;
        RECT 105.255 40.885 105.425 41.645 ;
        RECT 105.595 41.225 105.765 41.890 ;
        RECT 105.935 41.905 106.125 43.265 ;
        RECT 106.295 42.415 106.570 43.265 ;
        RECT 106.760 42.900 107.290 43.265 ;
        RECT 107.715 43.035 108.045 43.435 ;
        RECT 107.115 42.865 107.290 42.900 ;
        RECT 106.295 42.245 106.575 42.415 ;
        RECT 106.295 42.105 106.570 42.245 ;
        RECT 106.775 41.905 106.945 42.705 ;
        RECT 105.935 41.735 106.945 41.905 ;
        RECT 107.115 42.695 108.045 42.865 ;
        RECT 108.215 42.695 108.470 43.265 ;
        RECT 108.645 42.710 108.935 43.435 ;
        RECT 109.110 42.885 109.365 43.175 ;
        RECT 109.535 43.055 109.865 43.435 ;
        RECT 109.110 42.715 109.860 42.885 ;
        RECT 107.115 41.565 107.285 42.695 ;
        RECT 107.875 42.525 108.045 42.695 ;
        RECT 106.160 41.395 107.285 41.565 ;
        RECT 107.455 42.195 107.650 42.525 ;
        RECT 107.875 42.195 108.130 42.525 ;
        RECT 107.455 41.225 107.625 42.195 ;
        RECT 108.300 42.025 108.470 42.695 ;
        RECT 105.595 41.055 107.625 41.225 ;
        RECT 107.795 40.885 107.965 42.025 ;
        RECT 108.135 41.055 108.470 42.025 ;
        RECT 108.645 40.885 108.935 42.050 ;
        RECT 109.110 41.895 109.460 42.545 ;
        RECT 109.630 41.725 109.860 42.715 ;
        RECT 109.110 41.555 109.860 41.725 ;
        RECT 109.110 41.055 109.365 41.555 ;
        RECT 109.535 40.885 109.865 41.385 ;
        RECT 110.035 41.055 110.205 43.175 ;
        RECT 110.565 43.075 110.895 43.435 ;
        RECT 111.065 43.045 111.560 43.215 ;
        RECT 111.765 43.045 112.620 43.215 ;
        RECT 110.435 41.855 110.895 42.905 ;
        RECT 110.375 41.070 110.700 41.855 ;
        RECT 111.065 41.685 111.235 43.045 ;
        RECT 111.405 42.135 111.755 42.755 ;
        RECT 111.925 42.535 112.280 42.755 ;
        RECT 111.925 41.945 112.095 42.535 ;
        RECT 112.450 42.335 112.620 43.045 ;
        RECT 113.495 42.975 113.825 43.435 ;
        RECT 114.035 43.075 114.385 43.245 ;
        RECT 112.825 42.505 113.615 42.755 ;
        RECT 114.035 42.685 114.295 43.075 ;
        RECT 114.605 42.985 115.555 43.265 ;
        RECT 115.725 42.995 115.915 43.435 ;
        RECT 116.085 43.055 117.155 43.225 ;
        RECT 113.785 42.335 113.955 42.515 ;
        RECT 111.065 41.515 111.460 41.685 ;
        RECT 111.630 41.555 112.095 41.945 ;
        RECT 112.265 42.165 113.955 42.335 ;
        RECT 111.290 41.385 111.460 41.515 ;
        RECT 112.265 41.385 112.435 42.165 ;
        RECT 114.125 41.995 114.295 42.685 ;
        RECT 112.795 41.825 114.295 41.995 ;
        RECT 114.485 42.025 114.695 42.815 ;
        RECT 114.865 42.195 115.215 42.815 ;
        RECT 115.385 42.205 115.555 42.985 ;
        RECT 116.085 42.825 116.255 43.055 ;
        RECT 115.725 42.655 116.255 42.825 ;
        RECT 115.725 42.375 115.945 42.655 ;
        RECT 116.425 42.485 116.665 42.885 ;
        RECT 115.385 42.035 115.790 42.205 ;
        RECT 116.125 42.115 116.665 42.485 ;
        RECT 116.835 42.700 117.155 43.055 ;
        RECT 117.400 42.975 117.705 43.435 ;
        RECT 117.875 42.725 118.130 43.255 ;
        RECT 116.835 42.525 117.160 42.700 ;
        RECT 116.835 42.225 117.750 42.525 ;
        RECT 117.010 42.195 117.750 42.225 ;
        RECT 114.485 41.865 115.160 42.025 ;
        RECT 115.620 41.945 115.790 42.035 ;
        RECT 114.485 41.855 115.450 41.865 ;
        RECT 114.125 41.685 114.295 41.825 ;
        RECT 110.870 40.885 111.120 41.345 ;
        RECT 111.290 41.055 111.540 41.385 ;
        RECT 111.755 41.055 112.435 41.385 ;
        RECT 112.605 41.485 113.680 41.655 ;
        RECT 114.125 41.515 114.685 41.685 ;
        RECT 114.990 41.565 115.450 41.855 ;
        RECT 115.620 41.775 116.840 41.945 ;
        RECT 112.605 41.145 112.775 41.485 ;
        RECT 113.010 40.885 113.340 41.315 ;
        RECT 113.510 41.145 113.680 41.485 ;
        RECT 113.975 40.885 114.345 41.345 ;
        RECT 114.515 41.055 114.685 41.515 ;
        RECT 115.620 41.395 115.790 41.775 ;
        RECT 117.010 41.605 117.180 42.195 ;
        RECT 117.920 42.075 118.130 42.725 ;
        RECT 118.305 42.665 121.815 43.435 ;
        RECT 122.445 42.685 123.655 43.435 ;
        RECT 118.305 42.145 119.955 42.665 ;
        RECT 114.920 41.055 115.790 41.395 ;
        RECT 116.380 41.435 117.180 41.605 ;
        RECT 115.960 40.885 116.210 41.345 ;
        RECT 116.380 41.145 116.550 41.435 ;
        RECT 116.730 40.885 117.060 41.265 ;
        RECT 117.400 40.885 117.705 42.025 ;
        RECT 117.875 41.195 118.130 42.075 ;
        RECT 120.125 41.975 121.815 42.495 ;
        RECT 118.305 40.885 121.815 41.975 ;
        RECT 122.445 41.975 122.965 42.515 ;
        RECT 123.135 42.145 123.655 42.685 ;
        RECT 122.445 40.885 123.655 41.975 ;
        RECT 5.520 40.715 123.740 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 6.985 40.280 12.330 40.715 ;
        RECT 12.505 40.280 17.850 40.715 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 8.570 38.710 8.910 39.540 ;
        RECT 10.390 39.030 10.740 40.280 ;
        RECT 14.090 38.710 14.430 39.540 ;
        RECT 15.910 39.030 16.260 40.280 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.945 40.280 24.290 40.715 ;
        RECT 6.985 38.165 12.330 38.710 ;
        RECT 12.505 38.165 17.850 38.710 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 20.530 38.710 20.870 39.540 ;
        RECT 22.350 39.030 22.700 40.280 ;
        RECT 25.390 40.045 25.645 40.545 ;
        RECT 25.815 40.215 26.145 40.715 ;
        RECT 25.390 39.875 26.140 40.045 ;
        RECT 25.390 39.055 25.740 39.705 ;
        RECT 25.910 38.885 26.140 39.875 ;
        RECT 25.390 38.715 26.140 38.885 ;
        RECT 18.945 38.165 24.290 38.710 ;
        RECT 25.390 38.425 25.645 38.715 ;
        RECT 25.815 38.165 26.145 38.545 ;
        RECT 26.315 38.425 26.485 40.545 ;
        RECT 26.655 39.745 26.980 40.530 ;
        RECT 27.150 40.255 27.400 40.715 ;
        RECT 27.570 40.215 27.820 40.545 ;
        RECT 28.035 40.215 28.715 40.545 ;
        RECT 27.570 40.085 27.740 40.215 ;
        RECT 27.345 39.915 27.740 40.085 ;
        RECT 26.715 38.695 27.175 39.745 ;
        RECT 27.345 38.555 27.515 39.915 ;
        RECT 27.910 39.655 28.375 40.045 ;
        RECT 27.685 38.845 28.035 39.465 ;
        RECT 28.205 39.065 28.375 39.655 ;
        RECT 28.545 39.435 28.715 40.215 ;
        RECT 28.885 40.115 29.055 40.455 ;
        RECT 29.290 40.285 29.620 40.715 ;
        RECT 29.790 40.115 29.960 40.455 ;
        RECT 30.255 40.255 30.625 40.715 ;
        RECT 28.885 39.945 29.960 40.115 ;
        RECT 30.795 40.085 30.965 40.545 ;
        RECT 31.200 40.205 32.070 40.545 ;
        RECT 32.240 40.255 32.490 40.715 ;
        RECT 30.405 39.915 30.965 40.085 ;
        RECT 30.405 39.775 30.575 39.915 ;
        RECT 29.075 39.605 30.575 39.775 ;
        RECT 31.270 39.745 31.730 40.035 ;
        RECT 28.545 39.265 30.235 39.435 ;
        RECT 28.205 38.845 28.560 39.065 ;
        RECT 28.730 38.555 28.900 39.265 ;
        RECT 29.105 38.845 29.895 39.095 ;
        RECT 30.065 39.085 30.235 39.265 ;
        RECT 30.405 38.915 30.575 39.605 ;
        RECT 26.845 38.165 27.175 38.525 ;
        RECT 27.345 38.385 27.840 38.555 ;
        RECT 28.045 38.385 28.900 38.555 ;
        RECT 29.775 38.165 30.105 38.625 ;
        RECT 30.315 38.525 30.575 38.915 ;
        RECT 30.765 39.735 31.730 39.745 ;
        RECT 31.900 39.825 32.070 40.205 ;
        RECT 32.660 40.165 32.830 40.455 ;
        RECT 33.010 40.335 33.340 40.715 ;
        RECT 32.660 39.995 33.460 40.165 ;
        RECT 30.765 39.575 31.440 39.735 ;
        RECT 31.900 39.655 33.120 39.825 ;
        RECT 30.765 38.785 30.975 39.575 ;
        RECT 31.900 39.565 32.070 39.655 ;
        RECT 31.145 38.785 31.495 39.405 ;
        RECT 31.665 39.395 32.070 39.565 ;
        RECT 31.665 38.615 31.835 39.395 ;
        RECT 32.005 38.945 32.225 39.225 ;
        RECT 32.405 39.115 32.945 39.485 ;
        RECT 33.290 39.405 33.460 39.995 ;
        RECT 33.680 39.575 33.985 40.715 ;
        RECT 34.155 39.525 34.410 40.405 ;
        RECT 34.645 39.575 34.855 40.715 ;
        RECT 33.290 39.375 34.030 39.405 ;
        RECT 32.005 38.775 32.535 38.945 ;
        RECT 30.315 38.355 30.665 38.525 ;
        RECT 30.885 38.335 31.835 38.615 ;
        RECT 32.005 38.165 32.195 38.605 ;
        RECT 32.365 38.545 32.535 38.775 ;
        RECT 32.705 38.715 32.945 39.115 ;
        RECT 33.115 39.075 34.030 39.375 ;
        RECT 33.115 38.900 33.440 39.075 ;
        RECT 33.115 38.545 33.435 38.900 ;
        RECT 34.200 38.875 34.410 39.525 ;
        RECT 35.025 39.565 35.355 40.545 ;
        RECT 35.525 39.575 35.755 40.715 ;
        RECT 35.965 39.625 39.475 40.715 ;
        RECT 32.365 38.375 33.435 38.545 ;
        RECT 33.680 38.165 33.985 38.625 ;
        RECT 34.155 38.345 34.410 38.875 ;
        RECT 34.645 38.165 34.855 38.985 ;
        RECT 35.025 38.965 35.275 39.565 ;
        RECT 35.445 39.155 35.775 39.405 ;
        RECT 35.025 38.335 35.355 38.965 ;
        RECT 35.525 38.165 35.755 38.985 ;
        RECT 35.965 38.935 37.615 39.455 ;
        RECT 37.785 39.105 39.475 39.625 ;
        RECT 39.645 39.640 39.915 40.545 ;
        RECT 40.085 39.955 40.415 40.715 ;
        RECT 40.595 39.785 40.765 40.545 ;
        RECT 35.965 38.165 39.475 38.935 ;
        RECT 39.645 38.840 39.815 39.640 ;
        RECT 40.100 39.615 40.765 39.785 ;
        RECT 41.025 39.625 43.615 40.715 ;
        RECT 40.100 39.470 40.270 39.615 ;
        RECT 39.985 39.140 40.270 39.470 ;
        RECT 40.100 38.885 40.270 39.140 ;
        RECT 40.505 39.065 40.835 39.435 ;
        RECT 41.025 38.935 42.235 39.455 ;
        RECT 42.405 39.105 43.615 39.625 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.705 40.280 50.050 40.715 ;
        RECT 39.645 38.335 39.905 38.840 ;
        RECT 40.100 38.715 40.765 38.885 ;
        RECT 40.085 38.165 40.415 38.545 ;
        RECT 40.595 38.335 40.765 38.715 ;
        RECT 41.025 38.165 43.615 38.935 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 46.290 38.710 46.630 39.540 ;
        RECT 48.110 39.030 48.460 40.280 ;
        RECT 50.225 39.625 51.435 40.715 ;
        RECT 51.610 40.045 51.865 40.545 ;
        RECT 52.035 40.215 52.365 40.715 ;
        RECT 51.610 39.875 52.360 40.045 ;
        RECT 50.225 38.915 50.745 39.455 ;
        RECT 50.915 39.085 51.435 39.625 ;
        RECT 51.610 39.055 51.960 39.705 ;
        RECT 44.705 38.165 50.050 38.710 ;
        RECT 50.225 38.165 51.435 38.915 ;
        RECT 52.130 38.885 52.360 39.875 ;
        RECT 51.610 38.715 52.360 38.885 ;
        RECT 51.610 38.425 51.865 38.715 ;
        RECT 52.035 38.165 52.365 38.545 ;
        RECT 52.535 38.425 52.705 40.545 ;
        RECT 52.875 39.745 53.200 40.530 ;
        RECT 53.370 40.255 53.620 40.715 ;
        RECT 53.790 40.215 54.040 40.545 ;
        RECT 54.255 40.215 54.935 40.545 ;
        RECT 53.790 40.085 53.960 40.215 ;
        RECT 53.565 39.915 53.960 40.085 ;
        RECT 52.935 38.695 53.395 39.745 ;
        RECT 53.565 38.555 53.735 39.915 ;
        RECT 54.130 39.655 54.595 40.045 ;
        RECT 53.905 38.845 54.255 39.465 ;
        RECT 54.425 39.065 54.595 39.655 ;
        RECT 54.765 39.435 54.935 40.215 ;
        RECT 55.105 40.115 55.275 40.455 ;
        RECT 55.510 40.285 55.840 40.715 ;
        RECT 56.010 40.115 56.180 40.455 ;
        RECT 56.475 40.255 56.845 40.715 ;
        RECT 55.105 39.945 56.180 40.115 ;
        RECT 57.015 40.085 57.185 40.545 ;
        RECT 57.420 40.205 58.290 40.545 ;
        RECT 58.460 40.255 58.710 40.715 ;
        RECT 56.625 39.915 57.185 40.085 ;
        RECT 56.625 39.775 56.795 39.915 ;
        RECT 55.295 39.605 56.795 39.775 ;
        RECT 57.490 39.745 57.950 40.035 ;
        RECT 54.765 39.265 56.455 39.435 ;
        RECT 54.425 38.845 54.780 39.065 ;
        RECT 54.950 38.555 55.120 39.265 ;
        RECT 55.325 38.845 56.115 39.095 ;
        RECT 56.285 39.085 56.455 39.265 ;
        RECT 56.625 38.915 56.795 39.605 ;
        RECT 53.065 38.165 53.395 38.525 ;
        RECT 53.565 38.385 54.060 38.555 ;
        RECT 54.265 38.385 55.120 38.555 ;
        RECT 55.995 38.165 56.325 38.625 ;
        RECT 56.535 38.525 56.795 38.915 ;
        RECT 56.985 39.735 57.950 39.745 ;
        RECT 58.120 39.825 58.290 40.205 ;
        RECT 58.880 40.165 59.050 40.455 ;
        RECT 59.230 40.335 59.560 40.715 ;
        RECT 58.880 39.995 59.680 40.165 ;
        RECT 56.985 39.575 57.660 39.735 ;
        RECT 58.120 39.655 59.340 39.825 ;
        RECT 56.985 38.785 57.195 39.575 ;
        RECT 58.120 39.565 58.290 39.655 ;
        RECT 57.365 38.785 57.715 39.405 ;
        RECT 57.885 39.395 58.290 39.565 ;
        RECT 57.885 38.615 58.055 39.395 ;
        RECT 58.225 38.945 58.445 39.225 ;
        RECT 58.625 39.115 59.165 39.485 ;
        RECT 59.510 39.405 59.680 39.995 ;
        RECT 59.900 39.575 60.205 40.715 ;
        RECT 60.375 39.525 60.630 40.405 ;
        RECT 60.805 40.280 66.150 40.715 ;
        RECT 59.510 39.375 60.250 39.405 ;
        RECT 58.225 38.775 58.755 38.945 ;
        RECT 56.535 38.355 56.885 38.525 ;
        RECT 57.105 38.335 58.055 38.615 ;
        RECT 58.225 38.165 58.415 38.605 ;
        RECT 58.585 38.545 58.755 38.775 ;
        RECT 58.925 38.715 59.165 39.115 ;
        RECT 59.335 39.075 60.250 39.375 ;
        RECT 59.335 38.900 59.660 39.075 ;
        RECT 59.335 38.545 59.655 38.900 ;
        RECT 60.420 38.875 60.630 39.525 ;
        RECT 58.585 38.375 59.655 38.545 ;
        RECT 59.900 38.165 60.205 38.625 ;
        RECT 60.375 38.345 60.630 38.875 ;
        RECT 62.390 38.710 62.730 39.540 ;
        RECT 64.210 39.030 64.560 40.280 ;
        RECT 66.325 39.625 69.835 40.715 ;
        RECT 66.325 38.935 67.975 39.455 ;
        RECT 68.145 39.105 69.835 39.625 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.465 40.280 75.810 40.715 ;
        RECT 60.805 38.165 66.150 38.710 ;
        RECT 66.325 38.165 69.835 38.935 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 72.050 38.710 72.390 39.540 ;
        RECT 73.870 39.030 74.220 40.280 ;
        RECT 75.985 39.625 79.495 40.715 ;
        RECT 79.665 39.625 80.875 40.715 ;
        RECT 81.050 40.045 81.305 40.545 ;
        RECT 81.475 40.215 81.805 40.715 ;
        RECT 81.050 39.875 81.800 40.045 ;
        RECT 75.985 38.935 77.635 39.455 ;
        RECT 77.805 39.105 79.495 39.625 ;
        RECT 70.465 38.165 75.810 38.710 ;
        RECT 75.985 38.165 79.495 38.935 ;
        RECT 79.665 38.915 80.185 39.455 ;
        RECT 80.355 39.085 80.875 39.625 ;
        RECT 81.050 39.055 81.400 39.705 ;
        RECT 79.665 38.165 80.875 38.915 ;
        RECT 81.570 38.885 81.800 39.875 ;
        RECT 81.050 38.715 81.800 38.885 ;
        RECT 81.050 38.425 81.305 38.715 ;
        RECT 81.475 38.165 81.805 38.545 ;
        RECT 81.975 38.425 82.145 40.545 ;
        RECT 82.315 39.745 82.640 40.530 ;
        RECT 82.810 40.255 83.060 40.715 ;
        RECT 83.230 40.215 83.480 40.545 ;
        RECT 83.695 40.215 84.375 40.545 ;
        RECT 83.230 40.085 83.400 40.215 ;
        RECT 83.005 39.915 83.400 40.085 ;
        RECT 82.375 38.695 82.835 39.745 ;
        RECT 83.005 38.555 83.175 39.915 ;
        RECT 83.570 39.655 84.035 40.045 ;
        RECT 83.345 38.845 83.695 39.465 ;
        RECT 83.865 39.065 84.035 39.655 ;
        RECT 84.205 39.435 84.375 40.215 ;
        RECT 84.545 40.115 84.715 40.455 ;
        RECT 84.950 40.285 85.280 40.715 ;
        RECT 85.450 40.115 85.620 40.455 ;
        RECT 85.915 40.255 86.285 40.715 ;
        RECT 84.545 39.945 85.620 40.115 ;
        RECT 86.455 40.085 86.625 40.545 ;
        RECT 86.860 40.205 87.730 40.545 ;
        RECT 87.900 40.255 88.150 40.715 ;
        RECT 86.065 39.915 86.625 40.085 ;
        RECT 86.065 39.775 86.235 39.915 ;
        RECT 84.735 39.605 86.235 39.775 ;
        RECT 86.930 39.745 87.390 40.035 ;
        RECT 84.205 39.265 85.895 39.435 ;
        RECT 83.865 38.845 84.220 39.065 ;
        RECT 84.390 38.555 84.560 39.265 ;
        RECT 84.765 38.845 85.555 39.095 ;
        RECT 85.725 39.085 85.895 39.265 ;
        RECT 86.065 38.915 86.235 39.605 ;
        RECT 82.505 38.165 82.835 38.525 ;
        RECT 83.005 38.385 83.500 38.555 ;
        RECT 83.705 38.385 84.560 38.555 ;
        RECT 85.435 38.165 85.765 38.625 ;
        RECT 85.975 38.525 86.235 38.915 ;
        RECT 86.425 39.735 87.390 39.745 ;
        RECT 87.560 39.825 87.730 40.205 ;
        RECT 88.320 40.165 88.490 40.455 ;
        RECT 88.670 40.335 89.000 40.715 ;
        RECT 88.320 39.995 89.120 40.165 ;
        RECT 86.425 39.575 87.100 39.735 ;
        RECT 87.560 39.655 88.780 39.825 ;
        RECT 86.425 38.785 86.635 39.575 ;
        RECT 87.560 39.565 87.730 39.655 ;
        RECT 86.805 38.785 87.155 39.405 ;
        RECT 87.325 39.395 87.730 39.565 ;
        RECT 87.325 38.615 87.495 39.395 ;
        RECT 87.665 38.945 87.885 39.225 ;
        RECT 88.065 39.115 88.605 39.485 ;
        RECT 88.950 39.405 89.120 39.995 ;
        RECT 89.340 39.575 89.645 40.715 ;
        RECT 89.815 39.525 90.070 40.405 ;
        RECT 90.245 40.280 95.590 40.715 ;
        RECT 88.950 39.375 89.690 39.405 ;
        RECT 87.665 38.775 88.195 38.945 ;
        RECT 85.975 38.355 86.325 38.525 ;
        RECT 86.545 38.335 87.495 38.615 ;
        RECT 87.665 38.165 87.855 38.605 ;
        RECT 88.025 38.545 88.195 38.775 ;
        RECT 88.365 38.715 88.605 39.115 ;
        RECT 88.775 39.075 89.690 39.375 ;
        RECT 88.775 38.900 89.100 39.075 ;
        RECT 88.775 38.545 89.095 38.900 ;
        RECT 89.860 38.875 90.070 39.525 ;
        RECT 88.025 38.375 89.095 38.545 ;
        RECT 89.340 38.165 89.645 38.625 ;
        RECT 89.815 38.345 90.070 38.875 ;
        RECT 91.830 38.710 92.170 39.540 ;
        RECT 93.650 39.030 94.000 40.280 ;
        RECT 95.765 39.550 96.055 40.715 ;
        RECT 96.285 39.575 96.495 40.715 ;
        RECT 96.665 39.565 96.995 40.545 ;
        RECT 97.165 39.575 97.395 40.715 ;
        RECT 97.605 39.625 101.115 40.715 ;
        RECT 102.210 40.045 102.465 40.545 ;
        RECT 102.635 40.215 102.965 40.715 ;
        RECT 102.210 39.875 102.960 40.045 ;
        RECT 90.245 38.165 95.590 38.710 ;
        RECT 95.765 38.165 96.055 38.890 ;
        RECT 96.285 38.165 96.495 38.985 ;
        RECT 96.665 38.965 96.915 39.565 ;
        RECT 97.085 39.155 97.415 39.405 ;
        RECT 96.665 38.335 96.995 38.965 ;
        RECT 97.165 38.165 97.395 38.985 ;
        RECT 97.605 38.935 99.255 39.455 ;
        RECT 99.425 39.105 101.115 39.625 ;
        RECT 102.210 39.055 102.560 39.705 ;
        RECT 97.605 38.165 101.115 38.935 ;
        RECT 102.730 38.885 102.960 39.875 ;
        RECT 102.210 38.715 102.960 38.885 ;
        RECT 102.210 38.425 102.465 38.715 ;
        RECT 102.635 38.165 102.965 38.545 ;
        RECT 103.135 38.425 103.305 40.545 ;
        RECT 103.475 39.745 103.800 40.530 ;
        RECT 103.970 40.255 104.220 40.715 ;
        RECT 104.390 40.215 104.640 40.545 ;
        RECT 104.855 40.215 105.535 40.545 ;
        RECT 104.390 40.085 104.560 40.215 ;
        RECT 104.165 39.915 104.560 40.085 ;
        RECT 103.535 38.695 103.995 39.745 ;
        RECT 104.165 38.555 104.335 39.915 ;
        RECT 104.730 39.655 105.195 40.045 ;
        RECT 104.505 38.845 104.855 39.465 ;
        RECT 105.025 39.065 105.195 39.655 ;
        RECT 105.365 39.435 105.535 40.215 ;
        RECT 105.705 40.115 105.875 40.455 ;
        RECT 106.110 40.285 106.440 40.715 ;
        RECT 106.610 40.115 106.780 40.455 ;
        RECT 107.075 40.255 107.445 40.715 ;
        RECT 105.705 39.945 106.780 40.115 ;
        RECT 107.615 40.085 107.785 40.545 ;
        RECT 108.020 40.205 108.890 40.545 ;
        RECT 109.060 40.255 109.310 40.715 ;
        RECT 107.225 39.915 107.785 40.085 ;
        RECT 107.225 39.775 107.395 39.915 ;
        RECT 105.895 39.605 107.395 39.775 ;
        RECT 108.090 39.745 108.550 40.035 ;
        RECT 105.365 39.265 107.055 39.435 ;
        RECT 105.025 38.845 105.380 39.065 ;
        RECT 105.550 38.555 105.720 39.265 ;
        RECT 105.925 38.845 106.715 39.095 ;
        RECT 106.885 39.085 107.055 39.265 ;
        RECT 107.225 38.915 107.395 39.605 ;
        RECT 103.665 38.165 103.995 38.525 ;
        RECT 104.165 38.385 104.660 38.555 ;
        RECT 104.865 38.385 105.720 38.555 ;
        RECT 106.595 38.165 106.925 38.625 ;
        RECT 107.135 38.525 107.395 38.915 ;
        RECT 107.585 39.735 108.550 39.745 ;
        RECT 108.720 39.825 108.890 40.205 ;
        RECT 109.480 40.165 109.650 40.455 ;
        RECT 109.830 40.335 110.160 40.715 ;
        RECT 109.480 39.995 110.280 40.165 ;
        RECT 107.585 39.575 108.260 39.735 ;
        RECT 108.720 39.655 109.940 39.825 ;
        RECT 107.585 38.785 107.795 39.575 ;
        RECT 108.720 39.565 108.890 39.655 ;
        RECT 107.965 38.785 108.315 39.405 ;
        RECT 108.485 39.395 108.890 39.565 ;
        RECT 108.485 38.615 108.655 39.395 ;
        RECT 108.825 38.945 109.045 39.225 ;
        RECT 109.225 39.115 109.765 39.485 ;
        RECT 110.110 39.405 110.280 39.995 ;
        RECT 110.500 39.575 110.805 40.715 ;
        RECT 110.975 39.525 111.230 40.405 ;
        RECT 111.445 39.575 111.675 40.715 ;
        RECT 111.845 39.565 112.175 40.545 ;
        RECT 112.345 39.575 112.555 40.715 ;
        RECT 112.785 40.280 118.130 40.715 ;
        RECT 110.110 39.375 110.850 39.405 ;
        RECT 108.825 38.775 109.355 38.945 ;
        RECT 107.135 38.355 107.485 38.525 ;
        RECT 107.705 38.335 108.655 38.615 ;
        RECT 108.825 38.165 109.015 38.605 ;
        RECT 109.185 38.545 109.355 38.775 ;
        RECT 109.525 38.715 109.765 39.115 ;
        RECT 109.935 39.075 110.850 39.375 ;
        RECT 109.935 38.900 110.260 39.075 ;
        RECT 109.935 38.545 110.255 38.900 ;
        RECT 111.020 38.875 111.230 39.525 ;
        RECT 111.425 39.155 111.755 39.405 ;
        RECT 109.185 38.375 110.255 38.545 ;
        RECT 110.500 38.165 110.805 38.625 ;
        RECT 110.975 38.345 111.230 38.875 ;
        RECT 111.445 38.165 111.675 38.985 ;
        RECT 111.925 38.965 112.175 39.565 ;
        RECT 111.845 38.335 112.175 38.965 ;
        RECT 112.345 38.165 112.555 38.985 ;
        RECT 114.370 38.710 114.710 39.540 ;
        RECT 116.190 39.030 116.540 40.280 ;
        RECT 118.305 39.625 120.895 40.715 ;
        RECT 118.305 38.935 119.515 39.455 ;
        RECT 119.685 39.105 120.895 39.625 ;
        RECT 121.525 39.550 121.815 40.715 ;
        RECT 122.445 39.625 123.655 40.715 ;
        RECT 122.445 39.085 122.965 39.625 ;
        RECT 112.785 38.165 118.130 38.710 ;
        RECT 118.305 38.165 120.895 38.935 ;
        RECT 123.135 38.915 123.655 39.455 ;
        RECT 121.525 38.165 121.815 38.890 ;
        RECT 122.445 38.165 123.655 38.915 ;
        RECT 5.520 37.995 123.740 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 6.985 37.450 12.330 37.995 ;
        RECT 12.505 37.450 17.850 37.995 ;
        RECT 18.025 37.450 23.370 37.995 ;
        RECT 23.545 37.450 28.890 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 8.570 36.620 8.910 37.450 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 10.390 35.880 10.740 37.130 ;
        RECT 14.090 36.620 14.430 37.450 ;
        RECT 15.910 35.880 16.260 37.130 ;
        RECT 19.610 36.620 19.950 37.450 ;
        RECT 21.430 35.880 21.780 37.130 ;
        RECT 25.130 36.620 25.470 37.450 ;
        RECT 29.065 37.225 30.735 37.995 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 31.825 37.450 37.170 37.995 ;
        RECT 26.950 35.880 27.300 37.130 ;
        RECT 29.065 36.705 29.815 37.225 ;
        RECT 29.985 36.535 30.735 37.055 ;
        RECT 33.410 36.620 33.750 37.450 ;
        RECT 37.810 37.445 38.065 37.735 ;
        RECT 38.235 37.615 38.565 37.995 ;
        RECT 37.810 37.275 38.560 37.445 ;
        RECT 6.985 35.445 12.330 35.880 ;
        RECT 12.505 35.445 17.850 35.880 ;
        RECT 18.025 35.445 23.370 35.880 ;
        RECT 23.545 35.445 28.890 35.880 ;
        RECT 29.065 35.445 30.735 36.535 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 35.230 35.880 35.580 37.130 ;
        RECT 37.810 36.455 38.160 37.105 ;
        RECT 38.330 36.285 38.560 37.275 ;
        RECT 37.810 36.115 38.560 36.285 ;
        RECT 31.825 35.445 37.170 35.880 ;
        RECT 37.810 35.615 38.065 36.115 ;
        RECT 38.235 35.445 38.565 35.945 ;
        RECT 38.735 35.615 38.905 37.735 ;
        RECT 39.265 37.635 39.595 37.995 ;
        RECT 39.765 37.605 40.260 37.775 ;
        RECT 40.465 37.605 41.320 37.775 ;
        RECT 39.135 36.415 39.595 37.465 ;
        RECT 39.075 35.630 39.400 36.415 ;
        RECT 39.765 36.245 39.935 37.605 ;
        RECT 40.105 36.695 40.455 37.315 ;
        RECT 40.625 37.095 40.980 37.315 ;
        RECT 40.625 36.505 40.795 37.095 ;
        RECT 41.150 36.895 41.320 37.605 ;
        RECT 42.195 37.535 42.525 37.995 ;
        RECT 42.735 37.635 43.085 37.805 ;
        RECT 41.525 37.065 42.315 37.315 ;
        RECT 42.735 37.245 42.995 37.635 ;
        RECT 43.305 37.545 44.255 37.825 ;
        RECT 44.425 37.555 44.615 37.995 ;
        RECT 44.785 37.615 45.855 37.785 ;
        RECT 42.485 36.895 42.655 37.075 ;
        RECT 39.765 36.075 40.160 36.245 ;
        RECT 40.330 36.115 40.795 36.505 ;
        RECT 40.965 36.725 42.655 36.895 ;
        RECT 39.990 35.945 40.160 36.075 ;
        RECT 40.965 35.945 41.135 36.725 ;
        RECT 42.825 36.555 42.995 37.245 ;
        RECT 41.495 36.385 42.995 36.555 ;
        RECT 43.185 36.585 43.395 37.375 ;
        RECT 43.565 36.755 43.915 37.375 ;
        RECT 44.085 36.765 44.255 37.545 ;
        RECT 44.785 37.385 44.955 37.615 ;
        RECT 44.425 37.215 44.955 37.385 ;
        RECT 44.425 36.935 44.645 37.215 ;
        RECT 45.125 37.045 45.365 37.445 ;
        RECT 44.085 36.595 44.490 36.765 ;
        RECT 44.825 36.675 45.365 37.045 ;
        RECT 45.535 37.260 45.855 37.615 ;
        RECT 46.100 37.535 46.405 37.995 ;
        RECT 46.575 37.285 46.830 37.815 ;
        RECT 45.535 37.085 45.860 37.260 ;
        RECT 45.535 36.785 46.450 37.085 ;
        RECT 45.710 36.755 46.450 36.785 ;
        RECT 43.185 36.425 43.860 36.585 ;
        RECT 44.320 36.505 44.490 36.595 ;
        RECT 43.185 36.415 44.150 36.425 ;
        RECT 42.825 36.245 42.995 36.385 ;
        RECT 39.570 35.445 39.820 35.905 ;
        RECT 39.990 35.615 40.240 35.945 ;
        RECT 40.455 35.615 41.135 35.945 ;
        RECT 41.305 36.045 42.380 36.215 ;
        RECT 42.825 36.075 43.385 36.245 ;
        RECT 43.690 36.125 44.150 36.415 ;
        RECT 44.320 36.335 45.540 36.505 ;
        RECT 41.305 35.705 41.475 36.045 ;
        RECT 41.710 35.445 42.040 35.875 ;
        RECT 42.210 35.705 42.380 36.045 ;
        RECT 42.675 35.445 43.045 35.905 ;
        RECT 43.215 35.615 43.385 36.075 ;
        RECT 44.320 35.955 44.490 36.335 ;
        RECT 45.710 36.165 45.880 36.755 ;
        RECT 46.620 36.635 46.830 37.285 ;
        RECT 43.620 35.615 44.490 35.955 ;
        RECT 45.080 35.995 45.880 36.165 ;
        RECT 44.660 35.445 44.910 35.905 ;
        RECT 45.080 35.705 45.250 35.995 ;
        RECT 45.430 35.445 45.760 35.825 ;
        RECT 46.100 35.445 46.405 36.585 ;
        RECT 46.575 35.755 46.830 36.635 ;
        RECT 47.010 37.255 47.265 37.825 ;
        RECT 47.435 37.595 47.765 37.995 ;
        RECT 48.190 37.460 48.720 37.825 ;
        RECT 48.190 37.425 48.365 37.460 ;
        RECT 47.435 37.255 48.365 37.425 ;
        RECT 47.010 36.585 47.180 37.255 ;
        RECT 47.435 37.085 47.605 37.255 ;
        RECT 47.350 36.755 47.605 37.085 ;
        RECT 47.830 36.755 48.025 37.085 ;
        RECT 47.010 35.615 47.345 36.585 ;
        RECT 47.515 35.445 47.685 36.585 ;
        RECT 47.855 35.785 48.025 36.755 ;
        RECT 48.195 36.125 48.365 37.255 ;
        RECT 48.535 36.465 48.705 37.265 ;
        RECT 48.910 36.975 49.185 37.825 ;
        RECT 48.905 36.805 49.185 36.975 ;
        RECT 48.910 36.665 49.185 36.805 ;
        RECT 49.355 36.465 49.545 37.825 ;
        RECT 49.725 37.460 50.235 37.995 ;
        RECT 50.455 37.185 50.700 37.790 ;
        RECT 51.145 37.225 54.655 37.995 ;
        RECT 49.745 37.015 50.975 37.185 ;
        RECT 48.535 36.295 49.545 36.465 ;
        RECT 49.715 36.450 50.465 36.640 ;
        RECT 48.195 35.955 49.320 36.125 ;
        RECT 49.715 35.785 49.885 36.450 ;
        RECT 50.635 36.205 50.975 37.015 ;
        RECT 51.145 36.705 52.795 37.225 ;
        RECT 55.785 37.175 56.015 37.995 ;
        RECT 56.185 37.195 56.515 37.825 ;
        RECT 52.965 36.535 54.655 37.055 ;
        RECT 55.765 36.755 56.095 37.005 ;
        RECT 56.265 36.595 56.515 37.195 ;
        RECT 56.685 37.175 56.895 37.995 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 57.585 37.320 57.845 37.825 ;
        RECT 58.025 37.615 58.355 37.995 ;
        RECT 58.535 37.445 58.705 37.825 ;
        RECT 47.855 35.615 49.885 35.785 ;
        RECT 50.055 35.445 50.225 36.205 ;
        RECT 50.460 35.795 50.975 36.205 ;
        RECT 51.145 35.445 54.655 36.535 ;
        RECT 55.785 35.445 56.015 36.585 ;
        RECT 56.185 35.615 56.515 36.595 ;
        RECT 56.685 35.445 56.895 36.585 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 57.585 36.520 57.755 37.320 ;
        RECT 58.040 37.275 58.705 37.445 ;
        RECT 58.040 37.020 58.210 37.275 ;
        RECT 58.965 37.225 62.475 37.995 ;
        RECT 62.680 37.255 63.295 37.825 ;
        RECT 63.465 37.485 63.680 37.995 ;
        RECT 63.910 37.485 64.190 37.815 ;
        RECT 64.370 37.485 64.610 37.995 ;
        RECT 57.925 36.690 58.210 37.020 ;
        RECT 58.445 36.725 58.775 37.095 ;
        RECT 58.965 36.705 60.615 37.225 ;
        RECT 58.040 36.545 58.210 36.690 ;
        RECT 57.585 35.615 57.855 36.520 ;
        RECT 58.040 36.375 58.705 36.545 ;
        RECT 60.785 36.535 62.475 37.055 ;
        RECT 58.025 35.445 58.355 36.205 ;
        RECT 58.535 35.615 58.705 36.375 ;
        RECT 58.965 35.445 62.475 36.535 ;
        RECT 62.680 36.235 62.995 37.255 ;
        RECT 63.165 36.585 63.335 37.085 ;
        RECT 63.585 36.755 63.850 37.315 ;
        RECT 64.020 36.585 64.190 37.485 ;
        RECT 64.360 36.755 64.715 37.315 ;
        RECT 64.945 37.225 66.615 37.995 ;
        RECT 66.785 37.320 67.060 37.665 ;
        RECT 67.250 37.595 67.625 37.995 ;
        RECT 67.795 37.425 67.965 37.775 ;
        RECT 68.135 37.595 68.465 37.995 ;
        RECT 68.635 37.425 68.895 37.825 ;
        RECT 64.945 36.705 65.695 37.225 ;
        RECT 63.165 36.415 64.590 36.585 ;
        RECT 65.865 36.535 66.615 37.055 ;
        RECT 62.680 35.615 63.215 36.235 ;
        RECT 63.385 35.445 63.715 36.245 ;
        RECT 64.200 36.240 64.590 36.415 ;
        RECT 64.945 35.445 66.615 36.535 ;
        RECT 66.785 36.585 66.955 37.320 ;
        RECT 67.230 37.255 68.895 37.425 ;
        RECT 67.230 37.085 67.400 37.255 ;
        RECT 69.075 37.175 69.405 37.595 ;
        RECT 69.575 37.175 69.835 37.995 ;
        RECT 70.015 37.270 70.345 37.780 ;
        RECT 70.515 37.595 70.845 37.995 ;
        RECT 71.895 37.425 72.225 37.765 ;
        RECT 72.395 37.595 72.725 37.995 ;
        RECT 73.225 37.450 78.570 37.995 ;
        RECT 69.075 37.085 69.325 37.175 ;
        RECT 67.125 36.755 67.400 37.085 ;
        RECT 67.570 36.755 68.395 37.085 ;
        RECT 68.610 36.755 69.325 37.085 ;
        RECT 69.495 36.755 69.830 37.005 ;
        RECT 67.230 36.585 67.400 36.755 ;
        RECT 66.785 35.615 67.060 36.585 ;
        RECT 67.230 36.415 67.890 36.585 ;
        RECT 68.150 36.465 68.395 36.755 ;
        RECT 67.720 36.295 67.890 36.415 ;
        RECT 68.565 36.295 68.895 36.585 ;
        RECT 67.270 35.445 67.550 36.245 ;
        RECT 67.720 36.125 68.895 36.295 ;
        RECT 69.155 36.195 69.325 36.755 ;
        RECT 67.720 35.625 69.335 35.955 ;
        RECT 69.575 35.445 69.835 36.585 ;
        RECT 70.015 36.505 70.205 37.270 ;
        RECT 70.515 37.255 72.880 37.425 ;
        RECT 70.515 37.085 70.685 37.255 ;
        RECT 70.375 36.755 70.685 37.085 ;
        RECT 70.855 36.755 71.160 37.085 ;
        RECT 70.015 35.655 70.345 36.505 ;
        RECT 70.515 35.445 70.765 36.585 ;
        RECT 70.945 36.425 71.160 36.755 ;
        RECT 71.335 36.425 71.620 37.085 ;
        RECT 71.815 36.425 72.080 37.085 ;
        RECT 72.295 36.425 72.540 37.085 ;
        RECT 72.710 36.255 72.880 37.255 ;
        RECT 74.810 36.620 75.150 37.450 ;
        RECT 78.745 37.225 82.255 37.995 ;
        RECT 82.885 37.270 83.175 37.995 ;
        RECT 83.345 37.320 83.605 37.825 ;
        RECT 83.785 37.615 84.115 37.995 ;
        RECT 84.295 37.445 84.465 37.825 ;
        RECT 70.955 36.085 72.245 36.255 ;
        RECT 70.955 35.665 71.205 36.085 ;
        RECT 71.435 35.445 71.765 35.915 ;
        RECT 71.995 35.665 72.245 36.085 ;
        RECT 72.425 36.085 72.880 36.255 ;
        RECT 72.425 35.655 72.755 36.085 ;
        RECT 76.630 35.880 76.980 37.130 ;
        RECT 78.745 36.705 80.395 37.225 ;
        RECT 80.565 36.535 82.255 37.055 ;
        RECT 73.225 35.445 78.570 35.880 ;
        RECT 78.745 35.445 82.255 36.535 ;
        RECT 82.885 35.445 83.175 36.610 ;
        RECT 83.345 36.520 83.515 37.320 ;
        RECT 83.800 37.275 84.465 37.445 ;
        RECT 83.800 37.020 83.970 37.275 ;
        RECT 84.765 37.175 84.995 37.995 ;
        RECT 85.165 37.195 85.495 37.825 ;
        RECT 83.685 36.690 83.970 37.020 ;
        RECT 84.205 36.725 84.535 37.095 ;
        RECT 84.745 36.755 85.075 37.005 ;
        RECT 83.800 36.545 83.970 36.690 ;
        RECT 85.245 36.595 85.495 37.195 ;
        RECT 85.665 37.175 85.875 37.995 ;
        RECT 86.105 37.450 91.450 37.995 ;
        RECT 91.625 37.450 96.970 37.995 ;
        RECT 87.690 36.620 88.030 37.450 ;
        RECT 83.345 35.615 83.615 36.520 ;
        RECT 83.800 36.375 84.465 36.545 ;
        RECT 83.785 35.445 84.115 36.205 ;
        RECT 84.295 35.615 84.465 36.375 ;
        RECT 84.765 35.445 84.995 36.585 ;
        RECT 85.165 35.615 85.495 36.595 ;
        RECT 85.665 35.445 85.875 36.585 ;
        RECT 89.510 35.880 89.860 37.130 ;
        RECT 93.210 36.620 93.550 37.450 ;
        RECT 97.645 37.175 97.875 37.995 ;
        RECT 98.045 37.195 98.375 37.825 ;
        RECT 95.030 35.880 95.380 37.130 ;
        RECT 97.625 36.755 97.955 37.005 ;
        RECT 98.125 36.595 98.375 37.195 ;
        RECT 98.545 37.175 98.755 37.995 ;
        RECT 98.985 37.225 101.575 37.995 ;
        RECT 102.295 37.445 102.465 37.825 ;
        RECT 102.645 37.615 102.975 37.995 ;
        RECT 102.295 37.275 102.960 37.445 ;
        RECT 103.155 37.320 103.415 37.825 ;
        RECT 98.985 36.705 100.195 37.225 ;
        RECT 86.105 35.445 91.450 35.880 ;
        RECT 91.625 35.445 96.970 35.880 ;
        RECT 97.645 35.445 97.875 36.585 ;
        RECT 98.045 35.615 98.375 36.595 ;
        RECT 98.545 35.445 98.755 36.585 ;
        RECT 100.365 36.535 101.575 37.055 ;
        RECT 102.225 36.725 102.555 37.095 ;
        RECT 102.790 37.020 102.960 37.275 ;
        RECT 102.790 36.690 103.075 37.020 ;
        RECT 102.790 36.545 102.960 36.690 ;
        RECT 98.985 35.445 101.575 36.535 ;
        RECT 102.295 36.375 102.960 36.545 ;
        RECT 103.245 36.520 103.415 37.320 ;
        RECT 102.295 35.615 102.465 36.375 ;
        RECT 102.645 35.445 102.975 36.205 ;
        RECT 103.145 35.615 103.415 36.520 ;
        RECT 103.590 37.255 103.845 37.825 ;
        RECT 104.015 37.595 104.345 37.995 ;
        RECT 104.770 37.460 105.300 37.825 ;
        RECT 105.490 37.655 105.765 37.825 ;
        RECT 105.485 37.485 105.765 37.655 ;
        RECT 104.770 37.425 104.945 37.460 ;
        RECT 104.015 37.255 104.945 37.425 ;
        RECT 103.590 36.585 103.760 37.255 ;
        RECT 104.015 37.085 104.185 37.255 ;
        RECT 103.930 36.755 104.185 37.085 ;
        RECT 104.410 36.755 104.605 37.085 ;
        RECT 103.590 35.615 103.925 36.585 ;
        RECT 104.095 35.445 104.265 36.585 ;
        RECT 104.435 35.785 104.605 36.755 ;
        RECT 104.775 36.125 104.945 37.255 ;
        RECT 105.115 36.465 105.285 37.265 ;
        RECT 105.490 36.665 105.765 37.485 ;
        RECT 105.935 36.465 106.125 37.825 ;
        RECT 106.305 37.460 106.815 37.995 ;
        RECT 107.035 37.185 107.280 37.790 ;
        RECT 108.645 37.270 108.935 37.995 ;
        RECT 106.325 37.015 107.555 37.185 ;
        RECT 109.165 37.175 109.375 37.995 ;
        RECT 109.545 37.195 109.875 37.825 ;
        RECT 105.115 36.295 106.125 36.465 ;
        RECT 106.295 36.450 107.045 36.640 ;
        RECT 104.775 35.955 105.900 36.125 ;
        RECT 106.295 35.785 106.465 36.450 ;
        RECT 107.215 36.205 107.555 37.015 ;
        RECT 104.435 35.615 106.465 35.785 ;
        RECT 106.635 35.445 106.805 36.205 ;
        RECT 107.040 35.795 107.555 36.205 ;
        RECT 108.645 35.445 108.935 36.610 ;
        RECT 109.545 36.595 109.795 37.195 ;
        RECT 110.045 37.175 110.275 37.995 ;
        RECT 110.485 37.450 115.830 37.995 ;
        RECT 116.005 37.450 121.350 37.995 ;
        RECT 109.965 36.755 110.295 37.005 ;
        RECT 112.070 36.620 112.410 37.450 ;
        RECT 109.165 35.445 109.375 36.585 ;
        RECT 109.545 35.615 109.875 36.595 ;
        RECT 110.045 35.445 110.275 36.585 ;
        RECT 113.890 35.880 114.240 37.130 ;
        RECT 117.590 36.620 117.930 37.450 ;
        RECT 122.445 37.245 123.655 37.995 ;
        RECT 119.410 35.880 119.760 37.130 ;
        RECT 122.445 36.535 122.965 37.075 ;
        RECT 123.135 36.705 123.655 37.245 ;
        RECT 110.485 35.445 115.830 35.880 ;
        RECT 116.005 35.445 121.350 35.880 ;
        RECT 122.445 35.445 123.655 36.535 ;
        RECT 5.520 35.275 123.740 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.840 12.330 35.275 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 8.570 33.270 8.910 34.100 ;
        RECT 10.390 33.590 10.740 34.840 ;
        RECT 12.505 34.185 15.095 35.275 ;
        RECT 12.505 33.495 13.715 34.015 ;
        RECT 13.885 33.665 15.095 34.185 ;
        RECT 15.265 34.200 15.535 35.105 ;
        RECT 15.705 34.515 16.035 35.275 ;
        RECT 16.215 34.345 16.385 35.105 ;
        RECT 6.985 32.725 12.330 33.270 ;
        RECT 12.505 32.725 15.095 33.495 ;
        RECT 15.265 33.400 15.435 34.200 ;
        RECT 15.720 34.175 16.385 34.345 ;
        RECT 16.645 34.185 18.315 35.275 ;
        RECT 15.720 34.030 15.890 34.175 ;
        RECT 15.605 33.700 15.890 34.030 ;
        RECT 15.720 33.445 15.890 33.700 ;
        RECT 16.125 33.625 16.455 33.995 ;
        RECT 16.645 33.495 17.395 34.015 ;
        RECT 17.565 33.665 18.315 34.185 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 18.950 34.135 19.285 35.105 ;
        RECT 19.455 34.135 19.625 35.275 ;
        RECT 19.795 34.935 21.825 35.105 ;
        RECT 15.265 32.895 15.525 33.400 ;
        RECT 15.720 33.275 16.385 33.445 ;
        RECT 15.705 32.725 16.035 33.105 ;
        RECT 16.215 32.895 16.385 33.275 ;
        RECT 16.645 32.725 18.315 33.495 ;
        RECT 18.950 33.465 19.120 34.135 ;
        RECT 19.795 33.965 19.965 34.935 ;
        RECT 19.290 33.635 19.545 33.965 ;
        RECT 19.770 33.635 19.965 33.965 ;
        RECT 20.135 34.595 21.260 34.765 ;
        RECT 19.375 33.465 19.545 33.635 ;
        RECT 20.135 33.465 20.305 34.595 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 18.950 32.895 19.205 33.465 ;
        RECT 19.375 33.295 20.305 33.465 ;
        RECT 20.475 34.255 21.485 34.425 ;
        RECT 20.475 33.455 20.645 34.255 ;
        RECT 20.850 33.575 21.125 34.055 ;
        RECT 20.845 33.405 21.125 33.575 ;
        RECT 20.130 33.260 20.305 33.295 ;
        RECT 19.375 32.725 19.705 33.125 ;
        RECT 20.130 32.895 20.660 33.260 ;
        RECT 20.850 32.895 21.125 33.405 ;
        RECT 21.295 32.895 21.485 34.255 ;
        RECT 21.655 34.270 21.825 34.935 ;
        RECT 21.995 34.515 22.165 35.275 ;
        RECT 22.400 34.515 22.915 34.925 ;
        RECT 21.655 34.080 22.405 34.270 ;
        RECT 22.575 33.705 22.915 34.515 ;
        RECT 21.685 33.535 22.915 33.705 ;
        RECT 23.090 34.135 23.425 35.105 ;
        RECT 23.595 34.135 23.765 35.275 ;
        RECT 23.935 34.935 25.965 35.105 ;
        RECT 21.665 32.725 22.175 33.260 ;
        RECT 22.395 32.930 22.640 33.535 ;
        RECT 23.090 33.465 23.260 34.135 ;
        RECT 23.935 33.965 24.105 34.935 ;
        RECT 23.430 33.635 23.685 33.965 ;
        RECT 23.910 33.635 24.105 33.965 ;
        RECT 24.275 34.595 25.400 34.765 ;
        RECT 23.515 33.465 23.685 33.635 ;
        RECT 24.275 33.465 24.445 34.595 ;
        RECT 23.090 32.895 23.345 33.465 ;
        RECT 23.515 33.295 24.445 33.465 ;
        RECT 24.615 34.255 25.625 34.425 ;
        RECT 24.615 33.455 24.785 34.255 ;
        RECT 24.990 33.915 25.265 34.055 ;
        RECT 24.985 33.745 25.265 33.915 ;
        RECT 24.270 33.260 24.445 33.295 ;
        RECT 23.515 32.725 23.845 33.125 ;
        RECT 24.270 32.895 24.800 33.260 ;
        RECT 24.990 32.895 25.265 33.745 ;
        RECT 25.435 32.895 25.625 34.255 ;
        RECT 25.795 34.270 25.965 34.935 ;
        RECT 26.135 34.515 26.305 35.275 ;
        RECT 26.540 34.515 27.055 34.925 ;
        RECT 27.225 34.840 32.570 35.275 ;
        RECT 32.745 34.840 38.090 35.275 ;
        RECT 25.795 34.080 26.545 34.270 ;
        RECT 26.715 33.705 27.055 34.515 ;
        RECT 25.825 33.535 27.055 33.705 ;
        RECT 25.805 32.725 26.315 33.260 ;
        RECT 26.535 32.930 26.780 33.535 ;
        RECT 28.810 33.270 29.150 34.100 ;
        RECT 30.630 33.590 30.980 34.840 ;
        RECT 34.330 33.270 34.670 34.100 ;
        RECT 36.150 33.590 36.500 34.840 ;
        RECT 38.265 34.185 40.855 35.275 ;
        RECT 38.265 33.495 39.475 34.015 ;
        RECT 39.645 33.665 40.855 34.185 ;
        RECT 41.025 34.200 41.295 35.105 ;
        RECT 41.465 34.515 41.795 35.275 ;
        RECT 41.975 34.345 42.145 35.105 ;
        RECT 27.225 32.725 32.570 33.270 ;
        RECT 32.745 32.725 38.090 33.270 ;
        RECT 38.265 32.725 40.855 33.495 ;
        RECT 41.025 33.400 41.195 34.200 ;
        RECT 41.480 34.175 42.145 34.345 ;
        RECT 41.480 34.030 41.650 34.175 ;
        RECT 42.445 34.135 42.675 35.275 ;
        RECT 42.845 34.125 43.175 35.105 ;
        RECT 43.345 34.135 43.555 35.275 ;
        RECT 41.365 33.700 41.650 34.030 ;
        RECT 41.480 33.445 41.650 33.700 ;
        RECT 41.885 33.625 42.215 33.995 ;
        RECT 42.425 33.715 42.755 33.965 ;
        RECT 41.025 32.895 41.285 33.400 ;
        RECT 41.480 33.275 42.145 33.445 ;
        RECT 41.465 32.725 41.795 33.105 ;
        RECT 41.975 32.895 42.145 33.275 ;
        RECT 42.445 32.725 42.675 33.545 ;
        RECT 42.925 33.525 43.175 34.125 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 44.765 34.135 44.975 35.275 ;
        RECT 45.145 34.125 45.475 35.105 ;
        RECT 45.645 34.135 45.875 35.275 ;
        RECT 46.085 34.840 51.430 35.275 ;
        RECT 51.605 34.840 56.950 35.275 ;
        RECT 42.845 32.895 43.175 33.525 ;
        RECT 43.345 32.725 43.555 33.545 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 44.765 32.725 44.975 33.545 ;
        RECT 45.145 33.525 45.395 34.125 ;
        RECT 45.565 33.715 45.895 33.965 ;
        RECT 45.145 32.895 45.475 33.525 ;
        RECT 45.645 32.725 45.875 33.545 ;
        RECT 47.670 33.270 48.010 34.100 ;
        RECT 49.490 33.590 49.840 34.840 ;
        RECT 53.190 33.270 53.530 34.100 ;
        RECT 55.010 33.590 55.360 34.840 ;
        RECT 57.125 34.185 58.795 35.275 ;
        RECT 57.125 33.495 57.875 34.015 ;
        RECT 58.045 33.665 58.795 34.185 ;
        RECT 59.425 34.135 59.705 35.275 ;
        RECT 59.875 34.125 60.205 35.105 ;
        RECT 60.375 34.135 60.635 35.275 ;
        RECT 60.805 34.405 61.080 35.105 ;
        RECT 61.250 34.730 61.505 35.275 ;
        RECT 61.675 34.765 62.155 35.105 ;
        RECT 62.330 34.720 62.935 35.275 ;
        RECT 62.320 34.620 62.935 34.720 ;
        RECT 62.320 34.595 62.505 34.620 ;
        RECT 59.435 33.695 59.770 33.965 ;
        RECT 59.940 33.575 60.110 34.125 ;
        RECT 60.280 33.715 60.615 33.965 ;
        RECT 59.940 33.525 60.115 33.575 ;
        RECT 46.085 32.725 51.430 33.270 ;
        RECT 51.605 32.725 56.950 33.270 ;
        RECT 57.125 32.725 58.795 33.495 ;
        RECT 59.425 32.725 59.735 33.525 ;
        RECT 59.940 32.895 60.635 33.525 ;
        RECT 60.805 33.375 60.975 34.405 ;
        RECT 61.250 34.275 62.005 34.525 ;
        RECT 62.175 34.350 62.505 34.595 ;
        RECT 61.250 34.240 62.020 34.275 ;
        RECT 61.250 34.230 62.035 34.240 ;
        RECT 61.145 34.215 62.040 34.230 ;
        RECT 61.145 34.200 62.060 34.215 ;
        RECT 61.145 34.190 62.080 34.200 ;
        RECT 61.145 34.180 62.105 34.190 ;
        RECT 61.145 34.150 62.175 34.180 ;
        RECT 61.145 34.120 62.195 34.150 ;
        RECT 61.145 34.090 62.215 34.120 ;
        RECT 61.145 34.065 62.245 34.090 ;
        RECT 61.145 34.030 62.280 34.065 ;
        RECT 61.145 34.025 62.310 34.030 ;
        RECT 61.145 33.630 61.375 34.025 ;
        RECT 61.920 34.020 62.310 34.025 ;
        RECT 61.945 34.010 62.310 34.020 ;
        RECT 61.960 34.005 62.310 34.010 ;
        RECT 61.975 34.000 62.310 34.005 ;
        RECT 62.675 34.000 62.935 34.450 ;
        RECT 63.105 34.135 63.365 35.275 ;
        RECT 63.535 34.305 63.865 35.105 ;
        RECT 64.035 34.475 64.205 35.275 ;
        RECT 64.405 34.305 64.735 35.105 ;
        RECT 64.935 34.475 65.215 35.275 ;
        RECT 63.535 34.135 64.815 34.305 ;
        RECT 61.975 33.995 62.935 34.000 ;
        RECT 61.985 33.985 62.935 33.995 ;
        RECT 61.995 33.980 62.935 33.985 ;
        RECT 62.005 33.970 62.935 33.980 ;
        RECT 62.010 33.960 62.935 33.970 ;
        RECT 62.015 33.955 62.935 33.960 ;
        RECT 62.025 33.940 62.935 33.955 ;
        RECT 62.030 33.925 62.935 33.940 ;
        RECT 62.040 33.900 62.935 33.925 ;
        RECT 61.545 33.430 61.875 33.855 ;
        RECT 60.805 32.895 61.065 33.375 ;
        RECT 61.235 32.725 61.485 33.265 ;
        RECT 61.655 32.945 61.875 33.430 ;
        RECT 62.045 33.830 62.935 33.900 ;
        RECT 62.045 33.105 62.215 33.830 ;
        RECT 62.385 33.275 62.935 33.660 ;
        RECT 63.130 33.635 63.415 33.965 ;
        RECT 63.615 33.635 63.995 33.965 ;
        RECT 64.165 33.635 64.475 33.965 ;
        RECT 62.045 32.935 62.935 33.105 ;
        RECT 63.110 32.725 63.445 33.465 ;
        RECT 63.615 32.940 63.830 33.635 ;
        RECT 64.165 33.465 64.370 33.635 ;
        RECT 64.645 33.465 64.815 34.135 ;
        RECT 64.995 33.635 65.235 34.305 ;
        RECT 65.405 34.135 65.665 35.275 ;
        RECT 65.905 34.765 67.520 35.095 ;
        RECT 65.915 33.965 66.085 34.525 ;
        RECT 66.345 34.425 67.520 34.595 ;
        RECT 67.690 34.475 67.970 35.275 ;
        RECT 66.345 34.135 66.675 34.425 ;
        RECT 67.350 34.305 67.520 34.425 ;
        RECT 66.845 33.965 67.090 34.255 ;
        RECT 67.350 34.135 68.010 34.305 ;
        RECT 68.180 34.135 68.455 35.105 ;
        RECT 68.625 34.185 69.835 35.275 ;
        RECT 67.840 33.965 68.010 34.135 ;
        RECT 65.410 33.715 65.745 33.965 ;
        RECT 65.915 33.635 66.630 33.965 ;
        RECT 66.845 33.635 67.670 33.965 ;
        RECT 67.840 33.635 68.115 33.965 ;
        RECT 65.915 33.545 66.165 33.635 ;
        RECT 64.020 32.940 64.370 33.465 ;
        RECT 64.540 32.895 65.235 33.465 ;
        RECT 65.405 32.725 65.665 33.545 ;
        RECT 65.835 33.125 66.165 33.545 ;
        RECT 67.840 33.465 68.010 33.635 ;
        RECT 66.345 33.295 68.010 33.465 ;
        RECT 68.285 33.400 68.455 34.135 ;
        RECT 66.345 32.895 66.605 33.295 ;
        RECT 66.775 32.725 67.105 33.125 ;
        RECT 67.275 32.945 67.445 33.295 ;
        RECT 67.615 32.725 67.990 33.125 ;
        RECT 68.180 33.055 68.455 33.400 ;
        RECT 68.625 33.475 69.145 34.015 ;
        RECT 69.315 33.645 69.835 34.185 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 70.465 34.405 70.740 35.105 ;
        RECT 70.910 34.730 71.165 35.275 ;
        RECT 71.335 34.765 71.815 35.105 ;
        RECT 71.990 34.720 72.595 35.275 ;
        RECT 72.765 34.840 78.110 35.275 ;
        RECT 78.285 34.840 83.630 35.275 ;
        RECT 83.805 34.840 89.150 35.275 ;
        RECT 71.980 34.620 72.595 34.720 ;
        RECT 71.980 34.595 72.165 34.620 ;
        RECT 68.625 32.725 69.835 33.475 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 70.465 33.375 70.635 34.405 ;
        RECT 70.910 34.275 71.665 34.525 ;
        RECT 71.835 34.350 72.165 34.595 ;
        RECT 70.910 34.240 71.680 34.275 ;
        RECT 70.910 34.230 71.695 34.240 ;
        RECT 70.805 34.215 71.700 34.230 ;
        RECT 70.805 34.200 71.720 34.215 ;
        RECT 70.805 34.190 71.740 34.200 ;
        RECT 70.805 34.180 71.765 34.190 ;
        RECT 70.805 34.150 71.835 34.180 ;
        RECT 70.805 34.120 71.855 34.150 ;
        RECT 70.805 34.090 71.875 34.120 ;
        RECT 70.805 34.065 71.905 34.090 ;
        RECT 70.805 34.030 71.940 34.065 ;
        RECT 70.805 34.025 71.970 34.030 ;
        RECT 70.805 33.630 71.035 34.025 ;
        RECT 71.580 34.020 71.970 34.025 ;
        RECT 71.605 34.010 71.970 34.020 ;
        RECT 71.620 34.005 71.970 34.010 ;
        RECT 71.635 34.000 71.970 34.005 ;
        RECT 72.335 34.000 72.595 34.450 ;
        RECT 71.635 33.995 72.595 34.000 ;
        RECT 71.645 33.985 72.595 33.995 ;
        RECT 71.655 33.980 72.595 33.985 ;
        RECT 71.665 33.970 72.595 33.980 ;
        RECT 71.670 33.960 72.595 33.970 ;
        RECT 71.675 33.955 72.595 33.960 ;
        RECT 71.685 33.940 72.595 33.955 ;
        RECT 71.690 33.925 72.595 33.940 ;
        RECT 71.700 33.900 72.595 33.925 ;
        RECT 71.205 33.430 71.535 33.855 ;
        RECT 70.465 32.895 70.725 33.375 ;
        RECT 70.895 32.725 71.145 33.265 ;
        RECT 71.315 32.945 71.535 33.430 ;
        RECT 71.705 33.830 72.595 33.900 ;
        RECT 71.705 33.105 71.875 33.830 ;
        RECT 72.045 33.275 72.595 33.660 ;
        RECT 74.350 33.270 74.690 34.100 ;
        RECT 76.170 33.590 76.520 34.840 ;
        RECT 79.870 33.270 80.210 34.100 ;
        RECT 81.690 33.590 82.040 34.840 ;
        RECT 85.390 33.270 85.730 34.100 ;
        RECT 87.210 33.590 87.560 34.840 ;
        RECT 90.250 34.135 90.585 35.105 ;
        RECT 90.755 34.135 90.925 35.275 ;
        RECT 91.095 34.935 93.125 35.105 ;
        RECT 90.250 33.465 90.420 34.135 ;
        RECT 91.095 33.965 91.265 34.935 ;
        RECT 90.590 33.635 90.845 33.965 ;
        RECT 91.070 33.635 91.265 33.965 ;
        RECT 91.435 34.595 92.560 34.765 ;
        RECT 90.675 33.465 90.845 33.635 ;
        RECT 91.435 33.465 91.605 34.595 ;
        RECT 71.705 32.935 72.595 33.105 ;
        RECT 72.765 32.725 78.110 33.270 ;
        RECT 78.285 32.725 83.630 33.270 ;
        RECT 83.805 32.725 89.150 33.270 ;
        RECT 90.250 32.895 90.505 33.465 ;
        RECT 90.675 33.295 91.605 33.465 ;
        RECT 91.775 34.255 92.785 34.425 ;
        RECT 91.775 33.455 91.945 34.255 ;
        RECT 91.430 33.260 91.605 33.295 ;
        RECT 90.675 32.725 91.005 33.125 ;
        RECT 91.430 32.895 91.960 33.260 ;
        RECT 92.150 33.235 92.425 34.055 ;
        RECT 92.145 33.065 92.425 33.235 ;
        RECT 92.150 32.895 92.425 33.065 ;
        RECT 92.595 32.895 92.785 34.255 ;
        RECT 92.955 34.270 93.125 34.935 ;
        RECT 93.295 34.515 93.465 35.275 ;
        RECT 93.700 34.515 94.215 34.925 ;
        RECT 92.955 34.080 93.705 34.270 ;
        RECT 93.875 33.705 94.215 34.515 ;
        RECT 94.475 34.345 94.645 35.105 ;
        RECT 94.825 34.515 95.155 35.275 ;
        RECT 94.475 34.175 95.140 34.345 ;
        RECT 95.325 34.200 95.595 35.105 ;
        RECT 94.970 34.030 95.140 34.175 ;
        RECT 92.985 33.535 94.215 33.705 ;
        RECT 94.405 33.625 94.735 33.995 ;
        RECT 94.970 33.700 95.255 34.030 ;
        RECT 92.965 32.725 93.475 33.260 ;
        RECT 93.695 32.930 93.940 33.535 ;
        RECT 94.970 33.445 95.140 33.700 ;
        RECT 94.475 33.275 95.140 33.445 ;
        RECT 95.425 33.400 95.595 34.200 ;
        RECT 95.765 34.110 96.055 35.275 ;
        RECT 96.315 34.605 96.485 35.105 ;
        RECT 96.655 34.775 96.985 35.275 ;
        RECT 96.315 34.435 96.980 34.605 ;
        RECT 96.230 33.615 96.580 34.265 ;
        RECT 94.475 32.895 94.645 33.275 ;
        RECT 94.825 32.725 95.155 33.105 ;
        RECT 95.335 32.895 95.595 33.400 ;
        RECT 95.765 32.725 96.055 33.450 ;
        RECT 96.750 33.445 96.980 34.435 ;
        RECT 96.315 33.275 96.980 33.445 ;
        RECT 96.315 32.985 96.485 33.275 ;
        RECT 96.655 32.725 96.985 33.105 ;
        RECT 97.155 32.985 97.380 35.105 ;
        RECT 97.595 34.775 97.925 35.275 ;
        RECT 98.095 34.605 98.265 35.105 ;
        RECT 98.500 34.890 99.330 35.060 ;
        RECT 99.570 34.895 99.950 35.275 ;
        RECT 97.570 34.435 98.265 34.605 ;
        RECT 97.570 33.465 97.740 34.435 ;
        RECT 97.910 33.645 98.320 34.265 ;
        RECT 98.490 34.215 98.990 34.595 ;
        RECT 97.570 33.275 98.265 33.465 ;
        RECT 98.490 33.345 98.710 34.215 ;
        RECT 99.160 34.045 99.330 34.890 ;
        RECT 100.130 34.725 100.300 35.015 ;
        RECT 100.470 34.895 100.800 35.275 ;
        RECT 101.270 34.805 101.900 35.055 ;
        RECT 102.080 34.895 102.500 35.275 ;
        RECT 101.730 34.725 101.900 34.805 ;
        RECT 102.700 34.725 102.940 35.015 ;
        RECT 99.500 34.475 100.870 34.725 ;
        RECT 99.500 34.215 99.750 34.475 ;
        RECT 100.260 34.045 100.510 34.205 ;
        RECT 99.160 33.875 100.510 34.045 ;
        RECT 99.160 33.835 99.580 33.875 ;
        RECT 98.890 33.285 99.240 33.655 ;
        RECT 97.595 32.725 97.925 33.105 ;
        RECT 98.095 32.945 98.265 33.275 ;
        RECT 99.410 33.105 99.580 33.835 ;
        RECT 100.680 33.705 100.870 34.475 ;
        RECT 99.750 33.375 100.160 33.705 ;
        RECT 100.450 33.365 100.870 33.705 ;
        RECT 101.040 34.295 101.560 34.605 ;
        RECT 101.730 34.555 102.940 34.725 ;
        RECT 103.170 34.585 103.500 35.275 ;
        RECT 101.040 33.535 101.210 34.295 ;
        RECT 101.380 33.705 101.560 34.115 ;
        RECT 101.730 34.045 101.900 34.555 ;
        RECT 103.670 34.405 103.840 35.015 ;
        RECT 104.110 34.555 104.440 35.065 ;
        RECT 103.670 34.385 103.990 34.405 ;
        RECT 102.070 34.215 103.990 34.385 ;
        RECT 101.730 33.875 103.630 34.045 ;
        RECT 101.960 33.535 102.290 33.655 ;
        RECT 101.040 33.365 102.290 33.535 ;
        RECT 98.565 32.905 99.580 33.105 ;
        RECT 99.750 32.725 100.160 33.165 ;
        RECT 100.450 32.935 100.700 33.365 ;
        RECT 100.900 32.725 101.220 33.185 ;
        RECT 102.460 33.115 102.630 33.875 ;
        RECT 103.300 33.815 103.630 33.875 ;
        RECT 102.820 33.645 103.150 33.705 ;
        RECT 102.820 33.375 103.480 33.645 ;
        RECT 103.800 33.320 103.990 34.215 ;
        RECT 101.780 32.945 102.630 33.115 ;
        RECT 102.830 32.725 103.490 33.205 ;
        RECT 103.670 32.990 103.990 33.320 ;
        RECT 104.190 33.965 104.440 34.555 ;
        RECT 104.620 34.475 104.905 35.275 ;
        RECT 105.085 34.295 105.340 34.965 ;
        RECT 105.885 34.840 111.230 35.275 ;
        RECT 111.405 34.840 116.750 35.275 ;
        RECT 105.160 34.255 105.340 34.295 ;
        RECT 105.160 34.085 105.425 34.255 ;
        RECT 104.190 33.635 104.990 33.965 ;
        RECT 104.190 32.985 104.440 33.635 ;
        RECT 105.160 33.435 105.340 34.085 ;
        RECT 104.620 32.725 104.905 33.185 ;
        RECT 105.085 32.905 105.340 33.435 ;
        RECT 107.470 33.270 107.810 34.100 ;
        RECT 109.290 33.590 109.640 34.840 ;
        RECT 112.990 33.270 113.330 34.100 ;
        RECT 114.810 33.590 115.160 34.840 ;
        RECT 116.925 34.185 120.435 35.275 ;
        RECT 116.925 33.495 118.575 34.015 ;
        RECT 118.745 33.665 120.435 34.185 ;
        RECT 121.525 34.110 121.815 35.275 ;
        RECT 122.445 34.185 123.655 35.275 ;
        RECT 122.445 33.645 122.965 34.185 ;
        RECT 105.885 32.725 111.230 33.270 ;
        RECT 111.405 32.725 116.750 33.270 ;
        RECT 116.925 32.725 120.435 33.495 ;
        RECT 123.135 33.475 123.655 34.015 ;
        RECT 121.525 32.725 121.815 33.450 ;
        RECT 122.445 32.725 123.655 33.475 ;
        RECT 5.520 32.555 123.740 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.985 31.785 8.655 32.555 ;
        RECT 9.290 32.005 9.545 32.295 ;
        RECT 9.715 32.175 10.045 32.555 ;
        RECT 9.290 31.835 10.040 32.005 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 6.985 31.265 7.735 31.785 ;
        RECT 7.905 31.095 8.655 31.615 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 6.985 30.005 8.655 31.095 ;
        RECT 9.290 31.015 9.640 31.665 ;
        RECT 9.810 30.845 10.040 31.835 ;
        RECT 9.290 30.675 10.040 30.845 ;
        RECT 9.290 30.175 9.545 30.675 ;
        RECT 9.715 30.005 10.045 30.505 ;
        RECT 10.215 30.175 10.385 32.295 ;
        RECT 10.745 32.195 11.075 32.555 ;
        RECT 11.245 32.165 11.740 32.335 ;
        RECT 11.945 32.165 12.800 32.335 ;
        RECT 10.615 30.975 11.075 32.025 ;
        RECT 10.555 30.190 10.880 30.975 ;
        RECT 11.245 30.805 11.415 32.165 ;
        RECT 11.585 31.255 11.935 31.875 ;
        RECT 12.105 31.655 12.460 31.875 ;
        RECT 12.105 31.065 12.275 31.655 ;
        RECT 12.630 31.455 12.800 32.165 ;
        RECT 13.675 32.095 14.005 32.555 ;
        RECT 14.215 32.195 14.565 32.365 ;
        RECT 13.005 31.625 13.795 31.875 ;
        RECT 14.215 31.805 14.475 32.195 ;
        RECT 14.785 32.105 15.735 32.385 ;
        RECT 15.905 32.115 16.095 32.555 ;
        RECT 16.265 32.175 17.335 32.345 ;
        RECT 13.965 31.455 14.135 31.635 ;
        RECT 11.245 30.635 11.640 30.805 ;
        RECT 11.810 30.675 12.275 31.065 ;
        RECT 12.445 31.285 14.135 31.455 ;
        RECT 11.470 30.505 11.640 30.635 ;
        RECT 12.445 30.505 12.615 31.285 ;
        RECT 14.305 31.115 14.475 31.805 ;
        RECT 12.975 30.945 14.475 31.115 ;
        RECT 14.665 31.145 14.875 31.935 ;
        RECT 15.045 31.315 15.395 31.935 ;
        RECT 15.565 31.325 15.735 32.105 ;
        RECT 16.265 31.945 16.435 32.175 ;
        RECT 15.905 31.775 16.435 31.945 ;
        RECT 15.905 31.495 16.125 31.775 ;
        RECT 16.605 31.605 16.845 32.005 ;
        RECT 15.565 31.155 15.970 31.325 ;
        RECT 16.305 31.235 16.845 31.605 ;
        RECT 17.015 31.820 17.335 32.175 ;
        RECT 17.580 32.095 17.885 32.555 ;
        RECT 18.055 31.845 18.310 32.375 ;
        RECT 17.015 31.645 17.340 31.820 ;
        RECT 17.015 31.345 17.930 31.645 ;
        RECT 17.190 31.315 17.930 31.345 ;
        RECT 14.665 30.985 15.340 31.145 ;
        RECT 15.800 31.065 15.970 31.155 ;
        RECT 14.665 30.975 15.630 30.985 ;
        RECT 14.305 30.805 14.475 30.945 ;
        RECT 11.050 30.005 11.300 30.465 ;
        RECT 11.470 30.175 11.720 30.505 ;
        RECT 11.935 30.175 12.615 30.505 ;
        RECT 12.785 30.605 13.860 30.775 ;
        RECT 14.305 30.635 14.865 30.805 ;
        RECT 15.170 30.685 15.630 30.975 ;
        RECT 15.800 30.895 17.020 31.065 ;
        RECT 12.785 30.265 12.955 30.605 ;
        RECT 13.190 30.005 13.520 30.435 ;
        RECT 13.690 30.265 13.860 30.605 ;
        RECT 14.155 30.005 14.525 30.465 ;
        RECT 14.695 30.175 14.865 30.635 ;
        RECT 15.800 30.515 15.970 30.895 ;
        RECT 17.190 30.725 17.360 31.315 ;
        RECT 18.100 31.195 18.310 31.845 ;
        RECT 18.490 32.005 18.745 32.295 ;
        RECT 18.915 32.175 19.245 32.555 ;
        RECT 18.490 31.835 19.240 32.005 ;
        RECT 15.100 30.175 15.970 30.515 ;
        RECT 16.560 30.555 17.360 30.725 ;
        RECT 16.140 30.005 16.390 30.465 ;
        RECT 16.560 30.265 16.730 30.555 ;
        RECT 16.910 30.005 17.240 30.385 ;
        RECT 17.580 30.005 17.885 31.145 ;
        RECT 18.055 30.315 18.310 31.195 ;
        RECT 18.490 31.015 18.840 31.665 ;
        RECT 19.010 30.845 19.240 31.835 ;
        RECT 18.490 30.675 19.240 30.845 ;
        RECT 18.490 30.175 18.745 30.675 ;
        RECT 18.915 30.005 19.245 30.505 ;
        RECT 19.415 30.175 19.585 32.295 ;
        RECT 19.945 32.195 20.275 32.555 ;
        RECT 20.445 32.165 20.940 32.335 ;
        RECT 21.145 32.165 22.000 32.335 ;
        RECT 19.815 30.975 20.275 32.025 ;
        RECT 19.755 30.190 20.080 30.975 ;
        RECT 20.445 30.805 20.615 32.165 ;
        RECT 20.785 31.255 21.135 31.875 ;
        RECT 21.305 31.655 21.660 31.875 ;
        RECT 21.305 31.065 21.475 31.655 ;
        RECT 21.830 31.455 22.000 32.165 ;
        RECT 22.875 32.095 23.205 32.555 ;
        RECT 23.415 32.195 23.765 32.365 ;
        RECT 22.205 31.625 22.995 31.875 ;
        RECT 23.415 31.805 23.675 32.195 ;
        RECT 23.985 32.105 24.935 32.385 ;
        RECT 25.105 32.115 25.295 32.555 ;
        RECT 25.465 32.175 26.535 32.345 ;
        RECT 23.165 31.455 23.335 31.635 ;
        RECT 20.445 30.635 20.840 30.805 ;
        RECT 21.010 30.675 21.475 31.065 ;
        RECT 21.645 31.285 23.335 31.455 ;
        RECT 20.670 30.505 20.840 30.635 ;
        RECT 21.645 30.505 21.815 31.285 ;
        RECT 23.505 31.115 23.675 31.805 ;
        RECT 22.175 30.945 23.675 31.115 ;
        RECT 23.865 31.145 24.075 31.935 ;
        RECT 24.245 31.315 24.595 31.935 ;
        RECT 24.765 31.325 24.935 32.105 ;
        RECT 25.465 31.945 25.635 32.175 ;
        RECT 25.105 31.775 25.635 31.945 ;
        RECT 25.105 31.495 25.325 31.775 ;
        RECT 25.805 31.605 26.045 32.005 ;
        RECT 24.765 31.155 25.170 31.325 ;
        RECT 25.505 31.235 26.045 31.605 ;
        RECT 26.215 31.820 26.535 32.175 ;
        RECT 26.780 32.095 27.085 32.555 ;
        RECT 27.255 31.845 27.510 32.375 ;
        RECT 26.215 31.645 26.540 31.820 ;
        RECT 26.215 31.345 27.130 31.645 ;
        RECT 26.390 31.315 27.130 31.345 ;
        RECT 23.865 30.985 24.540 31.145 ;
        RECT 25.000 31.065 25.170 31.155 ;
        RECT 23.865 30.975 24.830 30.985 ;
        RECT 23.505 30.805 23.675 30.945 ;
        RECT 20.250 30.005 20.500 30.465 ;
        RECT 20.670 30.175 20.920 30.505 ;
        RECT 21.135 30.175 21.815 30.505 ;
        RECT 21.985 30.605 23.060 30.775 ;
        RECT 23.505 30.635 24.065 30.805 ;
        RECT 24.370 30.685 24.830 30.975 ;
        RECT 25.000 30.895 26.220 31.065 ;
        RECT 21.985 30.265 22.155 30.605 ;
        RECT 22.390 30.005 22.720 30.435 ;
        RECT 22.890 30.265 23.060 30.605 ;
        RECT 23.355 30.005 23.725 30.465 ;
        RECT 23.895 30.175 24.065 30.635 ;
        RECT 25.000 30.515 25.170 30.895 ;
        RECT 26.390 30.725 26.560 31.315 ;
        RECT 27.300 31.195 27.510 31.845 ;
        RECT 24.300 30.175 25.170 30.515 ;
        RECT 25.760 30.555 26.560 30.725 ;
        RECT 25.340 30.005 25.590 30.465 ;
        RECT 25.760 30.265 25.930 30.555 ;
        RECT 26.110 30.005 26.440 30.385 ;
        RECT 26.780 30.005 27.085 31.145 ;
        RECT 27.255 30.315 27.510 31.195 ;
        RECT 28.145 31.880 28.405 32.385 ;
        RECT 28.585 32.175 28.915 32.555 ;
        RECT 29.095 32.005 29.265 32.385 ;
        RECT 28.145 31.080 28.315 31.880 ;
        RECT 28.600 31.835 29.265 32.005 ;
        RECT 28.600 31.580 28.770 31.835 ;
        RECT 29.525 31.785 31.195 32.555 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 31.830 31.815 32.085 32.385 ;
        RECT 32.255 32.155 32.585 32.555 ;
        RECT 33.010 32.020 33.540 32.385 ;
        RECT 33.010 31.985 33.185 32.020 ;
        RECT 32.255 31.815 33.185 31.985 ;
        RECT 33.730 31.875 34.005 32.385 ;
        RECT 28.485 31.250 28.770 31.580 ;
        RECT 29.005 31.285 29.335 31.655 ;
        RECT 29.525 31.265 30.275 31.785 ;
        RECT 28.600 31.105 28.770 31.250 ;
        RECT 28.145 30.175 28.415 31.080 ;
        RECT 28.600 30.935 29.265 31.105 ;
        RECT 30.445 31.095 31.195 31.615 ;
        RECT 28.585 30.005 28.915 30.765 ;
        RECT 29.095 30.175 29.265 30.935 ;
        RECT 29.525 30.005 31.195 31.095 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 31.830 31.145 32.000 31.815 ;
        RECT 32.255 31.645 32.425 31.815 ;
        RECT 32.170 31.315 32.425 31.645 ;
        RECT 32.650 31.315 32.845 31.645 ;
        RECT 31.830 30.175 32.165 31.145 ;
        RECT 32.335 30.005 32.505 31.145 ;
        RECT 32.675 30.345 32.845 31.315 ;
        RECT 33.015 30.685 33.185 31.815 ;
        RECT 33.355 31.025 33.525 31.825 ;
        RECT 33.725 31.705 34.005 31.875 ;
        RECT 33.730 31.225 34.005 31.705 ;
        RECT 34.175 31.025 34.365 32.385 ;
        RECT 34.545 32.020 35.055 32.555 ;
        RECT 35.275 31.745 35.520 32.350 ;
        RECT 35.965 31.785 38.555 32.555 ;
        RECT 38.815 32.005 38.985 32.295 ;
        RECT 39.155 32.175 39.485 32.555 ;
        RECT 38.815 31.835 39.480 32.005 ;
        RECT 34.565 31.575 35.795 31.745 ;
        RECT 33.355 30.855 34.365 31.025 ;
        RECT 34.535 31.010 35.285 31.200 ;
        RECT 33.015 30.515 34.140 30.685 ;
        RECT 34.535 30.345 34.705 31.010 ;
        RECT 35.455 30.765 35.795 31.575 ;
        RECT 35.965 31.265 37.175 31.785 ;
        RECT 37.345 31.095 38.555 31.615 ;
        RECT 32.675 30.175 34.705 30.345 ;
        RECT 34.875 30.005 35.045 30.765 ;
        RECT 35.280 30.355 35.795 30.765 ;
        RECT 35.965 30.005 38.555 31.095 ;
        RECT 38.730 31.015 39.080 31.665 ;
        RECT 39.250 30.845 39.480 31.835 ;
        RECT 38.815 30.675 39.480 30.845 ;
        RECT 38.815 30.175 38.985 30.675 ;
        RECT 39.155 30.005 39.485 30.505 ;
        RECT 39.655 30.175 39.880 32.295 ;
        RECT 40.095 32.175 40.425 32.555 ;
        RECT 40.595 32.005 40.765 32.335 ;
        RECT 41.065 32.175 42.080 32.375 ;
        RECT 40.070 31.815 40.765 32.005 ;
        RECT 40.070 30.845 40.240 31.815 ;
        RECT 40.410 31.015 40.820 31.635 ;
        RECT 40.990 31.065 41.210 31.935 ;
        RECT 41.390 31.625 41.740 31.995 ;
        RECT 41.910 31.445 42.080 32.175 ;
        RECT 42.250 32.115 42.660 32.555 ;
        RECT 42.950 31.915 43.200 32.345 ;
        RECT 43.400 32.095 43.720 32.555 ;
        RECT 44.280 32.165 45.130 32.335 ;
        RECT 42.250 31.575 42.660 31.905 ;
        RECT 42.950 31.575 43.370 31.915 ;
        RECT 41.660 31.405 42.080 31.445 ;
        RECT 41.660 31.235 43.010 31.405 ;
        RECT 40.070 30.675 40.765 30.845 ;
        RECT 40.990 30.685 41.490 31.065 ;
        RECT 40.095 30.005 40.425 30.505 ;
        RECT 40.595 30.175 40.765 30.675 ;
        RECT 41.660 30.390 41.830 31.235 ;
        RECT 42.760 31.075 43.010 31.235 ;
        RECT 42.000 30.805 42.250 31.065 ;
        RECT 43.180 30.805 43.370 31.575 ;
        RECT 42.000 30.555 43.370 30.805 ;
        RECT 43.540 31.745 44.790 31.915 ;
        RECT 43.540 30.985 43.710 31.745 ;
        RECT 44.460 31.625 44.790 31.745 ;
        RECT 43.880 31.165 44.060 31.575 ;
        RECT 44.960 31.405 45.130 32.165 ;
        RECT 45.330 32.075 45.990 32.555 ;
        RECT 46.170 31.960 46.490 32.290 ;
        RECT 45.320 31.635 45.980 31.905 ;
        RECT 45.320 31.575 45.650 31.635 ;
        RECT 45.800 31.405 46.130 31.465 ;
        RECT 44.230 31.235 46.130 31.405 ;
        RECT 43.540 30.675 44.060 30.985 ;
        RECT 44.230 30.725 44.400 31.235 ;
        RECT 46.300 31.065 46.490 31.960 ;
        RECT 44.570 30.895 46.490 31.065 ;
        RECT 46.170 30.875 46.490 30.895 ;
        RECT 46.690 31.645 46.940 32.295 ;
        RECT 47.120 32.095 47.405 32.555 ;
        RECT 47.585 32.215 47.840 32.375 ;
        RECT 47.585 32.045 47.925 32.215 ;
        RECT 47.585 31.845 47.840 32.045 ;
        RECT 48.385 32.010 53.730 32.555 ;
        RECT 46.690 31.315 47.490 31.645 ;
        RECT 44.230 30.555 45.440 30.725 ;
        RECT 41.000 30.220 41.830 30.390 ;
        RECT 42.070 30.005 42.450 30.385 ;
        RECT 42.630 30.265 42.800 30.555 ;
        RECT 44.230 30.475 44.400 30.555 ;
        RECT 42.970 30.005 43.300 30.385 ;
        RECT 43.770 30.225 44.400 30.475 ;
        RECT 44.580 30.005 45.000 30.385 ;
        RECT 45.200 30.265 45.440 30.555 ;
        RECT 45.670 30.005 46.000 30.695 ;
        RECT 46.170 30.265 46.340 30.875 ;
        RECT 46.690 30.725 46.940 31.315 ;
        RECT 47.660 30.985 47.840 31.845 ;
        RECT 49.970 31.180 50.310 32.010 ;
        RECT 53.905 31.785 56.495 32.555 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 57.585 31.815 57.905 32.295 ;
        RECT 58.075 31.985 58.305 32.385 ;
        RECT 58.475 32.165 58.825 32.555 ;
        RECT 58.075 31.905 58.585 31.985 ;
        RECT 58.995 31.905 59.325 32.385 ;
        RECT 58.075 31.815 59.325 31.905 ;
        RECT 46.610 30.215 46.940 30.725 ;
        RECT 47.120 30.005 47.405 30.805 ;
        RECT 47.585 30.315 47.840 30.985 ;
        RECT 51.790 30.440 52.140 31.690 ;
        RECT 53.905 31.265 55.115 31.785 ;
        RECT 55.285 31.095 56.495 31.615 ;
        RECT 48.385 30.005 53.730 30.440 ;
        RECT 53.905 30.005 56.495 31.095 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 57.585 30.885 57.755 31.815 ;
        RECT 58.415 31.735 59.325 31.815 ;
        RECT 59.495 31.735 59.665 32.555 ;
        RECT 60.170 31.815 60.635 32.360 ;
        RECT 57.925 31.225 58.095 31.645 ;
        RECT 58.325 31.395 58.925 31.565 ;
        RECT 57.925 31.055 58.585 31.225 ;
        RECT 57.585 30.685 58.245 30.885 ;
        RECT 58.415 30.855 58.585 31.055 ;
        RECT 58.755 31.195 58.925 31.395 ;
        RECT 59.095 31.365 59.790 31.565 ;
        RECT 60.050 31.195 60.295 31.645 ;
        RECT 58.755 31.025 60.295 31.195 ;
        RECT 60.465 30.855 60.635 31.815 ;
        RECT 60.810 31.715 61.070 32.555 ;
        RECT 61.245 31.810 61.500 32.385 ;
        RECT 61.670 32.175 62.000 32.555 ;
        RECT 62.215 32.005 62.385 32.385 ;
        RECT 61.670 31.835 62.385 32.005 ;
        RECT 58.415 30.685 60.635 30.855 ;
        RECT 58.075 30.515 58.245 30.685 ;
        RECT 57.605 30.005 57.905 30.515 ;
        RECT 58.075 30.345 58.455 30.515 ;
        RECT 59.035 30.005 59.665 30.515 ;
        RECT 59.835 30.175 60.165 30.685 ;
        RECT 60.335 30.005 60.635 30.515 ;
        RECT 60.810 30.005 61.070 31.155 ;
        RECT 61.245 31.080 61.415 31.810 ;
        RECT 61.670 31.645 61.840 31.835 ;
        RECT 62.645 31.785 65.235 32.555 ;
        RECT 65.955 32.005 66.125 32.385 ;
        RECT 66.305 32.175 66.635 32.555 ;
        RECT 65.955 31.835 66.620 32.005 ;
        RECT 66.815 31.880 67.075 32.385 ;
        RECT 61.585 31.315 61.840 31.645 ;
        RECT 61.670 31.105 61.840 31.315 ;
        RECT 62.120 31.285 62.475 31.655 ;
        RECT 62.645 31.265 63.855 31.785 ;
        RECT 61.245 30.175 61.500 31.080 ;
        RECT 61.670 30.935 62.385 31.105 ;
        RECT 64.025 31.095 65.235 31.615 ;
        RECT 65.885 31.285 66.215 31.655 ;
        RECT 66.450 31.580 66.620 31.835 ;
        RECT 66.450 31.250 66.735 31.580 ;
        RECT 66.450 31.105 66.620 31.250 ;
        RECT 61.670 30.005 62.000 30.765 ;
        RECT 62.215 30.175 62.385 30.935 ;
        RECT 62.645 30.005 65.235 31.095 ;
        RECT 65.955 30.935 66.620 31.105 ;
        RECT 66.905 31.080 67.075 31.880 ;
        RECT 67.250 32.005 67.505 32.295 ;
        RECT 67.675 32.175 68.005 32.555 ;
        RECT 67.250 31.835 68.000 32.005 ;
        RECT 65.955 30.175 66.125 30.935 ;
        RECT 66.305 30.005 66.635 30.765 ;
        RECT 66.805 30.175 67.075 31.080 ;
        RECT 67.250 31.015 67.600 31.665 ;
        RECT 67.770 30.845 68.000 31.835 ;
        RECT 67.250 30.675 68.000 30.845 ;
        RECT 67.250 30.175 67.505 30.675 ;
        RECT 67.675 30.005 68.005 30.505 ;
        RECT 68.175 30.175 68.345 32.295 ;
        RECT 68.705 32.195 69.035 32.555 ;
        RECT 69.205 32.165 69.700 32.335 ;
        RECT 69.905 32.165 70.760 32.335 ;
        RECT 68.575 30.975 69.035 32.025 ;
        RECT 68.515 30.190 68.840 30.975 ;
        RECT 69.205 30.805 69.375 32.165 ;
        RECT 69.545 31.255 69.895 31.875 ;
        RECT 70.065 31.655 70.420 31.875 ;
        RECT 70.065 31.065 70.235 31.655 ;
        RECT 70.590 31.455 70.760 32.165 ;
        RECT 71.635 32.095 71.965 32.555 ;
        RECT 72.175 32.195 72.525 32.365 ;
        RECT 70.965 31.625 71.755 31.875 ;
        RECT 72.175 31.805 72.435 32.195 ;
        RECT 72.745 32.105 73.695 32.385 ;
        RECT 73.865 32.115 74.055 32.555 ;
        RECT 74.225 32.175 75.295 32.345 ;
        RECT 71.925 31.455 72.095 31.635 ;
        RECT 69.205 30.635 69.600 30.805 ;
        RECT 69.770 30.675 70.235 31.065 ;
        RECT 70.405 31.285 72.095 31.455 ;
        RECT 69.430 30.505 69.600 30.635 ;
        RECT 70.405 30.505 70.575 31.285 ;
        RECT 72.265 31.115 72.435 31.805 ;
        RECT 70.935 30.945 72.435 31.115 ;
        RECT 72.625 31.145 72.835 31.935 ;
        RECT 73.005 31.315 73.355 31.935 ;
        RECT 73.525 31.325 73.695 32.105 ;
        RECT 74.225 31.945 74.395 32.175 ;
        RECT 73.865 31.775 74.395 31.945 ;
        RECT 73.865 31.495 74.085 31.775 ;
        RECT 74.565 31.605 74.805 32.005 ;
        RECT 73.525 31.155 73.930 31.325 ;
        RECT 74.265 31.235 74.805 31.605 ;
        RECT 74.975 31.820 75.295 32.175 ;
        RECT 74.975 31.565 75.300 31.820 ;
        RECT 75.495 31.745 75.665 32.555 ;
        RECT 75.835 31.905 76.165 32.385 ;
        RECT 76.335 32.085 76.505 32.555 ;
        RECT 76.675 31.905 77.005 32.385 ;
        RECT 77.175 32.085 77.345 32.555 ;
        RECT 75.835 31.735 77.600 31.905 ;
        RECT 74.975 31.355 77.005 31.565 ;
        RECT 74.975 31.345 75.320 31.355 ;
        RECT 72.625 30.985 73.300 31.145 ;
        RECT 73.760 31.065 73.930 31.155 ;
        RECT 72.625 30.975 73.590 30.985 ;
        RECT 72.265 30.805 72.435 30.945 ;
        RECT 69.010 30.005 69.260 30.465 ;
        RECT 69.430 30.175 69.680 30.505 ;
        RECT 69.895 30.175 70.575 30.505 ;
        RECT 70.745 30.605 71.820 30.775 ;
        RECT 72.265 30.635 72.825 30.805 ;
        RECT 73.130 30.685 73.590 30.975 ;
        RECT 73.760 30.895 74.980 31.065 ;
        RECT 70.745 30.265 70.915 30.605 ;
        RECT 71.150 30.005 71.480 30.435 ;
        RECT 71.650 30.265 71.820 30.605 ;
        RECT 72.115 30.005 72.485 30.465 ;
        RECT 72.655 30.175 72.825 30.635 ;
        RECT 73.760 30.515 73.930 30.895 ;
        RECT 75.150 30.725 75.320 31.345 ;
        RECT 77.190 31.185 77.600 31.735 ;
        RECT 77.825 31.785 79.495 32.555 ;
        RECT 79.665 31.880 79.925 32.385 ;
        RECT 80.105 32.175 80.435 32.555 ;
        RECT 80.615 32.005 80.785 32.385 ;
        RECT 77.825 31.265 78.575 31.785 ;
        RECT 73.060 30.175 73.930 30.515 ;
        RECT 74.520 30.555 75.320 30.725 ;
        RECT 74.100 30.005 74.350 30.465 ;
        RECT 74.520 30.265 74.690 30.555 ;
        RECT 74.870 30.005 75.200 30.385 ;
        RECT 75.495 30.005 75.665 31.065 ;
        RECT 75.875 31.015 77.600 31.185 ;
        RECT 78.745 31.095 79.495 31.615 ;
        RECT 75.875 30.175 76.165 31.015 ;
        RECT 76.335 30.005 76.505 30.845 ;
        RECT 76.715 30.175 76.965 31.015 ;
        RECT 77.175 30.005 77.345 30.845 ;
        RECT 77.825 30.005 79.495 31.095 ;
        RECT 79.665 31.080 79.835 31.880 ;
        RECT 80.120 31.835 80.785 32.005 ;
        RECT 80.120 31.580 80.290 31.835 ;
        RECT 81.545 31.735 81.775 32.555 ;
        RECT 81.945 31.755 82.275 32.385 ;
        RECT 80.005 31.250 80.290 31.580 ;
        RECT 80.525 31.285 80.855 31.655 ;
        RECT 81.525 31.315 81.855 31.565 ;
        RECT 80.120 31.105 80.290 31.250 ;
        RECT 82.025 31.155 82.275 31.755 ;
        RECT 82.445 31.735 82.655 32.555 ;
        RECT 82.885 31.830 83.175 32.555 ;
        RECT 83.350 31.815 83.605 32.385 ;
        RECT 83.775 32.155 84.105 32.555 ;
        RECT 84.530 32.020 85.060 32.385 ;
        RECT 84.530 31.985 84.705 32.020 ;
        RECT 83.775 31.815 84.705 31.985 ;
        RECT 85.250 31.875 85.525 32.385 ;
        RECT 79.665 30.175 79.935 31.080 ;
        RECT 80.120 30.935 80.785 31.105 ;
        RECT 80.105 30.005 80.435 30.765 ;
        RECT 80.615 30.175 80.785 30.935 ;
        RECT 81.545 30.005 81.775 31.145 ;
        RECT 81.945 30.175 82.275 31.155 ;
        RECT 82.445 30.005 82.655 31.145 ;
        RECT 82.885 30.005 83.175 31.170 ;
        RECT 83.350 31.145 83.520 31.815 ;
        RECT 83.775 31.645 83.945 31.815 ;
        RECT 83.690 31.315 83.945 31.645 ;
        RECT 84.170 31.315 84.365 31.645 ;
        RECT 83.350 30.175 83.685 31.145 ;
        RECT 83.855 30.005 84.025 31.145 ;
        RECT 84.195 30.345 84.365 31.315 ;
        RECT 84.535 30.685 84.705 31.815 ;
        RECT 84.875 31.025 85.045 31.825 ;
        RECT 85.245 31.705 85.525 31.875 ;
        RECT 85.250 31.225 85.525 31.705 ;
        RECT 85.695 31.025 85.885 32.385 ;
        RECT 86.065 32.020 86.575 32.555 ;
        RECT 86.795 31.745 87.040 32.350 ;
        RECT 86.085 31.575 87.315 31.745 ;
        RECT 87.525 31.735 87.755 32.555 ;
        RECT 87.925 31.755 88.255 32.385 ;
        RECT 84.875 30.855 85.885 31.025 ;
        RECT 86.055 31.010 86.805 31.200 ;
        RECT 84.535 30.515 85.660 30.685 ;
        RECT 86.055 30.345 86.225 31.010 ;
        RECT 86.975 30.765 87.315 31.575 ;
        RECT 87.505 31.315 87.835 31.565 ;
        RECT 88.005 31.155 88.255 31.755 ;
        RECT 88.425 31.735 88.635 32.555 ;
        RECT 88.955 32.005 89.125 32.385 ;
        RECT 89.305 32.175 89.635 32.555 ;
        RECT 88.955 31.835 89.620 32.005 ;
        RECT 89.815 31.880 90.075 32.385 ;
        RECT 88.885 31.285 89.215 31.655 ;
        RECT 89.450 31.580 89.620 31.835 ;
        RECT 84.195 30.175 86.225 30.345 ;
        RECT 86.395 30.005 86.565 30.765 ;
        RECT 86.800 30.355 87.315 30.765 ;
        RECT 87.525 30.005 87.755 31.145 ;
        RECT 87.925 30.175 88.255 31.155 ;
        RECT 89.450 31.250 89.735 31.580 ;
        RECT 88.425 30.005 88.635 31.145 ;
        RECT 89.450 31.105 89.620 31.250 ;
        RECT 88.955 30.935 89.620 31.105 ;
        RECT 89.905 31.080 90.075 31.880 ;
        RECT 90.245 31.785 93.755 32.555 ;
        RECT 94.850 31.815 95.105 32.385 ;
        RECT 95.275 32.155 95.605 32.555 ;
        RECT 96.030 32.020 96.560 32.385 ;
        RECT 96.030 31.985 96.205 32.020 ;
        RECT 95.275 31.815 96.205 31.985 ;
        RECT 96.750 31.875 97.025 32.385 ;
        RECT 90.245 31.265 91.895 31.785 ;
        RECT 92.065 31.095 93.755 31.615 ;
        RECT 88.955 30.175 89.125 30.935 ;
        RECT 89.305 30.005 89.635 30.765 ;
        RECT 89.805 30.175 90.075 31.080 ;
        RECT 90.245 30.005 93.755 31.095 ;
        RECT 94.850 31.145 95.020 31.815 ;
        RECT 95.275 31.645 95.445 31.815 ;
        RECT 95.190 31.315 95.445 31.645 ;
        RECT 95.670 31.315 95.865 31.645 ;
        RECT 94.850 30.175 95.185 31.145 ;
        RECT 95.355 30.005 95.525 31.145 ;
        RECT 95.695 30.345 95.865 31.315 ;
        RECT 96.035 30.685 96.205 31.815 ;
        RECT 96.375 31.025 96.545 31.825 ;
        RECT 96.745 31.705 97.025 31.875 ;
        RECT 96.750 31.225 97.025 31.705 ;
        RECT 97.195 31.025 97.385 32.385 ;
        RECT 97.565 32.020 98.075 32.555 ;
        RECT 98.295 31.745 98.540 32.350 ;
        RECT 98.985 32.010 104.330 32.555 ;
        RECT 97.585 31.575 98.815 31.745 ;
        RECT 96.375 30.855 97.385 31.025 ;
        RECT 97.555 31.010 98.305 31.200 ;
        RECT 96.035 30.515 97.160 30.685 ;
        RECT 97.555 30.345 97.725 31.010 ;
        RECT 98.475 30.765 98.815 31.575 ;
        RECT 100.570 31.180 100.910 32.010 ;
        RECT 104.505 31.785 108.015 32.555 ;
        RECT 108.645 31.830 108.935 32.555 ;
        RECT 109.105 32.010 114.450 32.555 ;
        RECT 114.625 32.010 119.970 32.555 ;
        RECT 95.695 30.175 97.725 30.345 ;
        RECT 97.895 30.005 98.065 30.765 ;
        RECT 98.300 30.355 98.815 30.765 ;
        RECT 102.390 30.440 102.740 31.690 ;
        RECT 104.505 31.265 106.155 31.785 ;
        RECT 106.325 31.095 108.015 31.615 ;
        RECT 110.690 31.180 111.030 32.010 ;
        RECT 98.985 30.005 104.330 30.440 ;
        RECT 104.505 30.005 108.015 31.095 ;
        RECT 108.645 30.005 108.935 31.170 ;
        RECT 112.510 30.440 112.860 31.690 ;
        RECT 116.210 31.180 116.550 32.010 ;
        RECT 120.145 31.785 121.815 32.555 ;
        RECT 122.445 31.805 123.655 32.555 ;
        RECT 118.030 30.440 118.380 31.690 ;
        RECT 120.145 31.265 120.895 31.785 ;
        RECT 121.065 31.095 121.815 31.615 ;
        RECT 109.105 30.005 114.450 30.440 ;
        RECT 114.625 30.005 119.970 30.440 ;
        RECT 120.145 30.005 121.815 31.095 ;
        RECT 122.445 31.095 122.965 31.635 ;
        RECT 123.135 31.265 123.655 31.805 ;
        RECT 122.445 30.005 123.655 31.095 ;
        RECT 5.520 29.835 123.740 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 6.985 29.400 12.330 29.835 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 8.570 27.830 8.910 28.660 ;
        RECT 10.390 28.150 10.740 29.400 ;
        RECT 12.505 28.745 16.015 29.835 ;
        RECT 12.505 28.055 14.155 28.575 ;
        RECT 14.325 28.225 16.015 28.745 ;
        RECT 16.705 28.695 16.915 29.835 ;
        RECT 17.085 28.685 17.415 29.665 ;
        RECT 17.585 28.695 17.815 29.835 ;
        RECT 6.985 27.285 12.330 27.830 ;
        RECT 12.505 27.285 16.015 28.055 ;
        RECT 16.705 27.285 16.915 28.105 ;
        RECT 17.085 28.085 17.335 28.685 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.945 28.745 20.615 29.835 ;
        RECT 17.505 28.275 17.835 28.525 ;
        RECT 17.085 27.455 17.415 28.085 ;
        RECT 17.585 27.285 17.815 28.105 ;
        RECT 18.945 28.055 19.695 28.575 ;
        RECT 19.865 28.225 20.615 28.745 ;
        RECT 21.245 28.760 21.515 29.665 ;
        RECT 21.685 29.075 22.015 29.835 ;
        RECT 22.195 28.905 22.365 29.665 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 18.945 27.285 20.615 28.055 ;
        RECT 21.245 27.960 21.415 28.760 ;
        RECT 21.700 28.735 22.365 28.905 ;
        RECT 21.700 28.590 21.870 28.735 ;
        RECT 23.585 28.695 23.815 29.835 ;
        RECT 23.985 28.685 24.315 29.665 ;
        RECT 24.485 28.695 24.695 29.835 ;
        RECT 25.390 29.165 25.645 29.665 ;
        RECT 25.815 29.335 26.145 29.835 ;
        RECT 25.390 28.995 26.140 29.165 ;
        RECT 21.585 28.260 21.870 28.590 ;
        RECT 21.700 28.005 21.870 28.260 ;
        RECT 22.105 28.185 22.435 28.555 ;
        RECT 23.565 28.275 23.895 28.525 ;
        RECT 21.245 27.455 21.505 27.960 ;
        RECT 21.700 27.835 22.365 28.005 ;
        RECT 21.685 27.285 22.015 27.665 ;
        RECT 22.195 27.455 22.365 27.835 ;
        RECT 23.585 27.285 23.815 28.105 ;
        RECT 24.065 28.085 24.315 28.685 ;
        RECT 25.390 28.175 25.740 28.825 ;
        RECT 23.985 27.455 24.315 28.085 ;
        RECT 24.485 27.285 24.695 28.105 ;
        RECT 25.910 28.005 26.140 28.995 ;
        RECT 25.390 27.835 26.140 28.005 ;
        RECT 25.390 27.545 25.645 27.835 ;
        RECT 25.815 27.285 26.145 27.665 ;
        RECT 26.315 27.545 26.485 29.665 ;
        RECT 26.655 28.865 26.980 29.650 ;
        RECT 27.150 29.375 27.400 29.835 ;
        RECT 27.570 29.335 27.820 29.665 ;
        RECT 28.035 29.335 28.715 29.665 ;
        RECT 27.570 29.205 27.740 29.335 ;
        RECT 27.345 29.035 27.740 29.205 ;
        RECT 26.715 27.815 27.175 28.865 ;
        RECT 27.345 27.675 27.515 29.035 ;
        RECT 27.910 28.775 28.375 29.165 ;
        RECT 27.685 27.965 28.035 28.585 ;
        RECT 28.205 28.185 28.375 28.775 ;
        RECT 28.545 28.555 28.715 29.335 ;
        RECT 28.885 29.235 29.055 29.575 ;
        RECT 29.290 29.405 29.620 29.835 ;
        RECT 29.790 29.235 29.960 29.575 ;
        RECT 30.255 29.375 30.625 29.835 ;
        RECT 28.885 29.065 29.960 29.235 ;
        RECT 30.795 29.205 30.965 29.665 ;
        RECT 31.200 29.325 32.070 29.665 ;
        RECT 32.240 29.375 32.490 29.835 ;
        RECT 30.405 29.035 30.965 29.205 ;
        RECT 30.405 28.895 30.575 29.035 ;
        RECT 29.075 28.725 30.575 28.895 ;
        RECT 31.270 28.865 31.730 29.155 ;
        RECT 28.545 28.385 30.235 28.555 ;
        RECT 28.205 27.965 28.560 28.185 ;
        RECT 28.730 27.675 28.900 28.385 ;
        RECT 29.105 27.965 29.895 28.215 ;
        RECT 30.065 28.205 30.235 28.385 ;
        RECT 30.405 28.035 30.575 28.725 ;
        RECT 26.845 27.285 27.175 27.645 ;
        RECT 27.345 27.505 27.840 27.675 ;
        RECT 28.045 27.505 28.900 27.675 ;
        RECT 29.775 27.285 30.105 27.745 ;
        RECT 30.315 27.645 30.575 28.035 ;
        RECT 30.765 28.855 31.730 28.865 ;
        RECT 31.900 28.945 32.070 29.325 ;
        RECT 32.660 29.285 32.830 29.575 ;
        RECT 33.010 29.455 33.340 29.835 ;
        RECT 32.660 29.115 33.460 29.285 ;
        RECT 30.765 28.695 31.440 28.855 ;
        RECT 31.900 28.775 33.120 28.945 ;
        RECT 30.765 27.905 30.975 28.695 ;
        RECT 31.900 28.685 32.070 28.775 ;
        RECT 31.145 27.905 31.495 28.525 ;
        RECT 31.665 28.515 32.070 28.685 ;
        RECT 31.665 27.735 31.835 28.515 ;
        RECT 32.005 28.065 32.225 28.345 ;
        RECT 32.405 28.235 32.945 28.605 ;
        RECT 33.290 28.525 33.460 29.115 ;
        RECT 33.680 28.695 33.985 29.835 ;
        RECT 34.155 28.645 34.410 29.525 ;
        RECT 34.645 28.695 34.855 29.835 ;
        RECT 33.290 28.495 34.030 28.525 ;
        RECT 32.005 27.895 32.535 28.065 ;
        RECT 30.315 27.475 30.665 27.645 ;
        RECT 30.885 27.455 31.835 27.735 ;
        RECT 32.005 27.285 32.195 27.725 ;
        RECT 32.365 27.665 32.535 27.895 ;
        RECT 32.705 27.835 32.945 28.235 ;
        RECT 33.115 28.195 34.030 28.495 ;
        RECT 33.115 28.020 33.440 28.195 ;
        RECT 33.115 27.665 33.435 28.020 ;
        RECT 34.200 27.995 34.410 28.645 ;
        RECT 35.025 28.685 35.355 29.665 ;
        RECT 35.525 28.695 35.755 29.835 ;
        RECT 35.965 28.745 39.475 29.835 ;
        RECT 32.365 27.495 33.435 27.665 ;
        RECT 33.680 27.285 33.985 27.745 ;
        RECT 34.155 27.465 34.410 27.995 ;
        RECT 34.645 27.285 34.855 28.105 ;
        RECT 35.025 28.085 35.275 28.685 ;
        RECT 35.445 28.275 35.775 28.525 ;
        RECT 35.025 27.455 35.355 28.085 ;
        RECT 35.525 27.285 35.755 28.105 ;
        RECT 35.965 28.055 37.615 28.575 ;
        RECT 37.785 28.225 39.475 28.745 ;
        RECT 40.565 28.760 40.835 29.665 ;
        RECT 41.005 29.075 41.335 29.835 ;
        RECT 41.515 28.905 41.685 29.665 ;
        RECT 35.965 27.285 39.475 28.055 ;
        RECT 40.565 27.960 40.735 28.760 ;
        RECT 41.020 28.735 41.685 28.905 ;
        RECT 41.020 28.590 41.190 28.735 ;
        RECT 42.905 28.695 43.135 29.835 ;
        RECT 43.305 28.685 43.635 29.665 ;
        RECT 43.805 28.695 44.015 29.835 ;
        RECT 40.905 28.260 41.190 28.590 ;
        RECT 41.020 28.005 41.190 28.260 ;
        RECT 41.425 28.185 41.755 28.555 ;
        RECT 42.885 28.275 43.215 28.525 ;
        RECT 40.565 27.455 40.825 27.960 ;
        RECT 41.020 27.835 41.685 28.005 ;
        RECT 41.005 27.285 41.335 27.665 ;
        RECT 41.515 27.455 41.685 27.835 ;
        RECT 42.905 27.285 43.135 28.105 ;
        RECT 43.385 28.085 43.635 28.685 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.710 28.695 45.045 29.665 ;
        RECT 45.215 28.695 45.385 29.835 ;
        RECT 45.555 29.495 47.585 29.665 ;
        RECT 43.305 27.455 43.635 28.085 ;
        RECT 43.805 27.285 44.015 28.105 ;
        RECT 44.710 28.025 44.880 28.695 ;
        RECT 45.555 28.525 45.725 29.495 ;
        RECT 45.050 28.195 45.305 28.525 ;
        RECT 45.530 28.195 45.725 28.525 ;
        RECT 45.895 29.155 47.020 29.325 ;
        RECT 45.135 28.025 45.305 28.195 ;
        RECT 45.895 28.025 46.065 29.155 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 44.710 27.455 44.965 28.025 ;
        RECT 45.135 27.855 46.065 28.025 ;
        RECT 46.235 28.815 47.245 28.985 ;
        RECT 46.235 28.015 46.405 28.815 ;
        RECT 46.610 28.475 46.885 28.615 ;
        RECT 46.605 28.305 46.885 28.475 ;
        RECT 45.890 27.820 46.065 27.855 ;
        RECT 45.135 27.285 45.465 27.685 ;
        RECT 45.890 27.455 46.420 27.820 ;
        RECT 46.610 27.455 46.885 28.305 ;
        RECT 47.055 27.455 47.245 28.815 ;
        RECT 47.415 28.830 47.585 29.495 ;
        RECT 47.755 29.075 47.925 29.835 ;
        RECT 48.160 29.075 48.675 29.485 ;
        RECT 47.415 28.640 48.165 28.830 ;
        RECT 48.335 28.265 48.675 29.075 ;
        RECT 48.845 28.745 51.435 29.835 ;
        RECT 51.610 29.165 51.865 29.665 ;
        RECT 52.035 29.335 52.365 29.835 ;
        RECT 51.610 28.995 52.360 29.165 ;
        RECT 47.445 28.095 48.675 28.265 ;
        RECT 47.425 27.285 47.935 27.820 ;
        RECT 48.155 27.490 48.400 28.095 ;
        RECT 48.845 28.055 50.055 28.575 ;
        RECT 50.225 28.225 51.435 28.745 ;
        RECT 51.610 28.175 51.960 28.825 ;
        RECT 48.845 27.285 51.435 28.055 ;
        RECT 52.130 28.005 52.360 28.995 ;
        RECT 51.610 27.835 52.360 28.005 ;
        RECT 51.610 27.545 51.865 27.835 ;
        RECT 52.035 27.285 52.365 27.665 ;
        RECT 52.535 27.545 52.705 29.665 ;
        RECT 52.875 28.865 53.200 29.650 ;
        RECT 53.370 29.375 53.620 29.835 ;
        RECT 53.790 29.335 54.040 29.665 ;
        RECT 54.255 29.335 54.935 29.665 ;
        RECT 53.790 29.205 53.960 29.335 ;
        RECT 53.565 29.035 53.960 29.205 ;
        RECT 52.935 27.815 53.395 28.865 ;
        RECT 53.565 27.675 53.735 29.035 ;
        RECT 54.130 28.775 54.595 29.165 ;
        RECT 53.905 27.965 54.255 28.585 ;
        RECT 54.425 28.185 54.595 28.775 ;
        RECT 54.765 28.555 54.935 29.335 ;
        RECT 55.105 29.235 55.275 29.575 ;
        RECT 55.510 29.405 55.840 29.835 ;
        RECT 56.010 29.235 56.180 29.575 ;
        RECT 56.475 29.375 56.845 29.835 ;
        RECT 55.105 29.065 56.180 29.235 ;
        RECT 57.015 29.205 57.185 29.665 ;
        RECT 57.420 29.325 58.290 29.665 ;
        RECT 58.460 29.375 58.710 29.835 ;
        RECT 56.625 29.035 57.185 29.205 ;
        RECT 56.625 28.895 56.795 29.035 ;
        RECT 55.295 28.725 56.795 28.895 ;
        RECT 57.490 28.865 57.950 29.155 ;
        RECT 54.765 28.385 56.455 28.555 ;
        RECT 54.425 27.965 54.780 28.185 ;
        RECT 54.950 27.675 55.120 28.385 ;
        RECT 55.325 27.965 56.115 28.215 ;
        RECT 56.285 28.205 56.455 28.385 ;
        RECT 56.625 28.035 56.795 28.725 ;
        RECT 53.065 27.285 53.395 27.645 ;
        RECT 53.565 27.505 54.060 27.675 ;
        RECT 54.265 27.505 55.120 27.675 ;
        RECT 55.995 27.285 56.325 27.745 ;
        RECT 56.535 27.645 56.795 28.035 ;
        RECT 56.985 28.855 57.950 28.865 ;
        RECT 58.120 28.945 58.290 29.325 ;
        RECT 58.880 29.285 59.050 29.575 ;
        RECT 59.230 29.455 59.560 29.835 ;
        RECT 58.880 29.115 59.680 29.285 ;
        RECT 56.985 28.695 57.660 28.855 ;
        RECT 58.120 28.775 59.340 28.945 ;
        RECT 56.985 27.905 57.195 28.695 ;
        RECT 58.120 28.685 58.290 28.775 ;
        RECT 57.365 27.905 57.715 28.525 ;
        RECT 57.885 28.515 58.290 28.685 ;
        RECT 57.885 27.735 58.055 28.515 ;
        RECT 58.225 28.065 58.445 28.345 ;
        RECT 58.625 28.235 59.165 28.605 ;
        RECT 59.510 28.525 59.680 29.115 ;
        RECT 59.900 28.695 60.205 29.835 ;
        RECT 60.375 28.645 60.630 29.525 ;
        RECT 60.805 29.400 66.150 29.835 ;
        RECT 59.510 28.495 60.250 28.525 ;
        RECT 58.225 27.895 58.755 28.065 ;
        RECT 56.535 27.475 56.885 27.645 ;
        RECT 57.105 27.455 58.055 27.735 ;
        RECT 58.225 27.285 58.415 27.725 ;
        RECT 58.585 27.665 58.755 27.895 ;
        RECT 58.925 27.835 59.165 28.235 ;
        RECT 59.335 28.195 60.250 28.495 ;
        RECT 59.335 28.020 59.660 28.195 ;
        RECT 59.335 27.665 59.655 28.020 ;
        RECT 60.420 27.995 60.630 28.645 ;
        RECT 58.585 27.495 59.655 27.665 ;
        RECT 59.900 27.285 60.205 27.745 ;
        RECT 60.375 27.465 60.630 27.995 ;
        RECT 62.390 27.830 62.730 28.660 ;
        RECT 64.210 28.150 64.560 29.400 ;
        RECT 66.325 28.745 69.835 29.835 ;
        RECT 66.325 28.055 67.975 28.575 ;
        RECT 68.145 28.225 69.835 28.745 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 70.965 28.695 71.195 29.835 ;
        RECT 71.365 28.685 71.695 29.665 ;
        RECT 71.865 28.695 72.075 29.835 ;
        RECT 72.305 28.745 75.815 29.835 ;
        RECT 76.910 29.165 77.165 29.665 ;
        RECT 77.335 29.335 77.665 29.835 ;
        RECT 76.910 28.995 77.660 29.165 ;
        RECT 70.945 28.275 71.275 28.525 ;
        RECT 60.805 27.285 66.150 27.830 ;
        RECT 66.325 27.285 69.835 28.055 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 70.965 27.285 71.195 28.105 ;
        RECT 71.445 28.085 71.695 28.685 ;
        RECT 71.365 27.455 71.695 28.085 ;
        RECT 71.865 27.285 72.075 28.105 ;
        RECT 72.305 28.055 73.955 28.575 ;
        RECT 74.125 28.225 75.815 28.745 ;
        RECT 76.910 28.175 77.260 28.825 ;
        RECT 72.305 27.285 75.815 28.055 ;
        RECT 77.430 28.005 77.660 28.995 ;
        RECT 76.910 27.835 77.660 28.005 ;
        RECT 76.910 27.545 77.165 27.835 ;
        RECT 77.335 27.285 77.665 27.665 ;
        RECT 77.835 27.545 78.005 29.665 ;
        RECT 78.175 28.865 78.500 29.650 ;
        RECT 78.670 29.375 78.920 29.835 ;
        RECT 79.090 29.335 79.340 29.665 ;
        RECT 79.555 29.335 80.235 29.665 ;
        RECT 79.090 29.205 79.260 29.335 ;
        RECT 78.865 29.035 79.260 29.205 ;
        RECT 78.235 27.815 78.695 28.865 ;
        RECT 78.865 27.675 79.035 29.035 ;
        RECT 79.430 28.775 79.895 29.165 ;
        RECT 79.205 27.965 79.555 28.585 ;
        RECT 79.725 28.185 79.895 28.775 ;
        RECT 80.065 28.555 80.235 29.335 ;
        RECT 80.405 29.235 80.575 29.575 ;
        RECT 80.810 29.405 81.140 29.835 ;
        RECT 81.310 29.235 81.480 29.575 ;
        RECT 81.775 29.375 82.145 29.835 ;
        RECT 80.405 29.065 81.480 29.235 ;
        RECT 82.315 29.205 82.485 29.665 ;
        RECT 82.720 29.325 83.590 29.665 ;
        RECT 83.760 29.375 84.010 29.835 ;
        RECT 81.925 29.035 82.485 29.205 ;
        RECT 81.925 28.895 82.095 29.035 ;
        RECT 80.595 28.725 82.095 28.895 ;
        RECT 82.790 28.865 83.250 29.155 ;
        RECT 80.065 28.385 81.755 28.555 ;
        RECT 79.725 27.965 80.080 28.185 ;
        RECT 80.250 27.675 80.420 28.385 ;
        RECT 80.625 27.965 81.415 28.215 ;
        RECT 81.585 28.205 81.755 28.385 ;
        RECT 81.925 28.035 82.095 28.725 ;
        RECT 78.365 27.285 78.695 27.645 ;
        RECT 78.865 27.505 79.360 27.675 ;
        RECT 79.565 27.505 80.420 27.675 ;
        RECT 81.295 27.285 81.625 27.745 ;
        RECT 81.835 27.645 82.095 28.035 ;
        RECT 82.285 28.855 83.250 28.865 ;
        RECT 83.420 28.945 83.590 29.325 ;
        RECT 84.180 29.285 84.350 29.575 ;
        RECT 84.530 29.455 84.860 29.835 ;
        RECT 84.180 29.115 84.980 29.285 ;
        RECT 82.285 28.695 82.960 28.855 ;
        RECT 83.420 28.775 84.640 28.945 ;
        RECT 82.285 27.905 82.495 28.695 ;
        RECT 83.420 28.685 83.590 28.775 ;
        RECT 82.665 27.905 83.015 28.525 ;
        RECT 83.185 28.515 83.590 28.685 ;
        RECT 83.185 27.735 83.355 28.515 ;
        RECT 83.525 28.065 83.745 28.345 ;
        RECT 83.925 28.235 84.465 28.605 ;
        RECT 84.810 28.525 84.980 29.115 ;
        RECT 85.200 28.695 85.505 29.835 ;
        RECT 85.675 28.645 85.930 29.525 ;
        RECT 84.810 28.495 85.550 28.525 ;
        RECT 83.525 27.895 84.055 28.065 ;
        RECT 81.835 27.475 82.185 27.645 ;
        RECT 82.405 27.455 83.355 27.735 ;
        RECT 83.525 27.285 83.715 27.725 ;
        RECT 83.885 27.665 84.055 27.895 ;
        RECT 84.225 27.835 84.465 28.235 ;
        RECT 84.635 28.195 85.550 28.495 ;
        RECT 84.635 28.020 84.960 28.195 ;
        RECT 84.635 27.665 84.955 28.020 ;
        RECT 85.720 27.995 85.930 28.645 ;
        RECT 83.885 27.495 84.955 27.665 ;
        RECT 85.200 27.285 85.505 27.745 ;
        RECT 85.675 27.465 85.930 27.995 ;
        RECT 86.110 28.645 86.365 29.525 ;
        RECT 86.535 28.695 86.840 29.835 ;
        RECT 87.180 29.455 87.510 29.835 ;
        RECT 87.690 29.285 87.860 29.575 ;
        RECT 88.030 29.375 88.280 29.835 ;
        RECT 87.060 29.115 87.860 29.285 ;
        RECT 88.450 29.325 89.320 29.665 ;
        RECT 86.110 27.995 86.320 28.645 ;
        RECT 87.060 28.525 87.230 29.115 ;
        RECT 88.450 28.945 88.620 29.325 ;
        RECT 89.555 29.205 89.725 29.665 ;
        RECT 89.895 29.375 90.265 29.835 ;
        RECT 90.560 29.235 90.730 29.575 ;
        RECT 90.900 29.405 91.230 29.835 ;
        RECT 91.465 29.235 91.635 29.575 ;
        RECT 87.400 28.775 88.620 28.945 ;
        RECT 88.790 28.865 89.250 29.155 ;
        RECT 89.555 29.035 90.115 29.205 ;
        RECT 90.560 29.065 91.635 29.235 ;
        RECT 91.805 29.335 92.485 29.665 ;
        RECT 92.700 29.335 92.950 29.665 ;
        RECT 93.120 29.375 93.370 29.835 ;
        RECT 89.945 28.895 90.115 29.035 ;
        RECT 88.790 28.855 89.755 28.865 ;
        RECT 88.450 28.685 88.620 28.775 ;
        RECT 89.080 28.695 89.755 28.855 ;
        RECT 86.490 28.495 87.230 28.525 ;
        RECT 86.490 28.195 87.405 28.495 ;
        RECT 87.080 28.020 87.405 28.195 ;
        RECT 86.110 27.465 86.365 27.995 ;
        RECT 86.535 27.285 86.840 27.745 ;
        RECT 87.085 27.665 87.405 28.020 ;
        RECT 87.575 28.235 88.115 28.605 ;
        RECT 88.450 28.515 88.855 28.685 ;
        RECT 87.575 27.835 87.815 28.235 ;
        RECT 88.295 28.065 88.515 28.345 ;
        RECT 87.985 27.895 88.515 28.065 ;
        RECT 87.985 27.665 88.155 27.895 ;
        RECT 88.685 27.735 88.855 28.515 ;
        RECT 89.025 27.905 89.375 28.525 ;
        RECT 89.545 27.905 89.755 28.695 ;
        RECT 89.945 28.725 91.445 28.895 ;
        RECT 89.945 28.035 90.115 28.725 ;
        RECT 91.805 28.555 91.975 29.335 ;
        RECT 92.780 29.205 92.950 29.335 ;
        RECT 90.285 28.385 91.975 28.555 ;
        RECT 92.145 28.775 92.610 29.165 ;
        RECT 92.780 29.035 93.175 29.205 ;
        RECT 90.285 28.205 90.455 28.385 ;
        RECT 87.085 27.495 88.155 27.665 ;
        RECT 88.325 27.285 88.515 27.725 ;
        RECT 88.685 27.455 89.635 27.735 ;
        RECT 89.945 27.645 90.205 28.035 ;
        RECT 90.625 27.965 91.415 28.215 ;
        RECT 89.855 27.475 90.205 27.645 ;
        RECT 90.415 27.285 90.745 27.745 ;
        RECT 91.620 27.675 91.790 28.385 ;
        RECT 92.145 28.185 92.315 28.775 ;
        RECT 91.960 27.965 92.315 28.185 ;
        RECT 92.485 27.965 92.835 28.585 ;
        RECT 93.005 27.675 93.175 29.035 ;
        RECT 93.540 28.865 93.865 29.650 ;
        RECT 93.345 27.815 93.805 28.865 ;
        RECT 91.620 27.505 92.475 27.675 ;
        RECT 92.680 27.505 93.175 27.675 ;
        RECT 93.345 27.285 93.675 27.645 ;
        RECT 94.035 27.545 94.205 29.665 ;
        RECT 94.375 29.335 94.705 29.835 ;
        RECT 94.875 29.165 95.130 29.665 ;
        RECT 94.380 28.995 95.130 29.165 ;
        RECT 94.380 28.005 94.610 28.995 ;
        RECT 94.780 28.175 95.130 28.825 ;
        RECT 95.765 28.670 96.055 29.835 ;
        RECT 96.225 29.400 101.570 29.835 ;
        RECT 101.745 29.400 107.090 29.835 ;
        RECT 107.265 29.400 112.610 29.835 ;
        RECT 112.785 29.400 118.130 29.835 ;
        RECT 94.380 27.835 95.130 28.005 ;
        RECT 94.375 27.285 94.705 27.665 ;
        RECT 94.875 27.545 95.130 27.835 ;
        RECT 95.765 27.285 96.055 28.010 ;
        RECT 97.810 27.830 98.150 28.660 ;
        RECT 99.630 28.150 99.980 29.400 ;
        RECT 103.330 27.830 103.670 28.660 ;
        RECT 105.150 28.150 105.500 29.400 ;
        RECT 108.850 27.830 109.190 28.660 ;
        RECT 110.670 28.150 111.020 29.400 ;
        RECT 114.370 27.830 114.710 28.660 ;
        RECT 116.190 28.150 116.540 29.400 ;
        RECT 118.305 28.745 120.895 29.835 ;
        RECT 118.305 28.055 119.515 28.575 ;
        RECT 119.685 28.225 120.895 28.745 ;
        RECT 121.525 28.670 121.815 29.835 ;
        RECT 122.445 28.745 123.655 29.835 ;
        RECT 122.445 28.205 122.965 28.745 ;
        RECT 96.225 27.285 101.570 27.830 ;
        RECT 101.745 27.285 107.090 27.830 ;
        RECT 107.265 27.285 112.610 27.830 ;
        RECT 112.785 27.285 118.130 27.830 ;
        RECT 118.305 27.285 120.895 28.055 ;
        RECT 123.135 28.035 123.655 28.575 ;
        RECT 121.525 27.285 121.815 28.010 ;
        RECT 122.445 27.285 123.655 28.035 ;
        RECT 5.520 27.115 123.740 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 6.985 26.570 12.330 27.115 ;
        RECT 12.505 26.570 17.850 27.115 ;
        RECT 18.025 26.570 23.370 27.115 ;
        RECT 23.545 26.570 28.890 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 8.570 25.740 8.910 26.570 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 10.390 25.000 10.740 26.250 ;
        RECT 14.090 25.740 14.430 26.570 ;
        RECT 15.910 25.000 16.260 26.250 ;
        RECT 19.610 25.740 19.950 26.570 ;
        RECT 21.430 25.000 21.780 26.250 ;
        RECT 25.130 25.740 25.470 26.570 ;
        RECT 29.065 26.345 30.735 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.825 26.570 37.170 27.115 ;
        RECT 26.950 25.000 27.300 26.250 ;
        RECT 29.065 25.825 29.815 26.345 ;
        RECT 29.985 25.655 30.735 26.175 ;
        RECT 33.410 25.740 33.750 26.570 ;
        RECT 38.355 26.565 38.525 26.855 ;
        RECT 38.695 26.735 39.025 27.115 ;
        RECT 38.355 26.395 39.020 26.565 ;
        RECT 6.985 24.565 12.330 25.000 ;
        RECT 12.505 24.565 17.850 25.000 ;
        RECT 18.025 24.565 23.370 25.000 ;
        RECT 23.545 24.565 28.890 25.000 ;
        RECT 29.065 24.565 30.735 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 35.230 25.000 35.580 26.250 ;
        RECT 38.270 25.575 38.620 26.225 ;
        RECT 38.790 25.405 39.020 26.395 ;
        RECT 38.355 25.235 39.020 25.405 ;
        RECT 31.825 24.565 37.170 25.000 ;
        RECT 38.355 24.735 38.525 25.235 ;
        RECT 38.695 24.565 39.025 25.065 ;
        RECT 39.195 24.735 39.420 26.855 ;
        RECT 39.635 26.735 39.965 27.115 ;
        RECT 40.135 26.565 40.305 26.895 ;
        RECT 40.605 26.735 41.620 26.935 ;
        RECT 39.610 26.375 40.305 26.565 ;
        RECT 39.610 25.405 39.780 26.375 ;
        RECT 39.950 25.575 40.360 26.195 ;
        RECT 40.530 25.625 40.750 26.495 ;
        RECT 40.930 26.185 41.280 26.555 ;
        RECT 41.450 26.005 41.620 26.735 ;
        RECT 41.790 26.675 42.200 27.115 ;
        RECT 42.490 26.475 42.740 26.905 ;
        RECT 42.940 26.655 43.260 27.115 ;
        RECT 43.820 26.725 44.670 26.895 ;
        RECT 41.790 26.135 42.200 26.465 ;
        RECT 42.490 26.135 42.910 26.475 ;
        RECT 41.200 25.965 41.620 26.005 ;
        RECT 41.200 25.795 42.550 25.965 ;
        RECT 39.610 25.235 40.305 25.405 ;
        RECT 40.530 25.245 41.030 25.625 ;
        RECT 39.635 24.565 39.965 25.065 ;
        RECT 40.135 24.735 40.305 25.235 ;
        RECT 41.200 24.950 41.370 25.795 ;
        RECT 42.300 25.635 42.550 25.795 ;
        RECT 41.540 25.365 41.790 25.625 ;
        RECT 42.720 25.365 42.910 26.135 ;
        RECT 41.540 25.115 42.910 25.365 ;
        RECT 43.080 26.305 44.330 26.475 ;
        RECT 43.080 25.545 43.250 26.305 ;
        RECT 44.000 26.185 44.330 26.305 ;
        RECT 43.420 25.725 43.600 26.135 ;
        RECT 44.500 25.965 44.670 26.725 ;
        RECT 44.870 26.635 45.530 27.115 ;
        RECT 45.710 26.520 46.030 26.850 ;
        RECT 44.860 26.195 45.520 26.465 ;
        RECT 44.860 26.135 45.190 26.195 ;
        RECT 45.340 25.965 45.670 26.025 ;
        RECT 43.770 25.795 45.670 25.965 ;
        RECT 43.080 25.235 43.600 25.545 ;
        RECT 43.770 25.285 43.940 25.795 ;
        RECT 45.840 25.625 46.030 26.520 ;
        RECT 44.110 25.455 46.030 25.625 ;
        RECT 45.710 25.435 46.030 25.455 ;
        RECT 46.230 26.205 46.480 26.855 ;
        RECT 46.660 26.655 46.945 27.115 ;
        RECT 47.125 26.775 47.380 26.935 ;
        RECT 47.125 26.605 47.465 26.775 ;
        RECT 47.125 26.405 47.380 26.605 ;
        RECT 47.925 26.570 53.270 27.115 ;
        RECT 46.230 25.875 47.030 26.205 ;
        RECT 43.770 25.115 44.980 25.285 ;
        RECT 40.540 24.780 41.370 24.950 ;
        RECT 41.610 24.565 41.990 24.945 ;
        RECT 42.170 24.825 42.340 25.115 ;
        RECT 43.770 25.035 43.940 25.115 ;
        RECT 42.510 24.565 42.840 24.945 ;
        RECT 43.310 24.785 43.940 25.035 ;
        RECT 44.120 24.565 44.540 24.945 ;
        RECT 44.740 24.825 44.980 25.115 ;
        RECT 45.210 24.565 45.540 25.255 ;
        RECT 45.710 24.825 45.880 25.435 ;
        RECT 46.230 25.285 46.480 25.875 ;
        RECT 47.200 25.545 47.380 26.405 ;
        RECT 49.510 25.740 49.850 26.570 ;
        RECT 53.445 26.345 55.115 27.115 ;
        RECT 46.150 24.775 46.480 25.285 ;
        RECT 46.660 24.565 46.945 25.365 ;
        RECT 47.125 24.875 47.380 25.545 ;
        RECT 51.330 25.000 51.680 26.250 ;
        RECT 53.445 25.825 54.195 26.345 ;
        RECT 55.785 26.295 56.015 27.115 ;
        RECT 56.185 26.315 56.515 26.945 ;
        RECT 54.365 25.655 55.115 26.175 ;
        RECT 55.765 25.875 56.095 26.125 ;
        RECT 56.265 25.715 56.515 26.315 ;
        RECT 56.685 26.295 56.895 27.115 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 57.585 26.570 62.930 27.115 ;
        RECT 59.170 25.740 59.510 26.570 ;
        RECT 63.105 26.375 63.570 26.920 ;
        RECT 47.925 24.565 53.270 25.000 ;
        RECT 53.445 24.565 55.115 25.655 ;
        RECT 55.785 24.565 56.015 25.705 ;
        RECT 56.185 24.735 56.515 25.715 ;
        RECT 56.685 24.565 56.895 25.705 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 60.990 25.000 61.340 26.250 ;
        RECT 63.105 25.415 63.275 26.375 ;
        RECT 64.075 26.295 64.245 27.115 ;
        RECT 64.415 26.465 64.745 26.945 ;
        RECT 64.915 26.725 65.265 27.115 ;
        RECT 65.435 26.545 65.665 26.945 ;
        RECT 65.155 26.465 65.665 26.545 ;
        RECT 64.415 26.375 65.665 26.465 ;
        RECT 65.835 26.375 66.155 26.855 ;
        RECT 64.415 26.295 65.325 26.375 ;
        RECT 63.445 25.755 63.690 26.205 ;
        RECT 63.950 25.925 64.645 26.125 ;
        RECT 64.815 25.955 65.415 26.125 ;
        RECT 64.815 25.755 64.985 25.955 ;
        RECT 65.645 25.785 65.815 26.205 ;
        RECT 63.445 25.585 64.985 25.755 ;
        RECT 65.155 25.615 65.815 25.785 ;
        RECT 65.155 25.415 65.325 25.615 ;
        RECT 65.985 25.445 66.155 26.375 ;
        RECT 66.375 26.360 66.625 27.115 ;
        RECT 66.795 26.405 67.045 26.935 ;
        RECT 67.215 26.655 67.520 27.115 ;
        RECT 67.765 26.735 68.835 26.905 ;
        RECT 66.795 25.755 67.000 26.405 ;
        RECT 67.765 26.380 68.085 26.735 ;
        RECT 67.760 26.205 68.085 26.380 ;
        RECT 67.170 25.905 68.085 26.205 ;
        RECT 68.255 26.165 68.495 26.565 ;
        RECT 68.665 26.505 68.835 26.735 ;
        RECT 69.005 26.675 69.195 27.115 ;
        RECT 69.365 26.665 70.315 26.945 ;
        RECT 70.535 26.755 70.885 26.925 ;
        RECT 68.665 26.335 69.195 26.505 ;
        RECT 67.170 25.875 67.910 25.905 ;
        RECT 63.105 25.245 65.325 25.415 ;
        RECT 65.495 25.245 66.155 25.445 ;
        RECT 57.585 24.565 62.930 25.000 ;
        RECT 63.105 24.565 63.405 25.075 ;
        RECT 63.575 24.735 63.905 25.245 ;
        RECT 65.495 25.075 65.665 25.245 ;
        RECT 64.075 24.565 64.705 25.075 ;
        RECT 65.285 24.905 65.665 25.075 ;
        RECT 65.835 24.565 66.135 25.075 ;
        RECT 66.375 24.565 66.625 25.705 ;
        RECT 66.795 24.875 67.045 25.755 ;
        RECT 67.215 24.565 67.520 25.705 ;
        RECT 67.740 25.285 67.910 25.875 ;
        RECT 68.255 25.795 68.795 26.165 ;
        RECT 68.975 26.055 69.195 26.335 ;
        RECT 69.365 25.885 69.535 26.665 ;
        RECT 69.130 25.715 69.535 25.885 ;
        RECT 69.705 25.875 70.055 26.495 ;
        RECT 69.130 25.625 69.300 25.715 ;
        RECT 70.225 25.705 70.435 26.495 ;
        RECT 68.080 25.455 69.300 25.625 ;
        RECT 69.760 25.545 70.435 25.705 ;
        RECT 67.740 25.115 68.540 25.285 ;
        RECT 67.860 24.565 68.190 24.945 ;
        RECT 68.370 24.825 68.540 25.115 ;
        RECT 69.130 25.075 69.300 25.455 ;
        RECT 69.470 25.535 70.435 25.545 ;
        RECT 70.625 26.365 70.885 26.755 ;
        RECT 71.095 26.655 71.425 27.115 ;
        RECT 72.300 26.725 73.155 26.895 ;
        RECT 73.360 26.725 73.855 26.895 ;
        RECT 74.025 26.755 74.355 27.115 ;
        RECT 70.625 25.675 70.795 26.365 ;
        RECT 70.965 26.015 71.135 26.195 ;
        RECT 71.305 26.185 72.095 26.435 ;
        RECT 72.300 26.015 72.470 26.725 ;
        RECT 72.640 26.215 72.995 26.435 ;
        RECT 70.965 25.845 72.655 26.015 ;
        RECT 69.470 25.245 69.930 25.535 ;
        RECT 70.625 25.505 72.125 25.675 ;
        RECT 70.625 25.365 70.795 25.505 ;
        RECT 70.235 25.195 70.795 25.365 ;
        RECT 68.710 24.565 68.960 25.025 ;
        RECT 69.130 24.735 70.000 25.075 ;
        RECT 70.235 24.735 70.405 25.195 ;
        RECT 71.240 25.165 72.315 25.335 ;
        RECT 70.575 24.565 70.945 25.025 ;
        RECT 71.240 24.825 71.410 25.165 ;
        RECT 71.580 24.565 71.910 24.995 ;
        RECT 72.145 24.825 72.315 25.165 ;
        RECT 72.485 25.065 72.655 25.845 ;
        RECT 72.825 25.625 72.995 26.215 ;
        RECT 73.165 25.815 73.515 26.435 ;
        RECT 72.825 25.235 73.290 25.625 ;
        RECT 73.685 25.365 73.855 26.725 ;
        RECT 74.025 25.535 74.485 26.585 ;
        RECT 73.460 25.195 73.855 25.365 ;
        RECT 73.460 25.065 73.630 25.195 ;
        RECT 72.485 24.735 73.165 25.065 ;
        RECT 73.380 24.735 73.630 25.065 ;
        RECT 73.800 24.565 74.050 25.025 ;
        RECT 74.220 24.750 74.545 25.535 ;
        RECT 74.715 24.735 74.885 26.855 ;
        RECT 75.055 26.735 75.385 27.115 ;
        RECT 75.555 26.565 75.810 26.855 ;
        RECT 75.985 26.570 81.330 27.115 ;
        RECT 75.060 26.395 75.810 26.565 ;
        RECT 75.060 25.405 75.290 26.395 ;
        RECT 75.460 25.575 75.810 26.225 ;
        RECT 77.570 25.740 77.910 26.570 ;
        RECT 81.505 26.365 82.715 27.115 ;
        RECT 82.885 26.390 83.175 27.115 ;
        RECT 83.345 26.570 88.690 27.115 ;
        RECT 88.865 26.570 94.210 27.115 ;
        RECT 94.385 26.570 99.730 27.115 ;
        RECT 99.905 26.570 105.250 27.115 ;
        RECT 75.060 25.235 75.810 25.405 ;
        RECT 75.055 24.565 75.385 25.065 ;
        RECT 75.555 24.735 75.810 25.235 ;
        RECT 79.390 25.000 79.740 26.250 ;
        RECT 81.505 25.825 82.025 26.365 ;
        RECT 82.195 25.655 82.715 26.195 ;
        RECT 84.930 25.740 85.270 26.570 ;
        RECT 75.985 24.565 81.330 25.000 ;
        RECT 81.505 24.565 82.715 25.655 ;
        RECT 82.885 24.565 83.175 25.730 ;
        RECT 86.750 25.000 87.100 26.250 ;
        RECT 90.450 25.740 90.790 26.570 ;
        RECT 92.270 25.000 92.620 26.250 ;
        RECT 95.970 25.740 96.310 26.570 ;
        RECT 97.790 25.000 98.140 26.250 ;
        RECT 101.490 25.740 101.830 26.570 ;
        RECT 105.425 26.345 108.015 27.115 ;
        RECT 108.645 26.390 108.935 27.115 ;
        RECT 109.105 26.570 114.450 27.115 ;
        RECT 114.625 26.570 119.970 27.115 ;
        RECT 103.310 25.000 103.660 26.250 ;
        RECT 105.425 25.825 106.635 26.345 ;
        RECT 106.805 25.655 108.015 26.175 ;
        RECT 110.690 25.740 111.030 26.570 ;
        RECT 83.345 24.565 88.690 25.000 ;
        RECT 88.865 24.565 94.210 25.000 ;
        RECT 94.385 24.565 99.730 25.000 ;
        RECT 99.905 24.565 105.250 25.000 ;
        RECT 105.425 24.565 108.015 25.655 ;
        RECT 108.645 24.565 108.935 25.730 ;
        RECT 112.510 25.000 112.860 26.250 ;
        RECT 116.210 25.740 116.550 26.570 ;
        RECT 120.145 26.345 121.815 27.115 ;
        RECT 122.445 26.365 123.655 27.115 ;
        RECT 118.030 25.000 118.380 26.250 ;
        RECT 120.145 25.825 120.895 26.345 ;
        RECT 121.065 25.655 121.815 26.175 ;
        RECT 109.105 24.565 114.450 25.000 ;
        RECT 114.625 24.565 119.970 25.000 ;
        RECT 120.145 24.565 121.815 25.655 ;
        RECT 122.445 25.655 122.965 26.195 ;
        RECT 123.135 25.825 123.655 26.365 ;
        RECT 122.445 24.565 123.655 25.655 ;
        RECT 5.520 24.395 123.740 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 6.985 23.960 12.330 24.395 ;
        RECT 12.505 23.960 17.850 24.395 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 8.570 22.390 8.910 23.220 ;
        RECT 10.390 22.710 10.740 23.960 ;
        RECT 14.090 22.390 14.430 23.220 ;
        RECT 15.910 22.710 16.260 23.960 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 18.945 23.960 24.290 24.395 ;
        RECT 24.465 23.960 29.810 24.395 ;
        RECT 29.985 23.960 35.330 24.395 ;
        RECT 35.505 23.960 40.850 24.395 ;
        RECT 6.985 21.845 12.330 22.390 ;
        RECT 12.505 21.845 17.850 22.390 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 20.530 22.390 20.870 23.220 ;
        RECT 22.350 22.710 22.700 23.960 ;
        RECT 26.050 22.390 26.390 23.220 ;
        RECT 27.870 22.710 28.220 23.960 ;
        RECT 31.570 22.390 31.910 23.220 ;
        RECT 33.390 22.710 33.740 23.960 ;
        RECT 37.090 22.390 37.430 23.220 ;
        RECT 38.910 22.710 39.260 23.960 ;
        RECT 41.025 23.305 43.615 24.395 ;
        RECT 41.025 22.615 42.235 23.135 ;
        RECT 42.405 22.785 43.615 23.305 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.705 23.960 50.050 24.395 ;
        RECT 50.225 23.960 55.570 24.395 ;
        RECT 55.745 23.960 61.090 24.395 ;
        RECT 61.265 23.960 66.610 24.395 ;
        RECT 18.945 21.845 24.290 22.390 ;
        RECT 24.465 21.845 29.810 22.390 ;
        RECT 29.985 21.845 35.330 22.390 ;
        RECT 35.505 21.845 40.850 22.390 ;
        RECT 41.025 21.845 43.615 22.615 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 46.290 22.390 46.630 23.220 ;
        RECT 48.110 22.710 48.460 23.960 ;
        RECT 51.810 22.390 52.150 23.220 ;
        RECT 53.630 22.710 53.980 23.960 ;
        RECT 57.330 22.390 57.670 23.220 ;
        RECT 59.150 22.710 59.500 23.960 ;
        RECT 62.850 22.390 63.190 23.220 ;
        RECT 64.670 22.710 65.020 23.960 ;
        RECT 66.785 23.305 69.375 24.395 ;
        RECT 66.785 22.615 67.995 23.135 ;
        RECT 68.165 22.785 69.375 23.305 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.505 23.255 70.735 24.395 ;
        RECT 70.905 23.245 71.235 24.225 ;
        RECT 71.405 23.255 71.615 24.395 ;
        RECT 71.845 23.960 77.190 24.395 ;
        RECT 77.365 23.960 82.710 24.395 ;
        RECT 82.885 23.960 88.230 24.395 ;
        RECT 88.405 23.960 93.750 24.395 ;
        RECT 70.485 22.835 70.815 23.085 ;
        RECT 44.705 21.845 50.050 22.390 ;
        RECT 50.225 21.845 55.570 22.390 ;
        RECT 55.745 21.845 61.090 22.390 ;
        RECT 61.265 21.845 66.610 22.390 ;
        RECT 66.785 21.845 69.375 22.615 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 70.505 21.845 70.735 22.665 ;
        RECT 70.985 22.645 71.235 23.245 ;
        RECT 70.905 22.015 71.235 22.645 ;
        RECT 71.405 21.845 71.615 22.665 ;
        RECT 73.430 22.390 73.770 23.220 ;
        RECT 75.250 22.710 75.600 23.960 ;
        RECT 78.950 22.390 79.290 23.220 ;
        RECT 80.770 22.710 81.120 23.960 ;
        RECT 84.470 22.390 84.810 23.220 ;
        RECT 86.290 22.710 86.640 23.960 ;
        RECT 89.990 22.390 90.330 23.220 ;
        RECT 91.810 22.710 92.160 23.960 ;
        RECT 93.925 23.305 95.595 24.395 ;
        RECT 93.925 22.615 94.675 23.135 ;
        RECT 94.845 22.785 95.595 23.305 ;
        RECT 95.765 23.230 96.055 24.395 ;
        RECT 96.225 23.960 101.570 24.395 ;
        RECT 101.745 23.960 107.090 24.395 ;
        RECT 107.265 23.960 112.610 24.395 ;
        RECT 112.785 23.960 118.130 24.395 ;
        RECT 71.845 21.845 77.190 22.390 ;
        RECT 77.365 21.845 82.710 22.390 ;
        RECT 82.885 21.845 88.230 22.390 ;
        RECT 88.405 21.845 93.750 22.390 ;
        RECT 93.925 21.845 95.595 22.615 ;
        RECT 95.765 21.845 96.055 22.570 ;
        RECT 97.810 22.390 98.150 23.220 ;
        RECT 99.630 22.710 99.980 23.960 ;
        RECT 103.330 22.390 103.670 23.220 ;
        RECT 105.150 22.710 105.500 23.960 ;
        RECT 108.850 22.390 109.190 23.220 ;
        RECT 110.670 22.710 111.020 23.960 ;
        RECT 114.370 22.390 114.710 23.220 ;
        RECT 116.190 22.710 116.540 23.960 ;
        RECT 118.305 23.305 120.895 24.395 ;
        RECT 118.305 22.615 119.515 23.135 ;
        RECT 119.685 22.785 120.895 23.305 ;
        RECT 121.525 23.230 121.815 24.395 ;
        RECT 122.445 23.305 123.655 24.395 ;
        RECT 122.445 22.765 122.965 23.305 ;
        RECT 96.225 21.845 101.570 22.390 ;
        RECT 101.745 21.845 107.090 22.390 ;
        RECT 107.265 21.845 112.610 22.390 ;
        RECT 112.785 21.845 118.130 22.390 ;
        RECT 118.305 21.845 120.895 22.615 ;
        RECT 123.135 22.595 123.655 23.135 ;
        RECT 121.525 21.845 121.815 22.570 ;
        RECT 122.445 21.845 123.655 22.595 ;
        RECT 5.520 21.675 123.740 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 6.985 21.130 12.330 21.675 ;
        RECT 12.505 21.130 17.850 21.675 ;
        RECT 18.025 21.130 23.370 21.675 ;
        RECT 23.545 21.130 28.890 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 8.570 20.300 8.910 21.130 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 10.390 19.560 10.740 20.810 ;
        RECT 14.090 20.300 14.430 21.130 ;
        RECT 15.910 19.560 16.260 20.810 ;
        RECT 19.610 20.300 19.950 21.130 ;
        RECT 21.430 19.560 21.780 20.810 ;
        RECT 25.130 20.300 25.470 21.130 ;
        RECT 29.065 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 37.345 21.130 42.690 21.675 ;
        RECT 42.865 21.130 48.210 21.675 ;
        RECT 48.385 21.130 53.730 21.675 ;
        RECT 26.950 19.560 27.300 20.810 ;
        RECT 29.065 20.385 29.815 20.905 ;
        RECT 29.985 20.215 30.735 20.735 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 6.985 19.125 12.330 19.560 ;
        RECT 12.505 19.125 17.850 19.560 ;
        RECT 18.025 19.125 23.370 19.560 ;
        RECT 23.545 19.125 28.890 19.560 ;
        RECT 29.065 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 38.930 20.300 39.270 21.130 ;
        RECT 40.750 19.560 41.100 20.810 ;
        RECT 44.450 20.300 44.790 21.130 ;
        RECT 46.270 19.560 46.620 20.810 ;
        RECT 49.970 20.300 50.310 21.130 ;
        RECT 53.905 20.905 56.495 21.675 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 57.585 21.130 62.930 21.675 ;
        RECT 63.105 21.130 68.450 21.675 ;
        RECT 68.625 21.130 73.970 21.675 ;
        RECT 74.145 21.130 79.490 21.675 ;
        RECT 51.790 19.560 52.140 20.810 ;
        RECT 53.905 20.385 55.115 20.905 ;
        RECT 55.285 20.215 56.495 20.735 ;
        RECT 59.170 20.300 59.510 21.130 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.345 19.125 42.690 19.560 ;
        RECT 42.865 19.125 48.210 19.560 ;
        RECT 48.385 19.125 53.730 19.560 ;
        RECT 53.905 19.125 56.495 20.215 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 60.990 19.560 61.340 20.810 ;
        RECT 64.690 20.300 65.030 21.130 ;
        RECT 66.510 19.560 66.860 20.810 ;
        RECT 70.210 20.300 70.550 21.130 ;
        RECT 72.030 19.560 72.380 20.810 ;
        RECT 75.730 20.300 76.070 21.130 ;
        RECT 79.665 20.905 82.255 21.675 ;
        RECT 82.885 20.950 83.175 21.675 ;
        RECT 83.345 21.130 88.690 21.675 ;
        RECT 88.865 21.130 94.210 21.675 ;
        RECT 94.385 21.130 99.730 21.675 ;
        RECT 99.905 21.130 105.250 21.675 ;
        RECT 77.550 19.560 77.900 20.810 ;
        RECT 79.665 20.385 80.875 20.905 ;
        RECT 81.045 20.215 82.255 20.735 ;
        RECT 84.930 20.300 85.270 21.130 ;
        RECT 57.585 19.125 62.930 19.560 ;
        RECT 63.105 19.125 68.450 19.560 ;
        RECT 68.625 19.125 73.970 19.560 ;
        RECT 74.145 19.125 79.490 19.560 ;
        RECT 79.665 19.125 82.255 20.215 ;
        RECT 82.885 19.125 83.175 20.290 ;
        RECT 86.750 19.560 87.100 20.810 ;
        RECT 90.450 20.300 90.790 21.130 ;
        RECT 92.270 19.560 92.620 20.810 ;
        RECT 95.970 20.300 96.310 21.130 ;
        RECT 97.790 19.560 98.140 20.810 ;
        RECT 101.490 20.300 101.830 21.130 ;
        RECT 105.425 20.905 108.015 21.675 ;
        RECT 108.645 20.950 108.935 21.675 ;
        RECT 109.105 21.130 114.450 21.675 ;
        RECT 114.625 21.130 119.970 21.675 ;
        RECT 103.310 19.560 103.660 20.810 ;
        RECT 105.425 20.385 106.635 20.905 ;
        RECT 106.805 20.215 108.015 20.735 ;
        RECT 110.690 20.300 111.030 21.130 ;
        RECT 83.345 19.125 88.690 19.560 ;
        RECT 88.865 19.125 94.210 19.560 ;
        RECT 94.385 19.125 99.730 19.560 ;
        RECT 99.905 19.125 105.250 19.560 ;
        RECT 105.425 19.125 108.015 20.215 ;
        RECT 108.645 19.125 108.935 20.290 ;
        RECT 112.510 19.560 112.860 20.810 ;
        RECT 116.210 20.300 116.550 21.130 ;
        RECT 120.145 20.905 121.815 21.675 ;
        RECT 122.445 20.925 123.655 21.675 ;
        RECT 118.030 19.560 118.380 20.810 ;
        RECT 120.145 20.385 120.895 20.905 ;
        RECT 121.065 20.215 121.815 20.735 ;
        RECT 109.105 19.125 114.450 19.560 ;
        RECT 114.625 19.125 119.970 19.560 ;
        RECT 120.145 19.125 121.815 20.215 ;
        RECT 122.445 20.215 122.965 20.755 ;
        RECT 123.135 20.385 123.655 20.925 ;
        RECT 122.445 19.125 123.655 20.215 ;
        RECT 5.520 18.955 123.740 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 6.985 18.520 12.330 18.955 ;
        RECT 12.505 18.520 17.850 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 8.570 16.950 8.910 17.780 ;
        RECT 10.390 17.270 10.740 18.520 ;
        RECT 14.090 16.950 14.430 17.780 ;
        RECT 15.910 17.270 16.260 18.520 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 18.520 24.290 18.955 ;
        RECT 24.465 18.520 29.810 18.955 ;
        RECT 29.985 18.520 35.330 18.955 ;
        RECT 35.505 18.520 40.850 18.955 ;
        RECT 6.985 16.405 12.330 16.950 ;
        RECT 12.505 16.405 17.850 16.950 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 20.530 16.950 20.870 17.780 ;
        RECT 22.350 17.270 22.700 18.520 ;
        RECT 26.050 16.950 26.390 17.780 ;
        RECT 27.870 17.270 28.220 18.520 ;
        RECT 31.570 16.950 31.910 17.780 ;
        RECT 33.390 17.270 33.740 18.520 ;
        RECT 37.090 16.950 37.430 17.780 ;
        RECT 38.910 17.270 39.260 18.520 ;
        RECT 41.025 17.865 43.615 18.955 ;
        RECT 41.025 17.175 42.235 17.695 ;
        RECT 42.405 17.345 43.615 17.865 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 44.705 18.520 50.050 18.955 ;
        RECT 50.225 18.520 55.570 18.955 ;
        RECT 55.745 18.520 61.090 18.955 ;
        RECT 61.265 18.520 66.610 18.955 ;
        RECT 18.945 16.405 24.290 16.950 ;
        RECT 24.465 16.405 29.810 16.950 ;
        RECT 29.985 16.405 35.330 16.950 ;
        RECT 35.505 16.405 40.850 16.950 ;
        RECT 41.025 16.405 43.615 17.175 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 46.290 16.950 46.630 17.780 ;
        RECT 48.110 17.270 48.460 18.520 ;
        RECT 51.810 16.950 52.150 17.780 ;
        RECT 53.630 17.270 53.980 18.520 ;
        RECT 57.330 16.950 57.670 17.780 ;
        RECT 59.150 17.270 59.500 18.520 ;
        RECT 62.850 16.950 63.190 17.780 ;
        RECT 64.670 17.270 65.020 18.520 ;
        RECT 66.785 17.865 69.375 18.955 ;
        RECT 66.785 17.175 67.995 17.695 ;
        RECT 68.165 17.345 69.375 17.865 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 70.465 18.520 75.810 18.955 ;
        RECT 75.985 18.520 81.330 18.955 ;
        RECT 81.505 18.520 86.850 18.955 ;
        RECT 87.025 18.520 92.370 18.955 ;
        RECT 44.705 16.405 50.050 16.950 ;
        RECT 50.225 16.405 55.570 16.950 ;
        RECT 55.745 16.405 61.090 16.950 ;
        RECT 61.265 16.405 66.610 16.950 ;
        RECT 66.785 16.405 69.375 17.175 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 72.050 16.950 72.390 17.780 ;
        RECT 73.870 17.270 74.220 18.520 ;
        RECT 77.570 16.950 77.910 17.780 ;
        RECT 79.390 17.270 79.740 18.520 ;
        RECT 83.090 16.950 83.430 17.780 ;
        RECT 84.910 17.270 85.260 18.520 ;
        RECT 88.610 16.950 88.950 17.780 ;
        RECT 90.430 17.270 90.780 18.520 ;
        RECT 92.545 17.865 95.135 18.955 ;
        RECT 92.545 17.175 93.755 17.695 ;
        RECT 93.925 17.345 95.135 17.865 ;
        RECT 95.765 17.790 96.055 18.955 ;
        RECT 96.225 18.520 101.570 18.955 ;
        RECT 101.745 18.520 107.090 18.955 ;
        RECT 107.265 18.520 112.610 18.955 ;
        RECT 112.785 18.520 118.130 18.955 ;
        RECT 70.465 16.405 75.810 16.950 ;
        RECT 75.985 16.405 81.330 16.950 ;
        RECT 81.505 16.405 86.850 16.950 ;
        RECT 87.025 16.405 92.370 16.950 ;
        RECT 92.545 16.405 95.135 17.175 ;
        RECT 95.765 16.405 96.055 17.130 ;
        RECT 97.810 16.950 98.150 17.780 ;
        RECT 99.630 17.270 99.980 18.520 ;
        RECT 103.330 16.950 103.670 17.780 ;
        RECT 105.150 17.270 105.500 18.520 ;
        RECT 108.850 16.950 109.190 17.780 ;
        RECT 110.670 17.270 111.020 18.520 ;
        RECT 114.370 16.950 114.710 17.780 ;
        RECT 116.190 17.270 116.540 18.520 ;
        RECT 118.305 17.865 120.895 18.955 ;
        RECT 118.305 17.175 119.515 17.695 ;
        RECT 119.685 17.345 120.895 17.865 ;
        RECT 121.525 17.790 121.815 18.955 ;
        RECT 122.445 17.865 123.655 18.955 ;
        RECT 122.445 17.325 122.965 17.865 ;
        RECT 96.225 16.405 101.570 16.950 ;
        RECT 101.745 16.405 107.090 16.950 ;
        RECT 107.265 16.405 112.610 16.950 ;
        RECT 112.785 16.405 118.130 16.950 ;
        RECT 118.305 16.405 120.895 17.175 ;
        RECT 123.135 17.155 123.655 17.695 ;
        RECT 121.525 16.405 121.815 17.130 ;
        RECT 122.445 16.405 123.655 17.155 ;
        RECT 5.520 16.235 123.740 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 18.025 15.690 23.370 16.235 ;
        RECT 23.545 15.690 28.890 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 19.610 14.860 19.950 15.690 ;
        RECT 21.430 14.120 21.780 15.370 ;
        RECT 25.130 14.860 25.470 15.690 ;
        RECT 29.065 15.465 30.735 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.690 37.170 16.235 ;
        RECT 37.345 15.690 42.690 16.235 ;
        RECT 42.865 15.690 48.210 16.235 ;
        RECT 48.385 15.690 53.730 16.235 ;
        RECT 26.950 14.120 27.300 15.370 ;
        RECT 29.065 14.945 29.815 15.465 ;
        RECT 29.985 14.775 30.735 15.295 ;
        RECT 33.410 14.860 33.750 15.690 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 23.370 14.120 ;
        RECT 23.545 13.685 28.890 14.120 ;
        RECT 29.065 13.685 30.735 14.775 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 35.230 14.120 35.580 15.370 ;
        RECT 38.930 14.860 39.270 15.690 ;
        RECT 40.750 14.120 41.100 15.370 ;
        RECT 44.450 14.860 44.790 15.690 ;
        RECT 46.270 14.120 46.620 15.370 ;
        RECT 49.970 14.860 50.310 15.690 ;
        RECT 53.905 15.465 56.495 16.235 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 57.585 15.690 62.930 16.235 ;
        RECT 63.105 15.690 68.450 16.235 ;
        RECT 68.625 15.690 73.970 16.235 ;
        RECT 74.145 15.690 79.490 16.235 ;
        RECT 51.790 14.120 52.140 15.370 ;
        RECT 53.905 14.945 55.115 15.465 ;
        RECT 55.285 14.775 56.495 15.295 ;
        RECT 59.170 14.860 59.510 15.690 ;
        RECT 31.825 13.685 37.170 14.120 ;
        RECT 37.345 13.685 42.690 14.120 ;
        RECT 42.865 13.685 48.210 14.120 ;
        RECT 48.385 13.685 53.730 14.120 ;
        RECT 53.905 13.685 56.495 14.775 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 60.990 14.120 61.340 15.370 ;
        RECT 64.690 14.860 65.030 15.690 ;
        RECT 66.510 14.120 66.860 15.370 ;
        RECT 70.210 14.860 70.550 15.690 ;
        RECT 72.030 14.120 72.380 15.370 ;
        RECT 75.730 14.860 76.070 15.690 ;
        RECT 79.665 15.465 82.255 16.235 ;
        RECT 82.885 15.510 83.175 16.235 ;
        RECT 83.345 15.690 88.690 16.235 ;
        RECT 88.865 15.690 94.210 16.235 ;
        RECT 94.385 15.690 99.730 16.235 ;
        RECT 99.905 15.690 105.250 16.235 ;
        RECT 77.550 14.120 77.900 15.370 ;
        RECT 79.665 14.945 80.875 15.465 ;
        RECT 81.045 14.775 82.255 15.295 ;
        RECT 84.930 14.860 85.270 15.690 ;
        RECT 57.585 13.685 62.930 14.120 ;
        RECT 63.105 13.685 68.450 14.120 ;
        RECT 68.625 13.685 73.970 14.120 ;
        RECT 74.145 13.685 79.490 14.120 ;
        RECT 79.665 13.685 82.255 14.775 ;
        RECT 82.885 13.685 83.175 14.850 ;
        RECT 86.750 14.120 87.100 15.370 ;
        RECT 90.450 14.860 90.790 15.690 ;
        RECT 92.270 14.120 92.620 15.370 ;
        RECT 95.970 14.860 96.310 15.690 ;
        RECT 97.790 14.120 98.140 15.370 ;
        RECT 101.490 14.860 101.830 15.690 ;
        RECT 105.425 15.465 108.015 16.235 ;
        RECT 108.645 15.510 108.935 16.235 ;
        RECT 109.105 15.690 114.450 16.235 ;
        RECT 114.625 15.690 119.970 16.235 ;
        RECT 103.310 14.120 103.660 15.370 ;
        RECT 105.425 14.945 106.635 15.465 ;
        RECT 106.805 14.775 108.015 15.295 ;
        RECT 110.690 14.860 111.030 15.690 ;
        RECT 83.345 13.685 88.690 14.120 ;
        RECT 88.865 13.685 94.210 14.120 ;
        RECT 94.385 13.685 99.730 14.120 ;
        RECT 99.905 13.685 105.250 14.120 ;
        RECT 105.425 13.685 108.015 14.775 ;
        RECT 108.645 13.685 108.935 14.850 ;
        RECT 112.510 14.120 112.860 15.370 ;
        RECT 116.210 14.860 116.550 15.690 ;
        RECT 120.145 15.465 121.815 16.235 ;
        RECT 122.445 15.485 123.655 16.235 ;
        RECT 118.030 14.120 118.380 15.370 ;
        RECT 120.145 14.945 120.895 15.465 ;
        RECT 121.065 14.775 121.815 15.295 ;
        RECT 109.105 13.685 114.450 14.120 ;
        RECT 114.625 13.685 119.970 14.120 ;
        RECT 120.145 13.685 121.815 14.775 ;
        RECT 122.445 14.775 122.965 15.315 ;
        RECT 123.135 14.945 123.655 15.485 ;
        RECT 122.445 13.685 123.655 14.775 ;
        RECT 5.520 13.515 123.740 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 12.505 13.080 17.850 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 14.090 11.510 14.430 12.340 ;
        RECT 15.910 11.830 16.260 13.080 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 13.080 24.290 13.515 ;
        RECT 24.465 13.080 29.810 13.515 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 12.505 10.965 17.850 11.510 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 20.530 11.510 20.870 12.340 ;
        RECT 22.350 11.830 22.700 13.080 ;
        RECT 26.050 11.510 26.390 12.340 ;
        RECT 27.870 11.830 28.220 13.080 ;
        RECT 29.985 12.425 31.195 13.515 ;
        RECT 29.985 11.715 30.505 12.255 ;
        RECT 30.675 11.885 31.195 12.425 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 31.825 13.080 37.170 13.515 ;
        RECT 37.345 13.080 42.690 13.515 ;
        RECT 18.945 10.965 24.290 11.510 ;
        RECT 24.465 10.965 29.810 11.510 ;
        RECT 29.985 10.965 31.195 11.715 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 33.410 11.510 33.750 12.340 ;
        RECT 35.230 11.830 35.580 13.080 ;
        RECT 38.930 11.510 39.270 12.340 ;
        RECT 40.750 11.830 41.100 13.080 ;
        RECT 42.865 12.425 44.075 13.515 ;
        RECT 42.865 11.715 43.385 12.255 ;
        RECT 43.555 11.885 44.075 12.425 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 44.705 13.080 50.050 13.515 ;
        RECT 50.225 13.080 55.570 13.515 ;
        RECT 31.825 10.965 37.170 11.510 ;
        RECT 37.345 10.965 42.690 11.510 ;
        RECT 42.865 10.965 44.075 11.715 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 46.290 11.510 46.630 12.340 ;
        RECT 48.110 11.830 48.460 13.080 ;
        RECT 51.810 11.510 52.150 12.340 ;
        RECT 53.630 11.830 53.980 13.080 ;
        RECT 55.745 12.425 56.955 13.515 ;
        RECT 55.745 11.715 56.265 12.255 ;
        RECT 56.435 11.885 56.955 12.425 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 57.585 13.080 62.930 13.515 ;
        RECT 63.105 13.080 68.450 13.515 ;
        RECT 44.705 10.965 50.050 11.510 ;
        RECT 50.225 10.965 55.570 11.510 ;
        RECT 55.745 10.965 56.955 11.715 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 59.170 11.510 59.510 12.340 ;
        RECT 60.990 11.830 61.340 13.080 ;
        RECT 64.690 11.510 65.030 12.340 ;
        RECT 66.510 11.830 66.860 13.080 ;
        RECT 68.625 12.425 69.835 13.515 ;
        RECT 68.625 11.715 69.145 12.255 ;
        RECT 69.315 11.885 69.835 12.425 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 70.465 13.080 75.810 13.515 ;
        RECT 75.985 13.080 81.330 13.515 ;
        RECT 57.585 10.965 62.930 11.510 ;
        RECT 63.105 10.965 68.450 11.510 ;
        RECT 68.625 10.965 69.835 11.715 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 72.050 11.510 72.390 12.340 ;
        RECT 73.870 11.830 74.220 13.080 ;
        RECT 77.570 11.510 77.910 12.340 ;
        RECT 79.390 11.830 79.740 13.080 ;
        RECT 81.505 12.425 82.715 13.515 ;
        RECT 81.505 11.715 82.025 12.255 ;
        RECT 82.195 11.885 82.715 12.425 ;
        RECT 82.885 12.350 83.175 13.515 ;
        RECT 83.345 13.080 88.690 13.515 ;
        RECT 88.865 13.080 94.210 13.515 ;
        RECT 70.465 10.965 75.810 11.510 ;
        RECT 75.985 10.965 81.330 11.510 ;
        RECT 81.505 10.965 82.715 11.715 ;
        RECT 82.885 10.965 83.175 11.690 ;
        RECT 84.930 11.510 85.270 12.340 ;
        RECT 86.750 11.830 87.100 13.080 ;
        RECT 90.450 11.510 90.790 12.340 ;
        RECT 92.270 11.830 92.620 13.080 ;
        RECT 94.385 12.425 95.595 13.515 ;
        RECT 94.385 11.715 94.905 12.255 ;
        RECT 95.075 11.885 95.595 12.425 ;
        RECT 95.765 12.350 96.055 13.515 ;
        RECT 96.225 13.080 101.570 13.515 ;
        RECT 101.745 13.080 107.090 13.515 ;
        RECT 83.345 10.965 88.690 11.510 ;
        RECT 88.865 10.965 94.210 11.510 ;
        RECT 94.385 10.965 95.595 11.715 ;
        RECT 95.765 10.965 96.055 11.690 ;
        RECT 97.810 11.510 98.150 12.340 ;
        RECT 99.630 11.830 99.980 13.080 ;
        RECT 103.330 11.510 103.670 12.340 ;
        RECT 105.150 11.830 105.500 13.080 ;
        RECT 107.265 12.425 108.475 13.515 ;
        RECT 107.265 11.715 107.785 12.255 ;
        RECT 107.955 11.885 108.475 12.425 ;
        RECT 108.645 12.350 108.935 13.515 ;
        RECT 109.105 13.080 114.450 13.515 ;
        RECT 114.625 13.080 119.970 13.515 ;
        RECT 96.225 10.965 101.570 11.510 ;
        RECT 101.745 10.965 107.090 11.510 ;
        RECT 107.265 10.965 108.475 11.715 ;
        RECT 108.645 10.965 108.935 11.690 ;
        RECT 110.690 11.510 111.030 12.340 ;
        RECT 112.510 11.830 112.860 13.080 ;
        RECT 116.210 11.510 116.550 12.340 ;
        RECT 118.030 11.830 118.380 13.080 ;
        RECT 120.145 12.425 121.355 13.515 ;
        RECT 120.145 11.715 120.665 12.255 ;
        RECT 120.835 11.885 121.355 12.425 ;
        RECT 121.525 12.350 121.815 13.515 ;
        RECT 122.445 12.425 123.655 13.515 ;
        RECT 122.445 11.885 122.965 12.425 ;
        RECT 123.135 11.715 123.655 12.255 ;
        RECT 109.105 10.965 114.450 11.510 ;
        RECT 114.625 10.965 119.970 11.510 ;
        RECT 120.145 10.965 121.355 11.715 ;
        RECT 121.525 10.965 121.815 11.690 ;
        RECT 122.445 10.965 123.655 11.715 ;
        RECT 5.520 10.795 123.740 10.965 ;
      LAYER met1 ;
        RECT 5.520 127.600 123.740 128.080 ;
        RECT 121.065 127.400 121.355 127.445 ;
        RECT 125.650 127.400 125.970 127.460 ;
        RECT 121.065 127.260 125.970 127.400 ;
        RECT 121.065 127.215 121.355 127.260 ;
        RECT 125.650 127.200 125.970 127.260 ;
        RECT 113.195 127.060 113.485 127.105 ;
        RECT 115.085 127.060 115.375 127.105 ;
        RECT 118.205 127.060 118.495 127.105 ;
        RECT 113.195 126.920 118.495 127.060 ;
        RECT 113.195 126.875 113.485 126.920 ;
        RECT 115.085 126.875 115.375 126.920 ;
        RECT 118.205 126.875 118.495 126.920 ;
        RECT 111.850 126.380 112.170 126.440 ;
        RECT 112.325 126.380 112.615 126.425 ;
        RECT 111.850 126.240 112.615 126.380 ;
        RECT 111.850 126.180 112.170 126.240 ;
        RECT 112.325 126.195 112.615 126.240 ;
        RECT 112.790 126.380 113.080 126.425 ;
        RECT 114.625 126.380 114.915 126.425 ;
        RECT 118.205 126.380 118.495 126.425 ;
        RECT 112.790 126.240 118.495 126.380 ;
        RECT 112.790 126.195 113.080 126.240 ;
        RECT 114.625 126.195 114.915 126.240 ;
        RECT 118.205 126.195 118.495 126.240 ;
        RECT 113.690 125.840 114.010 126.100 ;
        RECT 115.985 126.040 116.635 126.085 ;
        RECT 117.370 126.040 117.690 126.100 ;
        RECT 119.285 126.085 119.575 126.400 ;
        RECT 119.285 126.040 119.875 126.085 ;
        RECT 115.985 125.900 119.875 126.040 ;
        RECT 115.985 125.855 116.635 125.900 ;
        RECT 117.370 125.840 117.690 125.900 ;
        RECT 119.585 125.855 119.875 125.900 ;
        RECT 5.520 124.880 123.740 125.360 ;
        RECT 111.850 124.680 112.170 124.740 ;
        RECT 111.850 124.540 117.140 124.680 ;
        RECT 111.850 124.480 112.170 124.540 ;
        RECT 17.550 124.385 17.870 124.400 ;
        RECT 61.710 124.385 62.030 124.400 ;
        RECT 13.985 124.340 14.275 124.385 ;
        RECT 17.225 124.340 17.875 124.385 ;
        RECT 13.985 124.200 17.875 124.340 ;
        RECT 13.985 124.155 14.575 124.200 ;
        RECT 17.225 124.155 17.875 124.200 ;
        RECT 42.385 124.340 43.035 124.385 ;
        RECT 45.985 124.340 46.275 124.385 ;
        RECT 42.385 124.200 46.275 124.340 ;
        RECT 42.385 124.155 43.035 124.200 ;
        RECT 45.685 124.155 46.275 124.200 ;
        RECT 51.585 124.340 52.235 124.385 ;
        RECT 55.185 124.340 55.475 124.385 ;
        RECT 51.585 124.200 55.475 124.340 ;
        RECT 51.585 124.155 52.235 124.200 ;
        RECT 54.885 124.155 55.475 124.200 ;
        RECT 61.245 124.340 62.030 124.385 ;
        RECT 64.845 124.340 65.135 124.385 ;
        RECT 61.245 124.200 65.135 124.340 ;
        RECT 61.245 124.155 62.030 124.200 ;
        RECT 3.750 124.000 4.070 124.060 ;
        RECT 6.985 124.000 7.275 124.045 ;
        RECT 3.750 123.860 7.275 124.000 ;
        RECT 3.750 123.800 4.070 123.860 ;
        RECT 6.985 123.815 7.275 123.860 ;
        RECT 14.285 123.840 14.575 124.155 ;
        RECT 17.550 124.140 17.870 124.155 ;
        RECT 45.685 124.060 45.975 124.155 ;
        RECT 15.365 124.000 15.655 124.045 ;
        RECT 18.945 124.000 19.235 124.045 ;
        RECT 20.780 124.000 21.070 124.045 ;
        RECT 15.365 123.860 21.070 124.000 ;
        RECT 15.365 123.815 15.655 123.860 ;
        RECT 18.945 123.815 19.235 123.860 ;
        RECT 20.780 123.815 21.070 123.860 ;
        RECT 21.690 124.000 22.010 124.060 ;
        RECT 25.845 124.000 26.135 124.045 ;
        RECT 29.525 124.000 29.815 124.045 ;
        RECT 33.650 124.000 33.970 124.060 ;
        RECT 21.690 123.860 33.970 124.000 ;
        RECT 21.690 123.800 22.010 123.860 ;
        RECT 25.845 123.815 26.135 123.860 ;
        RECT 29.525 123.815 29.815 123.860 ;
        RECT 33.650 123.800 33.970 123.860 ;
        RECT 39.190 124.000 39.480 124.045 ;
        RECT 41.025 124.000 41.315 124.045 ;
        RECT 44.605 124.000 44.895 124.045 ;
        RECT 39.190 123.860 44.895 124.000 ;
        RECT 39.190 123.815 39.480 123.860 ;
        RECT 41.025 123.815 41.315 123.860 ;
        RECT 44.605 123.815 44.895 123.860 ;
        RECT 45.610 123.840 45.975 124.060 ;
        RECT 48.390 124.000 48.680 124.045 ;
        RECT 50.225 124.000 50.515 124.045 ;
        RECT 53.805 124.000 54.095 124.045 ;
        RECT 48.390 123.860 54.095 124.000 ;
        RECT 45.610 123.800 45.930 123.840 ;
        RECT 48.390 123.815 48.680 123.860 ;
        RECT 50.225 123.815 50.515 123.860 ;
        RECT 53.805 123.815 54.095 123.860 ;
        RECT 54.885 124.000 55.175 124.155 ;
        RECT 61.710 124.140 62.030 124.155 ;
        RECT 64.545 124.155 65.135 124.200 ;
        RECT 70.905 124.340 71.555 124.385 ;
        RECT 74.505 124.340 74.795 124.385 ;
        RECT 70.905 124.200 74.795 124.340 ;
        RECT 70.905 124.155 71.555 124.200 ;
        RECT 74.205 124.155 74.795 124.200 ;
        RECT 87.005 124.340 87.655 124.385 ;
        RECT 90.605 124.340 90.895 124.385 ;
        RECT 87.005 124.200 90.895 124.340 ;
        RECT 87.005 124.155 87.655 124.200 ;
        RECT 90.305 124.155 90.895 124.200 ;
        RECT 94.025 124.340 94.315 124.385 ;
        RECT 97.265 124.340 97.915 124.385 ;
        RECT 94.025 124.200 97.915 124.340 ;
        RECT 94.025 124.155 94.615 124.200 ;
        RECT 97.265 124.155 97.915 124.200 ;
        RECT 110.585 124.340 110.875 124.385 ;
        RECT 113.825 124.340 114.475 124.385 ;
        RECT 110.585 124.200 114.475 124.340 ;
        RECT 117.000 124.340 117.140 124.540 ;
        RECT 117.000 124.200 118.060 124.340 ;
        RECT 110.585 124.155 111.175 124.200 ;
        RECT 113.825 124.155 114.475 124.200 ;
        RECT 57.110 124.000 57.430 124.060 ;
        RECT 54.885 123.860 57.430 124.000 ;
        RECT 54.885 123.840 55.175 123.860 ;
        RECT 57.110 123.800 57.430 123.860 ;
        RECT 58.050 124.000 58.340 124.045 ;
        RECT 59.885 124.000 60.175 124.045 ;
        RECT 63.465 124.000 63.755 124.045 ;
        RECT 58.050 123.860 63.755 124.000 ;
        RECT 58.050 123.815 58.340 123.860 ;
        RECT 59.885 123.815 60.175 123.860 ;
        RECT 63.465 123.815 63.755 123.860 ;
        RECT 64.545 123.840 64.835 124.155 ;
        RECT 74.205 124.060 74.495 124.155 ;
        RECT 67.710 124.000 68.000 124.045 ;
        RECT 69.545 124.000 69.835 124.045 ;
        RECT 73.125 124.000 73.415 124.045 ;
        RECT 67.710 123.860 73.415 124.000 ;
        RECT 67.710 123.815 68.000 123.860 ;
        RECT 69.545 123.815 69.835 123.860 ;
        RECT 73.125 123.815 73.415 123.860 ;
        RECT 74.130 123.840 74.495 124.060 ;
        RECT 83.810 124.000 84.100 124.045 ;
        RECT 85.645 124.000 85.935 124.045 ;
        RECT 89.225 124.000 89.515 124.045 ;
        RECT 83.810 123.860 89.515 124.000 ;
        RECT 74.130 123.800 74.450 123.840 ;
        RECT 83.810 123.815 84.100 123.860 ;
        RECT 85.645 123.815 85.935 123.860 ;
        RECT 89.225 123.815 89.515 123.860 ;
        RECT 89.770 124.000 90.090 124.060 ;
        RECT 90.305 124.000 90.595 124.155 ;
        RECT 89.770 123.860 90.595 124.000 ;
        RECT 89.770 123.800 90.090 123.860 ;
        RECT 90.305 123.840 90.595 123.860 ;
        RECT 92.990 124.000 93.310 124.060 ;
        RECT 94.325 124.000 94.615 124.155 ;
        RECT 92.990 123.860 94.615 124.000 ;
        RECT 92.990 123.800 93.310 123.860 ;
        RECT 94.325 123.840 94.615 123.860 ;
        RECT 95.405 124.000 95.695 124.045 ;
        RECT 98.985 124.000 99.275 124.045 ;
        RECT 100.820 124.000 101.110 124.045 ;
        RECT 95.405 123.860 101.110 124.000 ;
        RECT 95.405 123.815 95.695 123.860 ;
        RECT 98.985 123.815 99.275 123.860 ;
        RECT 100.820 123.815 101.110 123.860 ;
        RECT 105.870 124.000 106.190 124.060 ;
        RECT 110.885 124.000 111.175 124.155 ;
        RECT 117.920 124.045 118.060 124.200 ;
        RECT 105.870 123.860 111.175 124.000 ;
        RECT 105.870 123.800 106.190 123.860 ;
        RECT 110.885 123.840 111.175 123.860 ;
        RECT 111.965 124.000 112.255 124.045 ;
        RECT 115.545 124.000 115.835 124.045 ;
        RECT 117.380 124.000 117.670 124.045 ;
        RECT 111.965 123.860 117.670 124.000 ;
        RECT 111.965 123.815 112.255 123.860 ;
        RECT 115.545 123.815 115.835 123.860 ;
        RECT 117.380 123.815 117.670 123.860 ;
        RECT 117.845 123.815 118.135 124.045 ;
        RECT 12.505 123.660 12.795 123.705 ;
        RECT 16.170 123.660 16.490 123.720 ;
        RECT 12.505 123.520 16.490 123.660 ;
        RECT 12.505 123.475 12.795 123.520 ;
        RECT 16.170 123.460 16.490 123.520 ;
        RECT 19.850 123.460 20.170 123.720 ;
        RECT 21.245 123.660 21.535 123.705 ;
        RECT 20.860 123.520 21.535 123.660 ;
        RECT 15.365 123.320 15.655 123.365 ;
        RECT 18.485 123.320 18.775 123.365 ;
        RECT 20.375 123.320 20.665 123.365 ;
        RECT 15.365 123.180 20.665 123.320 ;
        RECT 15.365 123.135 15.655 123.180 ;
        RECT 18.485 123.135 18.775 123.180 ;
        RECT 20.375 123.135 20.665 123.180 ;
        RECT 20.860 123.040 21.000 123.520 ;
        RECT 21.245 123.475 21.535 123.520 ;
        RECT 38.710 123.460 39.030 123.720 ;
        RECT 40.105 123.660 40.395 123.705 ;
        RECT 46.070 123.660 46.390 123.720 ;
        RECT 40.105 123.520 46.390 123.660 ;
        RECT 40.105 123.475 40.395 123.520 ;
        RECT 46.070 123.460 46.390 123.520 ;
        RECT 47.925 123.475 48.215 123.705 ;
        RECT 39.595 123.320 39.885 123.365 ;
        RECT 41.485 123.320 41.775 123.365 ;
        RECT 44.605 123.320 44.895 123.365 ;
        RECT 39.595 123.180 44.895 123.320 ;
        RECT 39.595 123.135 39.885 123.180 ;
        RECT 41.485 123.135 41.775 123.180 ;
        RECT 44.605 123.135 44.895 123.180 ;
        RECT 47.450 123.120 47.770 123.380 ;
        RECT 7.905 122.980 8.195 123.025 ;
        RECT 18.930 122.980 19.250 123.040 ;
        RECT 7.905 122.840 19.250 122.980 ;
        RECT 7.905 122.795 8.195 122.840 ;
        RECT 18.930 122.780 19.250 122.840 ;
        RECT 20.770 122.780 21.090 123.040 ;
        RECT 26.305 122.980 26.595 123.025 ;
        RECT 26.750 122.980 27.070 123.040 ;
        RECT 26.305 122.840 27.070 122.980 ;
        RECT 26.305 122.795 26.595 122.840 ;
        RECT 26.750 122.780 27.070 122.840 ;
        RECT 29.510 122.980 29.830 123.040 ;
        RECT 29.985 122.980 30.275 123.025 ;
        RECT 29.510 122.840 30.275 122.980 ;
        RECT 29.510 122.780 29.830 122.840 ;
        RECT 29.985 122.795 30.275 122.840 ;
        RECT 39.170 122.980 39.490 123.040 ;
        RECT 48.000 122.980 48.140 123.475 ;
        RECT 49.290 123.460 49.610 123.720 ;
        RECT 57.585 123.475 57.875 123.705 ;
        RECT 48.795 123.320 49.085 123.365 ;
        RECT 50.685 123.320 50.975 123.365 ;
        RECT 53.805 123.320 54.095 123.365 ;
        RECT 48.795 123.180 54.095 123.320 ;
        RECT 48.795 123.135 49.085 123.180 ;
        RECT 50.685 123.135 50.975 123.180 ;
        RECT 53.805 123.135 54.095 123.180 ;
        RECT 54.810 123.320 55.130 123.380 ;
        RECT 56.665 123.320 56.955 123.365 ;
        RECT 54.810 123.180 56.955 123.320 ;
        RECT 54.810 123.120 55.130 123.180 ;
        RECT 56.665 123.135 56.955 123.180 ;
        RECT 57.660 122.980 57.800 123.475 ;
        RECT 58.950 123.460 59.270 123.720 ;
        RECT 61.250 123.660 61.570 123.720 ;
        RECT 66.325 123.660 66.615 123.705 ;
        RECT 61.250 123.520 66.615 123.660 ;
        RECT 61.250 123.460 61.570 123.520 ;
        RECT 66.325 123.475 66.615 123.520 ;
        RECT 67.230 123.460 67.550 123.720 ;
        RECT 68.625 123.660 68.915 123.705 ;
        RECT 69.070 123.660 69.390 123.720 ;
        RECT 68.625 123.520 69.390 123.660 ;
        RECT 68.625 123.475 68.915 123.520 ;
        RECT 69.070 123.460 69.390 123.520 ;
        RECT 74.590 123.660 74.910 123.720 ;
        RECT 75.985 123.660 76.275 123.705 ;
        RECT 74.590 123.520 76.275 123.660 ;
        RECT 74.590 123.460 74.910 123.520 ;
        RECT 75.985 123.475 76.275 123.520 ;
        RECT 83.330 123.460 83.650 123.720 ;
        RECT 84.725 123.660 85.015 123.705 ;
        RECT 87.930 123.660 88.250 123.720 ;
        RECT 84.725 123.520 88.250 123.660 ;
        RECT 84.725 123.475 85.015 123.520 ;
        RECT 87.930 123.460 88.250 123.520 ;
        RECT 88.390 123.660 88.710 123.720 ;
        RECT 92.085 123.660 92.375 123.705 ;
        RECT 88.390 123.520 92.375 123.660 ;
        RECT 88.390 123.460 88.710 123.520 ;
        RECT 92.085 123.475 92.375 123.520 ;
        RECT 92.530 123.460 92.850 123.720 ;
        RECT 93.450 123.660 93.770 123.720 ;
        RECT 99.905 123.660 100.195 123.705 ;
        RECT 93.450 123.520 100.195 123.660 ;
        RECT 93.450 123.460 93.770 123.520 ;
        RECT 99.905 123.475 100.195 123.520 ;
        RECT 101.285 123.475 101.575 123.705 ;
        RECT 106.330 123.660 106.650 123.720 ;
        RECT 109.105 123.660 109.395 123.705 ;
        RECT 116.465 123.660 116.755 123.705 ;
        RECT 106.330 123.520 109.395 123.660 ;
        RECT 58.455 123.320 58.745 123.365 ;
        RECT 60.345 123.320 60.635 123.365 ;
        RECT 63.465 123.320 63.755 123.365 ;
        RECT 58.455 123.180 63.755 123.320 ;
        RECT 58.455 123.135 58.745 123.180 ;
        RECT 60.345 123.135 60.635 123.180 ;
        RECT 63.465 123.135 63.755 123.180 ;
        RECT 68.115 123.320 68.405 123.365 ;
        RECT 70.005 123.320 70.295 123.365 ;
        RECT 73.125 123.320 73.415 123.365 ;
        RECT 68.115 123.180 73.415 123.320 ;
        RECT 68.115 123.135 68.405 123.180 ;
        RECT 70.005 123.135 70.295 123.180 ;
        RECT 73.125 123.135 73.415 123.180 ;
        RECT 84.215 123.320 84.505 123.365 ;
        RECT 86.105 123.320 86.395 123.365 ;
        RECT 89.225 123.320 89.515 123.365 ;
        RECT 84.215 123.180 89.515 123.320 ;
        RECT 84.215 123.135 84.505 123.180 ;
        RECT 86.105 123.135 86.395 123.180 ;
        RECT 89.225 123.135 89.515 123.180 ;
        RECT 95.405 123.320 95.695 123.365 ;
        RECT 98.525 123.320 98.815 123.365 ;
        RECT 100.415 123.320 100.705 123.365 ;
        RECT 95.405 123.180 100.705 123.320 ;
        RECT 95.405 123.135 95.695 123.180 ;
        RECT 98.525 123.135 98.815 123.180 ;
        RECT 100.415 123.135 100.705 123.180 ;
        RECT 39.170 122.840 57.800 122.980 ;
        RECT 96.210 122.980 96.530 123.040 ;
        RECT 101.360 122.980 101.500 123.475 ;
        RECT 106.330 123.460 106.650 123.520 ;
        RECT 109.105 123.475 109.395 123.520 ;
        RECT 109.640 123.520 116.755 123.660 ;
        RECT 103.110 123.320 103.430 123.380 ;
        RECT 109.640 123.320 109.780 123.520 ;
        RECT 116.465 123.475 116.755 123.520 ;
        RECT 103.110 123.180 109.780 123.320 ;
        RECT 111.965 123.320 112.255 123.365 ;
        RECT 115.085 123.320 115.375 123.365 ;
        RECT 116.975 123.320 117.265 123.365 ;
        RECT 111.965 123.180 117.265 123.320 ;
        RECT 103.110 123.120 103.430 123.180 ;
        RECT 111.965 123.135 112.255 123.180 ;
        RECT 115.085 123.135 115.375 123.180 ;
        RECT 116.975 123.135 117.265 123.180 ;
        RECT 96.210 122.840 101.500 122.980 ;
        RECT 39.170 122.780 39.490 122.840 ;
        RECT 96.210 122.780 96.530 122.840 ;
        RECT 5.520 122.160 123.740 122.640 ;
        RECT 11.570 121.960 11.890 122.020 ;
        RECT 15.725 121.960 16.015 122.005 ;
        RECT 11.570 121.820 16.015 121.960 ;
        RECT 11.570 121.760 11.890 121.820 ;
        RECT 15.725 121.775 16.015 121.820 ;
        RECT 17.550 121.960 17.870 122.020 ;
        RECT 19.405 121.960 19.695 122.005 ;
        RECT 17.550 121.820 19.695 121.960 ;
        RECT 17.550 121.760 17.870 121.820 ;
        RECT 19.405 121.775 19.695 121.820 ;
        RECT 29.050 121.960 29.370 122.020 ;
        RECT 33.205 121.960 33.495 122.005 ;
        RECT 41.930 121.960 42.250 122.020 ;
        RECT 43.785 121.960 44.075 122.005 ;
        RECT 29.050 121.820 33.495 121.960 ;
        RECT 29.050 121.760 29.370 121.820 ;
        RECT 33.205 121.775 33.495 121.820 ;
        RECT 34.430 121.820 41.700 121.960 ;
        RECT 7.855 121.620 8.145 121.665 ;
        RECT 9.745 121.620 10.035 121.665 ;
        RECT 12.865 121.620 13.155 121.665 ;
        RECT 7.855 121.480 13.155 121.620 ;
        RECT 7.855 121.435 8.145 121.480 ;
        RECT 9.745 121.435 10.035 121.480 ;
        RECT 12.865 121.435 13.155 121.480 ;
        RECT 18.930 121.620 19.250 121.680 ;
        RECT 25.335 121.620 25.625 121.665 ;
        RECT 27.225 121.620 27.515 121.665 ;
        RECT 30.345 121.620 30.635 121.665 ;
        RECT 18.930 121.480 25.140 121.620 ;
        RECT 18.930 121.420 19.250 121.480 ;
        RECT 20.310 121.280 20.630 121.340 ;
        RECT 24.465 121.280 24.755 121.325 ;
        RECT 20.310 121.140 24.755 121.280 ;
        RECT 25.000 121.280 25.140 121.480 ;
        RECT 25.335 121.480 30.635 121.620 ;
        RECT 25.335 121.435 25.625 121.480 ;
        RECT 27.225 121.435 27.515 121.480 ;
        RECT 30.345 121.435 30.635 121.480 ;
        RECT 34.430 121.280 34.570 121.820 ;
        RECT 35.915 121.620 36.205 121.665 ;
        RECT 37.805 121.620 38.095 121.665 ;
        RECT 40.925 121.620 41.215 121.665 ;
        RECT 35.915 121.480 41.215 121.620 ;
        RECT 35.915 121.435 36.205 121.480 ;
        RECT 37.805 121.435 38.095 121.480 ;
        RECT 40.925 121.435 41.215 121.480 ;
        RECT 25.000 121.140 34.570 121.280 ;
        RECT 35.045 121.280 35.335 121.325 ;
        RECT 39.170 121.280 39.490 121.340 ;
        RECT 35.045 121.140 39.490 121.280 ;
        RECT 41.560 121.280 41.700 121.820 ;
        RECT 41.930 121.820 44.075 121.960 ;
        RECT 41.930 121.760 42.250 121.820 ;
        RECT 43.785 121.775 44.075 121.820 ;
        RECT 46.070 121.960 46.390 122.020 ;
        RECT 47.005 121.960 47.295 122.005 ;
        RECT 46.070 121.820 47.295 121.960 ;
        RECT 46.070 121.760 46.390 121.820 ;
        RECT 47.005 121.775 47.295 121.820 ;
        RECT 49.290 121.960 49.610 122.020 ;
        RECT 53.445 121.960 53.735 122.005 ;
        RECT 49.290 121.820 53.735 121.960 ;
        RECT 49.290 121.760 49.610 121.820 ;
        RECT 53.445 121.775 53.735 121.820 ;
        RECT 56.665 121.960 56.955 122.005 ;
        RECT 61.710 121.960 62.030 122.020 ;
        RECT 56.665 121.820 62.030 121.960 ;
        RECT 56.665 121.775 56.955 121.820 ;
        RECT 61.710 121.760 62.030 121.820 ;
        RECT 73.225 121.960 73.515 122.005 ;
        RECT 74.130 121.960 74.450 122.020 ;
        RECT 73.225 121.820 74.450 121.960 ;
        RECT 73.225 121.775 73.515 121.820 ;
        RECT 74.130 121.760 74.450 121.820 ;
        RECT 81.030 121.960 81.350 122.020 ;
        RECT 83.345 121.960 83.635 122.005 ;
        RECT 81.030 121.820 83.635 121.960 ;
        RECT 81.030 121.760 81.350 121.820 ;
        RECT 83.345 121.775 83.635 121.820 ;
        RECT 87.930 121.760 88.250 122.020 ;
        RECT 89.770 121.760 90.090 122.020 ;
        RECT 92.990 121.760 93.310 122.020 ;
        RECT 105.870 121.760 106.190 122.020 ;
        RECT 114.150 121.960 114.470 122.020 ;
        RECT 115.545 121.960 115.835 122.005 ;
        RECT 114.150 121.820 115.835 121.960 ;
        RECT 114.150 121.760 114.470 121.820 ;
        RECT 115.545 121.775 115.835 121.820 ;
        RECT 117.370 121.960 117.690 122.020 ;
        RECT 117.845 121.960 118.135 122.005 ;
        RECT 117.370 121.820 118.135 121.960 ;
        RECT 117.370 121.760 117.690 121.820 ;
        RECT 117.845 121.775 118.135 121.820 ;
        RECT 45.610 121.620 45.930 121.680 ;
        RECT 48.845 121.620 49.135 121.665 ;
        RECT 45.610 121.480 49.135 121.620 ;
        RECT 45.610 121.420 45.930 121.480 ;
        RECT 48.845 121.435 49.135 121.480 ;
        RECT 55.745 121.620 56.035 121.665 ;
        RECT 58.950 121.620 59.270 121.680 ;
        RECT 55.745 121.480 59.270 121.620 ;
        RECT 55.745 121.435 56.035 121.480 ;
        RECT 58.950 121.420 59.270 121.480 ;
        RECT 75.475 121.620 75.765 121.665 ;
        RECT 77.365 121.620 77.655 121.665 ;
        RECT 80.485 121.620 80.775 121.665 ;
        RECT 75.475 121.480 80.775 121.620 ;
        RECT 75.475 121.435 75.765 121.480 ;
        RECT 77.365 121.435 77.655 121.480 ;
        RECT 80.485 121.435 80.775 121.480 ;
        RECT 97.095 121.620 97.385 121.665 ;
        RECT 98.985 121.620 99.275 121.665 ;
        RECT 102.105 121.620 102.395 121.665 ;
        RECT 97.095 121.480 102.395 121.620 ;
        RECT 97.095 121.435 97.385 121.480 ;
        RECT 98.985 121.435 99.275 121.480 ;
        RECT 102.105 121.435 102.395 121.480 ;
        RECT 107.675 121.620 107.965 121.665 ;
        RECT 109.565 121.620 109.855 121.665 ;
        RECT 112.685 121.620 112.975 121.665 ;
        RECT 107.675 121.480 112.975 121.620 ;
        RECT 107.675 121.435 107.965 121.480 ;
        RECT 109.565 121.435 109.855 121.480 ;
        RECT 112.685 121.435 112.975 121.480 ;
        RECT 52.050 121.280 52.370 121.340 ;
        RECT 41.560 121.140 52.370 121.280 ;
        RECT 20.310 121.080 20.630 121.140 ;
        RECT 24.465 121.095 24.755 121.140 ;
        RECT 35.045 121.095 35.335 121.140 ;
        RECT 39.170 121.080 39.490 121.140 ;
        RECT 52.050 121.080 52.370 121.140 ;
        RECT 57.110 121.280 57.430 121.340 ;
        RECT 58.045 121.280 58.335 121.325 ;
        RECT 106.805 121.280 107.095 121.325 ;
        RECT 108.630 121.280 108.950 121.340 ;
        RECT 111.850 121.280 112.170 121.340 ;
        RECT 57.110 121.140 58.335 121.280 ;
        RECT 57.110 121.080 57.430 121.140 ;
        RECT 58.045 121.095 58.335 121.140 ;
        RECT 92.620 121.140 105.640 121.280 ;
        RECT 92.620 121.000 92.760 121.140 ;
        RECT 6.985 120.755 7.275 120.985 ;
        RECT 7.450 120.940 7.740 120.985 ;
        RECT 9.285 120.940 9.575 120.985 ;
        RECT 12.865 120.940 13.155 120.985 ;
        RECT 7.450 120.800 13.155 120.940 ;
        RECT 7.450 120.755 7.740 120.800 ;
        RECT 9.285 120.755 9.575 120.800 ;
        RECT 12.865 120.755 13.155 120.800 ;
        RECT 7.060 120.600 7.200 120.755 ;
        RECT 7.890 120.600 8.210 120.660 ;
        RECT 7.060 120.460 8.210 120.600 ;
        RECT 7.890 120.400 8.210 120.460 ;
        RECT 8.350 120.400 8.670 120.660 ;
        RECT 13.945 120.645 14.235 120.960 ;
        RECT 17.105 120.940 17.395 120.985 ;
        RECT 18.010 120.940 18.330 121.000 ;
        RECT 19.865 120.940 20.155 120.985 ;
        RECT 21.690 120.940 22.010 121.000 ;
        RECT 17.105 120.800 22.010 120.940 ;
        RECT 17.105 120.755 17.395 120.800 ;
        RECT 18.010 120.740 18.330 120.800 ;
        RECT 19.865 120.755 20.155 120.800 ;
        RECT 21.690 120.740 22.010 120.800 ;
        RECT 24.930 120.940 25.220 120.985 ;
        RECT 26.765 120.940 27.055 120.985 ;
        RECT 30.345 120.940 30.635 120.985 ;
        RECT 24.930 120.800 30.635 120.940 ;
        RECT 24.930 120.755 25.220 120.800 ;
        RECT 26.765 120.755 27.055 120.800 ;
        RECT 30.345 120.755 30.635 120.800 ;
        RECT 10.645 120.600 11.295 120.645 ;
        RECT 13.945 120.600 14.535 120.645 ;
        RECT 16.645 120.600 16.935 120.645 ;
        RECT 10.645 120.460 16.935 120.600 ;
        RECT 10.645 120.415 11.295 120.460 ;
        RECT 14.245 120.415 14.535 120.460 ;
        RECT 16.645 120.415 16.935 120.460 ;
        RECT 25.845 120.415 26.135 120.645 ;
        RECT 28.125 120.600 28.775 120.645 ;
        RECT 29.510 120.600 29.830 120.660 ;
        RECT 31.425 120.645 31.715 120.960 ;
        RECT 33.650 120.940 33.970 121.000 ;
        RECT 35.510 120.940 35.800 120.985 ;
        RECT 37.345 120.940 37.635 120.985 ;
        RECT 40.925 120.940 41.215 120.985 ;
        RECT 33.650 120.800 34.570 120.940 ;
        RECT 33.650 120.740 33.970 120.800 ;
        RECT 31.425 120.600 32.015 120.645 ;
        RECT 28.125 120.460 32.015 120.600 ;
        RECT 34.430 120.600 34.570 120.800 ;
        RECT 35.510 120.800 41.215 120.940 ;
        RECT 35.510 120.755 35.800 120.800 ;
        RECT 37.345 120.755 37.635 120.800 ;
        RECT 40.925 120.755 41.215 120.800 ;
        RECT 34.430 120.460 36.180 120.600 ;
        RECT 28.125 120.415 28.775 120.460 ;
        RECT 25.920 120.260 26.060 120.415 ;
        RECT 29.510 120.400 29.830 120.460 ;
        RECT 31.725 120.415 32.015 120.460 ;
        RECT 29.970 120.260 30.290 120.320 ;
        RECT 25.920 120.120 30.290 120.260 ;
        RECT 29.970 120.060 30.290 120.120 ;
        RECT 34.125 120.260 34.415 120.305 ;
        RECT 35.490 120.260 35.810 120.320 ;
        RECT 34.125 120.120 35.810 120.260 ;
        RECT 36.040 120.260 36.180 120.460 ;
        RECT 36.410 120.400 36.730 120.660 ;
        RECT 42.005 120.645 42.295 120.960 ;
        RECT 45.625 120.755 45.915 120.985 ;
        RECT 47.925 120.940 48.215 120.985 ;
        RECT 48.830 120.940 49.150 121.000 ;
        RECT 47.925 120.800 49.150 120.940 ;
        RECT 47.925 120.755 48.215 120.800 ;
        RECT 38.705 120.600 39.355 120.645 ;
        RECT 42.005 120.600 42.595 120.645 ;
        RECT 45.165 120.600 45.455 120.645 ;
        RECT 38.705 120.460 45.455 120.600 ;
        RECT 38.705 120.415 39.355 120.460 ;
        RECT 42.305 120.415 42.595 120.460 ;
        RECT 45.165 120.415 45.455 120.460 ;
        RECT 45.700 120.600 45.840 120.755 ;
        RECT 48.830 120.740 49.150 120.800 ;
        RECT 49.305 120.755 49.595 120.985 ;
        RECT 51.590 120.940 51.910 121.000 ;
        RECT 54.365 120.940 54.655 120.985 ;
        RECT 51.590 120.800 54.655 120.940 ;
        RECT 49.380 120.600 49.520 120.755 ;
        RECT 51.590 120.740 51.910 120.800 ;
        RECT 54.365 120.755 54.655 120.800 ;
        RECT 54.825 120.940 55.115 120.985 ;
        RECT 55.730 120.940 56.050 121.000 ;
        RECT 54.825 120.800 56.050 120.940 ;
        RECT 54.825 120.755 55.115 120.800 ;
        RECT 55.730 120.740 56.050 120.800 ;
        RECT 56.205 120.940 56.495 120.985 ;
        RECT 57.585 120.940 57.875 120.985 ;
        RECT 56.205 120.800 57.875 120.940 ;
        RECT 56.205 120.755 56.495 120.800 ;
        RECT 57.585 120.755 57.875 120.800 ;
        RECT 72.305 120.940 72.595 120.985 ;
        RECT 73.685 120.940 73.975 120.985 ;
        RECT 74.130 120.940 74.450 121.000 ;
        RECT 72.305 120.800 74.450 120.940 ;
        RECT 72.305 120.755 72.595 120.800 ;
        RECT 73.685 120.755 73.975 120.800 ;
        RECT 49.750 120.600 50.070 120.660 ;
        RECT 56.280 120.600 56.420 120.755 ;
        RECT 74.130 120.740 74.450 120.800 ;
        RECT 74.605 120.755 74.895 120.985 ;
        RECT 75.070 120.940 75.360 120.985 ;
        RECT 76.905 120.940 77.195 120.985 ;
        RECT 80.485 120.940 80.775 120.985 ;
        RECT 75.070 120.800 80.775 120.940 ;
        RECT 75.070 120.755 75.360 120.800 ;
        RECT 76.905 120.755 77.195 120.800 ;
        RECT 80.485 120.755 80.775 120.800 ;
        RECT 45.700 120.460 56.420 120.600 ;
        RECT 67.230 120.600 67.550 120.660 ;
        RECT 74.680 120.600 74.820 120.755 ;
        RECT 75.510 120.600 75.830 120.660 ;
        RECT 67.230 120.460 75.830 120.600 ;
        RECT 45.700 120.260 45.840 120.460 ;
        RECT 49.750 120.400 50.070 120.460 ;
        RECT 67.230 120.400 67.550 120.460 ;
        RECT 75.510 120.400 75.830 120.460 ;
        RECT 75.970 120.400 76.290 120.660 ;
        RECT 81.565 120.645 81.855 120.960 ;
        RECT 84.725 120.755 85.015 120.985 ;
        RECT 88.865 120.940 89.155 120.985 ;
        RECT 89.770 120.940 90.090 121.000 ;
        RECT 88.865 120.800 90.090 120.940 ;
        RECT 88.865 120.755 89.155 120.800 ;
        RECT 78.265 120.600 78.915 120.645 ;
        RECT 81.565 120.600 82.155 120.645 ;
        RECT 84.265 120.600 84.555 120.645 ;
        RECT 78.265 120.460 84.555 120.600 ;
        RECT 78.265 120.415 78.915 120.460 ;
        RECT 81.865 120.415 82.155 120.460 ;
        RECT 84.265 120.415 84.555 120.460 ;
        RECT 84.800 120.600 84.940 120.755 ;
        RECT 89.770 120.740 90.090 120.800 ;
        RECT 90.245 120.940 90.535 120.985 ;
        RECT 92.530 120.940 92.850 121.000 ;
        RECT 90.245 120.800 92.850 120.940 ;
        RECT 90.245 120.755 90.535 120.800 ;
        RECT 90.320 120.600 90.460 120.755 ;
        RECT 92.530 120.740 92.850 120.800 ;
        RECT 96.210 120.740 96.530 121.000 ;
        RECT 105.500 120.985 105.640 121.140 ;
        RECT 106.805 121.140 112.170 121.280 ;
        RECT 106.805 121.095 107.095 121.140 ;
        RECT 108.630 121.080 108.950 121.140 ;
        RECT 111.850 121.080 112.170 121.140 ;
        RECT 96.690 120.940 96.980 120.985 ;
        RECT 98.525 120.940 98.815 120.985 ;
        RECT 102.105 120.940 102.395 120.985 ;
        RECT 96.690 120.800 102.395 120.940 ;
        RECT 96.690 120.755 96.980 120.800 ;
        RECT 98.525 120.755 98.815 120.800 ;
        RECT 102.105 120.755 102.395 120.800 ;
        RECT 84.800 120.460 90.460 120.600 ;
        RECT 36.040 120.120 45.840 120.260 ;
        RECT 55.730 120.260 56.050 120.320 ;
        RECT 60.790 120.260 61.110 120.320 ;
        RECT 55.730 120.120 61.110 120.260 ;
        RECT 34.125 120.075 34.415 120.120 ;
        RECT 35.490 120.060 35.810 120.120 ;
        RECT 55.730 120.060 56.050 120.120 ;
        RECT 60.790 120.060 61.110 120.120 ;
        RECT 71.830 120.060 72.150 120.320 ;
        RECT 75.050 120.260 75.370 120.320 ;
        RECT 84.800 120.260 84.940 120.460 ;
        RECT 97.590 120.400 97.910 120.660 ;
        RECT 99.890 120.645 100.210 120.660 ;
        RECT 103.185 120.645 103.475 120.960 ;
        RECT 105.425 120.755 105.715 120.985 ;
        RECT 107.270 120.940 107.560 120.985 ;
        RECT 109.105 120.940 109.395 120.985 ;
        RECT 112.685 120.940 112.975 120.985 ;
        RECT 107.270 120.800 112.975 120.940 ;
        RECT 107.270 120.755 107.560 120.800 ;
        RECT 109.105 120.755 109.395 120.800 ;
        RECT 112.685 120.755 112.975 120.800 ;
        RECT 99.885 120.600 100.535 120.645 ;
        RECT 103.185 120.600 103.775 120.645 ;
        RECT 99.885 120.460 103.775 120.600 ;
        RECT 99.885 120.415 100.535 120.460 ;
        RECT 103.485 120.415 103.775 120.460 ;
        RECT 99.890 120.400 100.210 120.415 ;
        RECT 75.050 120.120 84.940 120.260 ;
        RECT 101.730 120.260 102.050 120.320 ;
        RECT 104.965 120.260 105.255 120.305 ;
        RECT 101.730 120.120 105.255 120.260 ;
        RECT 105.500 120.260 105.640 120.755 ;
        RECT 106.790 120.600 107.110 120.660 ;
        RECT 113.765 120.645 114.055 120.960 ;
        RECT 116.925 120.940 117.215 120.985 ;
        RECT 117.385 120.940 117.675 120.985 ;
        RECT 116.925 120.800 117.675 120.940 ;
        RECT 116.925 120.755 117.215 120.800 ;
        RECT 117.385 120.755 117.675 120.800 ;
        RECT 108.185 120.600 108.475 120.645 ;
        RECT 106.790 120.460 108.475 120.600 ;
        RECT 106.790 120.400 107.110 120.460 ;
        RECT 108.185 120.415 108.475 120.460 ;
        RECT 110.465 120.600 111.115 120.645 ;
        RECT 113.765 120.600 114.355 120.645 ;
        RECT 116.465 120.600 116.755 120.645 ;
        RECT 110.465 120.460 116.755 120.600 ;
        RECT 110.465 120.415 111.115 120.460 ;
        RECT 114.065 120.415 114.355 120.460 ;
        RECT 116.465 120.415 116.755 120.460 ;
        RECT 113.230 120.260 113.550 120.320 ;
        RECT 117.000 120.260 117.140 120.755 ;
        RECT 105.500 120.120 117.140 120.260 ;
        RECT 75.050 120.060 75.370 120.120 ;
        RECT 101.730 120.060 102.050 120.120 ;
        RECT 104.965 120.075 105.255 120.120 ;
        RECT 113.230 120.060 113.550 120.120 ;
        RECT 5.520 119.440 123.740 119.920 ;
        RECT 29.970 119.040 30.290 119.300 ;
        RECT 36.410 119.240 36.730 119.300 ;
        RECT 41.485 119.240 41.775 119.285 ;
        RECT 36.410 119.100 41.775 119.240 ;
        RECT 36.410 119.040 36.730 119.100 ;
        RECT 41.485 119.055 41.775 119.100 ;
        RECT 64.485 119.240 64.775 119.285 ;
        RECT 67.690 119.240 68.010 119.300 ;
        RECT 64.485 119.100 68.010 119.240 ;
        RECT 64.485 119.055 64.775 119.100 ;
        RECT 67.690 119.040 68.010 119.100 ;
        RECT 75.970 119.240 76.290 119.300 ;
        RECT 79.205 119.240 79.495 119.285 ;
        RECT 75.970 119.100 79.495 119.240 ;
        RECT 75.970 119.040 76.290 119.100 ;
        RECT 79.205 119.055 79.495 119.100 ;
        RECT 92.085 119.240 92.375 119.285 ;
        RECT 93.450 119.240 93.770 119.300 ;
        RECT 92.085 119.100 93.770 119.240 ;
        RECT 92.085 119.055 92.375 119.100 ;
        RECT 93.450 119.040 93.770 119.100 ;
        RECT 96.685 119.240 96.975 119.285 ;
        RECT 97.590 119.240 97.910 119.300 ;
        RECT 96.685 119.100 97.910 119.240 ;
        RECT 96.685 119.055 96.975 119.100 ;
        RECT 97.590 119.040 97.910 119.100 ;
        RECT 99.445 119.240 99.735 119.285 ;
        RECT 99.890 119.240 100.210 119.300 ;
        RECT 99.445 119.100 100.210 119.240 ;
        RECT 99.445 119.055 99.735 119.100 ;
        RECT 99.890 119.040 100.210 119.100 ;
        RECT 103.110 119.040 103.430 119.300 ;
        RECT 106.790 119.040 107.110 119.300 ;
        RECT 108.185 119.240 108.475 119.285 ;
        RECT 113.690 119.240 114.010 119.300 ;
        RECT 108.185 119.100 114.010 119.240 ;
        RECT 108.185 119.055 108.475 119.100 ;
        RECT 113.690 119.040 114.010 119.100 ;
        RECT 117.830 119.040 118.150 119.300 ;
        RECT 9.385 118.900 9.675 118.945 ;
        RECT 12.625 118.900 13.275 118.945 ;
        RECT 17.565 118.900 17.855 118.945 ;
        RECT 9.385 118.760 17.855 118.900 ;
        RECT 9.385 118.715 9.975 118.760 ;
        RECT 12.625 118.715 13.275 118.760 ;
        RECT 17.565 118.715 17.855 118.760 ;
        RECT 22.265 118.900 22.555 118.945 ;
        RECT 25.505 118.900 26.155 118.945 ;
        RECT 26.750 118.900 27.070 118.960 ;
        RECT 35.490 118.945 35.810 118.960 ;
        RECT 22.265 118.760 27.070 118.900 ;
        RECT 22.265 118.715 22.855 118.760 ;
        RECT 25.505 118.715 26.155 118.760 ;
        RECT 9.685 118.400 9.975 118.715 ;
        RECT 10.765 118.560 11.055 118.605 ;
        RECT 14.345 118.560 14.635 118.605 ;
        RECT 16.180 118.560 16.470 118.605 ;
        RECT 10.765 118.420 16.470 118.560 ;
        RECT 10.765 118.375 11.055 118.420 ;
        RECT 14.345 118.375 14.635 118.420 ;
        RECT 16.180 118.375 16.470 118.420 ;
        RECT 16.645 118.375 16.935 118.605 ;
        RECT 3.290 118.220 3.610 118.280 ;
        RECT 7.905 118.220 8.195 118.265 ;
        RECT 3.290 118.080 8.195 118.220 ;
        RECT 3.290 118.020 3.610 118.080 ;
        RECT 7.905 118.035 8.195 118.080 ;
        RECT 15.250 118.020 15.570 118.280 ;
        RECT 10.765 117.880 11.055 117.925 ;
        RECT 13.885 117.880 14.175 117.925 ;
        RECT 15.775 117.880 16.065 117.925 ;
        RECT 10.765 117.740 16.065 117.880 ;
        RECT 10.765 117.695 11.055 117.740 ;
        RECT 13.885 117.695 14.175 117.740 ;
        RECT 15.775 117.695 16.065 117.740 ;
        RECT 7.890 117.540 8.210 117.600 ;
        RECT 16.720 117.540 16.860 118.375 ;
        RECT 18.010 118.360 18.330 118.620 ;
        RECT 19.390 118.560 19.710 118.620 ;
        RECT 20.325 118.560 20.615 118.605 ;
        RECT 19.390 118.420 20.615 118.560 ;
        RECT 19.390 118.360 19.710 118.420 ;
        RECT 20.325 118.375 20.615 118.420 ;
        RECT 22.565 118.400 22.855 118.715 ;
        RECT 26.750 118.700 27.070 118.760 ;
        RECT 35.485 118.900 36.135 118.945 ;
        RECT 39.085 118.900 39.375 118.945 ;
        RECT 35.485 118.760 39.375 118.900 ;
        RECT 35.485 118.715 36.135 118.760 ;
        RECT 38.785 118.715 39.375 118.760 ;
        RECT 35.490 118.700 35.810 118.715 ;
        RECT 23.645 118.560 23.935 118.605 ;
        RECT 27.225 118.560 27.515 118.605 ;
        RECT 29.060 118.560 29.350 118.605 ;
        RECT 23.645 118.420 29.350 118.560 ;
        RECT 23.645 118.375 23.935 118.420 ;
        RECT 27.225 118.375 27.515 118.420 ;
        RECT 29.060 118.375 29.350 118.420 ;
        RECT 29.525 118.375 29.815 118.605 ;
        RECT 20.785 118.220 21.075 118.265 ;
        RECT 21.230 118.220 21.550 118.280 ;
        RECT 20.785 118.080 21.550 118.220 ;
        RECT 20.785 118.035 21.075 118.080 ;
        RECT 21.230 118.020 21.550 118.080 ;
        RECT 28.130 118.020 28.450 118.280 ;
        RECT 29.600 118.220 29.740 118.375 ;
        RECT 30.890 118.360 31.210 118.620 ;
        RECT 32.290 118.560 32.580 118.605 ;
        RECT 34.125 118.560 34.415 118.605 ;
        RECT 37.705 118.560 37.995 118.605 ;
        RECT 32.290 118.420 37.995 118.560 ;
        RECT 32.290 118.375 32.580 118.420 ;
        RECT 34.125 118.375 34.415 118.420 ;
        RECT 37.705 118.375 37.995 118.420 ;
        RECT 38.785 118.400 39.075 118.715 ;
        RECT 49.750 118.700 50.070 118.960 ;
        RECT 65.965 118.900 66.255 118.945 ;
        RECT 69.205 118.900 69.855 118.945 ;
        RECT 71.830 118.900 72.150 118.960 ;
        RECT 65.965 118.760 72.150 118.900 ;
        RECT 65.965 118.715 66.555 118.760 ;
        RECT 69.205 118.715 69.855 118.760 ;
        RECT 42.405 118.560 42.695 118.605 ;
        RECT 46.530 118.560 46.850 118.620 ;
        RECT 42.405 118.420 46.850 118.560 ;
        RECT 42.405 118.375 42.695 118.420 ;
        RECT 46.530 118.360 46.850 118.420 ;
        RECT 51.145 118.375 51.435 118.605 ;
        RECT 52.050 118.560 52.370 118.620 ;
        RECT 58.965 118.560 59.255 118.605 ;
        RECT 52.050 118.420 59.255 118.560 ;
        RECT 31.825 118.220 32.115 118.265 ;
        RECT 29.600 118.080 32.115 118.220 ;
        RECT 19.405 117.880 19.695 117.925 ;
        RECT 19.850 117.880 20.170 117.940 ;
        RECT 19.405 117.740 20.170 117.880 ;
        RECT 19.405 117.695 19.695 117.740 ;
        RECT 19.850 117.680 20.170 117.740 ;
        RECT 23.645 117.880 23.935 117.925 ;
        RECT 26.765 117.880 27.055 117.925 ;
        RECT 28.655 117.880 28.945 117.925 ;
        RECT 23.645 117.740 28.945 117.880 ;
        RECT 23.645 117.695 23.935 117.740 ;
        RECT 26.765 117.695 27.055 117.740 ;
        RECT 28.655 117.695 28.945 117.740 ;
        RECT 20.310 117.540 20.630 117.600 ;
        RECT 29.600 117.540 29.740 118.080 ;
        RECT 31.825 118.035 32.115 118.080 ;
        RECT 33.190 118.020 33.510 118.280 ;
        RECT 35.950 118.220 36.270 118.280 ;
        RECT 40.565 118.220 40.855 118.265 ;
        RECT 35.950 118.080 40.855 118.220 ;
        RECT 35.950 118.020 36.270 118.080 ;
        RECT 40.565 118.035 40.855 118.080 ;
        RECT 32.695 117.880 32.985 117.925 ;
        RECT 34.585 117.880 34.875 117.925 ;
        RECT 37.705 117.880 37.995 117.925 ;
        RECT 32.695 117.740 37.995 117.880 ;
        RECT 51.220 117.880 51.360 118.375 ;
        RECT 52.050 118.360 52.370 118.420 ;
        RECT 58.965 118.375 59.255 118.420 ;
        RECT 66.265 118.400 66.555 118.715 ;
        RECT 71.830 118.700 72.150 118.760 ;
        RECT 75.050 118.700 75.370 118.960 ;
        RECT 92.530 118.900 92.850 118.960 ;
        RECT 112.765 118.900 113.415 118.945 ;
        RECT 114.150 118.900 114.470 118.960 ;
        RECT 116.365 118.900 116.655 118.945 ;
        RECT 92.530 118.760 99.200 118.900 ;
        RECT 92.530 118.700 92.850 118.760 ;
        RECT 67.345 118.560 67.635 118.605 ;
        RECT 70.925 118.560 71.215 118.605 ;
        RECT 72.760 118.560 73.050 118.605 ;
        RECT 67.345 118.420 73.050 118.560 ;
        RECT 67.345 118.375 67.635 118.420 ;
        RECT 70.925 118.375 71.215 118.420 ;
        RECT 72.760 118.375 73.050 118.420 ;
        RECT 73.670 118.360 73.990 118.620 ;
        RECT 80.125 118.560 80.415 118.605 ;
        RECT 90.690 118.560 91.010 118.620 ;
        RECT 80.125 118.420 91.010 118.560 ;
        RECT 80.125 118.375 80.415 118.420 ;
        RECT 90.690 118.360 91.010 118.420 ;
        RECT 91.150 118.360 91.470 118.620 ;
        RECT 95.765 118.560 96.055 118.605 ;
        RECT 98.510 118.560 98.830 118.620 ;
        RECT 99.060 118.605 99.200 118.760 ;
        RECT 112.765 118.760 116.655 118.900 ;
        RECT 112.765 118.715 113.415 118.760 ;
        RECT 114.150 118.700 114.470 118.760 ;
        RECT 116.065 118.715 116.655 118.760 ;
        RECT 95.765 118.420 98.830 118.560 ;
        RECT 95.765 118.375 96.055 118.420 ;
        RECT 98.510 118.360 98.830 118.420 ;
        RECT 98.985 118.375 99.275 118.605 ;
        RECT 102.205 118.560 102.495 118.605 ;
        RECT 103.110 118.560 103.430 118.620 ;
        RECT 102.205 118.420 103.430 118.560 ;
        RECT 102.205 118.375 102.495 118.420 ;
        RECT 103.110 118.360 103.430 118.420 ;
        RECT 105.870 118.360 106.190 118.620 ;
        RECT 107.265 118.375 107.555 118.605 ;
        RECT 109.570 118.560 109.860 118.605 ;
        RECT 111.405 118.560 111.695 118.605 ;
        RECT 114.985 118.560 115.275 118.605 ;
        RECT 109.570 118.420 115.275 118.560 ;
        RECT 109.570 118.375 109.860 118.420 ;
        RECT 111.405 118.375 111.695 118.420 ;
        RECT 114.985 118.375 115.275 118.420 ;
        RECT 116.065 118.400 116.355 118.715 ;
        RECT 71.830 118.020 72.150 118.280 ;
        RECT 73.225 118.220 73.515 118.265 ;
        RECT 75.510 118.220 75.830 118.280 ;
        RECT 73.225 118.080 75.830 118.220 ;
        RECT 73.225 118.035 73.515 118.080 ;
        RECT 75.510 118.020 75.830 118.080 ;
        RECT 104.490 118.220 104.810 118.280 ;
        RECT 107.340 118.220 107.480 118.375 ;
        RECT 104.490 118.080 107.480 118.220 ;
        RECT 104.490 118.020 104.810 118.080 ;
        RECT 109.090 118.020 109.410 118.280 ;
        RECT 110.470 118.020 110.790 118.280 ;
        RECT 67.345 117.880 67.635 117.925 ;
        RECT 70.465 117.880 70.755 117.925 ;
        RECT 72.355 117.880 72.645 117.925 ;
        RECT 51.220 117.740 67.000 117.880 ;
        RECT 32.695 117.695 32.985 117.740 ;
        RECT 34.585 117.695 34.875 117.740 ;
        RECT 37.705 117.695 37.995 117.740 ;
        RECT 7.890 117.400 29.740 117.540 ;
        RECT 59.425 117.540 59.715 117.585 ;
        RECT 66.310 117.540 66.630 117.600 ;
        RECT 59.425 117.400 66.630 117.540 ;
        RECT 66.860 117.540 67.000 117.740 ;
        RECT 67.345 117.740 72.645 117.880 ;
        RECT 67.345 117.695 67.635 117.740 ;
        RECT 70.465 117.695 70.755 117.740 ;
        RECT 72.355 117.695 72.645 117.740 ;
        RECT 109.975 117.880 110.265 117.925 ;
        RECT 111.865 117.880 112.155 117.925 ;
        RECT 114.985 117.880 115.275 117.925 ;
        RECT 109.975 117.740 115.275 117.880 ;
        RECT 109.975 117.695 110.265 117.740 ;
        RECT 111.865 117.695 112.155 117.740 ;
        RECT 114.985 117.695 115.275 117.740 ;
        RECT 73.670 117.540 73.990 117.600 ;
        RECT 66.860 117.400 73.990 117.540 ;
        RECT 7.890 117.340 8.210 117.400 ;
        RECT 20.310 117.340 20.630 117.400 ;
        RECT 59.425 117.355 59.715 117.400 ;
        RECT 66.310 117.340 66.630 117.400 ;
        RECT 73.670 117.340 73.990 117.400 ;
        RECT 5.520 116.720 123.740 117.200 ;
        RECT 8.350 116.520 8.670 116.580 ;
        RECT 10.205 116.520 10.495 116.565 ;
        RECT 8.350 116.380 10.495 116.520 ;
        RECT 8.350 116.320 8.670 116.380 ;
        RECT 10.205 116.335 10.495 116.380 ;
        RECT 11.585 116.520 11.875 116.565 ;
        RECT 15.250 116.520 15.570 116.580 ;
        RECT 11.585 116.380 15.570 116.520 ;
        RECT 11.585 116.335 11.875 116.380 ;
        RECT 15.250 116.320 15.570 116.380 ;
        RECT 24.005 116.520 24.295 116.565 ;
        RECT 28.130 116.520 28.450 116.580 ;
        RECT 24.005 116.380 28.450 116.520 ;
        RECT 24.005 116.335 24.295 116.380 ;
        RECT 28.130 116.320 28.450 116.380 ;
        RECT 33.190 116.520 33.510 116.580 ;
        RECT 33.665 116.520 33.955 116.565 ;
        RECT 33.190 116.380 33.955 116.520 ;
        RECT 33.190 116.320 33.510 116.380 ;
        RECT 33.665 116.335 33.955 116.380 ;
        RECT 68.625 116.520 68.915 116.565 ;
        RECT 71.830 116.520 72.150 116.580 ;
        RECT 68.625 116.380 72.150 116.520 ;
        RECT 68.625 116.335 68.915 116.380 ;
        RECT 71.830 116.320 72.150 116.380 ;
        RECT 114.150 116.320 114.470 116.580 ;
        RECT 69.070 116.180 69.390 116.240 ;
        RECT 71.385 116.180 71.675 116.225 ;
        RECT 69.070 116.040 71.675 116.180 ;
        RECT 69.070 115.980 69.390 116.040 ;
        RECT 71.385 115.995 71.675 116.040 ;
        RECT 76.450 116.180 76.740 116.225 ;
        RECT 78.310 116.180 78.600 116.225 ;
        RECT 81.090 116.180 81.380 116.225 ;
        RECT 76.450 116.040 81.380 116.180 ;
        RECT 76.450 115.995 76.740 116.040 ;
        RECT 78.310 115.995 78.600 116.040 ;
        RECT 81.090 115.995 81.380 116.040 ;
        RECT 11.125 115.500 11.415 115.545 ;
        RECT 12.030 115.500 12.350 115.560 ;
        RECT 11.125 115.360 12.350 115.500 ;
        RECT 11.125 115.315 11.415 115.360 ;
        RECT 12.030 115.300 12.350 115.360 ;
        RECT 12.490 115.300 12.810 115.560 ;
        RECT 24.925 115.500 25.215 115.545 ;
        RECT 26.750 115.500 27.070 115.560 ;
        RECT 24.925 115.360 27.070 115.500 ;
        RECT 24.925 115.315 25.215 115.360 ;
        RECT 26.750 115.300 27.070 115.360 ;
        RECT 34.585 115.500 34.875 115.545 ;
        RECT 36.410 115.500 36.730 115.560 ;
        RECT 34.585 115.360 36.730 115.500 ;
        RECT 34.585 115.315 34.875 115.360 ;
        RECT 36.410 115.300 36.730 115.360 ;
        RECT 69.545 115.315 69.835 115.545 ;
        RECT 69.620 114.820 69.760 115.315 ;
        RECT 72.290 115.300 72.610 115.560 ;
        RECT 75.510 115.500 75.830 115.560 ;
        RECT 75.985 115.500 76.275 115.545 ;
        RECT 75.510 115.360 76.275 115.500 ;
        RECT 75.510 115.300 75.830 115.360 ;
        RECT 75.985 115.315 76.275 115.360 ;
        RECT 77.810 115.300 78.130 115.560 ;
        RECT 81.090 115.500 81.380 115.545 ;
        RECT 78.845 115.360 81.380 115.500 ;
        RECT 78.845 115.205 79.060 115.360 ;
        RECT 81.090 115.315 81.380 115.360 ;
        RECT 113.230 115.500 113.550 115.560 ;
        RECT 113.705 115.500 113.995 115.545 ;
        RECT 113.230 115.360 113.995 115.500 ;
        RECT 113.230 115.300 113.550 115.360 ;
        RECT 113.705 115.315 113.995 115.360 ;
        RECT 76.910 115.160 77.200 115.205 ;
        RECT 78.770 115.160 79.060 115.205 ;
        RECT 76.910 115.020 79.060 115.160 ;
        RECT 76.910 114.975 77.200 115.020 ;
        RECT 78.770 114.975 79.060 115.020 ;
        RECT 79.690 115.160 79.980 115.205 ;
        RECT 80.570 115.160 80.890 115.220 ;
        RECT 82.950 115.160 83.240 115.205 ;
        RECT 92.990 115.160 93.310 115.220 ;
        RECT 79.690 115.020 83.240 115.160 ;
        RECT 79.690 114.975 79.980 115.020 ;
        RECT 80.570 114.960 80.890 115.020 ;
        RECT 82.950 114.975 83.240 115.020 ;
        RECT 83.420 115.020 93.310 115.160 ;
        RECT 83.420 114.820 83.560 115.020 ;
        RECT 92.990 114.960 93.310 115.020 ;
        RECT 69.620 114.680 83.560 114.820 ;
        RECT 83.790 114.820 84.110 114.880 ;
        RECT 84.955 114.820 85.245 114.865 ;
        RECT 83.790 114.680 85.245 114.820 ;
        RECT 83.790 114.620 84.110 114.680 ;
        RECT 84.955 114.635 85.245 114.680 ;
        RECT 5.520 114.000 123.740 114.480 ;
        RECT 77.810 113.600 78.130 113.860 ;
        RECT 80.570 113.800 80.890 113.860 ;
        RECT 81.045 113.800 81.335 113.845 ;
        RECT 80.570 113.660 81.335 113.800 ;
        RECT 80.570 113.600 80.890 113.660 ;
        RECT 81.045 113.615 81.335 113.660 ;
        RECT 83.790 113.800 84.110 113.860 ;
        RECT 85.185 113.800 85.475 113.845 ;
        RECT 92.070 113.800 92.390 113.860 ;
        RECT 83.790 113.660 92.390 113.800 ;
        RECT 83.790 113.600 84.110 113.660 ;
        RECT 85.185 113.615 85.475 113.660 ;
        RECT 92.070 113.600 92.390 113.660 ;
        RECT 93.465 113.800 93.755 113.845 ;
        RECT 101.730 113.800 102.050 113.860 ;
        RECT 93.465 113.660 102.050 113.800 ;
        RECT 93.465 113.615 93.755 113.660 ;
        RECT 101.730 113.600 102.050 113.660 ;
        RECT 105.885 113.800 106.175 113.845 ;
        RECT 110.470 113.800 110.790 113.860 ;
        RECT 105.885 113.660 110.790 113.800 ;
        RECT 105.885 113.615 106.175 113.660 ;
        RECT 110.470 113.600 110.790 113.660 ;
        RECT 11.590 113.460 11.880 113.505 ;
        RECT 13.450 113.460 13.740 113.505 ;
        RECT 11.590 113.320 13.740 113.460 ;
        RECT 11.590 113.275 11.880 113.320 ;
        RECT 13.450 113.275 13.740 113.320 ;
        RECT 14.370 113.460 14.660 113.505 ;
        RECT 16.170 113.460 16.490 113.520 ;
        RECT 17.630 113.460 17.920 113.505 ;
        RECT 14.370 113.320 17.920 113.460 ;
        RECT 14.370 113.275 14.660 113.320 ;
        RECT 13.525 113.120 13.740 113.275 ;
        RECT 16.170 113.260 16.490 113.320 ;
        RECT 17.630 113.275 17.920 113.320 ;
        RECT 27.670 113.460 27.990 113.520 ;
        RECT 40.570 113.460 40.860 113.505 ;
        RECT 42.430 113.460 42.720 113.505 ;
        RECT 27.670 113.320 32.960 113.460 ;
        RECT 27.670 113.260 27.990 113.320 ;
        RECT 32.820 113.165 32.960 113.320 ;
        RECT 40.570 113.320 42.720 113.460 ;
        RECT 40.570 113.275 40.860 113.320 ;
        RECT 42.430 113.275 42.720 113.320 ;
        RECT 43.350 113.460 43.640 113.505 ;
        RECT 45.150 113.460 45.470 113.520 ;
        RECT 46.610 113.460 46.900 113.505 ;
        RECT 43.350 113.320 46.900 113.460 ;
        RECT 43.350 113.275 43.640 113.320 ;
        RECT 15.770 113.120 16.060 113.165 ;
        RECT 13.525 112.980 16.060 113.120 ;
        RECT 15.770 112.935 16.060 112.980 ;
        RECT 30.445 112.935 30.735 113.165 ;
        RECT 32.745 112.935 33.035 113.165 ;
        RECT 41.485 113.120 41.775 113.165 ;
        RECT 41.930 113.120 42.250 113.180 ;
        RECT 41.485 112.980 42.250 113.120 ;
        RECT 42.505 113.120 42.720 113.275 ;
        RECT 45.150 113.260 45.470 113.320 ;
        RECT 46.610 113.275 46.900 113.320 ;
        RECT 58.950 113.460 59.270 113.520 ;
        RECT 59.820 113.460 60.110 113.505 ;
        RECT 63.080 113.460 63.370 113.505 ;
        RECT 58.950 113.320 63.370 113.460 ;
        RECT 58.950 113.260 59.270 113.320 ;
        RECT 59.820 113.275 60.110 113.320 ;
        RECT 63.080 113.275 63.370 113.320 ;
        RECT 64.000 113.460 64.290 113.505 ;
        RECT 65.860 113.460 66.150 113.505 ;
        RECT 86.550 113.460 86.870 113.520 ;
        RECT 102.190 113.505 102.510 113.520 ;
        RECT 96.230 113.460 96.520 113.505 ;
        RECT 98.090 113.460 98.380 113.505 ;
        RECT 64.000 113.320 66.150 113.460 ;
        RECT 64.000 113.275 64.290 113.320 ;
        RECT 65.860 113.275 66.150 113.320 ;
        RECT 82.730 113.320 94.140 113.460 ;
        RECT 44.750 113.120 45.040 113.165 ;
        RECT 42.505 112.980 45.040 113.120 ;
        RECT 41.485 112.935 41.775 112.980 ;
        RECT 7.890 112.780 8.210 112.840 ;
        RECT 10.665 112.780 10.955 112.825 ;
        RECT 7.890 112.640 10.955 112.780 ;
        RECT 7.890 112.580 8.210 112.640 ;
        RECT 10.665 112.595 10.955 112.640 ;
        RECT 12.505 112.780 12.795 112.825 ;
        RECT 14.330 112.780 14.650 112.840 ;
        RECT 12.505 112.640 14.650 112.780 ;
        RECT 30.520 112.780 30.660 112.935 ;
        RECT 41.930 112.920 42.250 112.980 ;
        RECT 44.750 112.935 45.040 112.980 ;
        RECT 61.680 113.120 61.970 113.165 ;
        RECT 64.000 113.120 64.215 113.275 ;
        RECT 61.680 112.980 64.215 113.120 ;
        RECT 61.680 112.935 61.970 112.980 ;
        RECT 78.745 112.935 79.035 113.165 ;
        RECT 80.585 113.120 80.875 113.165 ;
        RECT 82.730 113.120 82.870 113.320 ;
        RECT 86.550 113.260 86.870 113.320 ;
        RECT 80.585 112.980 82.870 113.120 ;
        RECT 87.010 113.120 87.330 113.180 ;
        RECT 89.860 113.165 90.000 113.320 ;
        RECT 88.405 113.120 88.695 113.165 ;
        RECT 87.010 112.980 88.695 113.120 ;
        RECT 80.585 112.935 80.875 112.980 ;
        RECT 35.950 112.780 36.270 112.840 ;
        RECT 30.520 112.640 36.270 112.780 ;
        RECT 12.505 112.595 12.795 112.640 ;
        RECT 14.330 112.580 14.650 112.640 ;
        RECT 35.950 112.580 36.270 112.640 ;
        RECT 39.170 112.780 39.490 112.840 ;
        RECT 39.645 112.780 39.935 112.825 ;
        RECT 39.170 112.640 39.935 112.780 ;
        RECT 39.170 112.580 39.490 112.640 ;
        RECT 39.645 112.595 39.935 112.640 ;
        RECT 55.270 112.780 55.590 112.840 ;
        RECT 64.945 112.780 65.235 112.825 ;
        RECT 55.270 112.640 65.235 112.780 ;
        RECT 55.270 112.580 55.590 112.640 ;
        RECT 64.945 112.595 65.235 112.640 ;
        RECT 66.785 112.780 67.075 112.825 ;
        RECT 75.510 112.780 75.830 112.840 ;
        RECT 66.785 112.640 75.830 112.780 ;
        RECT 66.785 112.595 67.075 112.640 ;
        RECT 75.510 112.580 75.830 112.640 ;
        RECT 11.130 112.440 11.420 112.485 ;
        RECT 12.990 112.440 13.280 112.485 ;
        RECT 15.770 112.440 16.060 112.485 ;
        RECT 11.130 112.300 16.060 112.440 ;
        RECT 11.130 112.255 11.420 112.300 ;
        RECT 12.990 112.255 13.280 112.300 ;
        RECT 15.770 112.255 16.060 112.300 ;
        RECT 40.110 112.440 40.400 112.485 ;
        RECT 41.970 112.440 42.260 112.485 ;
        RECT 44.750 112.440 45.040 112.485 ;
        RECT 40.110 112.300 45.040 112.440 ;
        RECT 40.110 112.255 40.400 112.300 ;
        RECT 41.970 112.255 42.260 112.300 ;
        RECT 44.750 112.255 45.040 112.300 ;
        RECT 61.680 112.440 61.970 112.485 ;
        RECT 64.460 112.440 64.750 112.485 ;
        RECT 66.320 112.440 66.610 112.485 ;
        RECT 61.680 112.300 66.610 112.440 ;
        RECT 78.820 112.440 78.960 112.935 ;
        RECT 87.010 112.920 87.330 112.980 ;
        RECT 88.405 112.935 88.695 112.980 ;
        RECT 89.785 112.935 90.075 113.165 ;
        RECT 92.530 112.920 92.850 113.180 ;
        RECT 94.000 113.165 94.140 113.320 ;
        RECT 96.230 113.320 98.380 113.460 ;
        RECT 96.230 113.275 96.520 113.320 ;
        RECT 98.090 113.275 98.380 113.320 ;
        RECT 99.010 113.460 99.300 113.505 ;
        RECT 102.190 113.460 102.560 113.505 ;
        RECT 99.010 113.320 102.560 113.460 ;
        RECT 99.010 113.275 99.300 113.320 ;
        RECT 102.190 113.275 102.560 113.320 ;
        RECT 93.925 112.935 94.215 113.165 ;
        RECT 98.165 113.120 98.380 113.275 ;
        RECT 102.190 113.260 102.510 113.275 ;
        RECT 100.410 113.120 100.700 113.165 ;
        RECT 98.165 112.980 100.700 113.120 ;
        RECT 100.410 112.935 100.700 112.980 ;
        RECT 104.950 112.920 105.270 113.180 ;
        RECT 85.630 112.580 85.950 112.840 ;
        RECT 86.565 112.780 86.855 112.825 ;
        RECT 87.930 112.780 88.250 112.840 ;
        RECT 86.565 112.640 88.250 112.780 ;
        RECT 86.565 112.595 86.855 112.640 ;
        RECT 87.930 112.580 88.250 112.640 ;
        RECT 95.305 112.780 95.595 112.825 ;
        RECT 96.210 112.780 96.530 112.840 ;
        RECT 95.305 112.640 96.530 112.780 ;
        RECT 95.305 112.595 95.595 112.640 ;
        RECT 96.210 112.580 96.530 112.640 ;
        RECT 97.130 112.580 97.450 112.840 ;
        RECT 83.345 112.440 83.635 112.485 ;
        RECT 78.820 112.300 83.635 112.440 ;
        RECT 61.680 112.255 61.970 112.300 ;
        RECT 64.460 112.255 64.750 112.300 ;
        RECT 66.320 112.255 66.610 112.300 ;
        RECT 83.345 112.255 83.635 112.300 ;
        RECT 95.770 112.440 96.060 112.485 ;
        RECT 97.630 112.440 97.920 112.485 ;
        RECT 100.410 112.440 100.700 112.485 ;
        RECT 95.770 112.300 100.700 112.440 ;
        RECT 95.770 112.255 96.060 112.300 ;
        RECT 97.630 112.255 97.920 112.300 ;
        RECT 100.410 112.255 100.700 112.300 ;
        RECT 19.635 112.100 19.925 112.145 ;
        RECT 20.770 112.100 21.090 112.160 ;
        RECT 19.635 111.960 21.090 112.100 ;
        RECT 19.635 111.915 19.925 111.960 ;
        RECT 20.770 111.900 21.090 111.960 ;
        RECT 29.510 111.900 29.830 112.160 ;
        RECT 32.270 111.900 32.590 112.160 ;
        RECT 48.615 112.100 48.905 112.145 ;
        RECT 49.750 112.100 50.070 112.160 ;
        RECT 48.615 111.960 50.070 112.100 ;
        RECT 48.615 111.915 48.905 111.960 ;
        RECT 49.750 111.900 50.070 111.960 ;
        RECT 55.730 112.100 56.050 112.160 ;
        RECT 57.815 112.100 58.105 112.145 ;
        RECT 61.250 112.100 61.570 112.160 ;
        RECT 55.730 111.960 61.570 112.100 ;
        RECT 55.730 111.900 56.050 111.960 ;
        RECT 57.815 111.915 58.105 111.960 ;
        RECT 61.250 111.900 61.570 111.960 ;
        RECT 82.870 112.100 83.190 112.160 ;
        RECT 87.485 112.100 87.775 112.145 ;
        RECT 82.870 111.960 87.775 112.100 ;
        RECT 82.870 111.900 83.190 111.960 ;
        RECT 87.485 111.915 87.775 111.960 ;
        RECT 89.310 111.900 89.630 112.160 ;
        RECT 94.385 112.100 94.675 112.145 ;
        RECT 96.670 112.100 96.990 112.160 ;
        RECT 94.385 111.960 96.990 112.100 ;
        RECT 94.385 111.915 94.675 111.960 ;
        RECT 96.670 111.900 96.990 111.960 ;
        RECT 104.030 112.145 104.350 112.160 ;
        RECT 104.030 111.915 104.565 112.145 ;
        RECT 104.030 111.900 104.350 111.915 ;
        RECT 5.520 111.280 123.740 111.760 ;
        RECT 14.330 110.880 14.650 111.140 ;
        RECT 41.485 111.080 41.775 111.125 ;
        RECT 41.930 111.080 42.250 111.140 ;
        RECT 41.485 110.940 42.250 111.080 ;
        RECT 41.485 110.895 41.775 110.940 ;
        RECT 41.930 110.880 42.250 110.940 ;
        RECT 53.445 111.080 53.735 111.125 ;
        RECT 55.270 111.080 55.590 111.140 ;
        RECT 53.445 110.940 55.590 111.080 ;
        RECT 53.445 110.895 53.735 110.940 ;
        RECT 55.270 110.880 55.590 110.940 ;
        RECT 82.885 111.080 83.175 111.125 ;
        RECT 83.330 111.080 83.650 111.140 ;
        RECT 82.885 110.940 83.650 111.080 ;
        RECT 82.885 110.895 83.175 110.940 ;
        RECT 83.330 110.880 83.650 110.940 ;
        RECT 92.530 111.080 92.850 111.140 ;
        RECT 94.385 111.080 94.675 111.125 ;
        RECT 92.530 110.940 94.675 111.080 ;
        RECT 92.530 110.880 92.850 110.940 ;
        RECT 94.385 110.895 94.675 110.940 ;
        RECT 97.130 111.080 97.450 111.140 ;
        RECT 100.365 111.080 100.655 111.125 ;
        RECT 97.130 110.940 100.655 111.080 ;
        RECT 97.130 110.880 97.450 110.940 ;
        RECT 100.365 110.895 100.655 110.940 ;
        RECT 26.770 110.740 27.060 110.785 ;
        RECT 28.630 110.740 28.920 110.785 ;
        RECT 31.410 110.740 31.700 110.785 ;
        RECT 26.770 110.600 31.700 110.740 ;
        RECT 26.770 110.555 27.060 110.600 ;
        RECT 28.630 110.555 28.920 110.600 ;
        RECT 31.410 110.555 31.700 110.600 ;
        RECT 59.890 110.740 60.180 110.785 ;
        RECT 61.750 110.740 62.040 110.785 ;
        RECT 64.530 110.740 64.820 110.785 ;
        RECT 59.890 110.600 64.820 110.740 ;
        RECT 59.890 110.555 60.180 110.600 ;
        RECT 61.750 110.555 62.040 110.600 ;
        RECT 64.530 110.555 64.820 110.600 ;
        RECT 71.390 110.740 71.680 110.785 ;
        RECT 73.250 110.740 73.540 110.785 ;
        RECT 76.030 110.740 76.320 110.785 ;
        RECT 71.390 110.600 76.320 110.740 ;
        RECT 71.390 110.555 71.680 110.600 ;
        RECT 73.250 110.555 73.540 110.600 ;
        RECT 76.030 110.555 76.320 110.600 ;
        RECT 87.930 110.740 88.250 110.800 ;
        RECT 108.190 110.740 108.480 110.785 ;
        RECT 110.050 110.740 110.340 110.785 ;
        RECT 112.830 110.740 113.120 110.785 ;
        RECT 87.930 110.600 107.940 110.740 ;
        RECT 87.930 110.540 88.250 110.600 ;
        RECT 16.170 110.200 16.490 110.460 ;
        RECT 22.150 110.200 22.470 110.460 ;
        RECT 27.670 110.400 27.990 110.460 ;
        RECT 25.000 110.260 27.990 110.400 ;
        RECT 15.265 109.875 15.555 110.105 ;
        RECT 16.630 110.060 16.950 110.120 ;
        RECT 25.000 110.105 25.140 110.260 ;
        RECT 27.670 110.200 27.990 110.260 ;
        RECT 28.145 110.400 28.435 110.445 ;
        RECT 29.510 110.400 29.830 110.460 ;
        RECT 28.145 110.260 29.830 110.400 ;
        RECT 28.145 110.215 28.435 110.260 ;
        RECT 29.510 110.200 29.830 110.260 ;
        RECT 45.150 110.200 45.470 110.460 ;
        RECT 50.670 110.400 50.990 110.460 ;
        RECT 56.205 110.400 56.495 110.445 ;
        RECT 45.700 110.260 50.440 110.400 ;
        RECT 24.925 110.060 25.215 110.105 ;
        RECT 26.305 110.070 26.595 110.105 ;
        RECT 25.920 110.060 26.595 110.070 ;
        RECT 31.410 110.060 31.700 110.105 ;
        RECT 16.630 109.920 25.215 110.060 ;
        RECT 15.340 109.380 15.480 109.875 ;
        RECT 16.630 109.860 16.950 109.920 ;
        RECT 24.925 109.875 25.215 109.920 ;
        RECT 25.460 109.930 26.595 110.060 ;
        RECT 25.460 109.920 26.060 109.930 ;
        RECT 20.310 109.720 20.630 109.780 ;
        RECT 25.460 109.720 25.600 109.920 ;
        RECT 26.305 109.875 26.595 109.930 ;
        RECT 29.165 109.920 31.700 110.060 ;
        RECT 29.165 109.765 29.380 109.920 ;
        RECT 31.410 109.875 31.700 109.920 ;
        RECT 42.390 109.860 42.710 110.120 ;
        RECT 45.700 110.105 45.840 110.260 ;
        RECT 45.625 109.875 45.915 110.105 ;
        RECT 49.290 109.860 49.610 110.120 ;
        RECT 50.300 110.105 50.440 110.260 ;
        RECT 50.670 110.260 56.495 110.400 ;
        RECT 50.670 110.200 50.990 110.260 ;
        RECT 56.205 110.215 56.495 110.260 ;
        RECT 57.110 110.200 57.430 110.460 ;
        RECT 70.925 110.400 71.215 110.445 ;
        RECT 75.510 110.400 75.830 110.460 ;
        RECT 70.925 110.260 75.830 110.400 ;
        RECT 70.925 110.215 71.215 110.260 ;
        RECT 75.510 110.200 75.830 110.260 ;
        RECT 79.650 110.445 79.970 110.460 ;
        RECT 79.650 110.400 80.185 110.445 ;
        RECT 85.630 110.400 85.950 110.460 ;
        RECT 91.700 110.445 91.840 110.600 ;
        RECT 97.220 110.445 97.360 110.600 ;
        RECT 79.650 110.260 85.950 110.400 ;
        RECT 79.650 110.215 80.185 110.260 ;
        RECT 79.650 110.200 79.970 110.215 ;
        RECT 85.630 110.200 85.950 110.260 ;
        RECT 91.625 110.400 91.915 110.445 ;
        RECT 97.145 110.400 97.435 110.445 ;
        RECT 98.050 110.400 98.370 110.460 ;
        RECT 91.625 110.260 92.025 110.400 ;
        RECT 97.145 110.260 97.545 110.400 ;
        RECT 98.050 110.260 101.960 110.400 ;
        RECT 91.625 110.215 91.915 110.260 ;
        RECT 97.145 110.215 97.435 110.260 ;
        RECT 98.050 110.200 98.370 110.260 ;
        RECT 50.225 110.060 50.515 110.105 ;
        RECT 51.590 110.060 51.910 110.120 ;
        RECT 50.225 109.920 51.910 110.060 ;
        RECT 50.225 109.875 50.515 109.920 ;
        RECT 51.590 109.860 51.910 109.920 ;
        RECT 52.525 109.875 52.815 110.105 ;
        RECT 20.310 109.580 25.600 109.720 ;
        RECT 27.230 109.720 27.520 109.765 ;
        RECT 29.090 109.720 29.380 109.765 ;
        RECT 27.230 109.580 29.380 109.720 ;
        RECT 20.310 109.520 20.630 109.580 ;
        RECT 27.230 109.535 27.520 109.580 ;
        RECT 29.090 109.535 29.380 109.580 ;
        RECT 30.010 109.720 30.300 109.765 ;
        RECT 32.270 109.720 32.590 109.780 ;
        RECT 33.270 109.720 33.560 109.765 ;
        RECT 30.010 109.580 33.560 109.720 ;
        RECT 30.010 109.535 30.300 109.580 ;
        RECT 32.270 109.520 32.590 109.580 ;
        RECT 33.270 109.535 33.560 109.580 ;
        RECT 18.945 109.380 19.235 109.425 ;
        RECT 15.340 109.240 19.235 109.380 ;
        RECT 18.945 109.195 19.235 109.240 ;
        RECT 20.770 109.180 21.090 109.440 ;
        RECT 21.230 109.180 21.550 109.440 ;
        RECT 23.990 109.380 24.310 109.440 ;
        RECT 25.385 109.380 25.675 109.425 ;
        RECT 23.990 109.240 25.675 109.380 ;
        RECT 23.990 109.180 24.310 109.240 ;
        RECT 25.385 109.195 25.675 109.240 ;
        RECT 27.670 109.380 27.990 109.440 ;
        RECT 35.275 109.380 35.565 109.425 ;
        RECT 27.670 109.240 35.565 109.380 ;
        RECT 27.670 109.180 27.990 109.240 ;
        RECT 35.275 109.195 35.565 109.240 ;
        RECT 47.450 109.380 47.770 109.440 ;
        RECT 48.385 109.380 48.675 109.425 ;
        RECT 47.450 109.240 48.675 109.380 ;
        RECT 47.450 109.180 47.770 109.240 ;
        RECT 48.385 109.195 48.675 109.240 ;
        RECT 50.210 109.380 50.530 109.440 ;
        RECT 50.685 109.380 50.975 109.425 ;
        RECT 50.210 109.240 50.975 109.380 ;
        RECT 52.600 109.380 52.740 109.875 ;
        RECT 55.730 109.860 56.050 110.120 ;
        RECT 58.030 109.860 58.350 110.120 ;
        RECT 59.425 109.875 59.715 110.105 ;
        RECT 61.265 110.060 61.555 110.105 ;
        RECT 64.530 110.060 64.820 110.105 ;
        RECT 59.960 109.920 61.555 110.060 ;
        RECT 56.650 109.720 56.970 109.780 ;
        RECT 59.500 109.720 59.640 109.875 ;
        RECT 56.650 109.580 59.640 109.720 ;
        RECT 56.650 109.520 56.970 109.580 ;
        RECT 53.905 109.380 54.195 109.425 ;
        RECT 52.600 109.240 54.195 109.380 ;
        RECT 50.210 109.180 50.530 109.240 ;
        RECT 50.685 109.195 50.975 109.240 ;
        RECT 53.905 109.195 54.195 109.240 ;
        RECT 58.965 109.380 59.255 109.425 ;
        RECT 59.960 109.380 60.100 109.920 ;
        RECT 61.265 109.875 61.555 109.920 ;
        RECT 62.285 109.920 64.820 110.060 ;
        RECT 62.285 109.765 62.500 109.920 ;
        RECT 64.530 109.875 64.820 109.920 ;
        RECT 72.750 109.860 73.070 110.120 ;
        RECT 76.030 110.060 76.320 110.105 ;
        RECT 73.785 109.920 76.320 110.060 ;
        RECT 60.350 109.720 60.640 109.765 ;
        RECT 62.210 109.720 62.500 109.765 ;
        RECT 60.350 109.580 62.500 109.720 ;
        RECT 60.350 109.535 60.640 109.580 ;
        RECT 62.210 109.535 62.500 109.580 ;
        RECT 63.130 109.720 63.420 109.765 ;
        RECT 64.930 109.720 65.250 109.780 ;
        RECT 73.785 109.765 74.000 109.920 ;
        RECT 76.030 109.875 76.320 109.920 ;
        RECT 101.285 109.875 101.575 110.105 ;
        RECT 66.390 109.720 66.680 109.765 ;
        RECT 63.130 109.580 66.680 109.720 ;
        RECT 63.130 109.535 63.420 109.580 ;
        RECT 64.930 109.520 65.250 109.580 ;
        RECT 66.390 109.535 66.680 109.580 ;
        RECT 71.850 109.720 72.140 109.765 ;
        RECT 73.710 109.720 74.000 109.765 ;
        RECT 71.850 109.580 74.000 109.720 ;
        RECT 71.850 109.535 72.140 109.580 ;
        RECT 73.710 109.535 74.000 109.580 ;
        RECT 74.630 109.720 74.920 109.765 ;
        RECT 76.430 109.720 76.750 109.780 ;
        RECT 77.890 109.720 78.180 109.765 ;
        RECT 74.630 109.580 78.180 109.720 ;
        RECT 74.630 109.535 74.920 109.580 ;
        RECT 76.430 109.520 76.750 109.580 ;
        RECT 77.890 109.535 78.180 109.580 ;
        RECT 90.230 109.520 90.550 109.780 ;
        RECT 58.965 109.240 60.100 109.380 ;
        RECT 61.710 109.380 62.030 109.440 ;
        RECT 68.395 109.380 68.685 109.425 ;
        RECT 61.710 109.240 68.685 109.380 ;
        RECT 58.965 109.195 59.255 109.240 ;
        RECT 61.710 109.180 62.030 109.240 ;
        RECT 68.395 109.195 68.685 109.240 ;
        RECT 92.070 109.180 92.390 109.440 ;
        RECT 92.545 109.380 92.835 109.425 ;
        RECT 93.450 109.380 93.770 109.440 ;
        RECT 97.605 109.380 97.895 109.425 ;
        RECT 92.545 109.240 97.895 109.380 ;
        RECT 92.545 109.195 92.835 109.240 ;
        RECT 93.450 109.180 93.770 109.240 ;
        RECT 97.605 109.195 97.895 109.240 ;
        RECT 98.050 109.180 98.370 109.440 ;
        RECT 99.905 109.380 100.195 109.425 ;
        RECT 101.360 109.380 101.500 109.875 ;
        RECT 101.820 109.720 101.960 110.260 ;
        RECT 102.190 110.200 102.510 110.460 ;
        RECT 104.580 110.445 104.720 110.600 ;
        RECT 104.505 110.400 104.795 110.445 ;
        RECT 107.800 110.400 107.940 110.600 ;
        RECT 108.190 110.600 113.120 110.740 ;
        RECT 108.190 110.555 108.480 110.600 ;
        RECT 110.050 110.555 110.340 110.600 ;
        RECT 112.830 110.555 113.120 110.600 ;
        RECT 113.230 110.400 113.550 110.460 ;
        RECT 104.505 110.260 104.905 110.400 ;
        RECT 107.800 110.260 113.550 110.400 ;
        RECT 104.505 110.215 104.795 110.260 ;
        RECT 113.230 110.200 113.550 110.260 ;
        RECT 102.650 109.860 102.970 110.120 ;
        RECT 107.725 110.060 108.015 110.105 ;
        RECT 109.090 110.060 109.410 110.120 ;
        RECT 107.725 109.920 109.410 110.060 ;
        RECT 107.725 109.875 108.015 109.920 ;
        RECT 109.090 109.860 109.410 109.920 ;
        RECT 109.550 109.860 109.870 110.120 ;
        RECT 112.830 110.060 113.120 110.105 ;
        RECT 110.585 109.920 113.120 110.060 ;
        RECT 104.030 109.720 104.350 109.780 ;
        RECT 110.585 109.765 110.800 109.920 ;
        RECT 112.830 109.875 113.120 109.920 ;
        RECT 117.370 109.860 117.690 110.120 ;
        RECT 104.965 109.720 105.255 109.765 ;
        RECT 108.650 109.720 108.940 109.765 ;
        RECT 110.510 109.720 110.800 109.765 ;
        RECT 101.820 109.580 105.255 109.720 ;
        RECT 104.030 109.520 104.350 109.580 ;
        RECT 104.965 109.535 105.255 109.580 ;
        RECT 105.500 109.580 107.940 109.720 ;
        RECT 105.500 109.440 105.640 109.580 ;
        RECT 99.905 109.240 101.500 109.380 ;
        RECT 99.905 109.195 100.195 109.240 ;
        RECT 105.410 109.180 105.730 109.440 ;
        RECT 107.250 109.180 107.570 109.440 ;
        RECT 107.800 109.380 107.940 109.580 ;
        RECT 108.650 109.580 110.800 109.720 ;
        RECT 108.650 109.535 108.940 109.580 ;
        RECT 110.510 109.535 110.800 109.580 ;
        RECT 111.430 109.720 111.720 109.765 ;
        RECT 114.690 109.720 114.980 109.765 ;
        RECT 117.845 109.720 118.135 109.765 ;
        RECT 111.430 109.580 118.135 109.720 ;
        RECT 111.430 109.535 111.720 109.580 ;
        RECT 114.690 109.535 114.980 109.580 ;
        RECT 117.845 109.535 118.135 109.580 ;
        RECT 116.695 109.380 116.985 109.425 ;
        RECT 107.800 109.240 116.985 109.380 ;
        RECT 116.695 109.195 116.985 109.240 ;
        RECT 5.520 108.560 123.740 109.040 ;
        RECT 19.865 108.175 20.155 108.405 ;
        RECT 18.930 107.480 19.250 107.740 ;
        RECT 19.940 107.680 20.080 108.175 ;
        RECT 58.950 108.160 59.270 108.420 ;
        RECT 59.885 108.175 60.175 108.405 ;
        RECT 23.990 108.065 24.310 108.080 ;
        RECT 21.250 108.020 21.540 108.065 ;
        RECT 23.110 108.020 23.400 108.065 ;
        RECT 21.250 107.880 23.400 108.020 ;
        RECT 21.250 107.835 21.540 107.880 ;
        RECT 23.110 107.835 23.400 107.880 ;
        RECT 22.165 107.680 22.455 107.725 ;
        RECT 19.940 107.540 22.455 107.680 ;
        RECT 23.185 107.680 23.400 107.835 ;
        RECT 23.990 108.020 24.320 108.065 ;
        RECT 27.290 108.020 27.580 108.065 ;
        RECT 23.990 107.880 27.580 108.020 ;
        RECT 23.990 107.835 24.320 107.880 ;
        RECT 27.290 107.835 27.580 107.880 ;
        RECT 35.050 108.020 35.340 108.065 ;
        RECT 36.910 108.020 37.200 108.065 ;
        RECT 35.050 107.880 37.200 108.020 ;
        RECT 35.050 107.835 35.340 107.880 ;
        RECT 36.910 107.835 37.200 107.880 ;
        RECT 37.830 108.020 38.120 108.065 ;
        RECT 41.090 108.020 41.380 108.065 ;
        RECT 44.245 108.020 44.535 108.065 ;
        RECT 37.830 107.880 44.535 108.020 ;
        RECT 37.830 107.835 38.120 107.880 ;
        RECT 41.090 107.835 41.380 107.880 ;
        RECT 44.245 107.835 44.535 107.880 ;
        RECT 46.550 108.020 46.840 108.065 ;
        RECT 48.410 108.020 48.700 108.065 ;
        RECT 46.550 107.880 48.700 108.020 ;
        RECT 46.550 107.835 46.840 107.880 ;
        RECT 48.410 107.835 48.700 107.880 ;
        RECT 49.330 108.020 49.620 108.065 ;
        RECT 50.210 108.020 50.530 108.080 ;
        RECT 52.590 108.020 52.880 108.065 ;
        RECT 49.330 107.880 52.880 108.020 ;
        RECT 49.330 107.835 49.620 107.880 ;
        RECT 23.990 107.820 24.310 107.835 ;
        RECT 25.430 107.680 25.720 107.725 ;
        RECT 23.185 107.540 25.720 107.680 ;
        RECT 22.165 107.495 22.455 107.540 ;
        RECT 25.430 107.495 25.720 107.540 ;
        RECT 32.730 107.480 33.050 107.740 ;
        RECT 34.125 107.680 34.415 107.725 ;
        RECT 36.985 107.680 37.200 107.835 ;
        RECT 39.230 107.680 39.520 107.725 ;
        RECT 34.125 107.540 36.640 107.680 ;
        RECT 36.985 107.540 39.520 107.680 ;
        RECT 34.125 107.495 34.415 107.540 ;
        RECT 20.310 107.140 20.630 107.400 ;
        RECT 35.965 107.340 36.255 107.385 ;
        RECT 33.740 107.200 36.255 107.340 ;
        RECT 36.500 107.340 36.640 107.540 ;
        RECT 39.230 107.495 39.520 107.540 ;
        RECT 44.705 107.680 44.995 107.725 ;
        RECT 44.705 107.540 47.220 107.680 ;
        RECT 44.705 107.495 44.995 107.540 ;
        RECT 39.630 107.340 39.950 107.400 ;
        RECT 45.625 107.340 45.915 107.385 ;
        RECT 36.500 107.200 45.915 107.340 ;
        RECT 47.080 107.340 47.220 107.540 ;
        RECT 47.450 107.480 47.770 107.740 ;
        RECT 48.485 107.680 48.700 107.835 ;
        RECT 50.210 107.820 50.530 107.880 ;
        RECT 52.590 107.835 52.880 107.880 ;
        RECT 58.030 108.020 58.350 108.080 ;
        RECT 59.960 108.020 60.100 108.175 ;
        RECT 61.710 108.160 62.030 108.420 ;
        RECT 64.930 108.160 65.250 108.420 ;
        RECT 72.750 108.160 73.070 108.420 ;
        RECT 79.650 108.160 79.970 108.420 ;
        RECT 107.725 108.360 108.015 108.405 ;
        RECT 109.550 108.360 109.870 108.420 ;
        RECT 107.725 108.220 109.870 108.360 ;
        RECT 107.725 108.175 108.015 108.220 ;
        RECT 109.550 108.160 109.870 108.220 ;
        RECT 111.405 108.175 111.695 108.405 ;
        RECT 58.030 107.880 60.100 108.020 ;
        RECT 60.790 108.020 61.110 108.080 ;
        RECT 62.185 108.020 62.475 108.065 ;
        RECT 77.350 108.020 77.670 108.080 ;
        RECT 96.670 108.065 96.990 108.080 ;
        RECT 60.790 107.880 62.475 108.020 ;
        RECT 58.030 107.820 58.350 107.880 ;
        RECT 60.790 107.820 61.110 107.880 ;
        RECT 62.185 107.835 62.475 107.880 ;
        RECT 65.480 107.880 77.670 108.020 ;
        RECT 50.730 107.680 51.020 107.725 ;
        RECT 48.485 107.540 51.020 107.680 ;
        RECT 50.730 107.495 51.020 107.540 ;
        RECT 51.590 107.680 51.910 107.740 ;
        RECT 65.480 107.725 65.620 107.880 ;
        RECT 77.350 107.820 77.670 107.880 ;
        RECT 96.620 108.020 96.990 108.065 ;
        RECT 99.880 108.020 100.170 108.065 ;
        RECT 96.620 107.880 100.170 108.020 ;
        RECT 96.620 107.835 96.990 107.880 ;
        RECT 99.880 107.835 100.170 107.880 ;
        RECT 100.800 108.020 101.090 108.065 ;
        RECT 102.660 108.020 102.950 108.065 ;
        RECT 100.800 107.880 102.950 108.020 ;
        RECT 100.800 107.835 101.090 107.880 ;
        RECT 102.660 107.835 102.950 107.880 ;
        RECT 96.670 107.820 96.990 107.835 ;
        RECT 58.505 107.680 58.795 107.725 ;
        RECT 65.405 107.680 65.695 107.725 ;
        RECT 51.590 107.540 65.695 107.680 ;
        RECT 51.590 107.480 51.910 107.540 ;
        RECT 58.505 107.495 58.795 107.540 ;
        RECT 65.405 107.495 65.695 107.540 ;
        RECT 73.685 107.495 73.975 107.725 ;
        RECT 74.130 107.680 74.450 107.740 ;
        RECT 75.050 107.680 75.370 107.740 ;
        RECT 74.130 107.540 75.370 107.680 ;
        RECT 51.680 107.340 51.820 107.480 ;
        RECT 47.080 107.200 51.820 107.340 ;
        RECT 57.110 107.340 57.430 107.400 ;
        RECT 62.630 107.340 62.950 107.400 ;
        RECT 57.110 107.200 62.950 107.340 ;
        RECT 33.740 107.045 33.880 107.200 ;
        RECT 35.965 107.155 36.255 107.200 ;
        RECT 39.630 107.140 39.950 107.200 ;
        RECT 45.625 107.155 45.915 107.200 ;
        RECT 57.110 107.140 57.430 107.200 ;
        RECT 62.630 107.140 62.950 107.200 ;
        RECT 20.790 107.000 21.080 107.045 ;
        RECT 22.650 107.000 22.940 107.045 ;
        RECT 25.430 107.000 25.720 107.045 ;
        RECT 20.790 106.860 25.720 107.000 ;
        RECT 20.790 106.815 21.080 106.860 ;
        RECT 22.650 106.815 22.940 106.860 ;
        RECT 25.430 106.815 25.720 106.860 ;
        RECT 33.665 106.815 33.955 107.045 ;
        RECT 34.590 107.000 34.880 107.045 ;
        RECT 36.450 107.000 36.740 107.045 ;
        RECT 39.230 107.000 39.520 107.045 ;
        RECT 34.590 106.860 39.520 107.000 ;
        RECT 34.590 106.815 34.880 106.860 ;
        RECT 36.450 106.815 36.740 106.860 ;
        RECT 39.230 106.815 39.520 106.860 ;
        RECT 46.090 107.000 46.380 107.045 ;
        RECT 47.950 107.000 48.240 107.045 ;
        RECT 50.730 107.000 51.020 107.045 ;
        RECT 46.090 106.860 51.020 107.000 ;
        RECT 73.760 107.000 73.900 107.495 ;
        RECT 74.130 107.480 74.450 107.540 ;
        RECT 75.050 107.480 75.370 107.540 ;
        RECT 83.790 107.480 84.110 107.740 ;
        RECT 98.480 107.680 98.770 107.725 ;
        RECT 100.800 107.680 101.015 107.835 ;
        RECT 98.480 107.540 101.015 107.680 ;
        RECT 98.480 107.495 98.770 107.540 ;
        RECT 101.730 107.480 102.050 107.740 ;
        RECT 106.805 107.680 107.095 107.725 ;
        RECT 107.250 107.680 107.570 107.740 ;
        RECT 106.805 107.540 107.570 107.680 ;
        RECT 106.805 107.495 107.095 107.540 ;
        RECT 107.250 107.480 107.570 107.540 ;
        RECT 110.470 107.480 110.790 107.740 ;
        RECT 111.480 107.680 111.620 108.175 ;
        RECT 112.790 108.020 113.080 108.065 ;
        RECT 114.650 108.020 114.940 108.065 ;
        RECT 112.790 107.880 114.940 108.020 ;
        RECT 112.790 107.835 113.080 107.880 ;
        RECT 114.650 107.835 114.940 107.880 ;
        RECT 115.570 108.020 115.860 108.065 ;
        RECT 116.450 108.020 116.770 108.080 ;
        RECT 118.830 108.020 119.120 108.065 ;
        RECT 115.570 107.880 119.120 108.020 ;
        RECT 115.570 107.835 115.860 107.880 ;
        RECT 113.705 107.680 113.995 107.725 ;
        RECT 111.480 107.540 113.995 107.680 ;
        RECT 114.725 107.680 114.940 107.835 ;
        RECT 116.450 107.820 116.770 107.880 ;
        RECT 118.830 107.835 119.120 107.880 ;
        RECT 116.970 107.680 117.260 107.725 ;
        RECT 114.725 107.540 117.260 107.680 ;
        RECT 113.705 107.495 113.995 107.540 ;
        RECT 116.970 107.495 117.260 107.540 ;
        RECT 75.525 107.340 75.815 107.385 ;
        RECT 76.890 107.340 77.210 107.400 ;
        RECT 75.525 107.200 77.210 107.340 ;
        RECT 75.525 107.155 75.815 107.200 ;
        RECT 76.890 107.140 77.210 107.200 ;
        RECT 80.125 107.155 80.415 107.385 ;
        RECT 80.570 107.340 80.890 107.400 ;
        RECT 87.930 107.340 88.250 107.400 ;
        RECT 80.570 107.200 88.250 107.340 ;
        RECT 77.825 107.000 78.115 107.045 ;
        RECT 73.760 106.860 78.115 107.000 ;
        RECT 80.200 107.000 80.340 107.155 ;
        RECT 80.570 107.140 80.890 107.200 ;
        RECT 87.930 107.140 88.250 107.200 ;
        RECT 103.585 107.340 103.875 107.385 ;
        RECT 109.090 107.340 109.410 107.400 ;
        RECT 111.865 107.340 112.155 107.385 ;
        RECT 103.585 107.200 112.155 107.340 ;
        RECT 103.585 107.155 103.875 107.200 ;
        RECT 109.090 107.140 109.410 107.200 ;
        RECT 111.865 107.155 112.155 107.200 ;
        RECT 83.330 107.000 83.650 107.060 ;
        RECT 80.200 106.860 83.650 107.000 ;
        RECT 46.090 106.815 46.380 106.860 ;
        RECT 47.950 106.815 48.240 106.860 ;
        RECT 50.730 106.815 51.020 106.860 ;
        RECT 77.825 106.815 78.115 106.860 ;
        RECT 83.330 106.800 83.650 106.860 ;
        RECT 93.450 107.000 93.770 107.060 ;
        RECT 94.615 107.000 94.905 107.045 ;
        RECT 93.450 106.860 94.905 107.000 ;
        RECT 93.450 106.800 93.770 106.860 ;
        RECT 94.615 106.815 94.905 106.860 ;
        RECT 98.480 107.000 98.770 107.045 ;
        RECT 101.260 107.000 101.550 107.045 ;
        RECT 103.120 107.000 103.410 107.045 ;
        RECT 98.480 106.860 103.410 107.000 ;
        RECT 98.480 106.815 98.770 106.860 ;
        RECT 101.260 106.815 101.550 106.860 ;
        RECT 103.120 106.815 103.410 106.860 ;
        RECT 112.330 107.000 112.620 107.045 ;
        RECT 114.190 107.000 114.480 107.045 ;
        RECT 116.970 107.000 117.260 107.045 ;
        RECT 112.330 106.860 117.260 107.000 ;
        RECT 112.330 106.815 112.620 106.860 ;
        RECT 114.190 106.815 114.480 106.860 ;
        RECT 116.970 106.815 117.260 106.860 ;
        RECT 27.670 106.660 27.990 106.720 ;
        RECT 29.295 106.660 29.585 106.705 ;
        RECT 27.670 106.520 29.585 106.660 ;
        RECT 27.670 106.460 27.990 106.520 ;
        RECT 29.295 106.475 29.585 106.520 ;
        RECT 43.095 106.660 43.385 106.705 ;
        RECT 46.990 106.660 47.310 106.720 ;
        RECT 43.095 106.520 47.310 106.660 ;
        RECT 43.095 106.475 43.385 106.520 ;
        RECT 46.990 106.460 47.310 106.520 ;
        RECT 52.970 106.660 53.290 106.720 ;
        RECT 54.595 106.660 54.885 106.705 ;
        RECT 52.970 106.520 54.885 106.660 ;
        RECT 52.970 106.460 53.290 106.520 ;
        RECT 54.595 106.475 54.885 106.520 ;
        RECT 114.610 106.660 114.930 106.720 ;
        RECT 120.835 106.660 121.125 106.705 ;
        RECT 114.610 106.520 121.125 106.660 ;
        RECT 114.610 106.460 114.930 106.520 ;
        RECT 120.835 106.475 121.125 106.520 ;
        RECT 5.520 105.840 123.740 106.320 ;
        RECT 18.930 105.640 19.250 105.700 ;
        RECT 21.245 105.640 21.535 105.685 ;
        RECT 18.930 105.500 21.535 105.640 ;
        RECT 18.930 105.440 19.250 105.500 ;
        RECT 21.245 105.455 21.535 105.500 ;
        RECT 35.950 105.440 36.270 105.700 ;
        RECT 49.290 105.640 49.610 105.700 ;
        RECT 53.905 105.640 54.195 105.685 ;
        RECT 57.110 105.640 57.430 105.700 ;
        RECT 49.290 105.500 54.195 105.640 ;
        RECT 49.290 105.440 49.610 105.500 ;
        RECT 53.905 105.455 54.195 105.500 ;
        RECT 56.740 105.500 57.430 105.640 ;
        RECT 17.565 104.960 17.855 105.005 ;
        RECT 18.930 104.960 19.250 105.020 ;
        RECT 22.150 104.960 22.470 105.020 ;
        RECT 24.465 104.960 24.755 105.005 ;
        RECT 35.030 104.960 35.350 105.020 ;
        RECT 39.185 104.960 39.475 105.005 ;
        RECT 47.910 104.960 48.230 105.020 ;
        RECT 56.740 105.005 56.880 105.500 ;
        RECT 57.110 105.440 57.430 105.500 ;
        RECT 62.630 105.640 62.950 105.700 ;
        RECT 66.325 105.640 66.615 105.685 ;
        RECT 62.630 105.500 66.615 105.640 ;
        RECT 62.630 105.440 62.950 105.500 ;
        RECT 66.325 105.455 66.615 105.500 ;
        RECT 76.430 105.440 76.750 105.700 ;
        RECT 86.550 105.440 86.870 105.700 ;
        RECT 89.770 105.640 90.090 105.700 ;
        RECT 92.530 105.640 92.850 105.700 ;
        RECT 89.770 105.500 92.850 105.640 ;
        RECT 89.770 105.440 90.090 105.500 ;
        RECT 92.530 105.440 92.850 105.500 ;
        RECT 110.470 105.640 110.790 105.700 ;
        RECT 112.325 105.640 112.615 105.685 ;
        RECT 110.470 105.500 112.615 105.640 ;
        RECT 110.470 105.440 110.790 105.500 ;
        RECT 112.325 105.455 112.615 105.500 ;
        RECT 116.450 105.640 116.770 105.700 ;
        RECT 116.925 105.640 117.215 105.685 ;
        RECT 116.450 105.500 117.215 105.640 ;
        RECT 116.450 105.440 116.770 105.500 ;
        RECT 116.925 105.455 117.215 105.500 ;
        RECT 73.685 105.300 73.975 105.345 ;
        RECT 80.570 105.300 80.890 105.360 ;
        RECT 73.685 105.160 80.890 105.300 ;
        RECT 73.685 105.115 73.975 105.160 ;
        RECT 80.570 105.100 80.890 105.160 ;
        RECT 81.510 105.300 81.800 105.345 ;
        RECT 83.370 105.300 83.660 105.345 ;
        RECT 86.150 105.300 86.440 105.345 ;
        RECT 81.510 105.160 86.440 105.300 ;
        RECT 86.640 105.300 86.780 105.440 ;
        RECT 86.640 105.160 99.200 105.300 ;
        RECT 81.510 105.115 81.800 105.160 ;
        RECT 83.370 105.115 83.660 105.160 ;
        RECT 86.150 105.115 86.440 105.160 ;
        RECT 56.665 104.960 56.955 105.005 ;
        RECT 59.885 104.960 60.175 105.005 ;
        RECT 61.710 104.960 62.030 105.020 ;
        RECT 17.565 104.820 56.955 104.960 ;
        RECT 17.565 104.775 17.855 104.820 ;
        RECT 18.930 104.760 19.250 104.820 ;
        RECT 22.150 104.760 22.470 104.820 ;
        RECT 24.465 104.775 24.755 104.820 ;
        RECT 35.030 104.760 35.350 104.820 ;
        RECT 39.185 104.775 39.475 104.820 ;
        RECT 47.910 104.760 48.230 104.820 ;
        RECT 56.665 104.775 56.955 104.820 ;
        RECT 58.580 104.820 62.030 104.960 ;
        RECT 12.505 104.435 12.795 104.665 ;
        RECT 13.885 104.620 14.175 104.665 ;
        RECT 16.630 104.620 16.950 104.680 ;
        RECT 21.690 104.620 22.010 104.680 ;
        RECT 13.885 104.480 22.010 104.620 ;
        RECT 13.885 104.435 14.175 104.480 ;
        RECT 12.580 104.280 12.720 104.435 ;
        RECT 16.630 104.420 16.950 104.480 ;
        RECT 21.690 104.420 22.010 104.480 ;
        RECT 23.085 104.620 23.375 104.665 ;
        RECT 27.670 104.620 27.990 104.680 ;
        RECT 23.085 104.480 27.990 104.620 ;
        RECT 23.085 104.435 23.375 104.480 ;
        RECT 27.670 104.420 27.990 104.480 ;
        RECT 38.265 104.620 38.555 104.665 ;
        RECT 52.970 104.620 53.290 104.680 ;
        RECT 55.745 104.620 56.035 104.665 ;
        RECT 38.265 104.480 56.035 104.620 ;
        RECT 38.265 104.435 38.555 104.480 ;
        RECT 52.970 104.420 53.290 104.480 ;
        RECT 55.745 104.435 56.035 104.480 ;
        RECT 56.205 104.620 56.495 104.665 ;
        RECT 58.580 104.620 58.720 104.820 ;
        RECT 59.885 104.775 60.175 104.820 ;
        RECT 61.710 104.760 62.030 104.820 ;
        RECT 75.510 104.960 75.830 105.020 ;
        RECT 81.045 104.960 81.335 105.005 ;
        RECT 83.790 104.960 84.110 105.020 ;
        RECT 75.510 104.820 84.110 104.960 ;
        RECT 75.510 104.760 75.830 104.820 ;
        RECT 81.045 104.775 81.335 104.820 ;
        RECT 83.790 104.760 84.110 104.820 ;
        RECT 89.770 104.960 90.090 105.020 ;
        RECT 90.705 104.960 90.995 105.005 ;
        RECT 89.770 104.820 90.995 104.960 ;
        RECT 89.770 104.760 90.090 104.820 ;
        RECT 90.705 104.775 90.995 104.820 ;
        RECT 56.205 104.480 58.720 104.620 ;
        RECT 56.205 104.435 56.495 104.480 ;
        RECT 58.950 104.420 59.270 104.680 ;
        RECT 76.890 104.420 77.210 104.680 ;
        RECT 78.730 104.420 79.050 104.680 ;
        RECT 79.650 104.420 79.970 104.680 ;
        RECT 82.870 104.420 83.190 104.680 ;
        RECT 86.150 104.620 86.440 104.665 ;
        RECT 83.905 104.480 86.440 104.620 ;
        RECT 18.010 104.280 18.330 104.340 ;
        RECT 12.580 104.140 18.330 104.280 ;
        RECT 18.010 104.080 18.330 104.140 ;
        RECT 25.370 104.080 25.690 104.340 ;
        RECT 27.210 104.280 27.530 104.340 ;
        RECT 37.805 104.280 38.095 104.325 ;
        RECT 27.210 104.140 38.095 104.280 ;
        RECT 27.210 104.080 27.530 104.140 ;
        RECT 37.805 104.095 38.095 104.140 ;
        RECT 39.170 104.280 39.490 104.340 ;
        RECT 41.945 104.280 42.235 104.325 ;
        RECT 39.170 104.140 42.235 104.280 ;
        RECT 39.170 104.080 39.490 104.140 ;
        RECT 41.945 104.095 42.235 104.140 ;
        RECT 11.570 103.740 11.890 104.000 ;
        RECT 13.425 103.940 13.715 103.985 ;
        RECT 13.870 103.940 14.190 104.000 ;
        RECT 13.425 103.800 14.190 103.940 ;
        RECT 13.425 103.755 13.715 103.800 ;
        RECT 13.870 103.740 14.190 103.800 ;
        RECT 14.330 103.740 14.650 104.000 ;
        RECT 16.170 103.740 16.490 104.000 ;
        RECT 16.645 103.940 16.935 103.985 ;
        RECT 19.850 103.940 20.170 104.000 ;
        RECT 16.645 103.800 20.170 103.940 ;
        RECT 16.645 103.755 16.935 103.800 ;
        RECT 19.850 103.740 20.170 103.800 ;
        RECT 23.530 103.740 23.850 104.000 ;
        RECT 31.350 103.940 31.670 104.000 ;
        RECT 31.825 103.940 32.115 103.985 ;
        RECT 31.350 103.800 32.115 103.940 ;
        RECT 42.020 103.940 42.160 104.095 ;
        RECT 44.690 104.080 45.010 104.340 ;
        RECT 67.705 104.280 67.995 104.325 ;
        RECT 68.150 104.280 68.470 104.340 ;
        RECT 72.305 104.280 72.595 104.325 ;
        RECT 67.705 104.140 72.595 104.280 ;
        RECT 76.980 104.280 77.120 104.420 ;
        RECT 83.905 104.325 84.120 104.480 ;
        RECT 86.150 104.435 86.440 104.480 ;
        RECT 90.230 104.420 90.550 104.680 ;
        RECT 91.610 104.420 91.930 104.680 ;
        RECT 92.070 104.420 92.390 104.680 ;
        RECT 99.060 104.665 99.200 105.160 ;
        RECT 113.230 104.960 113.550 105.020 ;
        RECT 115.085 104.960 115.375 105.005 ;
        RECT 113.230 104.820 115.375 104.960 ;
        RECT 113.230 104.760 113.550 104.820 ;
        RECT 115.085 104.775 115.375 104.820 ;
        RECT 98.985 104.620 99.275 104.665 ;
        RECT 102.650 104.620 102.970 104.680 ;
        RECT 113.690 104.620 114.010 104.680 ;
        RECT 114.165 104.620 114.455 104.665 ;
        RECT 114.610 104.620 114.930 104.680 ;
        RECT 98.985 104.480 113.460 104.620 ;
        RECT 98.985 104.435 99.275 104.480 ;
        RECT 102.650 104.420 102.970 104.480 ;
        RECT 81.970 104.280 82.260 104.325 ;
        RECT 83.830 104.280 84.120 104.325 ;
        RECT 76.980 104.140 81.260 104.280 ;
        RECT 67.705 104.095 67.995 104.140 ;
        RECT 68.150 104.080 68.470 104.140 ;
        RECT 72.305 104.095 72.595 104.140 ;
        RECT 51.145 103.940 51.435 103.985 ;
        RECT 56.650 103.940 56.970 104.000 ;
        RECT 42.020 103.800 56.970 103.940 ;
        RECT 31.350 103.740 31.670 103.800 ;
        RECT 31.825 103.755 32.115 103.800 ;
        RECT 51.145 103.755 51.435 103.800 ;
        RECT 56.650 103.740 56.970 103.800 ;
        RECT 57.110 103.940 57.430 104.000 ;
        RECT 58.045 103.940 58.335 103.985 ;
        RECT 57.110 103.800 58.335 103.940 ;
        RECT 57.110 103.740 57.430 103.800 ;
        RECT 58.045 103.755 58.335 103.800 ;
        RECT 80.570 103.740 80.890 104.000 ;
        RECT 81.120 103.940 81.260 104.140 ;
        RECT 81.970 104.140 84.120 104.280 ;
        RECT 81.970 104.095 82.260 104.140 ;
        RECT 83.830 104.095 84.120 104.140 ;
        RECT 84.750 104.280 85.040 104.325 ;
        RECT 88.010 104.280 88.300 104.325 ;
        RECT 89.310 104.280 89.630 104.340 ;
        RECT 84.750 104.140 89.630 104.280 ;
        RECT 90.320 104.280 90.460 104.420 ;
        RECT 100.365 104.280 100.655 104.325 ;
        RECT 90.320 104.140 100.655 104.280 ;
        RECT 84.750 104.095 85.040 104.140 ;
        RECT 88.010 104.095 88.300 104.140 ;
        RECT 89.310 104.080 89.630 104.140 ;
        RECT 100.365 104.095 100.655 104.140 ;
        RECT 109.090 104.080 109.410 104.340 ;
        RECT 113.320 104.280 113.460 104.480 ;
        RECT 113.690 104.480 114.930 104.620 ;
        RECT 113.690 104.420 114.010 104.480 ;
        RECT 114.165 104.435 114.455 104.480 ;
        RECT 114.610 104.420 114.930 104.480 ;
        RECT 116.465 104.620 116.755 104.665 ;
        RECT 117.370 104.620 117.690 104.680 ;
        RECT 116.465 104.480 117.690 104.620 ;
        RECT 116.465 104.435 116.755 104.480 ;
        RECT 116.540 104.280 116.680 104.435 ;
        RECT 117.370 104.420 117.690 104.480 ;
        RECT 113.320 104.140 116.680 104.280 ;
        RECT 86.550 103.940 86.870 104.000 ;
        RECT 81.120 103.800 86.870 103.940 ;
        RECT 86.550 103.740 86.870 103.800 ;
        RECT 88.850 103.940 89.170 104.000 ;
        RECT 90.015 103.940 90.305 103.985 ;
        RECT 88.850 103.800 90.305 103.940 ;
        RECT 88.850 103.740 89.170 103.800 ;
        RECT 90.015 103.755 90.305 103.800 ;
        RECT 99.445 103.940 99.735 103.985 ;
        RECT 100.810 103.940 101.130 104.000 ;
        RECT 99.445 103.800 101.130 103.940 ;
        RECT 99.445 103.755 99.735 103.800 ;
        RECT 100.810 103.740 101.130 103.800 ;
        RECT 105.410 103.940 105.730 104.000 ;
        RECT 114.625 103.940 114.915 103.985 ;
        RECT 105.410 103.800 114.915 103.940 ;
        RECT 105.410 103.740 105.730 103.800 ;
        RECT 114.625 103.755 114.915 103.800 ;
        RECT 5.520 103.120 123.740 103.600 ;
        RECT 7.905 102.735 8.195 102.965 ;
        RECT 6.985 102.240 7.275 102.285 ;
        RECT 7.980 102.240 8.120 102.735 ;
        RECT 18.010 102.720 18.330 102.980 ;
        RECT 31.825 102.920 32.115 102.965 ;
        RECT 32.730 102.920 33.050 102.980 ;
        RECT 31.825 102.780 33.050 102.920 ;
        RECT 31.825 102.735 32.115 102.780 ;
        RECT 32.730 102.720 33.050 102.780 ;
        RECT 42.390 102.920 42.710 102.980 ;
        RECT 44.705 102.920 44.995 102.965 ;
        RECT 42.390 102.780 44.995 102.920 ;
        RECT 42.390 102.720 42.710 102.780 ;
        RECT 44.705 102.735 44.995 102.780 ;
        RECT 46.990 102.720 47.310 102.980 ;
        RECT 68.150 102.720 68.470 102.980 ;
        RECT 86.565 102.920 86.855 102.965 ;
        RECT 87.010 102.920 87.330 102.980 ;
        RECT 86.565 102.780 87.330 102.920 ;
        RECT 86.565 102.735 86.855 102.780 ;
        RECT 87.010 102.720 87.330 102.780 ;
        RECT 87.470 102.920 87.790 102.980 ;
        RECT 102.650 102.920 102.970 102.980 ;
        RECT 111.405 102.920 111.695 102.965 ;
        RECT 87.470 102.780 91.840 102.920 ;
        RECT 87.470 102.720 87.790 102.780 ;
        RECT 9.290 102.580 9.580 102.625 ;
        RECT 11.150 102.580 11.440 102.625 ;
        RECT 9.290 102.440 11.440 102.580 ;
        RECT 9.290 102.395 9.580 102.440 ;
        RECT 11.150 102.395 11.440 102.440 ;
        RECT 12.070 102.580 12.360 102.625 ;
        RECT 13.870 102.580 14.190 102.640 ;
        RECT 15.330 102.580 15.620 102.625 ;
        RECT 12.070 102.440 15.620 102.580 ;
        RECT 12.070 102.395 12.360 102.440 ;
        RECT 10.205 102.240 10.495 102.285 ;
        RECT 6.985 102.100 7.660 102.240 ;
        RECT 7.980 102.100 10.495 102.240 ;
        RECT 11.225 102.240 11.440 102.395 ;
        RECT 13.870 102.380 14.190 102.440 ;
        RECT 15.330 102.395 15.620 102.440 ;
        RECT 20.325 102.580 20.615 102.625 ;
        RECT 20.770 102.580 21.090 102.640 ;
        RECT 26.290 102.580 26.610 102.640 ;
        RECT 29.510 102.580 29.830 102.640 ;
        RECT 20.325 102.440 26.610 102.580 ;
        RECT 20.325 102.395 20.615 102.440 ;
        RECT 20.770 102.380 21.090 102.440 ;
        RECT 26.290 102.380 26.610 102.440 ;
        RECT 27.300 102.440 29.830 102.580 ;
        RECT 13.470 102.240 13.760 102.285 ;
        RECT 11.225 102.100 13.760 102.240 ;
        RECT 6.985 102.055 7.275 102.100 ;
        RECT 7.520 101.220 7.660 102.100 ;
        RECT 10.205 102.055 10.495 102.100 ;
        RECT 13.470 102.055 13.760 102.100 ;
        RECT 19.850 102.040 20.170 102.300 ;
        RECT 21.690 102.240 22.010 102.300 ;
        RECT 23.085 102.240 23.375 102.285 ;
        RECT 27.300 102.240 27.440 102.440 ;
        RECT 29.510 102.380 29.830 102.440 ;
        RECT 33.665 102.580 33.955 102.625 ;
        RECT 35.950 102.580 36.270 102.640 ;
        RECT 47.080 102.580 47.220 102.720 ;
        RECT 91.700 102.640 91.840 102.780 ;
        RECT 102.650 102.780 111.695 102.920 ;
        RECT 102.650 102.720 102.970 102.780 ;
        RECT 111.405 102.735 111.695 102.780 ;
        RECT 88.405 102.580 88.695 102.625 ;
        RECT 88.850 102.580 89.170 102.640 ;
        RECT 33.665 102.440 47.220 102.580 ;
        RECT 84.340 102.440 89.170 102.580 ;
        RECT 33.665 102.395 33.955 102.440 ;
        RECT 35.950 102.380 36.270 102.440 ;
        RECT 21.690 102.100 27.440 102.240 ;
        RECT 27.685 102.240 27.975 102.285 ;
        RECT 28.130 102.240 28.450 102.300 ;
        RECT 27.685 102.100 28.450 102.240 ;
        RECT 21.690 102.040 22.010 102.100 ;
        RECT 23.085 102.055 23.375 102.100 ;
        RECT 27.685 102.055 27.975 102.100 ;
        RECT 28.130 102.040 28.450 102.100 ;
        RECT 46.545 102.240 46.835 102.285 ;
        RECT 50.670 102.240 50.990 102.300 ;
        RECT 46.545 102.100 50.990 102.240 ;
        RECT 46.545 102.055 46.835 102.100 ;
        RECT 50.670 102.040 50.990 102.100 ;
        RECT 51.605 102.240 51.895 102.285 ;
        RECT 53.905 102.240 54.195 102.285 ;
        RECT 58.505 102.240 58.795 102.285 ;
        RECT 58.950 102.240 59.270 102.300 ;
        RECT 51.605 102.100 59.270 102.240 ;
        RECT 51.605 102.055 51.895 102.100 ;
        RECT 53.905 102.055 54.195 102.100 ;
        RECT 58.505 102.055 58.795 102.100 ;
        RECT 7.890 101.900 8.210 101.960 ;
        RECT 8.365 101.900 8.655 101.945 ;
        RECT 7.890 101.760 8.655 101.900 ;
        RECT 7.890 101.700 8.210 101.760 ;
        RECT 8.365 101.715 8.655 101.760 ;
        RECT 18.930 101.900 19.250 101.960 ;
        RECT 20.785 101.900 21.075 101.945 ;
        RECT 18.930 101.760 21.075 101.900 ;
        RECT 18.930 101.700 19.250 101.760 ;
        RECT 20.785 101.715 21.075 101.760 ;
        RECT 21.230 101.900 21.550 101.960 ;
        RECT 26.765 101.900 27.055 101.945 ;
        RECT 27.210 101.900 27.530 101.960 ;
        RECT 21.230 101.760 27.530 101.900 ;
        RECT 21.230 101.700 21.550 101.760 ;
        RECT 26.765 101.715 27.055 101.760 ;
        RECT 27.210 101.700 27.530 101.760 ;
        RECT 34.125 101.715 34.415 101.945 ;
        RECT 8.830 101.560 9.120 101.605 ;
        RECT 10.690 101.560 10.980 101.605 ;
        RECT 13.470 101.560 13.760 101.605 ;
        RECT 8.830 101.420 13.760 101.560 ;
        RECT 8.830 101.375 9.120 101.420 ;
        RECT 10.690 101.375 10.980 101.420 ;
        RECT 13.470 101.375 13.760 101.420 ;
        RECT 16.170 101.560 16.490 101.620 ;
        RECT 17.335 101.560 17.625 101.605 ;
        RECT 23.530 101.560 23.850 101.620 ;
        RECT 16.170 101.420 23.850 101.560 ;
        RECT 16.170 101.360 16.490 101.420 ;
        RECT 17.335 101.375 17.625 101.420 ;
        RECT 23.530 101.360 23.850 101.420 ;
        RECT 27.670 101.560 27.990 101.620 ;
        RECT 34.200 101.560 34.340 101.715 ;
        RECT 35.030 101.700 35.350 101.960 ;
        RECT 47.910 101.700 48.230 101.960 ;
        RECT 52.970 101.700 53.290 101.960 ;
        RECT 27.670 101.420 34.340 101.560 ;
        RECT 53.430 101.560 53.750 101.620 ;
        RECT 54.825 101.560 55.115 101.605 ;
        RECT 53.430 101.420 55.115 101.560 ;
        RECT 58.580 101.560 58.720 102.055 ;
        RECT 58.950 102.040 59.270 102.100 ;
        RECT 59.425 102.240 59.715 102.285 ;
        RECT 60.790 102.240 61.110 102.300 ;
        RECT 59.425 102.100 61.110 102.240 ;
        RECT 59.425 102.055 59.715 102.100 ;
        RECT 60.790 102.040 61.110 102.100 ;
        RECT 67.230 102.240 67.550 102.300 ;
        RECT 69.085 102.240 69.375 102.285 ;
        RECT 67.230 102.100 69.375 102.240 ;
        RECT 67.230 102.040 67.550 102.100 ;
        RECT 69.085 102.055 69.375 102.100 ;
        RECT 83.330 102.240 83.650 102.300 ;
        RECT 84.340 102.285 84.480 102.440 ;
        RECT 88.405 102.395 88.695 102.440 ;
        RECT 88.850 102.380 89.170 102.440 ;
        RECT 91.610 102.580 91.930 102.640 ;
        RECT 96.210 102.580 96.530 102.640 ;
        RECT 100.810 102.625 101.130 102.640 ;
        RECT 98.070 102.580 98.360 102.625 ;
        RECT 99.930 102.580 100.220 102.625 ;
        RECT 91.610 102.440 95.520 102.580 ;
        RECT 91.610 102.380 91.930 102.440 ;
        RECT 84.265 102.240 84.555 102.285 ;
        RECT 83.330 102.100 84.555 102.240 ;
        RECT 83.330 102.040 83.650 102.100 ;
        RECT 84.265 102.055 84.555 102.100 ;
        RECT 85.185 102.055 85.475 102.285 ;
        RECT 86.105 102.240 86.395 102.285 ;
        RECT 92.070 102.240 92.390 102.300 ;
        RECT 92.620 102.285 92.760 102.440 ;
        RECT 95.380 102.300 95.520 102.440 ;
        RECT 96.210 102.440 97.360 102.580 ;
        RECT 96.210 102.380 96.530 102.440 ;
        RECT 86.105 102.100 92.390 102.240 ;
        RECT 86.105 102.055 86.395 102.100 ;
        RECT 66.310 101.700 66.630 101.960 ;
        RECT 70.005 101.900 70.295 101.945 ;
        RECT 79.650 101.900 79.970 101.960 ;
        RECT 85.260 101.900 85.400 102.055 ;
        RECT 92.070 102.040 92.390 102.100 ;
        RECT 92.545 102.055 92.835 102.285 ;
        RECT 93.450 102.040 93.770 102.300 ;
        RECT 95.290 102.040 95.610 102.300 ;
        RECT 97.220 102.285 97.360 102.440 ;
        RECT 98.070 102.440 100.220 102.580 ;
        RECT 98.070 102.395 98.360 102.440 ;
        RECT 99.930 102.395 100.220 102.440 ;
        RECT 97.145 102.240 97.435 102.285 ;
        RECT 100.005 102.240 100.220 102.395 ;
        RECT 100.810 102.580 101.140 102.625 ;
        RECT 104.110 102.580 104.400 102.625 ;
        RECT 100.810 102.440 104.400 102.580 ;
        RECT 100.810 102.395 101.140 102.440 ;
        RECT 104.110 102.395 104.400 102.440 ;
        RECT 100.810 102.380 101.130 102.395 ;
        RECT 102.250 102.240 102.540 102.285 ;
        RECT 97.145 102.100 99.660 102.240 ;
        RECT 100.005 102.100 102.540 102.240 ;
        RECT 97.145 102.055 97.435 102.100 ;
        RECT 87.470 101.900 87.790 101.960 ;
        RECT 70.005 101.760 87.790 101.900 ;
        RECT 70.005 101.715 70.295 101.760 ;
        RECT 70.080 101.560 70.220 101.715 ;
        RECT 79.650 101.700 79.970 101.760 ;
        RECT 87.470 101.700 87.790 101.760 ;
        RECT 88.865 101.715 89.155 101.945 ;
        RECT 58.580 101.420 70.220 101.560 ;
        RECT 88.940 101.560 89.080 101.715 ;
        RECT 89.310 101.700 89.630 101.960 ;
        RECT 96.225 101.900 96.515 101.945 ;
        RECT 98.050 101.900 98.370 101.960 ;
        RECT 96.225 101.760 98.370 101.900 ;
        RECT 96.225 101.715 96.515 101.760 ;
        RECT 98.050 101.700 98.370 101.760 ;
        RECT 98.970 101.700 99.290 101.960 ;
        RECT 99.520 101.900 99.660 102.100 ;
        RECT 102.250 102.055 102.540 102.100 ;
        RECT 114.625 102.240 114.915 102.285 ;
        RECT 117.370 102.240 117.690 102.300 ;
        RECT 114.625 102.100 117.690 102.240 ;
        RECT 114.625 102.055 114.915 102.100 ;
        RECT 117.370 102.040 117.690 102.100 ;
        RECT 109.090 101.900 109.410 101.960 ;
        RECT 99.520 101.760 109.410 101.900 ;
        RECT 109.090 101.700 109.410 101.760 ;
        RECT 111.850 101.700 112.170 101.960 ;
        RECT 112.785 101.900 113.075 101.945 ;
        RECT 113.230 101.900 113.550 101.960 ;
        RECT 112.785 101.760 113.550 101.900 ;
        RECT 112.785 101.715 113.075 101.760 ;
        RECT 113.230 101.700 113.550 101.760 ;
        RECT 97.130 101.560 97.450 101.620 ;
        RECT 88.940 101.420 97.450 101.560 ;
        RECT 27.670 101.360 27.990 101.420 ;
        RECT 53.430 101.360 53.750 101.420 ;
        RECT 54.825 101.375 55.115 101.420 ;
        RECT 97.130 101.360 97.450 101.420 ;
        RECT 97.610 101.560 97.900 101.605 ;
        RECT 99.470 101.560 99.760 101.605 ;
        RECT 102.250 101.560 102.540 101.605 ;
        RECT 97.610 101.420 102.540 101.560 ;
        RECT 97.610 101.375 97.900 101.420 ;
        RECT 99.470 101.375 99.760 101.420 ;
        RECT 102.250 101.375 102.540 101.420 ;
        RECT 14.330 101.220 14.650 101.280 ;
        RECT 7.520 101.080 14.650 101.220 ;
        RECT 14.330 101.020 14.650 101.080 ;
        RECT 18.470 101.220 18.790 101.280 ;
        RECT 22.625 101.220 22.915 101.265 ;
        RECT 18.470 101.080 22.915 101.220 ;
        RECT 18.470 101.020 18.790 101.080 ;
        RECT 22.625 101.035 22.915 101.080 ;
        RECT 28.590 101.020 28.910 101.280 ;
        RECT 52.525 101.220 52.815 101.265 ;
        RECT 53.890 101.220 54.210 101.280 ;
        RECT 52.525 101.080 54.210 101.220 ;
        RECT 52.525 101.035 52.815 101.080 ;
        RECT 53.890 101.020 54.210 101.080 ;
        RECT 57.570 101.020 57.890 101.280 ;
        RECT 91.610 101.020 91.930 101.280 ;
        RECT 94.370 101.020 94.690 101.280 ;
        RECT 97.220 101.220 97.360 101.360 ;
        RECT 106.115 101.220 106.405 101.265 ;
        RECT 97.220 101.080 106.405 101.220 ;
        RECT 106.115 101.035 106.405 101.080 ;
        RECT 109.565 101.220 109.855 101.265 ;
        RECT 110.010 101.220 110.330 101.280 ;
        RECT 109.565 101.080 110.330 101.220 ;
        RECT 109.565 101.035 109.855 101.080 ;
        RECT 110.010 101.020 110.330 101.080 ;
        RECT 114.150 101.020 114.470 101.280 ;
        RECT 5.520 100.400 123.740 100.880 ;
        RECT 16.875 100.200 17.165 100.245 ;
        RECT 19.850 100.200 20.170 100.260 ;
        RECT 16.875 100.060 20.170 100.200 ;
        RECT 16.875 100.015 17.165 100.060 ;
        RECT 19.850 100.000 20.170 100.060 ;
        RECT 98.970 100.000 99.290 100.260 ;
        RECT 105.410 100.200 105.730 100.260 ;
        RECT 99.980 100.060 105.730 100.200 ;
        RECT 8.370 99.860 8.660 99.905 ;
        RECT 10.230 99.860 10.520 99.905 ;
        RECT 13.010 99.860 13.300 99.905 ;
        RECT 8.370 99.720 13.300 99.860 ;
        RECT 8.370 99.675 8.660 99.720 ;
        RECT 10.230 99.675 10.520 99.720 ;
        RECT 13.010 99.675 13.300 99.720 ;
        RECT 23.530 99.660 23.850 99.920 ;
        RECT 99.980 99.860 100.120 100.060 ;
        RECT 105.410 100.000 105.730 100.060 ;
        RECT 98.140 99.720 100.120 99.860 ;
        RECT 9.745 99.520 10.035 99.565 ;
        RECT 11.570 99.520 11.890 99.580 ;
        RECT 9.745 99.380 11.890 99.520 ;
        RECT 9.745 99.335 10.035 99.380 ;
        RECT 11.570 99.320 11.890 99.380 ;
        RECT 22.625 99.520 22.915 99.565 ;
        RECT 23.620 99.520 23.760 99.660 ;
        RECT 22.625 99.380 23.760 99.520 ;
        RECT 35.950 99.520 36.270 99.580 ;
        RECT 36.425 99.520 36.715 99.565 ;
        RECT 68.165 99.520 68.455 99.565 ;
        RECT 97.590 99.520 97.910 99.580 ;
        RECT 98.140 99.565 98.280 99.720 ;
        RECT 100.365 99.675 100.655 99.905 ;
        RECT 108.190 99.860 108.480 99.905 ;
        RECT 110.050 99.860 110.340 99.905 ;
        RECT 112.830 99.860 113.120 99.905 ;
        RECT 108.190 99.720 113.120 99.860 ;
        RECT 108.190 99.675 108.480 99.720 ;
        RECT 110.050 99.675 110.340 99.720 ;
        RECT 112.830 99.675 113.120 99.720 ;
        RECT 35.950 99.380 36.715 99.520 ;
        RECT 22.625 99.335 22.915 99.380 ;
        RECT 35.950 99.320 36.270 99.380 ;
        RECT 36.425 99.335 36.715 99.380 ;
        RECT 36.960 99.380 97.910 99.520 ;
        RECT 7.890 98.980 8.210 99.240 ;
        RECT 13.010 99.180 13.300 99.225 ;
        RECT 10.765 99.040 13.300 99.180 ;
        RECT 10.765 98.885 10.980 99.040 ;
        RECT 13.010 98.995 13.300 99.040 ;
        RECT 22.150 99.180 22.470 99.240 ;
        RECT 23.545 99.180 23.835 99.225 ;
        RECT 25.845 99.180 26.135 99.225 ;
        RECT 22.150 99.040 26.135 99.180 ;
        RECT 22.150 98.980 22.470 99.040 ;
        RECT 23.545 98.995 23.835 99.040 ;
        RECT 25.845 98.995 26.135 99.040 ;
        RECT 8.830 98.840 9.120 98.885 ;
        RECT 10.690 98.840 10.980 98.885 ;
        RECT 8.830 98.700 10.980 98.840 ;
        RECT 8.830 98.655 9.120 98.700 ;
        RECT 10.690 98.655 10.980 98.700 ;
        RECT 11.610 98.840 11.900 98.885 ;
        RECT 14.870 98.840 15.160 98.885 ;
        RECT 18.470 98.840 18.790 98.900 ;
        RECT 11.610 98.700 18.790 98.840 ;
        RECT 11.610 98.655 11.900 98.700 ;
        RECT 14.870 98.655 15.160 98.700 ;
        RECT 18.470 98.640 18.790 98.700 ;
        RECT 21.690 98.840 22.010 98.900 ;
        RECT 24.925 98.840 25.215 98.885 ;
        RECT 21.690 98.700 25.215 98.840 ;
        RECT 25.920 98.840 26.060 98.995 ;
        RECT 26.290 98.980 26.610 99.240 ;
        RECT 27.670 98.980 27.990 99.240 ;
        RECT 28.130 99.180 28.450 99.240 ;
        RECT 35.505 99.180 35.795 99.225 ;
        RECT 36.960 99.180 37.100 99.380 ;
        RECT 68.165 99.335 68.455 99.380 ;
        RECT 97.590 99.320 97.910 99.380 ;
        RECT 98.065 99.335 98.355 99.565 ;
        RECT 28.130 99.040 37.100 99.180 ;
        RECT 43.770 99.180 44.090 99.240 ;
        RECT 44.705 99.180 44.995 99.225 ;
        RECT 43.770 99.040 44.995 99.180 ;
        RECT 28.130 98.980 28.450 99.040 ;
        RECT 35.505 98.995 35.795 99.040 ;
        RECT 43.770 98.980 44.090 99.040 ;
        RECT 44.705 98.995 44.995 99.040 ;
        RECT 71.385 98.995 71.675 99.225 ;
        RECT 74.605 99.180 74.895 99.225 ;
        RECT 76.890 99.180 77.210 99.240 ;
        RECT 74.605 99.040 77.210 99.180 ;
        RECT 74.605 98.995 74.895 99.040 ;
        RECT 28.220 98.840 28.360 98.980 ;
        RECT 25.920 98.700 28.360 98.840 ;
        RECT 29.510 98.840 29.830 98.900 ;
        RECT 43.860 98.840 44.000 98.980 ;
        RECT 29.510 98.700 44.000 98.840 ;
        RECT 21.690 98.640 22.010 98.700 ;
        RECT 24.925 98.655 25.215 98.700 ;
        RECT 29.510 98.640 29.830 98.700 ;
        RECT 67.230 98.640 67.550 98.900 ;
        RECT 71.460 98.840 71.600 98.995 ;
        RECT 76.890 98.980 77.210 99.040 ;
        RECT 95.290 99.180 95.610 99.240 ;
        RECT 97.145 99.180 97.435 99.225 ;
        RECT 95.290 99.040 97.435 99.180 ;
        RECT 95.290 98.980 95.610 99.040 ;
        RECT 97.145 98.995 97.435 99.040 ;
        RECT 99.905 99.180 100.195 99.225 ;
        RECT 100.440 99.180 100.580 99.675 ;
        RECT 103.125 99.520 103.415 99.565 ;
        RECT 113.230 99.520 113.550 99.580 ;
        RECT 103.125 99.380 113.550 99.520 ;
        RECT 103.125 99.335 103.415 99.380 ;
        RECT 113.230 99.320 113.550 99.380 ;
        RECT 99.905 99.040 100.580 99.180 ;
        RECT 107.725 99.180 108.015 99.225 ;
        RECT 109.090 99.180 109.410 99.240 ;
        RECT 107.725 99.040 109.410 99.180 ;
        RECT 99.905 98.995 100.195 99.040 ;
        RECT 107.725 98.995 108.015 99.040 ;
        RECT 109.090 98.980 109.410 99.040 ;
        RECT 109.550 98.980 109.870 99.240 ;
        RECT 112.830 99.180 113.120 99.225 ;
        RECT 110.585 99.040 113.120 99.180 ;
        RECT 75.050 98.840 75.370 98.900 ;
        RECT 110.585 98.885 110.800 99.040 ;
        RECT 112.830 98.995 113.120 99.040 ;
        RECT 117.370 98.980 117.690 99.240 ;
        RECT 71.460 98.700 75.370 98.840 ;
        RECT 75.050 98.640 75.370 98.700 ;
        RECT 108.650 98.840 108.940 98.885 ;
        RECT 110.510 98.840 110.800 98.885 ;
        RECT 108.650 98.700 110.800 98.840 ;
        RECT 108.650 98.655 108.940 98.700 ;
        RECT 110.510 98.655 110.800 98.700 ;
        RECT 111.430 98.840 111.720 98.885 ;
        RECT 114.150 98.840 114.470 98.900 ;
        RECT 114.690 98.840 114.980 98.885 ;
        RECT 111.430 98.700 114.980 98.840 ;
        RECT 111.430 98.655 111.720 98.700 ;
        RECT 114.150 98.640 114.470 98.700 ;
        RECT 114.690 98.655 114.980 98.700 ;
        RECT 23.990 98.500 24.310 98.560 ;
        RECT 24.465 98.500 24.755 98.545 ;
        RECT 23.990 98.360 24.755 98.500 ;
        RECT 23.990 98.300 24.310 98.360 ;
        RECT 24.465 98.315 24.755 98.360 ;
        RECT 29.050 98.300 29.370 98.560 ;
        RECT 34.570 98.300 34.890 98.560 ;
        RECT 45.150 98.300 45.470 98.560 ;
        RECT 68.150 98.500 68.470 98.560 ;
        RECT 70.925 98.500 71.215 98.545 ;
        RECT 68.150 98.360 71.215 98.500 ;
        RECT 68.150 98.300 68.470 98.360 ;
        RECT 70.925 98.315 71.215 98.360 ;
        RECT 71.830 98.500 72.150 98.560 ;
        RECT 73.685 98.500 73.975 98.545 ;
        RECT 71.830 98.360 73.975 98.500 ;
        RECT 71.830 98.300 72.150 98.360 ;
        RECT 73.685 98.315 73.975 98.360 ;
        RECT 96.225 98.500 96.515 98.545 ;
        RECT 96.670 98.500 96.990 98.560 ;
        RECT 96.225 98.360 96.990 98.500 ;
        RECT 96.225 98.315 96.515 98.360 ;
        RECT 96.670 98.300 96.990 98.360 ;
        RECT 97.130 98.500 97.450 98.560 ;
        RECT 102.205 98.500 102.495 98.545 ;
        RECT 97.130 98.360 102.495 98.500 ;
        RECT 97.130 98.300 97.450 98.360 ;
        RECT 102.205 98.315 102.495 98.360 ;
        RECT 102.650 98.500 102.970 98.560 ;
        RECT 116.695 98.500 116.985 98.545 ;
        RECT 102.650 98.360 116.985 98.500 ;
        RECT 102.650 98.300 102.970 98.360 ;
        RECT 116.695 98.315 116.985 98.360 ;
        RECT 117.830 98.300 118.150 98.560 ;
        RECT 5.520 97.680 123.740 98.160 ;
        RECT 40.105 97.295 40.395 97.525 ;
        RECT 48.830 97.480 49.150 97.540 ;
        RECT 53.445 97.480 53.735 97.525 ;
        RECT 75.510 97.480 75.830 97.540 ;
        RECT 48.830 97.340 53.735 97.480 ;
        RECT 29.510 97.140 29.830 97.200 ;
        RECT 26.380 97.000 37.560 97.140 ;
        RECT 20.770 96.600 21.090 96.860 ;
        RECT 21.705 96.800 21.995 96.845 ;
        RECT 22.150 96.800 22.470 96.860 ;
        RECT 21.705 96.660 22.470 96.800 ;
        RECT 21.705 96.615 21.995 96.660 ;
        RECT 22.150 96.600 22.470 96.660 ;
        RECT 23.070 96.800 23.390 96.860 ;
        RECT 26.380 96.845 26.520 97.000 ;
        RECT 29.510 96.940 29.830 97.000 ;
        RECT 24.005 96.800 24.295 96.845 ;
        RECT 23.070 96.660 24.295 96.800 ;
        RECT 23.070 96.600 23.390 96.660 ;
        RECT 24.005 96.615 24.295 96.660 ;
        RECT 26.305 96.615 26.595 96.845 ;
        RECT 26.765 96.800 27.055 96.845 ;
        RECT 27.210 96.800 27.530 96.860 ;
        RECT 26.765 96.660 27.530 96.800 ;
        RECT 26.765 96.615 27.055 96.660 ;
        RECT 27.210 96.600 27.530 96.660 ;
        RECT 32.730 96.600 33.050 96.860 ;
        RECT 37.420 96.845 37.560 97.000 ;
        RECT 37.345 96.615 37.635 96.845 ;
        RECT 39.185 96.800 39.475 96.845 ;
        RECT 38.800 96.660 39.475 96.800 ;
        RECT 40.180 96.800 40.320 97.295 ;
        RECT 48.830 97.280 49.150 97.340 ;
        RECT 53.445 97.295 53.735 97.340 ;
        RECT 70.080 97.340 75.830 97.480 ;
        RECT 41.490 97.140 41.780 97.185 ;
        RECT 43.350 97.140 43.640 97.185 ;
        RECT 41.490 97.000 43.640 97.140 ;
        RECT 41.490 96.955 41.780 97.000 ;
        RECT 43.350 96.955 43.640 97.000 ;
        RECT 44.270 97.140 44.560 97.185 ;
        RECT 45.150 97.140 45.470 97.200 ;
        RECT 47.530 97.140 47.820 97.185 ;
        RECT 58.490 97.140 58.810 97.200 ;
        RECT 44.270 97.000 47.820 97.140 ;
        RECT 44.270 96.955 44.560 97.000 ;
        RECT 42.405 96.800 42.695 96.845 ;
        RECT 40.180 96.660 42.695 96.800 ;
        RECT 43.425 96.800 43.640 96.955 ;
        RECT 45.150 96.940 45.470 97.000 ;
        RECT 47.530 96.955 47.820 97.000 ;
        RECT 54.440 97.000 58.810 97.140 ;
        RECT 54.440 96.845 54.580 97.000 ;
        RECT 58.490 96.940 58.810 97.000 ;
        RECT 61.270 97.140 61.560 97.185 ;
        RECT 63.130 97.140 63.420 97.185 ;
        RECT 61.270 97.000 63.420 97.140 ;
        RECT 61.270 96.955 61.560 97.000 ;
        RECT 63.130 96.955 63.420 97.000 ;
        RECT 64.050 97.140 64.340 97.185 ;
        RECT 67.310 97.140 67.600 97.185 ;
        RECT 68.150 97.140 68.470 97.200 ;
        RECT 64.050 97.000 68.470 97.140 ;
        RECT 64.050 96.955 64.340 97.000 ;
        RECT 67.310 96.955 67.600 97.000 ;
        RECT 45.670 96.800 45.960 96.845 ;
        RECT 43.425 96.660 45.960 96.800 ;
        RECT 19.850 96.460 20.170 96.520 ;
        RECT 22.625 96.460 22.915 96.505 ;
        RECT 19.850 96.320 22.915 96.460 ;
        RECT 19.850 96.260 20.170 96.320 ;
        RECT 22.625 96.275 22.915 96.320 ;
        RECT 23.085 95.780 23.375 95.825 ;
        RECT 23.530 95.780 23.850 95.840 ;
        RECT 23.085 95.640 23.850 95.780 ;
        RECT 23.085 95.595 23.375 95.640 ;
        RECT 23.530 95.580 23.850 95.640 ;
        RECT 33.190 95.780 33.510 95.840 ;
        RECT 33.665 95.780 33.955 95.825 ;
        RECT 33.190 95.640 33.955 95.780 ;
        RECT 33.190 95.580 33.510 95.640 ;
        RECT 33.665 95.595 33.955 95.640 ;
        RECT 36.870 95.580 37.190 95.840 ;
        RECT 38.800 95.780 38.940 96.660 ;
        RECT 39.185 96.615 39.475 96.660 ;
        RECT 42.405 96.615 42.695 96.660 ;
        RECT 45.670 96.615 45.960 96.660 ;
        RECT 54.365 96.615 54.655 96.845 ;
        RECT 54.810 96.600 55.130 96.860 ;
        RECT 55.730 96.600 56.050 96.860 ;
        RECT 56.650 96.800 56.970 96.860 ;
        RECT 60.345 96.800 60.635 96.845 ;
        RECT 56.650 96.660 60.635 96.800 ;
        RECT 63.205 96.800 63.420 96.955 ;
        RECT 68.150 96.940 68.470 97.000 ;
        RECT 70.080 96.845 70.220 97.340 ;
        RECT 75.510 97.280 75.830 97.340 ;
        RECT 111.405 97.480 111.695 97.525 ;
        RECT 111.405 97.340 112.540 97.480 ;
        RECT 111.405 97.295 111.695 97.340 ;
        RECT 70.930 97.140 71.220 97.185 ;
        RECT 72.790 97.140 73.080 97.185 ;
        RECT 70.930 97.000 73.080 97.140 ;
        RECT 70.930 96.955 71.220 97.000 ;
        RECT 72.790 96.955 73.080 97.000 ;
        RECT 73.710 97.140 74.000 97.185 ;
        RECT 74.590 97.140 74.910 97.200 ;
        RECT 76.970 97.140 77.260 97.185 ;
        RECT 73.710 97.000 77.260 97.140 ;
        RECT 73.710 96.955 74.000 97.000 ;
        RECT 65.450 96.800 65.740 96.845 ;
        RECT 63.205 96.660 65.740 96.800 ;
        RECT 56.650 96.600 56.970 96.660 ;
        RECT 60.345 96.615 60.635 96.660 ;
        RECT 65.450 96.615 65.740 96.660 ;
        RECT 70.005 96.615 70.295 96.845 ;
        RECT 71.830 96.600 72.150 96.860 ;
        RECT 72.865 96.800 73.080 96.955 ;
        RECT 74.590 96.940 74.910 97.000 ;
        RECT 76.970 96.955 77.260 97.000 ;
        RECT 97.590 97.140 97.910 97.200 ;
        RECT 102.190 97.140 102.510 97.200 ;
        RECT 97.590 97.000 102.510 97.140 ;
        RECT 97.590 96.940 97.910 97.000 ;
        RECT 75.110 96.800 75.400 96.845 ;
        RECT 72.865 96.660 75.400 96.800 ;
        RECT 75.110 96.615 75.400 96.660 ;
        RECT 97.130 96.800 97.450 96.860 ;
        RECT 100.440 96.845 100.580 97.000 ;
        RECT 102.190 96.940 102.510 97.000 ;
        RECT 109.090 97.140 109.410 97.200 ;
        RECT 109.090 97.000 112.080 97.140 ;
        RECT 109.090 96.940 109.410 97.000 ;
        RECT 99.445 96.800 99.735 96.845 ;
        RECT 97.130 96.660 99.735 96.800 ;
        RECT 97.130 96.600 97.450 96.660 ;
        RECT 99.445 96.615 99.735 96.660 ;
        RECT 100.365 96.615 100.655 96.845 ;
        RECT 101.285 96.800 101.575 96.845 ;
        RECT 101.730 96.800 102.050 96.860 ;
        RECT 109.550 96.800 109.870 96.860 ;
        RECT 101.285 96.660 102.050 96.800 ;
        RECT 101.285 96.615 101.575 96.660 ;
        RECT 101.730 96.600 102.050 96.660 ;
        RECT 109.180 96.660 109.870 96.800 ;
        RECT 40.565 96.275 40.855 96.505 ;
        RECT 39.170 96.120 39.490 96.180 ;
        RECT 40.640 96.120 40.780 96.275 ;
        RECT 62.170 96.260 62.490 96.520 ;
        RECT 109.180 96.165 109.320 96.660 ;
        RECT 109.550 96.600 109.870 96.660 ;
        RECT 110.010 96.600 110.330 96.860 ;
        RECT 110.470 96.600 110.790 96.860 ;
        RECT 111.940 96.845 112.080 97.000 ;
        RECT 111.865 96.615 112.155 96.845 ;
        RECT 112.400 96.800 112.540 97.340 ;
        RECT 112.790 97.140 113.080 97.185 ;
        RECT 114.650 97.140 114.940 97.185 ;
        RECT 112.790 97.000 114.940 97.140 ;
        RECT 112.790 96.955 113.080 97.000 ;
        RECT 114.650 96.955 114.940 97.000 ;
        RECT 115.570 97.140 115.860 97.185 ;
        RECT 117.830 97.140 118.150 97.200 ;
        RECT 118.830 97.140 119.120 97.185 ;
        RECT 115.570 97.000 119.120 97.140 ;
        RECT 115.570 96.955 115.860 97.000 ;
        RECT 113.705 96.800 113.995 96.845 ;
        RECT 112.400 96.660 113.995 96.800 ;
        RECT 114.725 96.800 114.940 96.955 ;
        RECT 117.830 96.940 118.150 97.000 ;
        RECT 118.830 96.955 119.120 97.000 ;
        RECT 116.970 96.800 117.260 96.845 ;
        RECT 120.835 96.800 121.125 96.845 ;
        RECT 114.725 96.660 117.260 96.800 ;
        RECT 113.705 96.615 113.995 96.660 ;
        RECT 116.970 96.615 117.260 96.660 ;
        RECT 117.460 96.660 121.125 96.800 ;
        RECT 117.460 96.460 117.600 96.660 ;
        RECT 120.835 96.615 121.125 96.660 ;
        RECT 111.940 96.320 117.600 96.460 ;
        RECT 111.940 96.180 112.080 96.320 ;
        RECT 39.170 95.980 40.780 96.120 ;
        RECT 41.030 96.120 41.320 96.165 ;
        RECT 42.890 96.120 43.180 96.165 ;
        RECT 45.670 96.120 45.960 96.165 ;
        RECT 41.030 95.980 45.960 96.120 ;
        RECT 39.170 95.920 39.490 95.980 ;
        RECT 41.030 95.935 41.320 95.980 ;
        RECT 42.890 95.935 43.180 95.980 ;
        RECT 45.670 95.935 45.960 95.980 ;
        RECT 60.810 96.120 61.100 96.165 ;
        RECT 62.670 96.120 62.960 96.165 ;
        RECT 65.450 96.120 65.740 96.165 ;
        RECT 60.810 95.980 65.740 96.120 ;
        RECT 60.810 95.935 61.100 95.980 ;
        RECT 62.670 95.935 62.960 95.980 ;
        RECT 65.450 95.935 65.740 95.980 ;
        RECT 70.470 96.120 70.760 96.165 ;
        RECT 72.330 96.120 72.620 96.165 ;
        RECT 75.110 96.120 75.400 96.165 ;
        RECT 70.470 95.980 75.400 96.120 ;
        RECT 70.470 95.935 70.760 95.980 ;
        RECT 72.330 95.935 72.620 95.980 ;
        RECT 75.110 95.935 75.400 95.980 ;
        RECT 109.105 95.935 109.395 96.165 ;
        RECT 111.850 95.920 112.170 96.180 ;
        RECT 112.330 96.120 112.620 96.165 ;
        RECT 114.190 96.120 114.480 96.165 ;
        RECT 116.970 96.120 117.260 96.165 ;
        RECT 112.330 95.980 117.260 96.120 ;
        RECT 112.330 95.935 112.620 95.980 ;
        RECT 114.190 95.935 114.480 95.980 ;
        RECT 116.970 95.935 117.260 95.980 ;
        RECT 44.690 95.780 45.010 95.840 ;
        RECT 38.800 95.640 45.010 95.780 ;
        RECT 44.690 95.580 45.010 95.640 ;
        RECT 47.450 95.780 47.770 95.840 ;
        RECT 49.535 95.780 49.825 95.825 ;
        RECT 47.450 95.640 49.825 95.780 ;
        RECT 47.450 95.580 47.770 95.640 ;
        RECT 49.535 95.595 49.825 95.640 ;
        RECT 55.745 95.780 56.035 95.825 ;
        RECT 57.570 95.780 57.890 95.840 ;
        RECT 55.745 95.640 57.890 95.780 ;
        RECT 55.745 95.595 56.035 95.640 ;
        RECT 57.570 95.580 57.890 95.640 ;
        RECT 64.930 95.780 65.250 95.840 ;
        RECT 69.315 95.780 69.605 95.825 ;
        RECT 72.750 95.780 73.070 95.840 ;
        RECT 79.190 95.825 79.510 95.840 ;
        RECT 64.930 95.640 73.070 95.780 ;
        RECT 64.930 95.580 65.250 95.640 ;
        RECT 69.315 95.595 69.605 95.640 ;
        RECT 72.750 95.580 73.070 95.640 ;
        RECT 78.975 95.595 79.510 95.825 ;
        RECT 79.190 95.580 79.510 95.595 ;
        RECT 5.520 94.960 123.740 95.440 ;
        RECT 30.675 94.760 30.965 94.805 ;
        RECT 32.270 94.760 32.590 94.820 ;
        RECT 30.675 94.620 32.590 94.760 ;
        RECT 30.675 94.575 30.965 94.620 ;
        RECT 32.270 94.560 32.590 94.620 ;
        RECT 44.690 94.560 45.010 94.820 ;
        RECT 54.365 94.760 54.655 94.805 ;
        RECT 55.730 94.760 56.050 94.820 ;
        RECT 54.365 94.620 56.050 94.760 ;
        RECT 54.365 94.575 54.655 94.620 ;
        RECT 55.730 94.560 56.050 94.620 ;
        RECT 62.170 94.760 62.490 94.820 ;
        RECT 67.705 94.760 67.995 94.805 ;
        RECT 62.170 94.620 67.995 94.760 ;
        RECT 62.170 94.560 62.490 94.620 ;
        RECT 67.705 94.575 67.995 94.620 ;
        RECT 74.590 94.760 74.910 94.820 ;
        RECT 75.065 94.760 75.355 94.805 ;
        RECT 74.590 94.620 75.355 94.760 ;
        RECT 74.590 94.560 74.910 94.620 ;
        RECT 75.065 94.575 75.355 94.620 ;
        RECT 76.890 94.560 77.210 94.820 ;
        RECT 86.105 94.760 86.395 94.805 ;
        RECT 91.150 94.760 91.470 94.820 ;
        RECT 92.545 94.760 92.835 94.805 ;
        RECT 86.105 94.620 90.920 94.760 ;
        RECT 86.105 94.575 86.395 94.620 ;
        RECT 22.170 94.420 22.460 94.465 ;
        RECT 24.030 94.420 24.320 94.465 ;
        RECT 26.810 94.420 27.100 94.465 ;
        RECT 22.170 94.280 27.100 94.420 ;
        RECT 22.170 94.235 22.460 94.280 ;
        RECT 24.030 94.235 24.320 94.280 ;
        RECT 26.810 94.235 27.100 94.280 ;
        RECT 31.830 94.420 32.120 94.465 ;
        RECT 33.690 94.420 33.980 94.465 ;
        RECT 36.470 94.420 36.760 94.465 ;
        RECT 31.830 94.280 36.760 94.420 ;
        RECT 31.830 94.235 32.120 94.280 ;
        RECT 33.690 94.235 33.980 94.280 ;
        RECT 36.470 94.235 36.760 94.280 ;
        RECT 57.130 94.420 57.420 94.465 ;
        RECT 58.990 94.420 59.280 94.465 ;
        RECT 61.770 94.420 62.060 94.465 ;
        RECT 57.130 94.280 62.060 94.420 ;
        RECT 57.130 94.235 57.420 94.280 ;
        RECT 58.990 94.235 59.280 94.280 ;
        RECT 61.770 94.235 62.060 94.280 ;
        RECT 66.325 94.235 66.615 94.465 ;
        RECT 70.465 94.235 70.755 94.465 ;
        RECT 84.250 94.420 84.570 94.480 ;
        RECT 84.250 94.280 88.160 94.420 ;
        RECT 20.310 94.080 20.630 94.140 ;
        RECT 21.705 94.080 21.995 94.125 ;
        RECT 31.350 94.080 31.670 94.140 ;
        RECT 20.310 93.940 31.670 94.080 ;
        RECT 20.310 93.880 20.630 93.940 ;
        RECT 21.705 93.895 21.995 93.940 ;
        RECT 31.350 93.880 31.670 93.940 ;
        RECT 33.190 93.880 33.510 94.140 ;
        RECT 46.070 94.080 46.390 94.140 ;
        RECT 47.465 94.080 47.755 94.125 ;
        RECT 46.070 93.940 47.755 94.080 ;
        RECT 46.070 93.880 46.390 93.940 ;
        RECT 47.465 93.895 47.755 93.940 ;
        RECT 56.650 93.880 56.970 94.140 ;
        RECT 58.505 94.080 58.795 94.125 ;
        RECT 66.400 94.080 66.540 94.235 ;
        RECT 58.505 93.940 66.540 94.080 ;
        RECT 58.505 93.895 58.795 93.940 ;
        RECT 23.530 93.540 23.850 93.800 ;
        RECT 26.810 93.740 27.100 93.785 ;
        RECT 36.470 93.740 36.760 93.785 ;
        RECT 24.565 93.600 27.100 93.740 ;
        RECT 24.565 93.445 24.780 93.600 ;
        RECT 26.810 93.555 27.100 93.600 ;
        RECT 34.225 93.600 36.760 93.740 ;
        RECT 22.630 93.400 22.920 93.445 ;
        RECT 24.490 93.400 24.780 93.445 ;
        RECT 22.630 93.260 24.780 93.400 ;
        RECT 22.630 93.215 22.920 93.260 ;
        RECT 24.490 93.215 24.780 93.260 ;
        RECT 25.410 93.400 25.700 93.445 ;
        RECT 27.210 93.400 27.530 93.460 ;
        RECT 34.225 93.445 34.440 93.600 ;
        RECT 36.470 93.555 36.760 93.600 ;
        RECT 50.210 93.740 50.530 93.800 ;
        RECT 51.145 93.740 51.435 93.785 ;
        RECT 50.210 93.600 51.435 93.740 ;
        RECT 50.210 93.540 50.530 93.600 ;
        RECT 51.145 93.555 51.435 93.600 ;
        RECT 52.065 93.555 52.355 93.785 ;
        RECT 28.670 93.400 28.960 93.445 ;
        RECT 25.410 93.260 28.960 93.400 ;
        RECT 25.410 93.215 25.700 93.260 ;
        RECT 27.210 93.200 27.530 93.260 ;
        RECT 28.670 93.215 28.960 93.260 ;
        RECT 32.290 93.400 32.580 93.445 ;
        RECT 34.150 93.400 34.440 93.445 ;
        RECT 32.290 93.260 34.440 93.400 ;
        RECT 32.290 93.215 32.580 93.260 ;
        RECT 34.150 93.215 34.440 93.260 ;
        RECT 35.070 93.400 35.360 93.445 ;
        RECT 36.870 93.400 37.190 93.460 ;
        RECT 38.330 93.400 38.620 93.445 ;
        RECT 52.140 93.400 52.280 93.555 ;
        RECT 52.510 93.540 52.830 93.800 ;
        RECT 52.970 93.540 53.290 93.800 ;
        RECT 61.770 93.740 62.060 93.785 ;
        RECT 59.525 93.600 62.060 93.740 ;
        RECT 59.525 93.445 59.740 93.600 ;
        RECT 61.770 93.555 62.060 93.600 ;
        RECT 66.770 93.740 67.090 93.800 ;
        RECT 67.245 93.740 67.535 93.785 ;
        RECT 66.770 93.600 67.535 93.740 ;
        RECT 66.770 93.540 67.090 93.600 ;
        RECT 67.245 93.555 67.535 93.600 ;
        RECT 68.625 93.740 68.915 93.785 ;
        RECT 70.540 93.740 70.680 94.235 ;
        RECT 84.250 94.220 84.570 94.280 ;
        RECT 72.750 93.880 73.070 94.140 ;
        RECT 73.225 94.080 73.515 94.125 ;
        RECT 79.665 94.080 79.955 94.125 ;
        RECT 73.225 93.940 79.955 94.080 ;
        RECT 73.225 93.895 73.515 93.940 ;
        RECT 79.665 93.895 79.955 93.940 ;
        RECT 82.960 93.940 85.400 94.080 ;
        RECT 68.625 93.600 70.680 93.740 ;
        RECT 71.830 93.740 72.150 93.800 ;
        RECT 73.300 93.740 73.440 93.895 ;
        RECT 71.830 93.600 73.440 93.740 ;
        RECT 74.605 93.740 74.895 93.785 ;
        RECT 75.050 93.740 75.370 93.800 ;
        RECT 74.605 93.600 75.370 93.740 ;
        RECT 68.625 93.555 68.915 93.600 ;
        RECT 71.830 93.540 72.150 93.600 ;
        RECT 74.605 93.555 74.895 93.600 ;
        RECT 75.050 93.540 75.370 93.600 ;
        RECT 78.730 93.740 79.050 93.800 ;
        RECT 82.960 93.785 83.100 93.940 ;
        RECT 82.885 93.740 83.175 93.785 ;
        RECT 78.730 93.600 83.175 93.740 ;
        RECT 78.730 93.540 79.050 93.600 ;
        RECT 82.885 93.555 83.175 93.600 ;
        RECT 83.805 93.555 84.095 93.785 ;
        RECT 35.070 93.260 38.620 93.400 ;
        RECT 35.070 93.215 35.360 93.260 ;
        RECT 36.870 93.200 37.190 93.260 ;
        RECT 38.330 93.215 38.620 93.260 ;
        RECT 47.540 93.260 52.280 93.400 ;
        RECT 57.590 93.400 57.880 93.445 ;
        RECT 59.450 93.400 59.740 93.445 ;
        RECT 57.590 93.260 59.740 93.400 ;
        RECT 47.540 93.120 47.680 93.260 ;
        RECT 57.590 93.215 57.880 93.260 ;
        RECT 59.450 93.215 59.740 93.260 ;
        RECT 60.370 93.400 60.660 93.445 ;
        RECT 61.250 93.400 61.570 93.460 ;
        RECT 63.630 93.400 63.920 93.445 ;
        RECT 60.370 93.260 63.920 93.400 ;
        RECT 60.370 93.215 60.660 93.260 ;
        RECT 61.250 93.200 61.570 93.260 ;
        RECT 63.630 93.215 63.920 93.260 ;
        RECT 72.305 93.400 72.595 93.445 ;
        RECT 79.190 93.400 79.510 93.460 ;
        RECT 83.880 93.400 84.020 93.555 ;
        RECT 84.250 93.540 84.570 93.800 ;
        RECT 84.725 93.555 85.015 93.785 ;
        RECT 85.260 93.740 85.400 93.940 ;
        RECT 86.550 93.740 86.870 93.800 ;
        RECT 88.020 93.785 88.160 94.280 ;
        RECT 90.780 94.080 90.920 94.620 ;
        RECT 91.150 94.620 92.835 94.760 ;
        RECT 91.150 94.560 91.470 94.620 ;
        RECT 92.545 94.575 92.835 94.620 ;
        RECT 94.370 94.560 94.690 94.820 ;
        RECT 96.670 94.560 96.990 94.820 ;
        RECT 98.510 94.560 98.830 94.820 ;
        RECT 110.470 94.760 110.790 94.820 ;
        RECT 112.785 94.760 113.075 94.805 ;
        RECT 110.470 94.620 113.075 94.760 ;
        RECT 110.470 94.560 110.790 94.620 ;
        RECT 112.785 94.575 113.075 94.620 ;
        RECT 113.230 94.420 113.550 94.480 ;
        RECT 113.230 94.280 115.760 94.420 ;
        RECT 113.230 94.220 113.550 94.280 ;
        RECT 97.145 94.080 97.435 94.125 ;
        RECT 98.970 94.080 99.290 94.140 ;
        RECT 90.780 93.940 96.440 94.080 ;
        RECT 88.390 93.785 88.710 93.800 ;
        RECT 87.485 93.740 87.775 93.785 ;
        RECT 85.260 93.600 86.870 93.740 ;
        RECT 72.305 93.260 84.020 93.400 ;
        RECT 84.800 93.400 84.940 93.555 ;
        RECT 86.550 93.540 86.870 93.600 ;
        RECT 87.100 93.600 87.775 93.740 ;
        RECT 86.090 93.400 86.410 93.460 ;
        RECT 84.800 93.260 86.410 93.400 ;
        RECT 72.305 93.215 72.595 93.260 ;
        RECT 79.190 93.200 79.510 93.260 ;
        RECT 86.090 93.200 86.410 93.260 ;
        RECT 39.630 93.060 39.950 93.120 ;
        RECT 40.335 93.060 40.625 93.105 ;
        RECT 46.530 93.060 46.850 93.120 ;
        RECT 39.630 92.920 46.850 93.060 ;
        RECT 39.630 92.860 39.950 92.920 ;
        RECT 40.335 92.875 40.625 92.920 ;
        RECT 46.530 92.860 46.850 92.920 ;
        RECT 47.005 93.060 47.295 93.105 ;
        RECT 47.450 93.060 47.770 93.120 ;
        RECT 47.005 92.920 47.770 93.060 ;
        RECT 47.005 92.875 47.295 92.920 ;
        RECT 47.450 92.860 47.770 92.920 ;
        RECT 64.470 93.060 64.790 93.120 ;
        RECT 65.635 93.060 65.925 93.105 ;
        RECT 64.470 92.920 65.925 93.060 ;
        RECT 64.470 92.860 64.790 92.920 ;
        RECT 65.635 92.875 65.925 92.920 ;
        RECT 78.745 93.060 79.035 93.105 ;
        RECT 83.790 93.060 84.110 93.120 ;
        RECT 87.100 93.060 87.240 93.600 ;
        RECT 87.485 93.555 87.775 93.600 ;
        RECT 87.945 93.555 88.235 93.785 ;
        RECT 88.390 93.555 88.795 93.785 ;
        RECT 88.390 93.540 88.710 93.555 ;
        RECT 93.450 93.540 93.770 93.800 ;
        RECT 93.925 93.740 94.215 93.785 ;
        RECT 94.370 93.740 94.690 93.800 ;
        RECT 96.300 93.785 96.440 93.940 ;
        RECT 97.145 93.940 99.290 94.080 ;
        RECT 97.145 93.895 97.435 93.940 ;
        RECT 98.970 93.880 99.290 93.940 ;
        RECT 100.825 94.080 101.115 94.125 ;
        RECT 102.650 94.080 102.970 94.140 ;
        RECT 100.825 93.940 102.970 94.080 ;
        RECT 100.825 93.895 101.115 93.940 ;
        RECT 102.650 93.880 102.970 93.940 ;
        RECT 104.965 94.080 105.255 94.125 ;
        RECT 111.850 94.080 112.170 94.140 ;
        RECT 115.620 94.125 115.760 94.280 ;
        RECT 104.965 93.940 114.840 94.080 ;
        RECT 104.965 93.895 105.255 93.940 ;
        RECT 111.850 93.880 112.170 93.940 ;
        RECT 93.925 93.600 94.690 93.740 ;
        RECT 93.925 93.555 94.215 93.600 ;
        RECT 94.370 93.540 94.690 93.600 ;
        RECT 96.225 93.555 96.515 93.785 ;
        RECT 97.605 93.555 97.895 93.785 ;
        RECT 101.745 93.740 102.035 93.785 ;
        RECT 102.190 93.740 102.510 93.800 ;
        RECT 114.700 93.785 114.840 93.940 ;
        RECT 115.545 93.895 115.835 94.125 ;
        RECT 104.045 93.740 104.335 93.785 ;
        RECT 106.345 93.740 106.635 93.785 ;
        RECT 101.745 93.600 106.635 93.740 ;
        RECT 101.745 93.555 102.035 93.600 ;
        RECT 89.785 93.400 90.075 93.445 ;
        RECT 94.845 93.400 95.135 93.445 ;
        RECT 89.785 93.260 95.135 93.400 ;
        RECT 89.785 93.215 90.075 93.260 ;
        RECT 94.845 93.215 95.135 93.260 ;
        RECT 95.750 93.400 96.070 93.460 ;
        RECT 97.680 93.400 97.820 93.555 ;
        RECT 102.190 93.540 102.510 93.600 ;
        RECT 104.045 93.555 104.335 93.600 ;
        RECT 106.345 93.555 106.635 93.600 ;
        RECT 107.265 93.740 107.555 93.785 ;
        RECT 107.265 93.600 113.920 93.740 ;
        RECT 107.265 93.555 107.555 93.600 ;
        RECT 113.780 93.460 113.920 93.600 ;
        RECT 114.625 93.555 114.915 93.785 ;
        RECT 95.750 93.260 97.820 93.400 ;
        RECT 113.690 93.400 114.010 93.460 ;
        RECT 115.085 93.400 115.375 93.445 ;
        RECT 113.690 93.260 115.375 93.400 ;
        RECT 95.750 93.200 96.070 93.260 ;
        RECT 113.690 93.200 114.010 93.260 ;
        RECT 115.085 93.215 115.375 93.260 ;
        RECT 78.745 92.920 87.240 93.060 ;
        RECT 78.745 92.875 79.035 92.920 ;
        RECT 83.790 92.860 84.110 92.920 ;
        RECT 102.650 92.860 102.970 93.120 ;
        RECT 103.125 93.060 103.415 93.105 ;
        RECT 103.570 93.060 103.890 93.120 ;
        RECT 103.125 92.920 103.890 93.060 ;
        RECT 103.125 92.875 103.415 92.920 ;
        RECT 103.570 92.860 103.890 92.920 ;
        RECT 104.030 93.060 104.350 93.120 ;
        RECT 105.425 93.060 105.715 93.105 ;
        RECT 104.030 92.920 105.715 93.060 ;
        RECT 104.030 92.860 104.350 92.920 ;
        RECT 105.425 92.875 105.715 92.920 ;
        RECT 5.520 92.240 123.740 92.720 ;
        RECT 14.345 92.040 14.635 92.085 ;
        RECT 13.730 91.900 14.635 92.040 ;
        RECT 12.505 91.360 12.795 91.405 ;
        RECT 13.730 91.360 13.870 91.900 ;
        RECT 14.345 91.855 14.635 91.900 ;
        RECT 23.070 92.040 23.390 92.100 ;
        RECT 23.545 92.040 23.835 92.085 ;
        RECT 23.070 91.900 23.835 92.040 ;
        RECT 23.070 91.840 23.390 91.900 ;
        RECT 23.545 91.855 23.835 91.900 ;
        RECT 32.730 91.840 33.050 92.100 ;
        RECT 35.045 92.040 35.335 92.085 ;
        RECT 39.630 92.040 39.950 92.100 ;
        RECT 35.045 91.900 39.950 92.040 ;
        RECT 35.045 91.855 35.335 91.900 ;
        RECT 39.630 91.840 39.950 91.900 ;
        RECT 40.105 92.040 40.395 92.085 ;
        RECT 46.530 92.040 46.850 92.100 ;
        RECT 61.250 92.040 61.570 92.100 ;
        RECT 61.725 92.040 62.015 92.085 ;
        RECT 40.105 91.900 41.240 92.040 ;
        RECT 40.105 91.855 40.395 91.900 ;
        RECT 25.845 91.700 26.135 91.745 ;
        RECT 32.270 91.700 32.590 91.760 ;
        RECT 34.585 91.700 34.875 91.745 ;
        RECT 25.845 91.560 34.875 91.700 ;
        RECT 25.845 91.515 26.135 91.560 ;
        RECT 32.270 91.500 32.590 91.560 ;
        RECT 34.585 91.515 34.875 91.560 ;
        RECT 38.710 91.700 39.030 91.760 ;
        RECT 38.710 91.560 40.780 91.700 ;
        RECT 38.710 91.500 39.030 91.560 ;
        RECT 12.505 91.220 13.870 91.360 ;
        RECT 12.505 91.175 12.795 91.220 ;
        RECT 16.170 91.160 16.490 91.420 ;
        RECT 25.385 91.360 25.675 91.405 ;
        RECT 16.720 91.220 25.675 91.360 ;
        RECT 16.720 91.080 16.860 91.220 ;
        RECT 25.385 91.175 25.675 91.220 ;
        RECT 39.185 91.360 39.475 91.405 ;
        RECT 40.090 91.360 40.410 91.420 ;
        RECT 40.640 91.405 40.780 91.560 ;
        RECT 39.185 91.220 40.410 91.360 ;
        RECT 39.185 91.175 39.475 91.220 ;
        RECT 40.090 91.160 40.410 91.220 ;
        RECT 40.565 91.175 40.855 91.405 ;
        RECT 41.100 91.360 41.240 91.900 ;
        RECT 46.530 91.900 50.900 92.040 ;
        RECT 46.530 91.840 46.850 91.900 ;
        RECT 44.230 91.745 44.550 91.760 ;
        RECT 41.490 91.700 41.780 91.745 ;
        RECT 43.350 91.700 43.640 91.745 ;
        RECT 41.490 91.560 43.640 91.700 ;
        RECT 41.490 91.515 41.780 91.560 ;
        RECT 43.350 91.515 43.640 91.560 ;
        RECT 42.405 91.360 42.695 91.405 ;
        RECT 41.100 91.220 42.695 91.360 ;
        RECT 43.425 91.360 43.640 91.515 ;
        RECT 44.230 91.700 44.560 91.745 ;
        RECT 47.530 91.700 47.820 91.745 ;
        RECT 44.230 91.560 47.820 91.700 ;
        RECT 44.230 91.515 44.560 91.560 ;
        RECT 47.530 91.515 47.820 91.560 ;
        RECT 44.230 91.500 44.550 91.515 ;
        RECT 45.670 91.360 45.960 91.405 ;
        RECT 43.425 91.220 45.960 91.360 ;
        RECT 42.405 91.175 42.695 91.220 ;
        RECT 45.670 91.175 45.960 91.220 ;
        RECT 50.210 91.160 50.530 91.420 ;
        RECT 50.760 91.390 50.900 91.900 ;
        RECT 61.250 91.900 62.015 92.040 ;
        RECT 61.250 91.840 61.570 91.900 ;
        RECT 61.725 91.855 62.015 91.900 ;
        RECT 64.930 91.840 65.250 92.100 ;
        RECT 66.770 91.840 67.090 92.100 ;
        RECT 83.345 91.855 83.635 92.085 ;
        RECT 83.790 92.040 84.110 92.100 ;
        RECT 85.630 92.040 85.950 92.100 ;
        RECT 83.790 91.900 85.950 92.040 ;
        RECT 53.445 91.700 53.735 91.745 ;
        RECT 53.905 91.700 54.195 91.745 ;
        RECT 75.050 91.700 75.370 91.760 ;
        RECT 53.445 91.560 54.195 91.700 ;
        RECT 53.445 91.515 53.735 91.560 ;
        RECT 53.905 91.515 54.195 91.560 ;
        RECT 62.030 91.560 75.370 91.700 ;
        RECT 51.040 91.390 51.330 91.435 ;
        RECT 50.760 91.250 51.330 91.390 ;
        RECT 51.040 91.205 51.330 91.250 ;
        RECT 51.605 91.175 51.895 91.405 ;
        RECT 52.065 91.350 52.355 91.405 ;
        RECT 54.350 91.360 54.670 91.420 ;
        RECT 55.285 91.360 55.575 91.405 ;
        RECT 52.065 91.175 52.380 91.350 ;
        RECT 16.630 90.820 16.950 91.080 ;
        RECT 17.565 91.020 17.855 91.065 ;
        RECT 20.310 91.020 20.630 91.080 ;
        RECT 26.765 91.020 27.055 91.065 ;
        RECT 35.965 91.020 36.255 91.065 ;
        RECT 46.070 91.020 46.390 91.080 ;
        RECT 17.565 90.880 46.390 91.020 ;
        RECT 17.565 90.835 17.855 90.880 ;
        RECT 20.310 90.820 20.630 90.880 ;
        RECT 26.765 90.835 27.055 90.880 ;
        RECT 35.965 90.835 36.255 90.880 ;
        RECT 46.070 90.820 46.390 90.880 ;
        RECT 41.030 90.680 41.320 90.725 ;
        RECT 42.890 90.680 43.180 90.725 ;
        RECT 45.670 90.680 45.960 90.725 ;
        RECT 41.030 90.540 45.960 90.680 ;
        RECT 41.030 90.495 41.320 90.540 ;
        RECT 42.890 90.495 43.180 90.540 ;
        RECT 45.670 90.495 45.960 90.540 ;
        RECT 46.990 90.680 47.310 90.740 ;
        RECT 51.680 90.680 51.820 91.175 ;
        RECT 52.240 91.020 52.380 91.175 ;
        RECT 54.350 91.220 55.575 91.360 ;
        RECT 54.350 91.160 54.670 91.220 ;
        RECT 55.285 91.175 55.575 91.220 ;
        RECT 61.250 91.360 61.570 91.420 ;
        RECT 62.030 91.360 62.170 91.560 ;
        RECT 75.050 91.500 75.370 91.560 ;
        RECT 61.250 91.220 62.170 91.360 ;
        RECT 81.505 91.360 81.795 91.405 ;
        RECT 83.420 91.360 83.560 91.855 ;
        RECT 83.790 91.840 84.110 91.900 ;
        RECT 85.630 91.840 85.950 91.900 ;
        RECT 87.010 92.040 87.330 92.100 ;
        RECT 88.390 92.040 88.710 92.100 ;
        RECT 92.530 92.040 92.850 92.100 ;
        RECT 93.465 92.040 93.755 92.085 ;
        RECT 87.010 91.900 89.540 92.040 ;
        RECT 87.010 91.840 87.330 91.900 ;
        RECT 88.390 91.840 88.710 91.900 ;
        RECT 85.260 91.560 88.620 91.700 ;
        RECT 81.505 91.220 83.560 91.360 ;
        RECT 83.790 91.360 84.110 91.420 ;
        RECT 85.260 91.405 85.400 91.560 ;
        RECT 85.185 91.360 85.475 91.405 ;
        RECT 83.790 91.220 85.475 91.360 ;
        RECT 61.250 91.160 61.570 91.220 ;
        RECT 81.505 91.175 81.795 91.220 ;
        RECT 83.790 91.160 84.110 91.220 ;
        RECT 85.185 91.175 85.475 91.220 ;
        RECT 86.090 91.360 86.410 91.420 ;
        RECT 88.480 91.405 88.620 91.560 ;
        RECT 89.400 91.405 89.540 91.900 ;
        RECT 92.530 91.900 93.755 92.040 ;
        RECT 92.530 91.840 92.850 91.900 ;
        RECT 93.465 91.855 93.755 91.900 ;
        RECT 90.705 91.700 90.995 91.745 ;
        RECT 91.165 91.700 91.455 91.745 ;
        RECT 90.705 91.560 91.455 91.700 ;
        RECT 90.705 91.515 90.995 91.560 ;
        RECT 91.165 91.515 91.455 91.560 ;
        RECT 87.485 91.360 87.775 91.405 ;
        RECT 86.090 91.220 87.775 91.360 ;
        RECT 86.090 91.160 86.410 91.220 ;
        RECT 87.485 91.175 87.775 91.220 ;
        RECT 88.405 91.175 88.695 91.405 ;
        RECT 88.865 91.175 89.155 91.405 ;
        RECT 89.325 91.175 89.615 91.405 ;
        RECT 92.545 91.360 92.835 91.405 ;
        RECT 97.590 91.360 97.910 91.420 ;
        RECT 92.545 91.220 97.910 91.360 ;
        RECT 92.545 91.175 92.835 91.220 ;
        RECT 52.970 91.020 53.290 91.080 ;
        RECT 52.240 90.880 53.290 91.020 ;
        RECT 52.970 90.820 53.290 90.880 ;
        RECT 54.810 90.820 55.130 91.080 ;
        RECT 63.565 90.835 63.855 91.065 ;
        RECT 64.010 91.020 64.330 91.080 ;
        RECT 64.485 91.020 64.775 91.065 ;
        RECT 64.010 90.880 64.775 91.020 ;
        RECT 52.510 90.680 52.830 90.740 ;
        RECT 56.205 90.680 56.495 90.725 ;
        RECT 46.990 90.540 51.360 90.680 ;
        RECT 51.680 90.540 52.830 90.680 ;
        RECT 46.990 90.480 47.310 90.540 ;
        RECT 11.570 90.140 11.890 90.400 ;
        RECT 40.090 90.340 40.410 90.400 ;
        RECT 45.150 90.340 45.470 90.400 ;
        RECT 40.090 90.200 45.470 90.340 ;
        RECT 40.090 90.140 40.410 90.200 ;
        RECT 45.150 90.140 45.470 90.200 ;
        RECT 47.910 90.340 48.230 90.400 ;
        RECT 49.535 90.340 49.825 90.385 ;
        RECT 47.910 90.200 49.825 90.340 ;
        RECT 51.220 90.340 51.360 90.540 ;
        RECT 52.510 90.480 52.830 90.540 ;
        RECT 53.060 90.540 56.495 90.680 ;
        RECT 63.640 90.680 63.780 90.835 ;
        RECT 64.010 90.820 64.330 90.880 ;
        RECT 64.485 90.835 64.775 90.880 ;
        RECT 86.550 90.820 86.870 91.080 ;
        RECT 71.830 90.680 72.150 90.740 ;
        RECT 63.640 90.540 72.150 90.680 ;
        RECT 53.060 90.340 53.200 90.540 ;
        RECT 56.205 90.495 56.495 90.540 ;
        RECT 71.830 90.480 72.150 90.540 ;
        RECT 82.870 90.680 83.190 90.740 ;
        RECT 88.940 90.680 89.080 91.175 ;
        RECT 97.590 91.160 97.910 91.220 ;
        RECT 90.690 91.020 91.010 91.080 ;
        RECT 91.625 91.020 91.915 91.065 ;
        RECT 90.690 90.880 91.915 91.020 ;
        RECT 90.690 90.820 91.010 90.880 ;
        RECT 91.625 90.835 91.915 90.880 ;
        RECT 82.870 90.540 89.080 90.680 ;
        RECT 82.870 90.480 83.190 90.540 ;
        RECT 51.220 90.200 53.200 90.340 ;
        RECT 47.910 90.140 48.230 90.200 ;
        RECT 49.535 90.155 49.825 90.200 ;
        RECT 53.890 90.140 54.210 90.400 ;
        RECT 80.110 90.340 80.430 90.400 ;
        RECT 80.585 90.340 80.875 90.385 ;
        RECT 80.110 90.200 80.875 90.340 ;
        RECT 80.110 90.140 80.430 90.200 ;
        RECT 80.585 90.155 80.875 90.200 ;
        RECT 91.610 90.140 91.930 90.400 ;
        RECT 5.520 89.520 123.740 90.000 ;
        RECT 16.630 89.320 16.950 89.380 ;
        RECT 17.795 89.320 18.085 89.365 ;
        RECT 16.630 89.180 18.085 89.320 ;
        RECT 16.630 89.120 16.950 89.180 ;
        RECT 17.795 89.135 18.085 89.180 ;
        RECT 23.990 89.320 24.310 89.380 ;
        RECT 24.465 89.320 24.755 89.365 ;
        RECT 23.990 89.180 24.755 89.320 ;
        RECT 23.990 89.120 24.310 89.180 ;
        RECT 24.465 89.135 24.755 89.180 ;
        RECT 26.750 89.120 27.070 89.380 ;
        RECT 34.570 89.120 34.890 89.380 ;
        RECT 36.410 89.120 36.730 89.380 ;
        RECT 43.325 89.320 43.615 89.365 ;
        RECT 44.230 89.320 44.550 89.380 ;
        RECT 43.325 89.180 44.550 89.320 ;
        RECT 43.325 89.135 43.615 89.180 ;
        RECT 44.230 89.120 44.550 89.180 ;
        RECT 45.150 89.320 45.470 89.380 ;
        RECT 45.625 89.320 45.915 89.365 ;
        RECT 69.545 89.320 69.835 89.365 ;
        RECT 45.150 89.180 45.915 89.320 ;
        RECT 45.150 89.120 45.470 89.180 ;
        RECT 45.625 89.135 45.915 89.180 ;
        RECT 62.030 89.180 66.540 89.320 ;
        RECT 9.290 88.980 9.580 89.025 ;
        RECT 11.150 88.980 11.440 89.025 ;
        RECT 13.930 88.980 14.220 89.025 ;
        RECT 9.290 88.840 14.220 88.980 ;
        RECT 9.290 88.795 9.580 88.840 ;
        RECT 11.150 88.795 11.440 88.840 ;
        RECT 13.930 88.795 14.220 88.840 ;
        RECT 27.210 88.980 27.530 89.040 ;
        RECT 31.810 88.980 32.130 89.040 ;
        RECT 62.030 88.980 62.170 89.180 ;
        RECT 27.210 88.840 62.170 88.980 ;
        RECT 27.210 88.780 27.530 88.840 ;
        RECT 31.810 88.780 32.130 88.840 ;
        RECT 10.665 88.640 10.955 88.685 ;
        RECT 11.570 88.640 11.890 88.700 ;
        RECT 10.665 88.500 11.890 88.640 ;
        RECT 10.665 88.455 10.955 88.500 ;
        RECT 11.570 88.440 11.890 88.500 ;
        RECT 23.070 88.640 23.390 88.700 ;
        RECT 24.925 88.640 25.215 88.685 ;
        RECT 23.070 88.500 25.215 88.640 ;
        RECT 23.070 88.440 23.390 88.500 ;
        RECT 24.925 88.455 25.215 88.500 ;
        RECT 35.045 88.640 35.335 88.685 ;
        RECT 35.950 88.640 36.270 88.700 ;
        RECT 35.045 88.500 36.270 88.640 ;
        RECT 35.045 88.455 35.335 88.500 ;
        RECT 35.950 88.440 36.270 88.500 ;
        RECT 47.910 88.440 48.230 88.700 ;
        RECT 48.385 88.455 48.675 88.685 ;
        RECT 66.400 88.640 66.540 89.180 ;
        RECT 69.545 89.180 101.500 89.320 ;
        RECT 69.545 89.135 69.835 89.180 ;
        RECT 78.750 88.980 79.040 89.025 ;
        RECT 80.610 88.980 80.900 89.025 ;
        RECT 83.390 88.980 83.680 89.025 ;
        RECT 78.750 88.840 83.680 88.980 ;
        RECT 78.750 88.795 79.040 88.840 ;
        RECT 80.610 88.795 80.900 88.840 ;
        RECT 83.390 88.795 83.680 88.840 ;
        RECT 85.630 88.980 85.950 89.040 ;
        RECT 87.255 88.980 87.545 89.025 ;
        RECT 85.630 88.840 87.545 88.980 ;
        RECT 85.630 88.780 85.950 88.840 ;
        RECT 87.255 88.795 87.545 88.840 ;
        RECT 69.070 88.640 69.390 88.700 ;
        RECT 66.400 88.500 69.390 88.640 ;
        RECT 7.890 88.300 8.210 88.360 ;
        RECT 8.825 88.300 9.115 88.345 ;
        RECT 13.930 88.300 14.220 88.345 ;
        RECT 7.890 88.160 9.115 88.300 ;
        RECT 7.890 88.100 8.210 88.160 ;
        RECT 8.825 88.115 9.115 88.160 ;
        RECT 11.685 88.160 14.220 88.300 ;
        RECT 11.685 88.005 11.900 88.160 ;
        RECT 13.930 88.115 14.220 88.160 ;
        RECT 23.530 88.300 23.850 88.360 ;
        RECT 25.845 88.300 26.135 88.345 ;
        RECT 23.530 88.160 26.135 88.300 ;
        RECT 23.530 88.100 23.850 88.160 ;
        RECT 25.845 88.115 26.135 88.160 ;
        RECT 35.490 88.100 35.810 88.360 ;
        RECT 42.865 88.300 43.155 88.345 ;
        RECT 44.230 88.300 44.550 88.360 ;
        RECT 42.865 88.160 44.550 88.300 ;
        RECT 42.865 88.115 43.155 88.160 ;
        RECT 44.230 88.100 44.550 88.160 ;
        RECT 47.450 88.100 47.770 88.360 ;
        RECT 48.460 88.300 48.600 88.455 ;
        RECT 48.000 88.160 48.600 88.300 ;
        RECT 60.345 88.300 60.635 88.345 ;
        RECT 62.630 88.300 62.950 88.360 ;
        RECT 66.400 88.345 66.540 88.500 ;
        RECT 69.070 88.440 69.390 88.500 ;
        RECT 80.110 88.440 80.430 88.700 ;
        RECT 81.950 88.640 82.270 88.700 ;
        RECT 101.360 88.640 101.500 89.180 ;
        RECT 101.745 89.135 102.035 89.365 ;
        RECT 102.665 89.320 102.955 89.365 ;
        RECT 103.110 89.320 103.430 89.380 ;
        RECT 102.665 89.180 103.430 89.320 ;
        RECT 102.665 89.135 102.955 89.180 ;
        RECT 101.820 88.980 101.960 89.135 ;
        RECT 103.110 89.120 103.430 89.180 ;
        RECT 103.570 89.120 103.890 89.380 ;
        RECT 105.425 89.320 105.715 89.365 ;
        RECT 105.870 89.320 106.190 89.380 ;
        RECT 105.425 89.180 106.190 89.320 ;
        RECT 105.425 89.135 105.715 89.180 ;
        RECT 105.870 89.120 106.190 89.180 ;
        RECT 104.030 88.980 104.350 89.040 ;
        RECT 101.820 88.840 104.350 88.980 ;
        RECT 104.030 88.780 104.350 88.840 ;
        RECT 104.490 88.780 104.810 89.040 ;
        RECT 81.950 88.500 89.080 88.640 ;
        RECT 101.360 88.500 103.340 88.640 ;
        RECT 81.950 88.440 82.270 88.500 ;
        RECT 60.345 88.160 62.950 88.300 ;
        RECT 9.750 87.960 10.040 88.005 ;
        RECT 11.610 87.960 11.900 88.005 ;
        RECT 9.750 87.820 11.900 87.960 ;
        RECT 9.750 87.775 10.040 87.820 ;
        RECT 11.610 87.775 11.900 87.820 ;
        RECT 12.530 87.960 12.820 88.005 ;
        RECT 14.790 87.960 15.110 88.020 ;
        RECT 15.790 87.960 16.080 88.005 ;
        RECT 12.530 87.820 16.080 87.960 ;
        RECT 12.530 87.775 12.820 87.820 ;
        RECT 14.790 87.760 15.110 87.820 ;
        RECT 15.790 87.775 16.080 87.820 ;
        RECT 23.990 87.960 24.310 88.020 ;
        RECT 24.465 87.960 24.755 88.005 ;
        RECT 23.990 87.820 24.755 87.960 ;
        RECT 23.990 87.760 24.310 87.820 ;
        RECT 24.465 87.775 24.755 87.820 ;
        RECT 34.125 87.960 34.415 88.005 ;
        RECT 35.030 87.960 35.350 88.020 ;
        RECT 34.125 87.820 35.350 87.960 ;
        RECT 34.125 87.775 34.415 87.820 ;
        RECT 35.030 87.760 35.350 87.820 ;
        RECT 46.070 87.960 46.390 88.020 ;
        RECT 48.000 87.960 48.140 88.160 ;
        RECT 60.345 88.115 60.635 88.160 ;
        RECT 62.630 88.100 62.950 88.160 ;
        RECT 66.325 88.115 66.615 88.345 ;
        RECT 67.245 88.115 67.535 88.345 ;
        RECT 67.705 88.115 67.995 88.345 ;
        RECT 46.070 87.820 48.140 87.960 ;
        RECT 64.010 87.960 64.330 88.020 ;
        RECT 67.320 87.960 67.460 88.115 ;
        RECT 64.010 87.820 67.460 87.960 ;
        RECT 67.780 87.960 67.920 88.115 ;
        RECT 68.150 88.100 68.470 88.360 ;
        RECT 75.510 88.300 75.830 88.360 ;
        RECT 78.270 88.300 78.590 88.360 ;
        RECT 88.940 88.345 89.080 88.500 ;
        RECT 83.390 88.300 83.680 88.345 ;
        RECT 75.510 88.160 78.590 88.300 ;
        RECT 75.510 88.100 75.830 88.160 ;
        RECT 78.270 88.100 78.590 88.160 ;
        RECT 81.145 88.160 83.680 88.300 ;
        RECT 68.610 87.960 68.930 88.020 ;
        RECT 81.145 88.005 81.360 88.160 ;
        RECT 83.390 88.115 83.680 88.160 ;
        RECT 88.865 88.300 89.155 88.345 ;
        RECT 95.290 88.300 95.610 88.360 ;
        RECT 88.865 88.160 95.610 88.300 ;
        RECT 88.865 88.115 89.155 88.160 ;
        RECT 95.290 88.100 95.610 88.160 ;
        RECT 101.285 88.115 101.575 88.345 ;
        RECT 67.780 87.820 68.930 87.960 ;
        RECT 46.070 87.760 46.390 87.820 ;
        RECT 47.540 87.680 47.680 87.820 ;
        RECT 64.010 87.760 64.330 87.820 ;
        RECT 68.610 87.760 68.930 87.820 ;
        RECT 79.210 87.960 79.500 88.005 ;
        RECT 81.070 87.960 81.360 88.005 ;
        RECT 79.210 87.820 81.360 87.960 ;
        RECT 79.210 87.775 79.500 87.820 ;
        RECT 81.070 87.775 81.360 87.820 ;
        RECT 81.990 87.960 82.280 88.005 ;
        RECT 85.250 87.960 85.540 88.005 ;
        RECT 88.405 87.960 88.695 88.005 ;
        RECT 81.990 87.820 88.695 87.960 ;
        RECT 81.990 87.775 82.280 87.820 ;
        RECT 85.250 87.775 85.540 87.820 ;
        RECT 88.405 87.775 88.695 87.820 ;
        RECT 100.350 87.760 100.670 88.020 ;
        RECT 101.360 87.960 101.500 88.115 ;
        RECT 101.730 88.100 102.050 88.360 ;
        RECT 103.200 88.345 103.340 88.500 ;
        RECT 103.570 88.440 103.890 88.700 ;
        RECT 104.580 88.640 104.720 88.780 ;
        RECT 104.120 88.500 104.720 88.640 ;
        RECT 104.120 88.360 104.260 88.500 ;
        RECT 103.125 88.115 103.415 88.345 ;
        RECT 104.030 88.100 104.350 88.360 ;
        RECT 104.490 88.100 104.810 88.360 ;
        RECT 112.310 88.300 112.630 88.360 ;
        RECT 112.785 88.300 113.075 88.345 ;
        RECT 115.085 88.300 115.375 88.345 ;
        RECT 116.910 88.300 117.230 88.360 ;
        RECT 112.310 88.160 113.075 88.300 ;
        RECT 112.310 88.100 112.630 88.160 ;
        RECT 112.785 88.115 113.075 88.160 ;
        RECT 113.320 88.160 117.230 88.300 ;
        RECT 101.360 87.820 103.340 87.960 ;
        RECT 103.200 87.680 103.340 87.820 ;
        RECT 47.450 87.420 47.770 87.680 ;
        RECT 51.130 87.620 51.450 87.680 ;
        RECT 54.810 87.620 55.130 87.680 ;
        RECT 51.130 87.480 55.130 87.620 ;
        RECT 51.130 87.420 51.450 87.480 ;
        RECT 54.810 87.420 55.130 87.480 ;
        RECT 59.410 87.420 59.730 87.680 ;
        RECT 103.110 87.420 103.430 87.680 ;
        RECT 105.410 87.620 105.730 87.680 ;
        RECT 113.320 87.620 113.460 88.160 ;
        RECT 115.085 88.115 115.375 88.160 ;
        RECT 116.910 88.100 117.230 88.160 ;
        RECT 105.410 87.480 113.460 87.620 ;
        RECT 105.410 87.420 105.730 87.480 ;
        RECT 113.690 87.420 114.010 87.680 ;
        RECT 114.150 87.620 114.470 87.680 ;
        RECT 114.625 87.620 114.915 87.665 ;
        RECT 114.150 87.480 114.915 87.620 ;
        RECT 114.150 87.420 114.470 87.480 ;
        RECT 114.625 87.435 114.915 87.480 ;
        RECT 5.520 86.800 123.740 87.280 ;
        RECT 30.445 86.600 30.735 86.645 ;
        RECT 30.890 86.600 31.210 86.660 ;
        RECT 25.920 86.460 28.820 86.600 ;
        RECT 8.830 86.260 9.120 86.305 ;
        RECT 10.690 86.260 10.980 86.305 ;
        RECT 8.830 86.120 10.980 86.260 ;
        RECT 8.830 86.075 9.120 86.120 ;
        RECT 10.690 86.075 10.980 86.120 ;
        RECT 11.610 86.260 11.900 86.305 ;
        RECT 13.410 86.260 13.730 86.320 ;
        RECT 14.870 86.260 15.160 86.305 ;
        RECT 11.610 86.120 15.160 86.260 ;
        RECT 11.610 86.075 11.900 86.120 ;
        RECT 7.890 85.720 8.210 85.980 ;
        RECT 10.765 85.920 10.980 86.075 ;
        RECT 13.410 86.060 13.730 86.120 ;
        RECT 14.870 86.075 15.160 86.120 ;
        RECT 16.630 86.260 16.950 86.320 ;
        RECT 16.630 86.120 25.600 86.260 ;
        RECT 16.630 86.060 16.950 86.120 ;
        RECT 13.010 85.920 13.300 85.965 ;
        RECT 10.765 85.780 13.300 85.920 ;
        RECT 13.010 85.735 13.300 85.780 ;
        RECT 18.930 85.920 19.250 85.980 ;
        RECT 25.460 85.965 25.600 86.120 ;
        RECT 25.920 85.980 26.060 86.460 ;
        RECT 27.685 86.260 27.975 86.305 ;
        RECT 28.145 86.260 28.435 86.305 ;
        RECT 27.685 86.120 28.435 86.260 ;
        RECT 28.680 86.260 28.820 86.460 ;
        RECT 30.445 86.460 31.210 86.600 ;
        RECT 30.445 86.415 30.735 86.460 ;
        RECT 30.890 86.400 31.210 86.460 ;
        RECT 35.030 86.400 35.350 86.660 ;
        RECT 70.925 86.600 71.215 86.645 ;
        RECT 100.350 86.600 100.670 86.660 ;
        RECT 48.230 86.460 68.380 86.600 ;
        RECT 34.110 86.260 34.430 86.320 ;
        RECT 28.680 86.120 34.430 86.260 ;
        RECT 27.685 86.075 27.975 86.120 ;
        RECT 28.145 86.075 28.435 86.120 ;
        RECT 19.405 85.920 19.695 85.965 ;
        RECT 18.930 85.780 19.695 85.920 ;
        RECT 18.930 85.720 19.250 85.780 ;
        RECT 19.405 85.735 19.695 85.780 ;
        RECT 24.465 85.735 24.755 85.965 ;
        RECT 25.385 85.735 25.675 85.965 ;
        RECT 9.745 85.580 10.035 85.625 ;
        RECT 11.570 85.580 11.890 85.640 ;
        RECT 9.745 85.440 11.890 85.580 ;
        RECT 9.745 85.395 10.035 85.440 ;
        RECT 11.570 85.380 11.890 85.440 ;
        RECT 16.170 85.580 16.490 85.640 ;
        RECT 16.875 85.580 17.165 85.625 ;
        RECT 19.850 85.580 20.170 85.640 ;
        RECT 16.170 85.440 20.170 85.580 ;
        RECT 16.170 85.380 16.490 85.440 ;
        RECT 16.875 85.395 17.165 85.440 ;
        RECT 19.850 85.380 20.170 85.440 ;
        RECT 20.310 85.380 20.630 85.640 ;
        RECT 22.150 85.580 22.470 85.640 ;
        RECT 24.540 85.580 24.680 85.735 ;
        RECT 25.830 85.720 26.150 85.980 ;
        RECT 26.290 85.920 26.610 85.980 ;
        RECT 29.525 85.920 29.815 85.965 ;
        RECT 30.890 85.920 31.210 85.980 ;
        RECT 26.290 85.780 29.280 85.920 ;
        RECT 26.290 85.720 26.610 85.780 ;
        RECT 27.210 85.580 27.530 85.640 ;
        RECT 22.150 85.440 27.530 85.580 ;
        RECT 22.150 85.380 22.470 85.440 ;
        RECT 27.210 85.380 27.530 85.440 ;
        RECT 28.605 85.395 28.895 85.625 ;
        RECT 29.140 85.580 29.280 85.780 ;
        RECT 29.525 85.780 31.210 85.920 ;
        RECT 29.525 85.735 29.815 85.780 ;
        RECT 30.890 85.720 31.210 85.780 ;
        RECT 31.810 85.720 32.130 85.980 ;
        RECT 32.270 85.920 32.590 85.980 ;
        RECT 33.280 85.965 33.420 86.120 ;
        RECT 34.110 86.060 34.430 86.120 ;
        RECT 32.745 85.920 33.035 85.965 ;
        RECT 32.270 85.780 33.035 85.920 ;
        RECT 32.270 85.720 32.590 85.780 ;
        RECT 32.745 85.735 33.035 85.780 ;
        RECT 33.205 85.735 33.495 85.965 ;
        RECT 33.665 85.920 33.955 85.965 ;
        RECT 48.230 85.920 48.370 86.460 ;
        RECT 68.240 86.320 68.380 86.460 ;
        RECT 70.925 86.460 100.670 86.600 ;
        RECT 70.925 86.415 71.215 86.460 ;
        RECT 100.350 86.400 100.670 86.460 ;
        RECT 102.205 86.600 102.495 86.645 ;
        RECT 104.030 86.600 104.350 86.660 ;
        RECT 102.205 86.460 104.350 86.600 ;
        RECT 102.205 86.415 102.495 86.460 ;
        RECT 104.030 86.400 104.350 86.460 ;
        RECT 104.950 86.400 105.270 86.660 ;
        RECT 58.510 86.260 58.800 86.305 ;
        RECT 60.370 86.260 60.660 86.305 ;
        RECT 58.510 86.120 60.660 86.260 ;
        RECT 58.510 86.075 58.800 86.120 ;
        RECT 60.370 86.075 60.660 86.120 ;
        RECT 61.290 86.260 61.580 86.305 ;
        RECT 62.170 86.260 62.490 86.320 ;
        RECT 64.550 86.260 64.840 86.305 ;
        RECT 61.290 86.120 64.840 86.260 ;
        RECT 61.290 86.075 61.580 86.120 ;
        RECT 33.665 85.780 48.370 85.920 ;
        RECT 56.650 85.920 56.970 85.980 ;
        RECT 57.585 85.920 57.875 85.965 ;
        RECT 56.650 85.780 57.875 85.920 ;
        RECT 33.665 85.735 33.955 85.780 ;
        RECT 33.740 85.580 33.880 85.735 ;
        RECT 56.650 85.720 56.970 85.780 ;
        RECT 57.585 85.735 57.875 85.780 ;
        RECT 59.410 85.720 59.730 85.980 ;
        RECT 60.445 85.920 60.660 86.075 ;
        RECT 62.170 86.060 62.490 86.120 ;
        RECT 64.550 86.075 64.840 86.120 ;
        RECT 68.150 86.260 68.470 86.320 ;
        RECT 78.270 86.260 78.590 86.320 ;
        RECT 85.650 86.260 85.940 86.305 ;
        RECT 87.510 86.260 87.800 86.305 ;
        RECT 68.150 86.120 69.760 86.260 ;
        RECT 68.150 86.060 68.470 86.120 ;
        RECT 62.690 85.920 62.980 85.965 ;
        RECT 60.445 85.780 62.980 85.920 ;
        RECT 62.690 85.735 62.980 85.780 ;
        RECT 67.690 85.720 68.010 85.980 ;
        RECT 69.620 85.965 69.760 86.120 ;
        RECT 78.270 86.120 84.940 86.260 ;
        RECT 78.270 86.060 78.590 86.120 ;
        RECT 68.625 85.735 68.915 85.965 ;
        RECT 69.085 85.735 69.375 85.965 ;
        RECT 69.545 85.735 69.835 85.965 ;
        RECT 29.140 85.440 33.880 85.580 ;
        RECT 34.110 85.580 34.430 85.640 ;
        RECT 64.930 85.580 65.250 85.640 ;
        RECT 68.700 85.580 68.840 85.735 ;
        RECT 34.110 85.440 64.700 85.580 ;
        RECT 8.370 85.240 8.660 85.285 ;
        RECT 10.230 85.240 10.520 85.285 ;
        RECT 13.010 85.240 13.300 85.285 ;
        RECT 8.370 85.100 13.300 85.240 ;
        RECT 28.680 85.240 28.820 85.395 ;
        RECT 34.110 85.380 34.430 85.440 ;
        RECT 29.510 85.240 29.830 85.300 ;
        RECT 28.680 85.100 29.830 85.240 ;
        RECT 8.370 85.055 8.660 85.100 ;
        RECT 10.230 85.055 10.520 85.100 ;
        RECT 13.010 85.055 13.300 85.100 ;
        RECT 29.510 85.040 29.830 85.100 ;
        RECT 58.050 85.240 58.340 85.285 ;
        RECT 59.910 85.240 60.200 85.285 ;
        RECT 62.690 85.240 62.980 85.285 ;
        RECT 58.050 85.100 62.980 85.240 ;
        RECT 64.560 85.240 64.700 85.440 ;
        RECT 64.930 85.440 68.840 85.580 ;
        RECT 64.930 85.380 65.250 85.440 ;
        RECT 68.610 85.240 68.930 85.300 ;
        RECT 69.160 85.240 69.300 85.735 ;
        RECT 83.330 85.720 83.650 85.980 ;
        RECT 84.800 85.965 84.940 86.120 ;
        RECT 85.650 86.120 87.800 86.260 ;
        RECT 85.650 86.075 85.940 86.120 ;
        RECT 87.510 86.075 87.800 86.120 ;
        RECT 88.430 86.260 88.720 86.305 ;
        RECT 91.690 86.260 91.980 86.305 ;
        RECT 94.845 86.260 95.135 86.305 ;
        RECT 88.430 86.120 95.135 86.260 ;
        RECT 88.430 86.075 88.720 86.120 ;
        RECT 91.690 86.075 91.980 86.120 ;
        RECT 94.845 86.075 95.135 86.120 ;
        RECT 98.050 86.260 98.370 86.320 ;
        RECT 102.665 86.260 102.955 86.305 ;
        RECT 105.410 86.260 105.730 86.320 ;
        RECT 98.050 86.120 102.955 86.260 ;
        RECT 84.725 85.735 85.015 85.965 ;
        RECT 87.585 85.920 87.800 86.075 ;
        RECT 98.050 86.060 98.370 86.120 ;
        RECT 102.665 86.075 102.955 86.120 ;
        RECT 103.200 86.120 105.730 86.260 ;
        RECT 89.830 85.920 90.120 85.965 ;
        RECT 87.585 85.780 90.120 85.920 ;
        RECT 89.830 85.735 90.120 85.780 ;
        RECT 95.290 85.720 95.610 85.980 ;
        RECT 96.670 85.920 96.990 85.980 ;
        RECT 99.905 85.920 100.195 85.965 ;
        RECT 96.670 85.780 100.195 85.920 ;
        RECT 96.670 85.720 96.990 85.780 ;
        RECT 99.905 85.735 100.195 85.780 ;
        RECT 101.285 85.920 101.575 85.965 ;
        RECT 102.190 85.920 102.510 85.980 ;
        RECT 101.285 85.780 102.510 85.920 ;
        RECT 101.285 85.735 101.575 85.780 ;
        RECT 102.190 85.720 102.510 85.780 ;
        RECT 86.565 85.580 86.855 85.625 ;
        RECT 84.340 85.440 86.855 85.580 ;
        RECT 84.340 85.285 84.480 85.440 ;
        RECT 86.565 85.395 86.855 85.440 ;
        RECT 64.560 85.100 69.300 85.240 ;
        RECT 58.050 85.055 58.340 85.100 ;
        RECT 59.910 85.055 60.200 85.100 ;
        RECT 62.690 85.055 62.980 85.100 ;
        RECT 68.610 85.040 68.930 85.100 ;
        RECT 84.265 85.055 84.555 85.285 ;
        RECT 85.190 85.240 85.480 85.285 ;
        RECT 87.050 85.240 87.340 85.285 ;
        RECT 89.830 85.240 90.120 85.285 ;
        RECT 85.190 85.100 90.120 85.240 ;
        RECT 95.380 85.240 95.520 85.720 ;
        RECT 98.510 85.580 98.830 85.640 ;
        RECT 100.365 85.580 100.655 85.625 ;
        RECT 98.510 85.440 100.655 85.580 ;
        RECT 98.510 85.380 98.830 85.440 ;
        RECT 100.365 85.395 100.655 85.440 ;
        RECT 103.200 85.240 103.340 86.120 ;
        RECT 105.410 86.060 105.730 86.120 ;
        RECT 110.030 86.260 110.320 86.305 ;
        RECT 111.890 86.260 112.180 86.305 ;
        RECT 110.030 86.120 112.180 86.260 ;
        RECT 110.030 86.075 110.320 86.120 ;
        RECT 111.890 86.075 112.180 86.120 ;
        RECT 112.810 86.260 113.100 86.305 ;
        RECT 114.610 86.260 114.930 86.320 ;
        RECT 116.070 86.260 116.360 86.305 ;
        RECT 112.810 86.120 116.360 86.260 ;
        RECT 112.810 86.075 113.100 86.120 ;
        RECT 104.045 85.920 104.335 85.965 ;
        RECT 104.950 85.920 105.270 85.980 ;
        RECT 104.045 85.780 105.270 85.920 ;
        RECT 111.965 85.920 112.180 86.075 ;
        RECT 114.610 86.060 114.930 86.120 ;
        RECT 116.070 86.075 116.360 86.120 ;
        RECT 114.210 85.920 114.500 85.965 ;
        RECT 111.965 85.780 114.500 85.920 ;
        RECT 104.045 85.735 104.335 85.780 ;
        RECT 104.950 85.720 105.270 85.780 ;
        RECT 114.210 85.735 114.500 85.780 ;
        RECT 116.910 85.920 117.230 85.980 ;
        RECT 118.765 85.920 119.055 85.965 ;
        RECT 116.910 85.780 119.055 85.920 ;
        RECT 116.910 85.720 117.230 85.780 ;
        RECT 118.765 85.735 119.055 85.780 ;
        RECT 103.585 85.395 103.875 85.625 ;
        RECT 95.380 85.100 103.340 85.240 ;
        RECT 103.660 85.240 103.800 85.395 ;
        RECT 109.090 85.380 109.410 85.640 ;
        RECT 110.930 85.380 111.250 85.640 ;
        RECT 104.030 85.240 104.350 85.300 ;
        RECT 103.660 85.100 104.350 85.240 ;
        RECT 85.190 85.055 85.480 85.100 ;
        RECT 87.050 85.055 87.340 85.100 ;
        RECT 89.830 85.055 90.120 85.100 ;
        RECT 104.030 85.040 104.350 85.100 ;
        RECT 109.570 85.240 109.860 85.285 ;
        RECT 111.430 85.240 111.720 85.285 ;
        RECT 114.210 85.240 114.500 85.285 ;
        RECT 109.570 85.100 114.500 85.240 ;
        RECT 109.570 85.055 109.860 85.100 ;
        RECT 111.430 85.055 111.720 85.100 ;
        RECT 114.210 85.055 114.500 85.100 ;
        RECT 17.550 84.700 17.870 84.960 ;
        RECT 29.050 84.700 29.370 84.960 ;
        RECT 66.555 84.900 66.845 84.945 ;
        RECT 67.230 84.900 67.550 84.960 ;
        RECT 66.555 84.760 67.550 84.900 ;
        RECT 66.555 84.715 66.845 84.760 ;
        RECT 67.230 84.700 67.550 84.760 ;
        RECT 67.690 84.900 68.010 84.960 ;
        RECT 69.070 84.900 69.390 84.960 ;
        RECT 67.690 84.760 69.390 84.900 ;
        RECT 67.690 84.700 68.010 84.760 ;
        RECT 69.070 84.700 69.390 84.760 ;
        RECT 83.790 84.900 84.110 84.960 ;
        RECT 93.695 84.900 93.985 84.945 ;
        RECT 83.790 84.760 93.985 84.900 ;
        RECT 83.790 84.700 84.110 84.760 ;
        RECT 93.695 84.715 93.985 84.760 ;
        RECT 101.270 84.700 101.590 84.960 ;
        RECT 102.650 84.700 102.970 84.960 ;
        RECT 116.910 84.900 117.230 84.960 ;
        RECT 118.075 84.900 118.365 84.945 ;
        RECT 116.910 84.760 118.365 84.900 ;
        RECT 116.910 84.700 117.230 84.760 ;
        RECT 118.075 84.715 118.365 84.760 ;
        RECT 118.750 84.900 119.070 84.960 ;
        RECT 119.225 84.900 119.515 84.945 ;
        RECT 118.750 84.760 119.515 84.900 ;
        RECT 118.750 84.700 119.070 84.760 ;
        RECT 119.225 84.715 119.515 84.760 ;
        RECT 5.520 84.080 123.740 84.560 ;
        RECT 10.665 83.880 10.955 83.925 ;
        RECT 11.570 83.880 11.890 83.940 ;
        RECT 10.665 83.740 11.890 83.880 ;
        RECT 10.665 83.695 10.955 83.740 ;
        RECT 11.570 83.680 11.890 83.740 ;
        RECT 23.990 83.880 24.310 83.940 ;
        RECT 25.385 83.880 25.675 83.925 ;
        RECT 23.990 83.740 25.675 83.880 ;
        RECT 23.990 83.680 24.310 83.740 ;
        RECT 25.385 83.695 25.675 83.740 ;
        RECT 57.110 83.680 57.430 83.940 ;
        RECT 62.185 83.880 62.475 83.925 ;
        RECT 62.630 83.880 62.950 83.940 ;
        RECT 82.425 83.880 82.715 83.925 ;
        RECT 83.330 83.880 83.650 83.940 ;
        RECT 62.185 83.740 62.950 83.880 ;
        RECT 62.185 83.695 62.475 83.740 ;
        RECT 62.630 83.680 62.950 83.740 ;
        RECT 65.020 83.740 82.180 83.880 ;
        RECT 65.020 83.260 65.160 83.740 ;
        RECT 71.830 83.540 72.150 83.600 ;
        RECT 74.130 83.540 74.450 83.600 ;
        RECT 65.480 83.400 74.450 83.540 ;
        RECT 82.040 83.540 82.180 83.740 ;
        RECT 82.425 83.740 83.650 83.880 ;
        RECT 82.425 83.695 82.715 83.740 ;
        RECT 83.330 83.680 83.650 83.740 ;
        RECT 101.730 83.880 102.050 83.940 ;
        RECT 103.125 83.880 103.415 83.925 ;
        RECT 113.230 83.880 113.550 83.940 ;
        RECT 101.730 83.740 103.415 83.880 ;
        RECT 101.730 83.680 102.050 83.740 ;
        RECT 103.125 83.695 103.415 83.740 ;
        RECT 104.580 83.740 106.100 83.880 ;
        RECT 104.580 83.540 104.720 83.740 ;
        RECT 82.040 83.400 104.720 83.540 ;
        RECT 25.830 83.200 26.150 83.260 ;
        RECT 13.960 83.060 15.480 83.200 ;
        RECT 13.960 82.920 14.100 83.060 ;
        RECT 11.585 82.675 11.875 82.905 ;
        RECT 11.660 82.520 11.800 82.675 ;
        RECT 13.410 82.660 13.730 82.920 ;
        RECT 13.870 82.660 14.190 82.920 ;
        RECT 14.790 82.660 15.110 82.920 ;
        RECT 15.340 82.905 15.480 83.060 ;
        RECT 23.620 83.060 26.150 83.200 ;
        RECT 15.265 82.675 15.555 82.905 ;
        RECT 22.150 82.660 22.470 82.920 ;
        RECT 23.620 82.905 23.760 83.060 ;
        RECT 25.830 83.000 26.150 83.060 ;
        RECT 26.290 83.000 26.610 83.260 ;
        RECT 43.325 83.200 43.615 83.245 ;
        RECT 47.450 83.200 47.770 83.260 ;
        RECT 43.325 83.060 47.770 83.200 ;
        RECT 43.325 83.015 43.615 83.060 ;
        RECT 47.450 83.000 47.770 83.060 ;
        RECT 47.910 83.000 48.230 83.260 ;
        RECT 50.210 83.200 50.530 83.260 ;
        RECT 56.665 83.200 56.955 83.245 ;
        RECT 58.030 83.200 58.350 83.260 ;
        RECT 61.250 83.200 61.570 83.260 ;
        RECT 50.210 83.060 51.360 83.200 ;
        RECT 50.210 83.000 50.530 83.060 ;
        RECT 23.085 82.675 23.375 82.905 ;
        RECT 23.545 82.675 23.835 82.905 ;
        RECT 24.005 82.860 24.295 82.905 ;
        RECT 26.380 82.860 26.520 83.000 ;
        RECT 27.210 82.860 27.530 82.920 ;
        RECT 24.005 82.720 27.530 82.860 ;
        RECT 24.005 82.675 24.295 82.720 ;
        RECT 17.550 82.520 17.870 82.580 ;
        RECT 11.660 82.380 17.870 82.520 ;
        RECT 17.550 82.320 17.870 82.380 ;
        RECT 19.850 82.520 20.170 82.580 ;
        RECT 23.160 82.520 23.300 82.675 ;
        RECT 27.210 82.660 27.530 82.720 ;
        RECT 46.545 82.860 46.835 82.905 ;
        RECT 48.000 82.860 48.140 83.000 ;
        RECT 51.220 82.905 51.360 83.060 ;
        RECT 56.665 83.060 58.350 83.200 ;
        RECT 56.665 83.015 56.955 83.060 ;
        RECT 58.030 83.000 58.350 83.060 ;
        RECT 60.420 83.060 61.570 83.200 ;
        RECT 46.545 82.720 50.900 82.860 ;
        RECT 46.545 82.675 46.835 82.720 ;
        RECT 19.850 82.380 23.300 82.520 ;
        RECT 41.945 82.520 42.235 82.565 ;
        RECT 47.005 82.520 47.295 82.565 ;
        RECT 47.910 82.520 48.230 82.580 ;
        RECT 41.945 82.380 48.230 82.520 ;
        RECT 50.760 82.520 50.900 82.720 ;
        RECT 51.145 82.675 51.435 82.905 ;
        RECT 52.065 82.675 52.355 82.905 ;
        RECT 52.140 82.520 52.280 82.675 ;
        RECT 52.510 82.660 52.830 82.920 ;
        RECT 52.970 82.660 53.290 82.920 ;
        RECT 55.730 82.660 56.050 82.920 ;
        RECT 60.420 82.905 60.560 83.060 ;
        RECT 61.250 83.000 61.570 83.060 ;
        RECT 64.930 83.000 65.250 83.260 ;
        RECT 65.480 83.245 65.620 83.400 ;
        RECT 71.830 83.340 72.150 83.400 ;
        RECT 74.130 83.340 74.450 83.400 ;
        RECT 65.405 83.015 65.695 83.245 ;
        RECT 68.610 83.200 68.930 83.260 ;
        RECT 67.780 83.060 68.930 83.200 ;
        RECT 60.345 82.675 60.635 82.905 ;
        RECT 62.170 82.660 62.490 82.920 ;
        RECT 64.010 82.660 64.330 82.920 ;
        RECT 65.020 82.860 65.160 83.000 ;
        RECT 66.325 82.860 66.615 82.905 ;
        RECT 65.020 82.720 66.615 82.860 ;
        RECT 66.325 82.675 66.615 82.720 ;
        RECT 67.230 82.660 67.550 82.920 ;
        RECT 67.780 82.905 67.920 83.060 ;
        RECT 68.610 83.000 68.930 83.060 ;
        RECT 69.545 83.015 69.835 83.245 ;
        RECT 83.790 83.200 84.110 83.260 ;
        RECT 84.725 83.200 85.015 83.245 ;
        RECT 83.790 83.060 85.015 83.200 ;
        RECT 67.705 82.675 67.995 82.905 ;
        RECT 68.150 82.660 68.470 82.920 ;
        RECT 69.620 82.860 69.760 83.015 ;
        RECT 83.790 83.000 84.110 83.060 ;
        RECT 84.725 83.015 85.015 83.060 ;
        RECT 85.185 83.015 85.475 83.245 ;
        RECT 71.385 82.860 71.675 82.905 ;
        RECT 69.620 82.720 72.980 82.860 ;
        RECT 71.385 82.675 71.675 82.720 ;
        RECT 50.760 82.380 52.280 82.520 ;
        RECT 54.365 82.520 54.655 82.565 ;
        RECT 57.125 82.520 57.415 82.565 ;
        RECT 54.365 82.380 57.415 82.520 ;
        RECT 19.850 82.320 20.170 82.380 ;
        RECT 41.945 82.335 42.235 82.380 ;
        RECT 47.005 82.335 47.295 82.380 ;
        RECT 47.910 82.320 48.230 82.380 ;
        RECT 54.365 82.335 54.655 82.380 ;
        RECT 57.125 82.335 57.415 82.380 ;
        RECT 60.805 82.520 61.095 82.565 ;
        RECT 62.260 82.520 62.400 82.660 ;
        RECT 60.805 82.380 62.400 82.520 ;
        RECT 64.485 82.520 64.775 82.565 ;
        RECT 67.320 82.520 67.460 82.660 ;
        RECT 64.485 82.380 67.460 82.520 ;
        RECT 67.780 82.380 70.680 82.520 ;
        RECT 60.805 82.335 61.095 82.380 ;
        RECT 64.485 82.335 64.775 82.380 ;
        RECT 67.780 82.240 67.920 82.380 ;
        RECT 22.150 82.180 22.470 82.240 ;
        RECT 23.990 82.180 24.310 82.240 ;
        RECT 22.150 82.040 24.310 82.180 ;
        RECT 22.150 81.980 22.470 82.040 ;
        RECT 23.990 81.980 24.310 82.040 ;
        RECT 37.790 82.180 38.110 82.240 ;
        RECT 40.105 82.180 40.395 82.225 ;
        RECT 37.790 82.040 40.395 82.180 ;
        RECT 37.790 81.980 38.110 82.040 ;
        RECT 40.105 81.995 40.395 82.040 ;
        RECT 42.405 82.180 42.695 82.225 ;
        RECT 43.770 82.180 44.090 82.240 ;
        RECT 42.405 82.040 44.090 82.180 ;
        RECT 42.405 81.995 42.695 82.040 ;
        RECT 43.770 81.980 44.090 82.040 ;
        RECT 44.690 81.980 45.010 82.240 ;
        RECT 52.050 82.180 52.370 82.240 ;
        RECT 54.825 82.180 55.115 82.225 ;
        RECT 52.050 82.040 55.115 82.180 ;
        RECT 52.050 81.980 52.370 82.040 ;
        RECT 54.825 81.995 55.115 82.040 ;
        RECT 67.690 81.980 68.010 82.240 ;
        RECT 70.540 82.225 70.680 82.380 ;
        RECT 71.830 82.320 72.150 82.580 ;
        RECT 72.305 82.335 72.595 82.565 ;
        RECT 72.840 82.520 72.980 82.720 ;
        RECT 73.210 82.660 73.530 82.920 ;
        RECT 74.130 82.860 74.450 82.920 ;
        RECT 85.260 82.860 85.400 83.015 ;
        RECT 99.520 82.920 99.660 83.400 ;
        RECT 104.950 83.340 105.270 83.600 ;
        RECT 105.040 83.200 105.180 83.340 ;
        RECT 99.980 83.060 105.180 83.200 ;
        RECT 86.550 82.860 86.870 82.920 ;
        RECT 88.850 82.860 89.170 82.920 ;
        RECT 74.130 82.720 89.170 82.860 ;
        RECT 74.130 82.660 74.450 82.720 ;
        RECT 86.550 82.660 86.870 82.720 ;
        RECT 88.850 82.660 89.170 82.720 ;
        RECT 99.430 82.660 99.750 82.920 ;
        RECT 99.980 82.520 100.120 83.060 ;
        RECT 100.350 82.660 100.670 82.920 ;
        RECT 100.810 82.660 101.130 82.920 ;
        RECT 101.270 82.860 101.590 82.920 ;
        RECT 104.405 82.870 104.695 82.905 ;
        RECT 104.120 82.860 104.720 82.870 ;
        RECT 101.270 82.730 104.720 82.860 ;
        RECT 101.270 82.720 104.260 82.730 ;
        RECT 104.405 82.720 104.720 82.730 ;
        RECT 101.270 82.660 101.590 82.720 ;
        RECT 104.405 82.675 104.695 82.720 ;
        RECT 104.950 82.660 105.270 82.920 ;
        RECT 105.425 82.675 105.715 82.905 ;
        RECT 105.960 82.870 106.100 83.740 ;
        RECT 110.330 83.740 113.550 83.880 ;
        RECT 110.330 83.540 110.470 83.740 ;
        RECT 113.230 83.680 113.550 83.740 ;
        RECT 108.720 83.400 110.470 83.540 ;
        RECT 112.330 83.540 112.620 83.585 ;
        RECT 114.190 83.540 114.480 83.585 ;
        RECT 116.970 83.540 117.260 83.585 ;
        RECT 112.330 83.400 117.260 83.540 ;
        RECT 108.720 83.245 108.860 83.400 ;
        RECT 112.330 83.355 112.620 83.400 ;
        RECT 114.190 83.355 114.480 83.400 ;
        RECT 116.970 83.355 117.260 83.400 ;
        RECT 108.645 83.015 108.935 83.245 ;
        RECT 109.090 83.200 109.410 83.260 ;
        RECT 111.865 83.200 112.155 83.245 ;
        RECT 109.090 83.060 112.155 83.200 ;
        RECT 109.090 83.000 109.410 83.060 ;
        RECT 111.865 83.015 112.155 83.060 ;
        RECT 113.690 83.000 114.010 83.260 ;
        RECT 120.835 83.200 121.125 83.245 ;
        RECT 114.240 83.060 121.125 83.200 ;
        RECT 114.240 82.920 114.380 83.060 ;
        RECT 120.835 83.015 121.125 83.060 ;
        RECT 106.345 82.870 106.635 82.905 ;
        RECT 105.960 82.730 106.635 82.870 ;
        RECT 106.345 82.675 106.635 82.730 ;
        RECT 106.790 82.860 107.110 82.920 ;
        RECT 114.150 82.860 114.470 82.920 ;
        RECT 116.970 82.860 117.260 82.905 ;
        RECT 106.790 82.720 114.470 82.860 ;
        RECT 72.840 82.380 100.120 82.520 ;
        RECT 105.500 82.520 105.640 82.675 ;
        RECT 106.790 82.660 107.110 82.720 ;
        RECT 114.150 82.660 114.470 82.720 ;
        RECT 114.725 82.720 117.260 82.860 ;
        RECT 114.725 82.565 114.940 82.720 ;
        RECT 116.970 82.675 117.260 82.720 ;
        RECT 118.750 82.565 119.070 82.580 ;
        RECT 109.105 82.520 109.395 82.565 ;
        RECT 112.790 82.520 113.080 82.565 ;
        RECT 114.650 82.520 114.940 82.565 ;
        RECT 105.500 82.380 112.080 82.520 ;
        RECT 109.105 82.335 109.395 82.380 ;
        RECT 70.465 81.995 70.755 82.225 ;
        RECT 72.380 82.180 72.520 82.335 ;
        RECT 74.130 82.180 74.450 82.240 ;
        RECT 72.380 82.040 74.450 82.180 ;
        RECT 74.130 81.980 74.450 82.040 ;
        RECT 83.790 82.180 84.110 82.240 ;
        RECT 84.265 82.180 84.555 82.225 ;
        RECT 83.790 82.040 84.555 82.180 ;
        RECT 83.790 81.980 84.110 82.040 ;
        RECT 84.265 81.995 84.555 82.040 ;
        RECT 102.665 82.180 102.955 82.225 ;
        RECT 104.490 82.180 104.810 82.240 ;
        RECT 102.665 82.040 104.810 82.180 ;
        RECT 102.665 81.995 102.955 82.040 ;
        RECT 104.490 81.980 104.810 82.040 ;
        RECT 109.565 82.180 109.855 82.225 ;
        RECT 110.470 82.180 110.790 82.240 ;
        RECT 109.565 82.040 110.790 82.180 ;
        RECT 109.565 81.995 109.855 82.040 ;
        RECT 110.470 81.980 110.790 82.040 ;
        RECT 111.390 81.980 111.710 82.240 ;
        RECT 111.940 82.180 112.080 82.380 ;
        RECT 112.790 82.380 114.940 82.520 ;
        RECT 112.790 82.335 113.080 82.380 ;
        RECT 114.650 82.335 114.940 82.380 ;
        RECT 115.570 82.520 115.860 82.565 ;
        RECT 118.750 82.520 119.120 82.565 ;
        RECT 115.570 82.380 119.120 82.520 ;
        RECT 115.570 82.335 115.860 82.380 ;
        RECT 118.750 82.335 119.120 82.380 ;
        RECT 118.750 82.320 119.070 82.335 ;
        RECT 116.910 82.180 117.230 82.240 ;
        RECT 111.940 82.040 117.230 82.180 ;
        RECT 116.910 81.980 117.230 82.040 ;
        RECT 5.520 81.360 123.740 81.840 ;
        RECT 18.945 81.160 19.235 81.205 ;
        RECT 19.390 81.160 19.710 81.220 ;
        RECT 27.210 81.160 27.530 81.220 ;
        RECT 44.690 81.160 45.010 81.220 ;
        RECT 18.945 81.020 19.710 81.160 ;
        RECT 18.945 80.975 19.235 81.020 ;
        RECT 19.390 80.960 19.710 81.020 ;
        RECT 23.160 81.020 27.530 81.160 ;
        RECT 21.245 80.820 21.535 80.865 ;
        RECT 21.705 80.820 21.995 80.865 ;
        RECT 21.245 80.680 21.995 80.820 ;
        RECT 21.245 80.635 21.535 80.680 ;
        RECT 21.705 80.635 21.995 80.680 ;
        RECT 19.865 80.480 20.155 80.525 ;
        RECT 22.610 80.480 22.930 80.540 ;
        RECT 23.160 80.525 23.300 81.020 ;
        RECT 27.210 80.960 27.530 81.020 ;
        RECT 38.340 81.020 45.010 81.160 ;
        RECT 23.620 80.680 26.980 80.820 ;
        RECT 23.620 80.525 23.760 80.680 ;
        RECT 26.840 80.540 26.980 80.680 ;
        RECT 19.865 80.340 22.930 80.480 ;
        RECT 19.865 80.295 20.155 80.340 ;
        RECT 22.610 80.280 22.930 80.340 ;
        RECT 23.085 80.295 23.375 80.525 ;
        RECT 23.545 80.295 23.835 80.525 ;
        RECT 24.005 80.295 24.295 80.525 ;
        RECT 24.450 80.480 24.770 80.540 ;
        RECT 24.925 80.480 25.215 80.525 ;
        RECT 25.370 80.480 25.690 80.540 ;
        RECT 26.305 80.480 26.595 80.525 ;
        RECT 24.450 80.340 25.690 80.480 ;
        RECT 20.785 80.140 21.075 80.185 ;
        RECT 21.230 80.140 21.550 80.200 ;
        RECT 20.785 80.000 21.550 80.140 ;
        RECT 20.785 79.955 21.075 80.000 ;
        RECT 21.230 79.940 21.550 80.000 ;
        RECT 15.710 79.800 16.030 79.860 ;
        RECT 18.930 79.800 19.250 79.860 ;
        RECT 24.080 79.800 24.220 80.295 ;
        RECT 24.450 80.280 24.770 80.340 ;
        RECT 24.925 80.295 25.215 80.340 ;
        RECT 25.370 80.280 25.690 80.340 ;
        RECT 25.920 80.340 26.595 80.480 ;
        RECT 15.710 79.660 24.220 79.800 ;
        RECT 25.920 79.800 26.060 80.340 ;
        RECT 26.305 80.295 26.595 80.340 ;
        RECT 26.750 80.280 27.070 80.540 ;
        RECT 27.210 80.280 27.530 80.540 ;
        RECT 37.790 80.280 38.110 80.540 ;
        RECT 38.340 80.525 38.480 81.020 ;
        RECT 44.690 80.960 45.010 81.020 ;
        RECT 47.910 81.160 48.230 81.220 ;
        RECT 48.615 81.160 48.905 81.205 ;
        RECT 47.910 81.020 48.905 81.160 ;
        RECT 47.910 80.960 48.230 81.020 ;
        RECT 48.615 80.975 48.905 81.020 ;
        RECT 56.665 81.160 56.955 81.205 ;
        RECT 60.330 81.160 60.650 81.220 ;
        RECT 56.665 81.020 60.650 81.160 ;
        RECT 56.665 80.975 56.955 81.020 ;
        RECT 40.570 80.820 40.860 80.865 ;
        RECT 42.430 80.820 42.720 80.865 ;
        RECT 40.570 80.680 42.720 80.820 ;
        RECT 40.570 80.635 40.860 80.680 ;
        RECT 42.430 80.635 42.720 80.680 ;
        RECT 43.350 80.820 43.640 80.865 ;
        RECT 45.150 80.820 45.470 80.880 ;
        RECT 46.610 80.820 46.900 80.865 ;
        RECT 43.350 80.680 46.900 80.820 ;
        RECT 48.690 80.820 48.830 80.975 ;
        RECT 60.330 80.960 60.650 81.020 ;
        RECT 62.170 81.160 62.490 81.220 ;
        RECT 66.310 81.160 66.630 81.220 ;
        RECT 71.830 81.160 72.150 81.220 ;
        RECT 62.170 81.020 72.150 81.160 ;
        RECT 62.170 80.960 62.490 81.020 ;
        RECT 66.310 80.960 66.630 81.020 ;
        RECT 71.830 80.960 72.150 81.020 ;
        RECT 83.790 80.960 84.110 81.220 ;
        RECT 89.785 81.160 90.075 81.205 ;
        RECT 90.230 81.160 90.550 81.220 ;
        RECT 89.785 81.020 90.550 81.160 ;
        RECT 89.785 80.975 90.075 81.020 ;
        RECT 90.230 80.960 90.550 81.020 ;
        RECT 95.750 80.960 96.070 81.220 ;
        RECT 100.810 81.160 101.130 81.220 ;
        RECT 97.680 81.020 101.130 81.160 ;
        RECT 53.905 80.820 54.195 80.865 ;
        RECT 54.365 80.820 54.655 80.865 ;
        RECT 65.390 80.820 65.710 80.880 ;
        RECT 48.690 80.680 51.820 80.820 ;
        RECT 43.350 80.635 43.640 80.680 ;
        RECT 38.265 80.295 38.555 80.525 ;
        RECT 39.170 80.480 39.490 80.540 ;
        RECT 39.645 80.480 39.935 80.525 ;
        RECT 39.170 80.340 39.935 80.480 ;
        RECT 42.505 80.480 42.720 80.635 ;
        RECT 45.150 80.620 45.470 80.680 ;
        RECT 46.610 80.635 46.900 80.680 ;
        RECT 44.750 80.480 45.040 80.525 ;
        RECT 42.505 80.340 45.040 80.480 ;
        RECT 39.170 80.280 39.490 80.340 ;
        RECT 39.645 80.295 39.935 80.340 ;
        RECT 44.750 80.295 45.040 80.340 ;
        RECT 50.210 80.480 50.530 80.540 ;
        RECT 51.680 80.525 51.820 80.680 ;
        RECT 53.905 80.680 54.655 80.820 ;
        RECT 53.905 80.635 54.195 80.680 ;
        RECT 54.365 80.635 54.655 80.680 ;
        RECT 55.360 80.680 65.710 80.820 ;
        RECT 50.685 80.480 50.975 80.525 ;
        RECT 50.210 80.340 50.975 80.480 ;
        RECT 50.210 80.280 50.530 80.340 ;
        RECT 50.685 80.295 50.975 80.340 ;
        RECT 51.605 80.295 51.895 80.525 ;
        RECT 41.485 80.140 41.775 80.185 ;
        RECT 39.260 80.000 41.775 80.140 ;
        RECT 39.260 79.845 39.400 80.000 ;
        RECT 41.485 79.955 41.775 80.000 ;
        RECT 25.920 79.660 38.940 79.800 ;
        RECT 15.710 79.600 16.030 79.660 ;
        RECT 18.930 79.600 19.250 79.660 ;
        RECT 20.770 79.260 21.090 79.520 ;
        RECT 22.150 79.460 22.470 79.520 ;
        RECT 25.920 79.460 26.060 79.660 ;
        RECT 22.150 79.320 26.060 79.460 ;
        RECT 28.605 79.460 28.895 79.505 ;
        RECT 29.510 79.460 29.830 79.520 ;
        RECT 28.605 79.320 29.830 79.460 ;
        RECT 22.150 79.260 22.470 79.320 ;
        RECT 28.605 79.275 28.895 79.320 ;
        RECT 29.510 79.260 29.830 79.320 ;
        RECT 36.410 79.460 36.730 79.520 ;
        RECT 36.885 79.460 37.175 79.505 ;
        RECT 36.410 79.320 37.175 79.460 ;
        RECT 38.800 79.460 38.940 79.660 ;
        RECT 39.185 79.615 39.475 79.845 ;
        RECT 40.110 79.800 40.400 79.845 ;
        RECT 41.970 79.800 42.260 79.845 ;
        RECT 44.750 79.800 45.040 79.845 ;
        RECT 40.110 79.660 45.040 79.800 ;
        RECT 50.760 79.800 50.900 80.295 ;
        RECT 52.050 80.280 52.370 80.540 ;
        RECT 52.525 80.480 52.815 80.525 ;
        RECT 52.970 80.480 53.290 80.540 ;
        RECT 55.360 80.480 55.500 80.680 ;
        RECT 65.390 80.620 65.710 80.680 ;
        RECT 66.790 80.820 67.080 80.865 ;
        RECT 68.650 80.820 68.940 80.865 ;
        RECT 66.790 80.680 68.940 80.820 ;
        RECT 66.790 80.635 67.080 80.680 ;
        RECT 68.650 80.635 68.940 80.680 ;
        RECT 69.570 80.820 69.860 80.865 ;
        RECT 72.830 80.820 73.120 80.865 ;
        RECT 75.985 80.820 76.275 80.865 ;
        RECT 69.570 80.680 76.275 80.820 ;
        RECT 83.880 80.820 84.020 80.960 ;
        RECT 87.025 80.820 87.315 80.865 ;
        RECT 87.485 80.820 87.775 80.865 ;
        RECT 83.880 80.680 84.940 80.820 ;
        RECT 69.570 80.635 69.860 80.680 ;
        RECT 72.830 80.635 73.120 80.680 ;
        RECT 75.985 80.635 76.275 80.680 ;
        RECT 52.525 80.340 55.500 80.480 ;
        RECT 55.745 80.480 56.035 80.525 ;
        RECT 56.650 80.480 56.970 80.540 ;
        RECT 55.745 80.340 56.970 80.480 ;
        RECT 52.525 80.295 52.815 80.340 ;
        RECT 52.970 80.280 53.290 80.340 ;
        RECT 55.745 80.295 56.035 80.340 ;
        RECT 56.650 80.280 56.970 80.340 ;
        RECT 65.865 80.480 66.155 80.525 ;
        RECT 68.725 80.480 68.940 80.635 ;
        RECT 70.970 80.480 71.260 80.525 ;
        RECT 65.865 80.340 68.380 80.480 ;
        RECT 68.725 80.340 71.260 80.480 ;
        RECT 65.865 80.295 66.155 80.340 ;
        RECT 55.285 80.140 55.575 80.185 ;
        RECT 57.570 80.140 57.890 80.200 ;
        RECT 55.285 80.000 57.890 80.140 ;
        RECT 55.285 79.955 55.575 80.000 ;
        RECT 57.570 79.940 57.890 80.000 ;
        RECT 67.690 79.940 68.010 80.200 ;
        RECT 68.240 80.140 68.380 80.340 ;
        RECT 70.970 80.295 71.260 80.340 ;
        RECT 75.510 80.280 75.830 80.540 ;
        RECT 79.190 80.280 79.510 80.540 ;
        RECT 81.950 80.280 82.270 80.540 ;
        RECT 83.330 80.480 83.650 80.540 ;
        RECT 84.800 80.525 84.940 80.680 ;
        RECT 87.025 80.680 87.775 80.820 ;
        RECT 87.025 80.635 87.315 80.680 ;
        RECT 87.485 80.635 87.775 80.680 ;
        RECT 96.210 80.820 96.530 80.880 ;
        RECT 97.680 80.820 97.820 81.020 ;
        RECT 100.810 80.960 101.130 81.020 ;
        RECT 102.190 81.160 102.510 81.220 ;
        RECT 102.665 81.160 102.955 81.205 ;
        RECT 102.190 81.020 102.955 81.160 ;
        RECT 102.190 80.960 102.510 81.020 ;
        RECT 102.665 80.975 102.955 81.020 ;
        RECT 110.025 81.160 110.315 81.205 ;
        RECT 110.930 81.160 111.250 81.220 ;
        RECT 110.025 81.020 111.250 81.160 ;
        RECT 110.025 80.975 110.315 81.020 ;
        RECT 110.930 80.960 111.250 81.020 ;
        RECT 111.865 81.160 112.155 81.205 ;
        RECT 112.310 81.160 112.630 81.220 ;
        RECT 111.865 81.020 112.630 81.160 ;
        RECT 111.865 80.975 112.155 81.020 ;
        RECT 112.310 80.960 112.630 81.020 ;
        RECT 113.705 81.160 113.995 81.205 ;
        RECT 116.910 81.160 117.230 81.220 ;
        RECT 113.705 81.020 117.230 81.160 ;
        RECT 113.705 80.975 113.995 81.020 ;
        RECT 116.910 80.960 117.230 81.020 ;
        RECT 110.470 80.820 110.790 80.880 ;
        RECT 113.230 80.820 113.550 80.880 ;
        RECT 96.210 80.680 97.820 80.820 ;
        RECT 96.210 80.620 96.530 80.680 ;
        RECT 83.805 80.480 84.095 80.525 ;
        RECT 83.330 80.340 84.095 80.480 ;
        RECT 83.330 80.280 83.650 80.340 ;
        RECT 83.805 80.295 84.095 80.340 ;
        RECT 84.725 80.295 85.015 80.525 ;
        RECT 85.185 80.295 85.475 80.525 ;
        RECT 85.645 80.480 85.935 80.525 ;
        RECT 86.550 80.480 86.870 80.540 ;
        RECT 85.645 80.340 86.870 80.480 ;
        RECT 85.645 80.295 85.935 80.340 ;
        RECT 75.970 80.140 76.290 80.200 ;
        RECT 68.240 80.000 76.290 80.140 ;
        RECT 75.970 79.940 76.290 80.000 ;
        RECT 82.870 80.140 83.190 80.200 ;
        RECT 85.260 80.140 85.400 80.295 ;
        RECT 86.550 80.280 86.870 80.340 ;
        RECT 88.865 80.480 89.155 80.525 ;
        RECT 93.910 80.480 94.230 80.540 ;
        RECT 88.865 80.340 94.230 80.480 ;
        RECT 88.865 80.295 89.155 80.340 ;
        RECT 93.910 80.280 94.230 80.340 ;
        RECT 94.830 80.480 95.150 80.540 ;
        RECT 97.680 80.525 97.820 80.680 ;
        RECT 98.140 80.680 113.550 80.820 ;
        RECT 98.140 80.525 98.280 80.680 ;
        RECT 110.470 80.620 110.790 80.680 ;
        RECT 113.230 80.620 113.550 80.680 ;
        RECT 97.145 80.480 97.435 80.525 ;
        RECT 94.830 80.340 97.435 80.480 ;
        RECT 94.830 80.280 95.150 80.340 ;
        RECT 82.870 80.000 85.400 80.140 ;
        RECT 82.870 79.940 83.190 80.000 ;
        RECT 88.390 79.940 88.710 80.200 ;
        RECT 66.330 79.800 66.620 79.845 ;
        RECT 68.190 79.800 68.480 79.845 ;
        RECT 70.970 79.800 71.260 79.845 ;
        RECT 50.760 79.660 66.080 79.800 ;
        RECT 40.110 79.615 40.400 79.660 ;
        RECT 41.970 79.615 42.260 79.660 ;
        RECT 44.750 79.615 45.040 79.660 ;
        RECT 43.770 79.460 44.090 79.520 ;
        RECT 38.800 79.320 44.090 79.460 ;
        RECT 36.410 79.260 36.730 79.320 ;
        RECT 36.885 79.275 37.175 79.320 ;
        RECT 43.770 79.260 44.090 79.320 ;
        RECT 53.430 79.460 53.750 79.520 ;
        RECT 54.365 79.460 54.655 79.505 ;
        RECT 53.430 79.320 54.655 79.460 ;
        RECT 65.940 79.460 66.080 79.660 ;
        RECT 66.330 79.660 71.260 79.800 ;
        RECT 66.330 79.615 66.620 79.660 ;
        RECT 68.190 79.615 68.480 79.660 ;
        RECT 70.970 79.615 71.260 79.660 ;
        RECT 67.690 79.460 68.010 79.520 ;
        RECT 65.940 79.320 68.010 79.460 ;
        RECT 53.430 79.260 53.750 79.320 ;
        RECT 54.365 79.275 54.655 79.320 ;
        RECT 67.690 79.260 68.010 79.320 ;
        RECT 73.210 79.460 73.530 79.520 ;
        RECT 74.835 79.460 75.125 79.505 ;
        RECT 73.210 79.320 75.125 79.460 ;
        RECT 73.210 79.260 73.530 79.320 ;
        RECT 74.835 79.275 75.125 79.320 ;
        RECT 77.810 79.460 78.130 79.520 ;
        RECT 78.285 79.460 78.575 79.505 ;
        RECT 77.810 79.320 78.575 79.460 ;
        RECT 77.810 79.260 78.130 79.320 ;
        RECT 78.285 79.275 78.575 79.320 ;
        RECT 81.490 79.260 81.810 79.520 ;
        RECT 88.865 79.460 89.155 79.505 ;
        RECT 89.770 79.460 90.090 79.520 ;
        RECT 88.865 79.320 90.090 79.460 ;
        RECT 96.760 79.460 96.900 80.340 ;
        RECT 97.145 80.295 97.435 80.340 ;
        RECT 97.605 80.295 97.895 80.525 ;
        RECT 98.065 80.295 98.355 80.525 ;
        RECT 98.985 80.295 99.275 80.525 ;
        RECT 99.060 80.140 99.200 80.295 ;
        RECT 99.430 80.280 99.750 80.540 ;
        RECT 100.365 80.295 100.655 80.525 ;
        RECT 97.220 80.000 99.200 80.140 ;
        RECT 100.440 80.140 100.580 80.295 ;
        RECT 100.810 80.280 101.130 80.540 ;
        RECT 101.270 80.280 101.590 80.540 ;
        RECT 109.105 80.480 109.395 80.525 ;
        RECT 111.390 80.480 111.710 80.540 ;
        RECT 109.105 80.340 111.710 80.480 ;
        RECT 109.105 80.295 109.395 80.340 ;
        RECT 111.390 80.280 111.710 80.340 ;
        RECT 113.690 80.480 114.010 80.540 ;
        RECT 116.910 80.480 117.230 80.540 ;
        RECT 113.690 80.340 117.230 80.480 ;
        RECT 113.690 80.280 114.010 80.340 ;
        RECT 116.910 80.280 117.230 80.340 ;
        RECT 102.650 80.140 102.970 80.200 ;
        RECT 100.440 80.000 102.970 80.140 ;
        RECT 97.220 79.860 97.360 80.000 ;
        RECT 102.650 79.940 102.970 80.000 ;
        RECT 114.150 79.940 114.470 80.200 ;
        RECT 114.625 79.955 114.915 80.185 ;
        RECT 97.130 79.600 97.450 79.860 ;
        RECT 100.350 79.800 100.670 79.860 ;
        RECT 106.790 79.800 107.110 79.860 ;
        RECT 100.350 79.660 107.110 79.800 ;
        RECT 100.350 79.600 100.670 79.660 ;
        RECT 106.790 79.600 107.110 79.660 ;
        RECT 112.310 79.800 112.630 79.860 ;
        RECT 114.700 79.800 114.840 79.955 ;
        RECT 112.310 79.660 114.840 79.800 ;
        RECT 112.310 79.600 112.630 79.660 ;
        RECT 101.270 79.460 101.590 79.520 ;
        RECT 96.760 79.320 101.590 79.460 ;
        RECT 88.865 79.275 89.155 79.320 ;
        RECT 89.770 79.260 90.090 79.320 ;
        RECT 101.270 79.260 101.590 79.320 ;
        RECT 116.450 79.260 116.770 79.520 ;
        RECT 5.520 78.640 123.740 79.120 ;
        RECT 12.030 78.440 12.350 78.500 ;
        RECT 19.405 78.440 19.695 78.485 ;
        RECT 12.030 78.300 19.695 78.440 ;
        RECT 12.030 78.240 12.350 78.300 ;
        RECT 19.405 78.255 19.695 78.300 ;
        RECT 21.690 78.240 22.010 78.500 ;
        RECT 27.225 78.440 27.515 78.485 ;
        RECT 22.240 78.300 27.515 78.440 ;
        RECT 12.490 78.100 12.810 78.160 ;
        RECT 22.240 78.100 22.380 78.300 ;
        RECT 27.225 78.255 27.515 78.300 ;
        RECT 28.590 78.240 28.910 78.500 ;
        RECT 43.770 78.240 44.090 78.500 ;
        RECT 45.150 78.240 45.470 78.500 ;
        RECT 79.190 78.440 79.510 78.500 ;
        RECT 85.645 78.440 85.935 78.485 ;
        RECT 79.190 78.300 85.935 78.440 ;
        RECT 79.190 78.240 79.510 78.300 ;
        RECT 85.645 78.255 85.935 78.300 ;
        RECT 12.490 77.960 22.380 78.100 ;
        RECT 35.915 78.100 36.205 78.145 ;
        RECT 37.805 78.100 38.095 78.145 ;
        RECT 40.925 78.100 41.215 78.145 ;
        RECT 35.915 77.960 41.215 78.100 ;
        RECT 12.490 77.900 12.810 77.960 ;
        RECT 35.915 77.915 36.205 77.960 ;
        RECT 37.805 77.915 38.095 77.960 ;
        RECT 40.925 77.915 41.215 77.960 ;
        RECT 65.865 78.100 66.155 78.145 ;
        RECT 68.150 78.100 68.470 78.160 ;
        RECT 76.450 78.100 76.740 78.145 ;
        RECT 78.310 78.100 78.600 78.145 ;
        RECT 81.090 78.100 81.380 78.145 ;
        RECT 65.865 77.960 72.520 78.100 ;
        RECT 65.865 77.915 66.155 77.960 ;
        RECT 68.150 77.900 68.470 77.960 ;
        RECT 16.645 77.575 16.935 77.805 ;
        RECT 26.750 77.760 27.070 77.820 ;
        RECT 24.080 77.620 27.070 77.760 ;
        RECT 16.720 77.420 16.860 77.575 ;
        RECT 19.850 77.420 20.170 77.480 ;
        RECT 16.720 77.280 20.170 77.420 ;
        RECT 19.850 77.220 20.170 77.280 ;
        RECT 20.325 77.235 20.615 77.465 ;
        RECT 20.400 77.080 20.540 77.235 ;
        RECT 20.770 77.220 21.090 77.480 ;
        RECT 24.080 77.465 24.220 77.620 ;
        RECT 26.750 77.560 27.070 77.620 ;
        RECT 36.410 77.560 36.730 77.820 ;
        RECT 62.630 77.760 62.950 77.820 ;
        RECT 68.610 77.760 68.930 77.820 ;
        RECT 62.630 77.620 72.060 77.760 ;
        RECT 62.630 77.560 62.950 77.620 ;
        RECT 68.610 77.560 68.930 77.620 ;
        RECT 23.545 77.235 23.835 77.465 ;
        RECT 24.005 77.235 24.295 77.465 ;
        RECT 21.230 77.080 21.550 77.140 ;
        RECT 20.400 76.940 21.550 77.080 ;
        RECT 21.230 76.880 21.550 76.940 ;
        RECT 21.705 77.080 21.995 77.125 ;
        RECT 22.165 77.080 22.455 77.125 ;
        RECT 21.705 76.940 22.455 77.080 ;
        RECT 23.620 77.080 23.760 77.235 ;
        RECT 24.450 77.220 24.770 77.480 ;
        RECT 25.370 77.220 25.690 77.480 ;
        RECT 28.130 77.220 28.450 77.480 ;
        RECT 28.605 77.235 28.895 77.465 ;
        RECT 27.210 77.080 27.530 77.140 ;
        RECT 23.620 76.940 27.530 77.080 ;
        RECT 21.705 76.895 21.995 76.940 ;
        RECT 22.165 76.895 22.455 76.940 ;
        RECT 27.210 76.880 27.530 76.940 ;
        RECT 11.110 76.740 11.430 76.800 ;
        RECT 13.425 76.740 13.715 76.785 ;
        RECT 11.110 76.600 13.715 76.740 ;
        RECT 11.110 76.540 11.430 76.600 ;
        RECT 13.425 76.555 13.715 76.600 ;
        RECT 15.250 76.540 15.570 76.800 ;
        RECT 15.710 76.540 16.030 76.800 ;
        RECT 28.680 76.740 28.820 77.235 ;
        RECT 29.510 77.220 29.830 77.480 ;
        RECT 34.570 77.420 34.890 77.480 ;
        RECT 35.045 77.420 35.335 77.465 ;
        RECT 34.570 77.280 35.335 77.420 ;
        RECT 34.570 77.220 34.890 77.280 ;
        RECT 35.045 77.235 35.335 77.280 ;
        RECT 35.510 77.420 35.800 77.465 ;
        RECT 37.345 77.420 37.635 77.465 ;
        RECT 40.925 77.420 41.215 77.465 ;
        RECT 35.510 77.280 41.215 77.420 ;
        RECT 35.510 77.235 35.800 77.280 ;
        RECT 37.345 77.235 37.635 77.280 ;
        RECT 40.925 77.235 41.215 77.280 ;
        RECT 38.705 77.080 39.355 77.125 ;
        RECT 41.470 77.080 41.790 77.140 ;
        RECT 42.005 77.125 42.295 77.440 ;
        RECT 44.690 77.220 45.010 77.480 ;
        RECT 66.770 77.220 67.090 77.480 ;
        RECT 69.070 77.420 69.390 77.480 ;
        RECT 71.920 77.465 72.060 77.620 ;
        RECT 72.380 77.465 72.520 77.960 ;
        RECT 76.450 77.960 81.380 78.100 ;
        RECT 76.450 77.915 76.740 77.960 ;
        RECT 78.310 77.915 78.600 77.960 ;
        RECT 81.090 77.915 81.380 77.960 ;
        RECT 83.790 78.100 84.110 78.160 ;
        RECT 84.955 78.100 85.245 78.145 ;
        RECT 83.790 77.960 88.160 78.100 ;
        RECT 83.790 77.900 84.110 77.960 ;
        RECT 84.955 77.915 85.245 77.960 ;
        RECT 75.970 77.560 76.290 77.820 ;
        RECT 77.810 77.560 78.130 77.820 ;
        RECT 88.020 77.805 88.160 77.960 ;
        RECT 110.485 77.915 110.775 78.145 ;
        RECT 111.410 78.100 111.700 78.145 ;
        RECT 113.270 78.100 113.560 78.145 ;
        RECT 116.050 78.100 116.340 78.145 ;
        RECT 111.410 77.960 116.340 78.100 ;
        RECT 111.410 77.915 111.700 77.960 ;
        RECT 113.270 77.915 113.560 77.960 ;
        RECT 116.050 77.915 116.340 77.960 ;
        RECT 87.945 77.575 88.235 77.805 ;
        RECT 88.850 77.560 89.170 77.820 ;
        RECT 110.560 77.760 110.700 77.915 ;
        RECT 112.785 77.760 113.075 77.805 ;
        RECT 110.560 77.620 113.075 77.760 ;
        RECT 112.785 77.575 113.075 77.620 ;
        RECT 70.465 77.420 70.755 77.465 ;
        RECT 69.070 77.280 70.755 77.420 ;
        RECT 69.070 77.220 69.390 77.280 ;
        RECT 70.465 77.235 70.755 77.280 ;
        RECT 71.385 77.235 71.675 77.465 ;
        RECT 71.845 77.235 72.135 77.465 ;
        RECT 72.305 77.235 72.595 77.465 ;
        RECT 81.090 77.420 81.380 77.465 ;
        RECT 78.845 77.280 81.380 77.420 ;
        RECT 42.005 77.080 42.595 77.125 ;
        RECT 38.705 76.940 42.595 77.080 ;
        RECT 71.460 77.080 71.600 77.235 ;
        RECT 73.210 77.080 73.530 77.140 ;
        RECT 78.845 77.125 79.060 77.280 ;
        RECT 81.090 77.235 81.380 77.280 ;
        RECT 109.565 77.420 109.855 77.465 ;
        RECT 110.470 77.420 110.790 77.480 ;
        RECT 109.565 77.280 110.790 77.420 ;
        RECT 109.565 77.235 109.855 77.280 ;
        RECT 110.470 77.220 110.790 77.280 ;
        RECT 110.930 77.220 111.250 77.480 ;
        RECT 116.050 77.420 116.340 77.465 ;
        RECT 113.805 77.280 116.340 77.420 ;
        RECT 71.460 76.940 73.530 77.080 ;
        RECT 38.705 76.895 39.355 76.940 ;
        RECT 41.470 76.880 41.790 76.940 ;
        RECT 42.305 76.895 42.595 76.940 ;
        RECT 73.210 76.880 73.530 76.940 ;
        RECT 76.910 77.080 77.200 77.125 ;
        RECT 78.770 77.080 79.060 77.125 ;
        RECT 76.910 76.940 79.060 77.080 ;
        RECT 76.910 76.895 77.200 76.940 ;
        RECT 78.770 76.895 79.060 76.940 ;
        RECT 79.690 77.080 79.980 77.125 ;
        RECT 81.490 77.080 81.810 77.140 ;
        RECT 82.950 77.080 83.240 77.125 ;
        RECT 96.670 77.080 96.990 77.140 ;
        RECT 113.805 77.125 114.020 77.280 ;
        RECT 116.050 77.235 116.340 77.280 ;
        RECT 79.690 76.940 83.240 77.080 ;
        RECT 79.690 76.895 79.980 76.940 ;
        RECT 81.490 76.880 81.810 76.940 ;
        RECT 82.950 76.895 83.240 76.940 ;
        RECT 83.420 76.940 96.990 77.080 ;
        RECT 29.510 76.740 29.830 76.800 ;
        RECT 28.680 76.600 29.830 76.740 ;
        RECT 29.510 76.540 29.830 76.600 ;
        RECT 52.510 76.740 52.830 76.800 ;
        RECT 66.310 76.740 66.630 76.800 ;
        RECT 52.510 76.600 66.630 76.740 ;
        RECT 52.510 76.540 52.830 76.600 ;
        RECT 66.310 76.540 66.630 76.600 ;
        RECT 73.685 76.740 73.975 76.785 ;
        RECT 83.420 76.740 83.560 76.940 ;
        RECT 96.670 76.880 96.990 76.940 ;
        RECT 111.870 77.080 112.160 77.125 ;
        RECT 113.730 77.080 114.020 77.125 ;
        RECT 111.870 76.940 114.020 77.080 ;
        RECT 111.870 76.895 112.160 76.940 ;
        RECT 113.730 76.895 114.020 76.940 ;
        RECT 114.650 77.080 114.940 77.125 ;
        RECT 116.450 77.080 116.770 77.140 ;
        RECT 117.910 77.080 118.200 77.125 ;
        RECT 114.650 76.940 118.200 77.080 ;
        RECT 114.650 76.895 114.940 76.940 ;
        RECT 116.450 76.880 116.770 76.940 ;
        RECT 117.910 76.895 118.200 76.940 ;
        RECT 73.685 76.600 83.560 76.740 ;
        RECT 83.790 76.740 84.110 76.800 ;
        RECT 87.485 76.740 87.775 76.785 ;
        RECT 83.790 76.600 87.775 76.740 ;
        RECT 73.685 76.555 73.975 76.600 ;
        RECT 83.790 76.540 84.110 76.600 ;
        RECT 87.485 76.555 87.775 76.600 ;
        RECT 113.230 76.740 113.550 76.800 ;
        RECT 119.915 76.740 120.205 76.785 ;
        RECT 113.230 76.600 120.205 76.740 ;
        RECT 113.230 76.540 113.550 76.600 ;
        RECT 119.915 76.555 120.205 76.600 ;
        RECT 5.520 75.920 123.740 76.400 ;
        RECT 22.610 75.720 22.930 75.780 ;
        RECT 23.085 75.720 23.375 75.765 ;
        RECT 22.610 75.580 23.375 75.720 ;
        RECT 22.610 75.520 22.930 75.580 ;
        RECT 23.085 75.535 23.375 75.580 ;
        RECT 26.765 75.720 27.055 75.765 ;
        RECT 28.130 75.720 28.450 75.780 ;
        RECT 26.765 75.580 28.450 75.720 ;
        RECT 26.765 75.535 27.055 75.580 ;
        RECT 28.130 75.520 28.450 75.580 ;
        RECT 40.105 75.720 40.395 75.765 ;
        RECT 41.470 75.720 41.790 75.780 ;
        RECT 40.105 75.580 41.790 75.720 ;
        RECT 40.105 75.535 40.395 75.580 ;
        RECT 41.470 75.520 41.790 75.580 ;
        RECT 47.450 75.720 47.770 75.780 ;
        RECT 55.270 75.720 55.590 75.780 ;
        RECT 47.450 75.580 55.590 75.720 ;
        RECT 47.450 75.520 47.770 75.580 ;
        RECT 55.270 75.520 55.590 75.580 ;
        RECT 56.205 75.720 56.495 75.765 ;
        RECT 56.650 75.720 56.970 75.780 ;
        RECT 56.205 75.580 56.970 75.720 ;
        RECT 56.205 75.535 56.495 75.580 ;
        RECT 56.650 75.520 56.970 75.580 ;
        RECT 62.630 75.520 62.950 75.780 ;
        RECT 82.425 75.720 82.715 75.765 ;
        RECT 92.085 75.720 92.375 75.765 ;
        RECT 92.990 75.720 93.310 75.780 ;
        RECT 82.425 75.580 90.000 75.720 ;
        RECT 82.425 75.535 82.715 75.580 ;
        RECT 16.645 75.380 16.935 75.425 ;
        RECT 22.150 75.380 22.470 75.440 ;
        RECT 16.645 75.240 22.470 75.380 ;
        RECT 16.645 75.195 16.935 75.240 ;
        RECT 22.150 75.180 22.470 75.240 ;
        RECT 26.380 75.240 30.200 75.380 ;
        RECT 11.110 74.840 11.430 75.100 ;
        RECT 12.505 74.855 12.795 75.085 ;
        RECT 12.580 74.700 12.720 74.855 ;
        RECT 13.870 74.840 14.190 75.100 ;
        RECT 15.250 75.040 15.570 75.100 ;
        RECT 17.090 75.040 17.410 75.100 ;
        RECT 23.990 75.040 24.310 75.100 ;
        RECT 15.250 74.900 24.310 75.040 ;
        RECT 15.250 74.840 15.570 74.900 ;
        RECT 17.090 74.840 17.410 74.900 ;
        RECT 23.990 74.840 24.310 74.900 ;
        RECT 24.450 74.840 24.770 75.100 ;
        RECT 24.925 74.855 25.215 75.085 ;
        RECT 18.025 74.700 18.315 74.745 ;
        RECT 20.310 74.700 20.630 74.760 ;
        RECT 12.580 74.560 13.870 74.700 ;
        RECT 13.730 74.360 13.870 74.560 ;
        RECT 18.025 74.560 20.630 74.700 ;
        RECT 18.025 74.515 18.315 74.560 ;
        RECT 20.310 74.500 20.630 74.560 ;
        RECT 14.805 74.360 15.095 74.405 ;
        RECT 13.730 74.220 15.095 74.360 ;
        RECT 14.805 74.175 15.095 74.220 ;
        RECT 8.810 74.020 9.130 74.080 ;
        RECT 10.205 74.020 10.495 74.065 ;
        RECT 8.810 73.880 10.495 74.020 ;
        RECT 8.810 73.820 9.130 73.880 ;
        RECT 10.205 73.835 10.495 73.880 ;
        RECT 11.570 73.820 11.890 74.080 ;
        RECT 13.410 73.820 13.730 74.080 ;
        RECT 25.000 74.020 25.140 74.855 ;
        RECT 25.370 74.840 25.690 75.100 ;
        RECT 26.380 75.085 26.520 75.240 ;
        RECT 26.305 74.855 26.595 75.085 ;
        RECT 27.670 75.040 27.990 75.100 ;
        RECT 28.145 75.040 28.435 75.085 ;
        RECT 27.670 74.900 28.435 75.040 ;
        RECT 27.670 74.840 27.990 74.900 ;
        RECT 28.145 74.855 28.435 74.900 ;
        RECT 28.590 74.840 28.910 75.100 ;
        RECT 30.060 75.085 30.200 75.240 ;
        RECT 64.010 75.180 64.330 75.440 ;
        RECT 66.310 75.380 66.630 75.440 ;
        RECT 82.870 75.380 83.190 75.440 ;
        RECT 89.860 75.425 90.000 75.580 ;
        RECT 92.085 75.580 93.310 75.720 ;
        RECT 92.085 75.535 92.375 75.580 ;
        RECT 92.990 75.520 93.310 75.580 ;
        RECT 93.450 75.720 93.770 75.780 ;
        RECT 93.925 75.720 94.215 75.765 ;
        RECT 96.670 75.720 96.990 75.780 ;
        RECT 93.450 75.580 94.215 75.720 ;
        RECT 93.450 75.520 93.770 75.580 ;
        RECT 93.925 75.535 94.215 75.580 ;
        RECT 95.380 75.580 96.990 75.720 ;
        RECT 86.565 75.380 86.855 75.425 ;
        RECT 87.025 75.380 87.315 75.425 ;
        RECT 66.310 75.240 84.940 75.380 ;
        RECT 66.310 75.180 66.630 75.240 ;
        RECT 29.065 74.855 29.355 75.085 ;
        RECT 29.985 75.040 30.275 75.085 ;
        RECT 33.190 75.040 33.510 75.100 ;
        RECT 29.985 74.900 33.510 75.040 ;
        RECT 29.985 74.855 30.275 74.900 ;
        RECT 29.140 74.700 29.280 74.855 ;
        RECT 33.190 74.840 33.510 74.900 ;
        RECT 38.250 75.040 38.570 75.100 ;
        RECT 39.645 75.040 39.935 75.085 ;
        RECT 38.250 74.900 39.935 75.040 ;
        RECT 38.250 74.840 38.570 74.900 ;
        RECT 39.645 74.855 39.935 74.900 ;
        RECT 52.050 75.040 52.370 75.100 ;
        RECT 52.985 75.040 53.275 75.085 ;
        RECT 52.050 74.900 53.275 75.040 ;
        RECT 52.050 74.840 52.370 74.900 ;
        RECT 52.985 74.855 53.275 74.900 ;
        RECT 53.905 74.855 54.195 75.085 ;
        RECT 31.350 74.700 31.670 74.760 ;
        RECT 29.140 74.560 31.670 74.700 ;
        RECT 31.350 74.500 31.670 74.560 ;
        RECT 52.510 74.700 52.830 74.760 ;
        RECT 53.980 74.700 54.120 74.855 ;
        RECT 54.350 74.840 54.670 75.100 ;
        RECT 54.825 75.040 55.115 75.085 ;
        RECT 55.730 75.040 56.050 75.100 ;
        RECT 54.825 74.900 56.050 75.040 ;
        RECT 54.825 74.855 55.115 74.900 ;
        RECT 55.730 74.840 56.050 74.900 ;
        RECT 59.410 74.840 59.730 75.100 ;
        RECT 63.565 75.040 63.855 75.085 ;
        RECT 65.850 75.040 66.170 75.100 ;
        RECT 63.565 74.900 66.170 75.040 ;
        RECT 63.565 74.855 63.855 74.900 ;
        RECT 65.850 74.840 66.170 74.900 ;
        RECT 67.690 75.040 68.010 75.100 ;
        RECT 78.730 75.040 79.050 75.100 ;
        RECT 79.205 75.040 79.495 75.085 ;
        RECT 80.020 75.055 80.310 75.100 ;
        RECT 80.660 75.085 80.800 75.240 ;
        RECT 82.870 75.180 83.190 75.240 ;
        RECT 67.690 74.900 79.495 75.040 ;
        RECT 67.690 74.840 68.010 74.900 ;
        RECT 78.730 74.840 79.050 74.900 ;
        RECT 79.205 74.855 79.495 74.900 ;
        RECT 79.740 74.915 80.310 75.055 ;
        RECT 52.510 74.560 54.120 74.700 ;
        RECT 55.270 74.700 55.590 74.760 ;
        RECT 58.045 74.700 58.335 74.745 ;
        RECT 55.270 74.560 58.335 74.700 ;
        RECT 52.510 74.500 52.830 74.560 ;
        RECT 55.270 74.500 55.590 74.560 ;
        RECT 58.045 74.515 58.335 74.560 ;
        RECT 78.270 74.700 78.590 74.760 ;
        RECT 79.740 74.700 79.880 74.915 ;
        RECT 80.020 74.870 80.310 74.915 ;
        RECT 80.585 74.855 80.875 75.085 ;
        RECT 81.030 74.840 81.350 75.100 ;
        RECT 83.330 74.840 83.650 75.100 ;
        RECT 83.790 75.040 84.110 75.100 ;
        RECT 84.800 75.085 84.940 75.240 ;
        RECT 86.565 75.240 87.315 75.380 ;
        RECT 86.565 75.195 86.855 75.240 ;
        RECT 87.025 75.195 87.315 75.240 ;
        RECT 89.785 75.195 90.075 75.425 ;
        RECT 90.230 75.380 90.550 75.440 ;
        RECT 95.380 75.380 95.520 75.580 ;
        RECT 96.670 75.520 96.990 75.580 ;
        RECT 97.590 75.520 97.910 75.780 ;
        RECT 110.470 75.720 110.790 75.780 ;
        RECT 112.325 75.720 112.615 75.765 ;
        RECT 110.470 75.580 112.615 75.720 ;
        RECT 110.470 75.520 110.790 75.580 ;
        RECT 112.325 75.535 112.615 75.580 ;
        RECT 113.230 75.720 113.550 75.780 ;
        RECT 114.625 75.720 114.915 75.765 ;
        RECT 113.230 75.580 114.915 75.720 ;
        RECT 113.230 75.520 113.550 75.580 ;
        RECT 114.625 75.535 114.915 75.580 ;
        RECT 90.230 75.240 95.520 75.380 ;
        RECT 95.840 75.240 99.660 75.380 ;
        RECT 90.230 75.180 90.550 75.240 ;
        RECT 84.265 75.040 84.555 75.085 ;
        RECT 83.790 74.900 84.555 75.040 ;
        RECT 83.790 74.840 84.110 74.900 ;
        RECT 84.265 74.855 84.555 74.900 ;
        RECT 84.725 74.855 85.015 75.085 ;
        RECT 85.185 74.855 85.475 75.085 ;
        RECT 88.405 75.040 88.695 75.085 ;
        RECT 89.310 75.040 89.630 75.100 ;
        RECT 88.405 74.900 89.630 75.040 ;
        RECT 88.405 74.855 88.695 74.900 ;
        RECT 78.270 74.560 79.880 74.700 ;
        RECT 85.260 74.700 85.400 74.855 ;
        RECT 89.310 74.840 89.630 74.900 ;
        RECT 91.165 75.040 91.455 75.085 ;
        RECT 92.070 75.040 92.390 75.100 ;
        RECT 91.165 74.900 92.390 75.040 ;
        RECT 91.165 74.855 91.455 74.900 ;
        RECT 92.070 74.840 92.390 74.900 ;
        RECT 95.290 74.840 95.610 75.100 ;
        RECT 95.840 75.085 95.980 75.240 ;
        RECT 95.765 74.855 96.055 75.085 ;
        RECT 96.225 74.855 96.515 75.085 ;
        RECT 97.145 75.040 97.435 75.085 ;
        RECT 97.590 75.040 97.910 75.100 ;
        RECT 99.520 75.085 99.660 75.240 ;
        RECT 97.145 74.900 97.910 75.040 ;
        RECT 97.145 74.855 97.435 74.900 ;
        RECT 86.550 74.700 86.870 74.760 ;
        RECT 85.260 74.560 86.870 74.700 ;
        RECT 78.270 74.500 78.590 74.560 ;
        RECT 65.390 74.360 65.710 74.420 ;
        RECT 81.030 74.360 81.350 74.420 ;
        RECT 85.260 74.360 85.400 74.560 ;
        RECT 86.550 74.500 86.870 74.560 ;
        RECT 87.470 74.500 87.790 74.760 ;
        RECT 90.705 74.700 90.995 74.745 ;
        RECT 91.610 74.700 91.930 74.760 ;
        RECT 90.705 74.560 91.930 74.700 ;
        RECT 90.705 74.515 90.995 74.560 ;
        RECT 91.610 74.500 91.930 74.560 ;
        RECT 92.530 74.700 92.850 74.760 ;
        RECT 95.840 74.700 95.980 74.855 ;
        RECT 92.530 74.560 95.980 74.700 ;
        RECT 92.530 74.500 92.850 74.560 ;
        RECT 65.390 74.220 85.400 74.360 ;
        RECT 88.850 74.360 89.170 74.420 ;
        RECT 89.325 74.360 89.615 74.405 ;
        RECT 88.850 74.220 89.615 74.360 ;
        RECT 96.300 74.360 96.440 74.855 ;
        RECT 97.590 74.840 97.910 74.900 ;
        RECT 98.985 74.855 99.275 75.085 ;
        RECT 99.445 74.855 99.735 75.085 ;
        RECT 99.905 74.855 100.195 75.085 ;
        RECT 96.670 74.700 96.990 74.760 ;
        RECT 99.060 74.700 99.200 74.855 ;
        RECT 96.670 74.560 99.200 74.700 ;
        RECT 99.980 74.700 100.120 74.855 ;
        RECT 100.810 74.840 101.130 75.100 ;
        RECT 102.190 74.840 102.510 75.100 ;
        RECT 114.165 75.040 114.455 75.085 ;
        RECT 113.320 74.900 114.455 75.040 ;
        RECT 112.770 74.700 113.090 74.760 ;
        RECT 99.980 74.560 113.090 74.700 ;
        RECT 96.670 74.500 96.990 74.560 ;
        RECT 112.770 74.500 113.090 74.560 ;
        RECT 113.320 74.420 113.460 74.900 ;
        RECT 114.165 74.855 114.455 74.900 ;
        RECT 115.070 74.500 115.390 74.760 ;
        RECT 113.230 74.360 113.550 74.420 ;
        RECT 96.300 74.220 113.550 74.360 ;
        RECT 65.390 74.160 65.710 74.220 ;
        RECT 81.030 74.160 81.350 74.220 ;
        RECT 88.850 74.160 89.170 74.220 ;
        RECT 89.325 74.175 89.615 74.220 ;
        RECT 113.230 74.160 113.550 74.220 ;
        RECT 28.130 74.020 28.450 74.080 ;
        RECT 25.000 73.880 28.450 74.020 ;
        RECT 28.130 73.820 28.450 73.880 ;
        RECT 35.030 74.020 35.350 74.080 ;
        RECT 63.090 74.020 63.410 74.080 ;
        RECT 35.030 73.880 63.410 74.020 ;
        RECT 35.030 73.820 35.350 73.880 ;
        RECT 63.090 73.820 63.410 73.880 ;
        RECT 71.385 74.020 71.675 74.065 ;
        RECT 71.830 74.020 72.150 74.080 ;
        RECT 71.385 73.880 72.150 74.020 ;
        RECT 71.385 73.835 71.675 73.880 ;
        RECT 71.830 73.820 72.150 73.880 ;
        RECT 80.570 74.020 80.890 74.080 ;
        RECT 87.025 74.020 87.315 74.065 ;
        RECT 80.570 73.880 87.315 74.020 ;
        RECT 80.570 73.820 80.890 73.880 ;
        RECT 87.025 73.835 87.315 73.880 ;
        RECT 91.150 73.820 91.470 74.080 ;
        RECT 97.590 74.020 97.910 74.080 ;
        RECT 100.810 74.020 101.130 74.080 ;
        RECT 97.590 73.880 101.130 74.020 ;
        RECT 97.590 73.820 97.910 73.880 ;
        RECT 100.810 73.820 101.130 73.880 ;
        RECT 101.285 74.020 101.575 74.065 ;
        RECT 101.730 74.020 102.050 74.080 ;
        RECT 101.285 73.880 102.050 74.020 ;
        RECT 101.285 73.835 101.575 73.880 ;
        RECT 101.730 73.820 102.050 73.880 ;
        RECT 5.520 73.200 123.740 73.680 ;
        RECT 15.710 73.000 16.030 73.060 ;
        RECT 16.415 73.000 16.705 73.045 ;
        RECT 15.710 72.860 16.705 73.000 ;
        RECT 15.710 72.800 16.030 72.860 ;
        RECT 16.415 72.815 16.705 72.860 ;
        RECT 23.530 73.000 23.850 73.060 ;
        RECT 24.005 73.000 24.295 73.045 ;
        RECT 23.530 72.860 24.295 73.000 ;
        RECT 23.530 72.800 23.850 72.860 ;
        RECT 24.005 72.815 24.295 72.860 ;
        RECT 30.890 72.800 31.210 73.060 ;
        RECT 35.490 73.000 35.810 73.060 ;
        RECT 36.425 73.000 36.715 73.045 ;
        RECT 35.490 72.860 36.715 73.000 ;
        RECT 35.490 72.800 35.810 72.860 ;
        RECT 36.425 72.815 36.715 72.860 ;
        RECT 53.430 72.800 53.750 73.060 ;
        RECT 53.980 72.860 55.040 73.000 ;
        RECT 7.910 72.660 8.200 72.705 ;
        RECT 9.770 72.660 10.060 72.705 ;
        RECT 12.550 72.660 12.840 72.705 ;
        RECT 7.910 72.520 12.840 72.660 ;
        RECT 7.910 72.475 8.200 72.520 ;
        RECT 9.770 72.475 10.060 72.520 ;
        RECT 12.550 72.475 12.840 72.520 ;
        RECT 24.450 72.660 24.770 72.720 ;
        RECT 27.670 72.660 27.990 72.720 ;
        RECT 52.050 72.660 52.370 72.720 ;
        RECT 53.980 72.660 54.120 72.860 ;
        RECT 24.450 72.520 29.740 72.660 ;
        RECT 24.450 72.460 24.770 72.520 ;
        RECT 7.445 72.320 7.735 72.365 ;
        RECT 8.350 72.320 8.670 72.380 ;
        RECT 7.445 72.180 8.670 72.320 ;
        RECT 7.445 72.135 7.735 72.180 ;
        RECT 8.350 72.120 8.670 72.180 ;
        RECT 8.810 72.320 9.130 72.380 ;
        RECT 9.285 72.320 9.575 72.365 ;
        RECT 8.810 72.180 9.575 72.320 ;
        RECT 8.810 72.120 9.130 72.180 ;
        RECT 9.285 72.135 9.575 72.180 ;
        RECT 12.550 71.980 12.840 72.025 ;
        RECT 10.305 71.840 12.840 71.980 ;
        RECT 10.305 71.685 10.520 71.840 ;
        RECT 12.550 71.795 12.840 71.840 ;
        RECT 13.870 71.980 14.190 72.040 ;
        RECT 25.460 72.025 25.600 72.520 ;
        RECT 27.670 72.460 27.990 72.520 ;
        RECT 28.130 72.320 28.450 72.380 ;
        RECT 29.600 72.320 29.740 72.520 ;
        RECT 50.300 72.520 54.120 72.660 ;
        RECT 25.920 72.180 29.280 72.320 ;
        RECT 25.920 72.025 26.060 72.180 ;
        RECT 28.130 72.120 28.450 72.180 ;
        RECT 18.025 71.980 18.315 72.025 ;
        RECT 13.870 71.840 18.315 71.980 ;
        RECT 13.870 71.780 14.190 71.840 ;
        RECT 18.025 71.795 18.315 71.840 ;
        RECT 25.385 71.795 25.675 72.025 ;
        RECT 25.830 71.795 26.120 72.025 ;
        RECT 26.305 71.980 26.595 72.025 ;
        RECT 26.750 71.980 27.070 72.040 ;
        RECT 26.305 71.840 27.070 71.980 ;
        RECT 26.305 71.795 26.595 71.840 ;
        RECT 26.750 71.780 27.070 71.840 ;
        RECT 27.210 71.980 27.530 72.040 ;
        RECT 27.685 71.980 27.975 72.025 ;
        RECT 27.210 71.840 27.975 71.980 ;
        RECT 27.210 71.780 27.530 71.840 ;
        RECT 27.685 71.795 27.975 71.840 ;
        RECT 28.590 71.780 28.910 72.040 ;
        RECT 29.140 72.025 29.280 72.180 ;
        RECT 29.600 72.180 35.260 72.320 ;
        RECT 29.600 72.025 29.740 72.180 ;
        RECT 35.120 72.040 35.260 72.180 ;
        RECT 29.065 71.795 29.355 72.025 ;
        RECT 29.525 71.795 29.815 72.025 ;
        RECT 8.370 71.640 8.660 71.685 ;
        RECT 10.230 71.640 10.520 71.685 ;
        RECT 8.370 71.500 10.520 71.640 ;
        RECT 8.370 71.455 8.660 71.500 ;
        RECT 10.230 71.455 10.520 71.500 ;
        RECT 11.150 71.640 11.440 71.685 ;
        RECT 13.410 71.640 13.730 71.700 ;
        RECT 14.410 71.640 14.700 71.685 ;
        RECT 11.150 71.500 14.700 71.640 ;
        RECT 11.150 71.455 11.440 71.500 ;
        RECT 13.410 71.440 13.730 71.500 ;
        RECT 14.410 71.455 14.700 71.500 ;
        RECT 21.690 71.640 22.010 71.700 ;
        RECT 23.990 71.640 24.310 71.700 ;
        RECT 21.690 71.500 24.310 71.640 ;
        RECT 29.140 71.640 29.280 71.795 ;
        RECT 33.190 71.780 33.510 72.040 ;
        RECT 34.110 71.780 34.430 72.040 ;
        RECT 34.585 71.795 34.875 72.025 ;
        RECT 34.660 71.640 34.800 71.795 ;
        RECT 35.030 71.780 35.350 72.040 ;
        RECT 38.250 71.980 38.570 72.040 ;
        RECT 50.300 72.025 50.440 72.520 ;
        RECT 52.050 72.460 52.370 72.520 ;
        RECT 51.680 72.180 53.660 72.320 ;
        RECT 48.845 71.980 49.135 72.025 ;
        RECT 38.250 71.840 49.135 71.980 ;
        RECT 38.250 71.780 38.570 71.840 ;
        RECT 48.845 71.795 49.135 71.840 ;
        RECT 50.225 71.795 50.515 72.025 ;
        RECT 50.670 71.980 50.990 72.040 ;
        RECT 51.680 72.025 51.820 72.180 ;
        RECT 51.145 71.980 51.435 72.025 ;
        RECT 50.670 71.840 51.435 71.980 ;
        RECT 50.670 71.780 50.990 71.840 ;
        RECT 51.145 71.795 51.435 71.840 ;
        RECT 51.605 71.795 51.895 72.025 ;
        RECT 52.065 71.980 52.355 72.025 ;
        RECT 52.065 71.795 52.380 71.980 ;
        RECT 35.490 71.640 35.810 71.700 ;
        RECT 29.140 71.500 35.810 71.640 ;
        RECT 21.690 71.440 22.010 71.500 ;
        RECT 23.990 71.440 24.310 71.500 ;
        RECT 35.490 71.440 35.810 71.500 ;
        RECT 17.550 71.100 17.870 71.360 ;
        RECT 22.150 71.300 22.470 71.360 ;
        RECT 25.370 71.300 25.690 71.360 ;
        RECT 22.150 71.160 25.690 71.300 ;
        RECT 22.150 71.100 22.470 71.160 ;
        RECT 25.370 71.100 25.690 71.160 ;
        RECT 49.290 71.100 49.610 71.360 ;
        RECT 52.240 71.300 52.380 71.795 ;
        RECT 53.520 71.640 53.660 72.180 ;
        RECT 53.980 72.025 54.120 72.520 ;
        RECT 54.350 72.460 54.670 72.720 ;
        RECT 54.900 72.660 55.040 72.860 ;
        RECT 57.110 72.800 57.430 73.060 ;
        RECT 57.585 73.000 57.875 73.045 ;
        RECT 58.490 73.000 58.810 73.060 ;
        RECT 57.585 72.860 58.810 73.000 ;
        RECT 57.585 72.815 57.875 72.860 ;
        RECT 58.490 72.800 58.810 72.860 ;
        RECT 64.945 73.000 65.235 73.045 ;
        RECT 74.130 73.000 74.450 73.060 ;
        RECT 64.945 72.860 74.450 73.000 ;
        RECT 64.945 72.815 65.235 72.860 ;
        RECT 74.130 72.800 74.450 72.860 ;
        RECT 92.070 72.800 92.390 73.060 ;
        RECT 61.250 72.660 61.570 72.720 ;
        RECT 54.900 72.520 61.570 72.660 ;
        RECT 61.250 72.460 61.570 72.520 ;
        RECT 99.910 72.660 100.200 72.705 ;
        RECT 101.770 72.660 102.060 72.705 ;
        RECT 104.550 72.660 104.840 72.705 ;
        RECT 99.910 72.520 104.840 72.660 ;
        RECT 99.910 72.475 100.200 72.520 ;
        RECT 101.770 72.475 102.060 72.520 ;
        RECT 104.550 72.475 104.840 72.520 ;
        RECT 54.440 72.320 54.580 72.460 ;
        RECT 68.150 72.320 68.470 72.380 ;
        RECT 54.440 72.180 68.470 72.320 ;
        RECT 53.905 71.795 54.195 72.025 ;
        RECT 54.350 71.980 54.670 72.040 ;
        RECT 55.360 72.025 55.500 72.180 ;
        RECT 54.825 71.980 55.115 72.025 ;
        RECT 54.350 71.840 55.115 71.980 ;
        RECT 54.350 71.780 54.670 71.840 ;
        RECT 54.825 71.795 55.115 71.840 ;
        RECT 55.285 71.795 55.575 72.025 ;
        RECT 55.730 71.980 56.050 72.040 ;
        RECT 58.950 71.980 59.270 72.040 ;
        RECT 55.730 71.840 59.270 71.980 ;
        RECT 55.360 71.640 55.500 71.795 ;
        RECT 55.730 71.780 56.050 71.840 ;
        RECT 58.950 71.780 59.270 71.840 ;
        RECT 59.425 71.780 59.715 72.010 ;
        RECT 59.870 71.780 60.190 72.040 ;
        RECT 53.520 71.500 55.500 71.640 ;
        RECT 55.820 71.300 55.960 71.780 ;
        RECT 59.500 71.640 59.640 71.780 ;
        RECT 60.420 71.640 60.560 72.180 ;
        RECT 68.150 72.120 68.470 72.180 ;
        RECT 74.130 72.120 74.450 72.380 ;
        RECT 99.445 72.320 99.735 72.365 ;
        RECT 110.930 72.320 111.250 72.380 ;
        RECT 99.445 72.180 111.250 72.320 ;
        RECT 99.445 72.135 99.735 72.180 ;
        RECT 110.930 72.120 111.250 72.180 ;
        RECT 112.310 72.320 112.630 72.380 ;
        RECT 113.245 72.320 113.535 72.365 ;
        RECT 115.070 72.320 115.390 72.380 ;
        RECT 112.310 72.180 115.390 72.320 ;
        RECT 112.310 72.120 112.630 72.180 ;
        RECT 113.245 72.135 113.535 72.180 ;
        RECT 115.070 72.120 115.390 72.180 ;
        RECT 60.805 71.980 61.095 72.025 ;
        RECT 61.250 71.980 61.570 72.040 ;
        RECT 60.805 71.840 61.570 71.980 ;
        RECT 60.805 71.795 61.095 71.840 ;
        RECT 61.250 71.780 61.570 71.840 ;
        RECT 64.010 71.980 64.330 72.040 ;
        RECT 66.770 71.980 67.090 72.040 ;
        RECT 67.245 71.980 67.535 72.025 ;
        RECT 64.010 71.840 67.535 71.980 ;
        RECT 64.010 71.780 64.330 71.840 ;
        RECT 66.770 71.780 67.090 71.840 ;
        RECT 67.245 71.795 67.535 71.840 ;
        RECT 59.500 71.500 60.560 71.640 ;
        RECT 63.565 71.455 63.855 71.685 ;
        RECT 68.240 71.640 68.380 72.120 ;
        RECT 73.210 71.780 73.530 72.040 ;
        RECT 76.430 71.980 76.750 72.040 ;
        RECT 88.850 71.980 89.170 72.040 ;
        RECT 76.430 71.840 89.170 71.980 ;
        RECT 76.430 71.780 76.750 71.840 ;
        RECT 88.850 71.780 89.170 71.840 ;
        RECT 89.770 71.780 90.090 72.040 ;
        RECT 90.245 71.795 90.535 72.025 ;
        RECT 90.705 71.980 90.995 72.025 ;
        RECT 91.150 71.980 91.470 72.040 ;
        RECT 95.290 71.980 95.610 72.040 ;
        RECT 90.705 71.840 95.610 71.980 ;
        RECT 90.705 71.795 90.995 71.840 ;
        RECT 90.320 71.640 90.460 71.795 ;
        RECT 91.150 71.780 91.470 71.840 ;
        RECT 95.290 71.780 95.610 71.840 ;
        RECT 101.285 71.980 101.575 72.025 ;
        RECT 101.730 71.980 102.050 72.040 ;
        RECT 104.550 71.980 104.840 72.025 ;
        RECT 101.285 71.840 102.050 71.980 ;
        RECT 101.285 71.795 101.575 71.840 ;
        RECT 101.730 71.780 102.050 71.840 ;
        RECT 102.305 71.840 104.840 71.980 ;
        RECT 92.530 71.640 92.850 71.700 ;
        RECT 102.305 71.685 102.520 71.840 ;
        RECT 104.550 71.795 104.840 71.840 ;
        RECT 110.025 71.980 110.315 72.025 ;
        RECT 110.470 71.980 110.790 72.040 ;
        RECT 113.690 71.980 114.010 72.040 ;
        RECT 110.025 71.840 114.010 71.980 ;
        RECT 110.025 71.795 110.315 71.840 ;
        RECT 110.470 71.780 110.790 71.840 ;
        RECT 113.690 71.780 114.010 71.840 ;
        RECT 114.150 71.980 114.470 72.040 ;
        RECT 114.625 71.980 114.915 72.025 ;
        RECT 117.845 71.980 118.135 72.025 ;
        RECT 114.150 71.840 114.915 71.980 ;
        RECT 114.150 71.780 114.470 71.840 ;
        RECT 114.625 71.795 114.915 71.840 ;
        RECT 116.540 71.840 118.135 71.980 ;
        RECT 68.240 71.500 92.850 71.640 ;
        RECT 52.240 71.160 55.960 71.300 ;
        RECT 59.410 71.300 59.730 71.360 ;
        RECT 63.640 71.300 63.780 71.455 ;
        RECT 92.530 71.440 92.850 71.500 ;
        RECT 100.370 71.640 100.660 71.685 ;
        RECT 102.230 71.640 102.520 71.685 ;
        RECT 100.370 71.500 102.520 71.640 ;
        RECT 100.370 71.455 100.660 71.500 ;
        RECT 102.230 71.455 102.520 71.500 ;
        RECT 103.150 71.640 103.440 71.685 ;
        RECT 106.410 71.640 106.700 71.685 ;
        RECT 109.565 71.640 109.855 71.685 ;
        RECT 103.150 71.500 109.855 71.640 ;
        RECT 103.150 71.455 103.440 71.500 ;
        RECT 106.410 71.455 106.700 71.500 ;
        RECT 109.565 71.455 109.855 71.500 ;
        RECT 59.410 71.160 63.780 71.300 ;
        RECT 65.390 71.300 65.710 71.360 ;
        RECT 68.165 71.300 68.455 71.345 ;
        RECT 65.390 71.160 68.455 71.300 ;
        RECT 59.410 71.100 59.730 71.160 ;
        RECT 65.390 71.100 65.710 71.160 ;
        RECT 68.165 71.115 68.455 71.160 ;
        RECT 71.370 71.100 71.690 71.360 ;
        RECT 73.685 71.300 73.975 71.345 ;
        RECT 78.270 71.300 78.590 71.360 ;
        RECT 73.685 71.160 78.590 71.300 ;
        RECT 73.685 71.115 73.975 71.160 ;
        RECT 78.270 71.100 78.590 71.160 ;
        RECT 102.650 71.300 102.970 71.360 ;
        RECT 104.490 71.300 104.810 71.360 ;
        RECT 108.415 71.300 108.705 71.345 ;
        RECT 102.650 71.160 108.705 71.300 ;
        RECT 102.650 71.100 102.970 71.160 ;
        RECT 104.490 71.100 104.810 71.160 ;
        RECT 108.415 71.115 108.705 71.160 ;
        RECT 113.690 71.300 114.010 71.360 ;
        RECT 116.540 71.345 116.680 71.840 ;
        RECT 117.845 71.795 118.135 71.840 ;
        RECT 114.165 71.300 114.455 71.345 ;
        RECT 113.690 71.160 114.455 71.300 ;
        RECT 113.690 71.100 114.010 71.160 ;
        RECT 114.165 71.115 114.455 71.160 ;
        RECT 116.465 71.115 116.755 71.345 ;
        RECT 116.910 71.100 117.230 71.360 ;
        RECT 5.520 70.480 123.740 70.960 ;
        RECT 17.090 70.080 17.410 70.340 ;
        RECT 21.230 70.280 21.550 70.340 ;
        RECT 24.005 70.280 24.295 70.325 ;
        RECT 35.490 70.280 35.810 70.340 ;
        RECT 59.410 70.280 59.730 70.340 ;
        RECT 60.805 70.280 61.095 70.325 ;
        RECT 21.230 70.140 24.295 70.280 ;
        RECT 21.230 70.080 21.550 70.140 ;
        RECT 24.005 70.095 24.295 70.140 ;
        RECT 25.000 70.140 35.260 70.280 ;
        RECT 12.025 69.940 12.675 69.985 ;
        RECT 15.625 69.940 15.915 69.985 ;
        RECT 17.550 69.940 17.870 70.000 ;
        RECT 25.000 69.940 25.140 70.140 ;
        RECT 27.670 69.940 27.990 70.000 ;
        RECT 12.025 69.800 17.870 69.940 ;
        RECT 12.025 69.755 12.675 69.800 ;
        RECT 15.325 69.755 15.915 69.800 ;
        RECT 8.830 69.600 9.120 69.645 ;
        RECT 10.665 69.600 10.955 69.645 ;
        RECT 14.245 69.600 14.535 69.645 ;
        RECT 8.830 69.460 14.535 69.600 ;
        RECT 8.830 69.415 9.120 69.460 ;
        RECT 10.665 69.415 10.955 69.460 ;
        RECT 14.245 69.415 14.535 69.460 ;
        RECT 15.325 69.440 15.615 69.755 ;
        RECT 17.550 69.740 17.870 69.800 ;
        RECT 22.700 69.800 25.140 69.940 ;
        RECT 25.460 69.800 27.990 69.940 ;
        RECT 35.120 69.940 35.260 70.140 ;
        RECT 35.490 70.140 52.280 70.280 ;
        RECT 35.490 70.080 35.810 70.140 ;
        RECT 44.690 69.940 45.010 70.000 ;
        RECT 35.120 69.800 45.010 69.940 ;
        RECT 18.470 69.600 18.790 69.660 ;
        RECT 19.865 69.600 20.155 69.645 ;
        RECT 18.470 69.460 20.155 69.600 ;
        RECT 18.470 69.400 18.790 69.460 ;
        RECT 19.865 69.415 20.155 69.460 ;
        RECT 8.350 69.060 8.670 69.320 ;
        RECT 9.745 69.260 10.035 69.305 ;
        RECT 11.570 69.260 11.890 69.320 ;
        RECT 9.745 69.120 11.890 69.260 ;
        RECT 9.745 69.075 10.035 69.120 ;
        RECT 11.570 69.060 11.890 69.120 ;
        RECT 18.945 69.260 19.235 69.305 ;
        RECT 22.700 69.260 22.840 69.800 ;
        RECT 25.460 69.645 25.600 69.800 ;
        RECT 27.670 69.740 27.990 69.800 ;
        RECT 44.690 69.740 45.010 69.800 ;
        RECT 45.630 69.940 45.920 69.985 ;
        RECT 47.490 69.940 47.780 69.985 ;
        RECT 45.630 69.800 47.780 69.940 ;
        RECT 45.630 69.755 45.920 69.800 ;
        RECT 47.490 69.755 47.780 69.800 ;
        RECT 48.410 69.940 48.700 69.985 ;
        RECT 49.290 69.940 49.610 70.000 ;
        RECT 51.670 69.940 51.960 69.985 ;
        RECT 48.410 69.800 51.960 69.940 ;
        RECT 52.140 69.940 52.280 70.140 ;
        RECT 59.410 70.140 61.095 70.280 ;
        RECT 59.410 70.080 59.730 70.140 ;
        RECT 60.805 70.095 61.095 70.140 ;
        RECT 61.250 70.280 61.570 70.340 ;
        RECT 64.485 70.280 64.775 70.325 ;
        RECT 76.430 70.280 76.750 70.340 ;
        RECT 61.250 70.140 76.750 70.280 ;
        RECT 61.250 70.080 61.570 70.140 ;
        RECT 64.485 70.095 64.775 70.140 ;
        RECT 76.430 70.080 76.750 70.140 ;
        RECT 78.745 70.280 79.035 70.325 ;
        RECT 82.410 70.280 82.730 70.340 ;
        RECT 83.790 70.280 84.110 70.340 ;
        RECT 78.745 70.140 84.110 70.280 ;
        RECT 78.745 70.095 79.035 70.140 ;
        RECT 82.410 70.080 82.730 70.140 ;
        RECT 83.790 70.080 84.110 70.140 ;
        RECT 89.310 70.280 89.630 70.340 ;
        RECT 90.705 70.280 90.995 70.325 ;
        RECT 89.310 70.140 90.995 70.280 ;
        RECT 89.310 70.080 89.630 70.140 ;
        RECT 90.705 70.095 90.995 70.140 ;
        RECT 93.910 70.280 94.230 70.340 ;
        RECT 94.385 70.280 94.675 70.325 ;
        RECT 99.890 70.280 100.210 70.340 ;
        RECT 93.910 70.140 94.675 70.280 ;
        RECT 93.910 70.080 94.230 70.140 ;
        RECT 94.385 70.095 94.675 70.140 ;
        RECT 95.840 70.140 100.210 70.280 ;
        RECT 90.230 69.940 90.550 70.000 ;
        RECT 52.140 69.800 61.020 69.940 ;
        RECT 48.410 69.755 48.700 69.800 ;
        RECT 25.385 69.415 25.675 69.645 ;
        RECT 25.830 69.400 26.150 69.660 ;
        RECT 26.305 69.415 26.595 69.645 ;
        RECT 18.945 69.120 22.840 69.260 ;
        RECT 23.070 69.260 23.390 69.320 ;
        RECT 26.380 69.260 26.520 69.415 ;
        RECT 27.210 69.400 27.530 69.660 ;
        RECT 37.790 69.400 38.110 69.660 ;
        RECT 38.250 69.600 38.570 69.660 ;
        RECT 41.025 69.600 41.315 69.645 ;
        RECT 47.565 69.600 47.780 69.755 ;
        RECT 49.290 69.740 49.610 69.800 ;
        RECT 51.670 69.755 51.960 69.800 ;
        RECT 53.430 69.645 53.750 69.660 ;
        RECT 49.810 69.600 50.100 69.645 ;
        RECT 38.250 69.460 41.315 69.600 ;
        RECT 38.250 69.400 38.570 69.460 ;
        RECT 41.025 69.415 41.315 69.460 ;
        RECT 42.480 69.460 47.220 69.600 ;
        RECT 47.565 69.460 50.100 69.600 ;
        RECT 23.070 69.120 26.520 69.260 ;
        RECT 27.300 69.260 27.440 69.400 ;
        RECT 33.190 69.260 33.510 69.320 ;
        RECT 42.480 69.260 42.620 69.460 ;
        RECT 27.300 69.120 42.620 69.260 ;
        RECT 42.850 69.260 43.170 69.320 ;
        RECT 44.705 69.260 44.995 69.305 ;
        RECT 42.850 69.120 44.995 69.260 ;
        RECT 18.945 69.075 19.235 69.120 ;
        RECT 23.070 69.060 23.390 69.120 ;
        RECT 33.190 69.060 33.510 69.120 ;
        RECT 42.850 69.060 43.170 69.120 ;
        RECT 44.705 69.075 44.995 69.120 ;
        RECT 46.530 69.060 46.850 69.320 ;
        RECT 47.080 69.260 47.220 69.460 ;
        RECT 49.810 69.415 50.100 69.460 ;
        RECT 53.430 69.600 53.965 69.645 ;
        RECT 59.870 69.600 60.190 69.660 ;
        RECT 53.430 69.460 60.190 69.600 ;
        RECT 53.430 69.415 53.965 69.460 ;
        RECT 53.430 69.400 53.750 69.415 ;
        RECT 59.870 69.400 60.190 69.460 ;
        RECT 60.330 69.260 60.650 69.320 ;
        RECT 47.080 69.120 60.650 69.260 ;
        RECT 60.880 69.260 61.020 69.800 ;
        RECT 61.340 69.800 67.920 69.940 ;
        RECT 61.340 69.645 61.480 69.800 ;
        RECT 65.480 69.660 65.620 69.800 ;
        RECT 61.265 69.415 61.555 69.645 ;
        RECT 61.725 69.600 62.015 69.645 ;
        RECT 62.170 69.600 62.490 69.660 ;
        RECT 61.725 69.460 62.490 69.600 ;
        RECT 61.725 69.415 62.015 69.460 ;
        RECT 62.170 69.400 62.490 69.460 ;
        RECT 63.105 69.600 63.395 69.645 ;
        RECT 64.010 69.600 64.330 69.660 ;
        RECT 63.105 69.460 64.330 69.600 ;
        RECT 63.105 69.415 63.395 69.460 ;
        RECT 64.010 69.400 64.330 69.460 ;
        RECT 65.390 69.400 65.710 69.660 ;
        RECT 65.850 69.400 66.170 69.660 ;
        RECT 67.780 69.645 67.920 69.800 ;
        RECT 70.540 69.800 90.550 69.940 ;
        RECT 67.705 69.415 67.995 69.645 ;
        RECT 68.610 69.600 68.930 69.660 ;
        RECT 69.545 69.600 69.835 69.645 ;
        RECT 68.610 69.460 69.835 69.600 ;
        RECT 68.610 69.400 68.930 69.460 ;
        RECT 69.545 69.415 69.835 69.460 ;
        RECT 62.645 69.260 62.935 69.305 ;
        RECT 65.940 69.260 66.080 69.400 ;
        RECT 60.880 69.120 62.400 69.260 ;
        RECT 60.330 69.060 60.650 69.120 ;
        RECT 9.235 68.920 9.525 68.965 ;
        RECT 11.125 68.920 11.415 68.965 ;
        RECT 14.245 68.920 14.535 68.965 ;
        RECT 9.235 68.780 14.535 68.920 ;
        RECT 9.235 68.735 9.525 68.780 ;
        RECT 11.125 68.735 11.415 68.780 ;
        RECT 14.245 68.735 14.535 68.780 ;
        RECT 25.830 68.920 26.150 68.980 ;
        RECT 28.130 68.920 28.450 68.980 ;
        RECT 25.830 68.780 28.450 68.920 ;
        RECT 25.830 68.720 26.150 68.780 ;
        RECT 28.130 68.720 28.450 68.780 ;
        RECT 45.170 68.920 45.460 68.965 ;
        RECT 47.030 68.920 47.320 68.965 ;
        RECT 49.810 68.920 50.100 68.965 ;
        RECT 45.170 68.780 50.100 68.920 ;
        RECT 62.260 68.920 62.400 69.120 ;
        RECT 62.645 69.120 66.080 69.260 ;
        RECT 62.645 69.075 62.935 69.120 ;
        RECT 67.690 68.920 68.010 68.980 ;
        RECT 68.625 68.920 68.915 68.965 ;
        RECT 62.260 68.780 67.460 68.920 ;
        RECT 45.170 68.735 45.460 68.780 ;
        RECT 47.030 68.735 47.320 68.780 ;
        RECT 49.810 68.735 50.100 68.780 ;
        RECT 36.410 68.580 36.730 68.640 ;
        RECT 36.885 68.580 37.175 68.625 ;
        RECT 36.410 68.440 37.175 68.580 ;
        RECT 36.410 68.380 36.730 68.440 ;
        RECT 36.885 68.395 37.175 68.440 ;
        RECT 39.170 68.580 39.490 68.640 ;
        RECT 40.565 68.580 40.855 68.625 ;
        RECT 39.170 68.440 40.855 68.580 ;
        RECT 39.170 68.380 39.490 68.440 ;
        RECT 40.565 68.395 40.855 68.440 ;
        RECT 62.170 68.580 62.490 68.640 ;
        RECT 64.930 68.580 65.250 68.640 ;
        RECT 62.170 68.440 65.250 68.580 ;
        RECT 62.170 68.380 62.490 68.440 ;
        RECT 64.930 68.380 65.250 68.440 ;
        RECT 66.310 68.580 66.630 68.640 ;
        RECT 66.785 68.580 67.075 68.625 ;
        RECT 66.310 68.440 67.075 68.580 ;
        RECT 67.320 68.580 67.460 68.780 ;
        RECT 67.690 68.780 68.915 68.920 ;
        RECT 67.690 68.720 68.010 68.780 ;
        RECT 68.625 68.735 68.915 68.780 ;
        RECT 70.540 68.625 70.680 69.800 ;
        RECT 90.230 69.740 90.550 69.800 ;
        RECT 92.620 69.800 94.600 69.940 ;
        RECT 92.620 69.660 92.760 69.800 ;
        RECT 71.370 69.400 71.690 69.660 ;
        RECT 78.270 69.400 78.590 69.660 ;
        RECT 81.505 69.600 81.795 69.645 ;
        RECT 81.950 69.600 82.270 69.660 ;
        RECT 81.505 69.460 82.270 69.600 ;
        RECT 81.505 69.415 81.795 69.460 ;
        RECT 81.950 69.400 82.270 69.460 ;
        RECT 91.150 69.600 91.470 69.660 ;
        RECT 92.085 69.600 92.375 69.645 ;
        RECT 91.150 69.460 92.375 69.600 ;
        RECT 91.150 69.400 91.470 69.460 ;
        RECT 92.085 69.415 92.375 69.460 ;
        RECT 92.530 69.400 92.850 69.660 ;
        RECT 93.005 69.600 93.295 69.645 ;
        RECT 93.450 69.600 93.770 69.660 ;
        RECT 93.005 69.460 93.770 69.600 ;
        RECT 93.005 69.415 93.295 69.460 ;
        RECT 93.450 69.400 93.770 69.460 ;
        RECT 93.910 69.400 94.230 69.660 ;
        RECT 79.205 69.075 79.495 69.305 ;
        RECT 94.460 69.260 94.600 69.800 ;
        RECT 95.290 69.600 95.610 69.660 ;
        RECT 95.840 69.645 95.980 70.140 ;
        RECT 99.890 70.080 100.210 70.140 ;
        RECT 101.745 70.280 102.035 70.325 ;
        RECT 102.190 70.280 102.510 70.340 ;
        RECT 101.745 70.140 102.510 70.280 ;
        RECT 101.745 70.095 102.035 70.140 ;
        RECT 102.190 70.080 102.510 70.140 ;
        RECT 103.585 70.280 103.875 70.325 ;
        RECT 113.690 70.280 114.010 70.340 ;
        RECT 120.375 70.280 120.665 70.325 ;
        RECT 103.585 70.140 120.665 70.280 ;
        RECT 103.585 70.095 103.875 70.140 ;
        RECT 103.660 69.940 103.800 70.095 ;
        RECT 113.690 70.080 114.010 70.140 ;
        RECT 120.375 70.095 120.665 70.140 ;
        RECT 96.300 69.800 98.740 69.940 ;
        RECT 96.300 69.645 96.440 69.800 ;
        RECT 95.765 69.600 96.055 69.645 ;
        RECT 95.290 69.460 96.055 69.600 ;
        RECT 95.290 69.400 95.610 69.460 ;
        RECT 95.765 69.415 96.055 69.460 ;
        RECT 96.225 69.415 96.515 69.645 ;
        RECT 96.300 69.260 96.440 69.415 ;
        RECT 96.670 69.400 96.990 69.660 ;
        RECT 97.590 69.400 97.910 69.660 ;
        RECT 98.065 69.415 98.355 69.645 ;
        RECT 94.460 69.120 96.440 69.260 ;
        RECT 97.130 69.260 97.450 69.320 ;
        RECT 98.140 69.260 98.280 69.415 ;
        RECT 97.130 69.120 98.280 69.260 ;
        RECT 98.600 69.260 98.740 69.800 ;
        RECT 99.060 69.800 103.800 69.940 ;
        RECT 99.060 69.645 99.200 69.800 ;
        RECT 104.030 69.740 104.350 70.000 ;
        RECT 112.330 69.940 112.620 69.985 ;
        RECT 114.190 69.940 114.480 69.985 ;
        RECT 112.330 69.800 114.480 69.940 ;
        RECT 112.330 69.755 112.620 69.800 ;
        RECT 114.190 69.755 114.480 69.800 ;
        RECT 115.110 69.940 115.400 69.985 ;
        RECT 117.370 69.940 117.690 70.000 ;
        RECT 118.370 69.940 118.660 69.985 ;
        RECT 115.110 69.800 118.660 69.940 ;
        RECT 115.110 69.755 115.400 69.800 ;
        RECT 98.985 69.415 99.275 69.645 ;
        RECT 99.445 69.415 99.735 69.645 ;
        RECT 99.520 69.260 99.660 69.415 ;
        RECT 99.890 69.400 100.210 69.660 ;
        RECT 104.120 69.600 104.260 69.740 ;
        RECT 101.360 69.460 104.260 69.600 ;
        RECT 110.930 69.600 111.250 69.660 ;
        RECT 111.405 69.600 111.695 69.645 ;
        RECT 110.930 69.460 111.695 69.600 ;
        RECT 114.265 69.600 114.480 69.755 ;
        RECT 117.370 69.740 117.690 69.800 ;
        RECT 118.370 69.755 118.660 69.800 ;
        RECT 116.510 69.600 116.800 69.645 ;
        RECT 114.265 69.460 116.800 69.600 ;
        RECT 101.360 69.305 101.500 69.460 ;
        RECT 110.930 69.400 111.250 69.460 ;
        RECT 111.405 69.415 111.695 69.460 ;
        RECT 116.510 69.415 116.800 69.460 ;
        RECT 98.600 69.120 99.660 69.260 ;
        RECT 74.130 68.920 74.450 68.980 ;
        RECT 79.280 68.920 79.420 69.075 ;
        RECT 97.130 69.060 97.450 69.120 ;
        RECT 101.285 69.075 101.575 69.305 ;
        RECT 103.110 69.260 103.430 69.320 ;
        RECT 104.045 69.260 104.335 69.305 ;
        RECT 104.490 69.260 104.810 69.320 ;
        RECT 103.110 69.120 104.810 69.260 ;
        RECT 103.110 69.060 103.430 69.120 ;
        RECT 104.045 69.075 104.335 69.120 ;
        RECT 104.490 69.060 104.810 69.120 ;
        RECT 104.965 69.075 105.255 69.305 ;
        RECT 113.245 69.260 113.535 69.305 ;
        RECT 116.910 69.260 117.230 69.320 ;
        RECT 113.245 69.120 117.230 69.260 ;
        RECT 113.245 69.075 113.535 69.120 ;
        RECT 74.130 68.780 79.420 68.920 ;
        RECT 88.850 68.920 89.170 68.980 ;
        RECT 93.910 68.920 94.230 68.980 ;
        RECT 97.590 68.920 97.910 68.980 ;
        RECT 88.850 68.780 97.910 68.920 ;
        RECT 105.040 68.920 105.180 69.075 ;
        RECT 116.910 69.060 117.230 69.120 ;
        RECT 105.410 68.920 105.730 68.980 ;
        RECT 105.040 68.780 105.730 68.920 ;
        RECT 74.130 68.720 74.450 68.780 ;
        RECT 88.850 68.720 89.170 68.780 ;
        RECT 93.910 68.720 94.230 68.780 ;
        RECT 97.590 68.720 97.910 68.780 ;
        RECT 105.410 68.720 105.730 68.780 ;
        RECT 111.870 68.920 112.160 68.965 ;
        RECT 113.730 68.920 114.020 68.965 ;
        RECT 116.510 68.920 116.800 68.965 ;
        RECT 111.870 68.780 116.800 68.920 ;
        RECT 111.870 68.735 112.160 68.780 ;
        RECT 113.730 68.735 114.020 68.780 ;
        RECT 116.510 68.735 116.800 68.780 ;
        RECT 70.465 68.580 70.755 68.625 ;
        RECT 67.320 68.440 70.755 68.580 ;
        RECT 66.310 68.380 66.630 68.440 ;
        RECT 66.785 68.395 67.075 68.440 ;
        RECT 70.465 68.395 70.755 68.440 ;
        RECT 72.290 68.380 72.610 68.640 ;
        RECT 76.430 68.380 76.750 68.640 ;
        RECT 80.570 68.580 80.890 68.640 ;
        RECT 81.045 68.580 81.335 68.625 ;
        RECT 80.570 68.440 81.335 68.580 ;
        RECT 80.570 68.380 80.890 68.440 ;
        RECT 81.045 68.395 81.335 68.440 ;
        RECT 5.520 67.760 123.740 68.240 ;
        RECT 38.710 67.560 39.030 67.620 ;
        RECT 33.280 67.420 39.030 67.560 ;
        RECT 28.590 66.880 28.910 66.940 ;
        RECT 32.745 66.880 33.035 66.925 ;
        RECT 33.280 66.880 33.420 67.420 ;
        RECT 38.710 67.360 39.030 67.420 ;
        RECT 46.530 67.560 46.850 67.620 ;
        RECT 47.465 67.560 47.755 67.605 ;
        RECT 46.530 67.420 47.755 67.560 ;
        RECT 46.530 67.360 46.850 67.420 ;
        RECT 47.465 67.375 47.755 67.420 ;
        RECT 58.950 67.560 59.270 67.620 ;
        RECT 63.105 67.560 63.395 67.605 ;
        RECT 58.950 67.420 63.395 67.560 ;
        RECT 58.950 67.360 59.270 67.420 ;
        RECT 63.105 67.375 63.395 67.420 ;
        RECT 64.945 67.375 65.235 67.605 ;
        RECT 35.050 67.220 35.340 67.265 ;
        RECT 36.910 67.220 37.200 67.265 ;
        RECT 39.690 67.220 39.980 67.265 ;
        RECT 35.050 67.080 39.980 67.220 ;
        RECT 35.050 67.035 35.340 67.080 ;
        RECT 36.910 67.035 37.200 67.080 ;
        RECT 39.690 67.035 39.980 67.080 ;
        RECT 48.845 67.035 49.135 67.265 ;
        RECT 62.170 67.220 62.490 67.280 ;
        RECT 65.020 67.220 65.160 67.375 ;
        RECT 68.150 67.360 68.470 67.620 ;
        RECT 76.430 67.560 76.750 67.620 ;
        RECT 72.840 67.420 76.750 67.560 ;
        RECT 62.170 67.080 65.160 67.220 ;
        RECT 28.590 66.740 31.580 66.880 ;
        RECT 28.590 66.680 28.910 66.740 ;
        RECT 31.440 66.585 31.580 66.740 ;
        RECT 32.745 66.740 33.420 66.880 ;
        RECT 32.745 66.695 33.035 66.740 ;
        RECT 34.570 66.680 34.890 66.940 ;
        RECT 36.410 66.680 36.730 66.940 ;
        RECT 29.065 66.540 29.355 66.585 ;
        RECT 29.065 66.400 29.740 66.540 ;
        RECT 29.065 66.355 29.355 66.400 ;
        RECT 28.130 65.660 28.450 65.920 ;
        RECT 29.600 65.905 29.740 66.400 ;
        RECT 31.365 66.355 31.655 66.585 ;
        RECT 31.825 66.540 32.115 66.585 ;
        RECT 34.110 66.540 34.430 66.600 ;
        RECT 39.690 66.540 39.980 66.585 ;
        RECT 31.825 66.400 34.430 66.540 ;
        RECT 31.825 66.355 32.115 66.400 ;
        RECT 34.110 66.340 34.430 66.400 ;
        RECT 37.445 66.400 39.980 66.540 ;
        RECT 37.445 66.245 37.660 66.400 ;
        RECT 39.690 66.355 39.980 66.400 ;
        RECT 48.385 66.540 48.675 66.585 ;
        RECT 48.920 66.540 49.060 67.035 ;
        RECT 62.170 67.020 62.490 67.080 ;
        RECT 52.050 66.680 52.370 66.940 ;
        RECT 48.385 66.400 49.060 66.540 ;
        RECT 48.385 66.355 48.675 66.400 ;
        RECT 50.670 66.340 50.990 66.600 ;
        RECT 51.145 66.540 51.435 66.585 ;
        RECT 53.430 66.540 53.750 66.600 ;
        RECT 51.145 66.400 53.750 66.540 ;
        RECT 51.145 66.355 51.435 66.400 ;
        RECT 53.430 66.340 53.750 66.400 ;
        RECT 64.010 66.340 64.330 66.600 ;
        RECT 65.390 66.540 65.710 66.600 ;
        RECT 65.865 66.540 66.155 66.585 ;
        RECT 65.390 66.400 66.155 66.540 ;
        RECT 65.390 66.340 65.710 66.400 ;
        RECT 65.865 66.355 66.155 66.400 ;
        RECT 69.085 66.355 69.375 66.585 ;
        RECT 72.305 66.540 72.595 66.585 ;
        RECT 72.840 66.540 72.980 67.420 ;
        RECT 76.430 67.360 76.750 67.420 ;
        RECT 82.410 67.605 82.730 67.620 ;
        RECT 82.410 67.375 82.945 67.605 ;
        RECT 82.410 67.360 82.730 67.375 ;
        RECT 117.370 67.360 117.690 67.620 ;
        RECT 74.150 67.220 74.440 67.265 ;
        RECT 76.010 67.220 76.300 67.265 ;
        RECT 78.790 67.220 79.080 67.265 ;
        RECT 74.150 67.080 79.080 67.220 ;
        RECT 74.150 67.035 74.440 67.080 ;
        RECT 76.010 67.035 76.300 67.080 ;
        RECT 78.790 67.035 79.080 67.080 ;
        RECT 73.685 66.880 73.975 66.925 ;
        RECT 81.950 66.880 82.270 66.940 ;
        RECT 84.265 66.880 84.555 66.925 ;
        RECT 73.685 66.740 76.200 66.880 ;
        RECT 73.685 66.695 73.975 66.740 ;
        RECT 76.060 66.600 76.200 66.740 ;
        RECT 81.950 66.740 84.555 66.880 ;
        RECT 81.950 66.680 82.270 66.740 ;
        RECT 84.265 66.695 84.555 66.740 ;
        RECT 89.770 66.880 90.090 66.940 ;
        RECT 92.530 66.880 92.850 66.940 ;
        RECT 89.770 66.740 92.850 66.880 ;
        RECT 89.770 66.680 90.090 66.740 ;
        RECT 92.530 66.680 92.850 66.740 ;
        RECT 92.990 66.880 93.310 66.940 ;
        RECT 93.465 66.880 93.755 66.925 ;
        RECT 105.410 66.880 105.730 66.940 ;
        RECT 112.310 66.880 112.630 66.940 ;
        RECT 113.245 66.880 113.535 66.925 ;
        RECT 92.990 66.740 113.535 66.880 ;
        RECT 92.990 66.680 93.310 66.740 ;
        RECT 93.465 66.695 93.755 66.740 ;
        RECT 105.410 66.680 105.730 66.740 ;
        RECT 112.310 66.680 112.630 66.740 ;
        RECT 113.245 66.695 113.535 66.740 ;
        RECT 75.525 66.540 75.815 66.585 ;
        RECT 72.305 66.400 72.980 66.540 ;
        RECT 73.300 66.400 75.815 66.540 ;
        RECT 72.305 66.355 72.595 66.400 ;
        RECT 35.510 66.200 35.800 66.245 ;
        RECT 37.370 66.200 37.660 66.245 ;
        RECT 35.510 66.060 37.660 66.200 ;
        RECT 35.510 66.015 35.800 66.060 ;
        RECT 37.370 66.015 37.660 66.060 ;
        RECT 38.290 66.200 38.580 66.245 ;
        RECT 39.170 66.200 39.490 66.260 ;
        RECT 41.550 66.200 41.840 66.245 ;
        RECT 38.290 66.060 41.840 66.200 ;
        RECT 38.290 66.015 38.580 66.060 ;
        RECT 39.170 66.000 39.490 66.060 ;
        RECT 41.550 66.015 41.840 66.060 ;
        RECT 42.390 66.200 42.710 66.260 ;
        RECT 43.555 66.200 43.845 66.245 ;
        RECT 50.760 66.200 50.900 66.340 ;
        RECT 42.390 66.060 50.900 66.200 ;
        RECT 64.470 66.200 64.790 66.260 ;
        RECT 68.610 66.200 68.930 66.260 ;
        RECT 69.160 66.200 69.300 66.355 ;
        RECT 64.470 66.060 69.300 66.200 ;
        RECT 42.390 66.000 42.710 66.060 ;
        RECT 43.555 66.015 43.845 66.060 ;
        RECT 64.470 66.000 64.790 66.060 ;
        RECT 68.610 66.000 68.930 66.060 ;
        RECT 73.300 65.905 73.440 66.400 ;
        RECT 75.525 66.355 75.815 66.400 ;
        RECT 75.970 66.340 76.290 66.600 ;
        RECT 78.790 66.540 79.080 66.585 ;
        RECT 76.545 66.400 79.080 66.540 ;
        RECT 76.545 66.245 76.760 66.400 ;
        RECT 78.790 66.355 79.080 66.400 ;
        RECT 83.330 66.340 83.650 66.600 ;
        RECT 92.085 66.540 92.375 66.585 ;
        RECT 103.110 66.540 103.430 66.600 ;
        RECT 92.085 66.400 103.430 66.540 ;
        RECT 92.085 66.355 92.375 66.400 ;
        RECT 103.110 66.340 103.430 66.400 ;
        RECT 110.470 66.540 110.790 66.600 ;
        RECT 117.845 66.540 118.135 66.585 ;
        RECT 110.470 66.400 118.135 66.540 ;
        RECT 110.470 66.340 110.790 66.400 ;
        RECT 117.845 66.355 118.135 66.400 ;
        RECT 80.570 66.245 80.890 66.260 ;
        RECT 74.610 66.200 74.900 66.245 ;
        RECT 76.470 66.200 76.760 66.245 ;
        RECT 74.610 66.060 76.760 66.200 ;
        RECT 74.610 66.015 74.900 66.060 ;
        RECT 76.470 66.015 76.760 66.060 ;
        RECT 77.390 66.200 77.680 66.245 ;
        RECT 80.570 66.200 80.940 66.245 ;
        RECT 77.390 66.060 80.940 66.200 ;
        RECT 77.390 66.015 77.680 66.060 ;
        RECT 80.570 66.015 80.940 66.060 ;
        RECT 113.230 66.200 113.550 66.260 ;
        RECT 114.165 66.200 114.455 66.245 ;
        RECT 116.910 66.200 117.230 66.260 ;
        RECT 113.230 66.060 114.455 66.200 ;
        RECT 80.570 66.000 80.890 66.015 ;
        RECT 113.230 66.000 113.550 66.060 ;
        RECT 114.165 66.015 114.455 66.060 ;
        RECT 114.700 66.060 117.230 66.200 ;
        RECT 29.525 65.675 29.815 65.905 ;
        RECT 73.225 65.675 73.515 65.905 ;
        RECT 87.930 65.860 88.250 65.920 ;
        RECT 90.245 65.860 90.535 65.905 ;
        RECT 87.930 65.720 90.535 65.860 ;
        RECT 87.930 65.660 88.250 65.720 ;
        RECT 90.245 65.675 90.535 65.720 ;
        RECT 112.770 65.860 113.090 65.920 ;
        RECT 114.700 65.905 114.840 66.060 ;
        RECT 116.910 66.000 117.230 66.060 ;
        RECT 114.625 65.860 114.915 65.905 ;
        RECT 112.770 65.720 114.915 65.860 ;
        RECT 112.770 65.660 113.090 65.720 ;
        RECT 114.625 65.675 114.915 65.720 ;
        RECT 116.465 65.860 116.755 65.905 ;
        RECT 119.670 65.860 119.990 65.920 ;
        RECT 116.465 65.720 119.990 65.860 ;
        RECT 116.465 65.675 116.755 65.720 ;
        RECT 119.670 65.660 119.990 65.720 ;
        RECT 5.520 65.040 123.740 65.520 ;
        RECT 23.070 64.640 23.390 64.900 ;
        RECT 26.750 64.840 27.070 64.900 ;
        RECT 27.685 64.840 27.975 64.885 ;
        RECT 26.750 64.700 27.975 64.840 ;
        RECT 26.750 64.640 27.070 64.700 ;
        RECT 27.685 64.655 27.975 64.700 ;
        RECT 28.145 64.840 28.435 64.885 ;
        RECT 28.590 64.840 28.910 64.900 ;
        RECT 28.145 64.700 28.910 64.840 ;
        RECT 28.145 64.655 28.435 64.700 ;
        RECT 28.590 64.640 28.910 64.700 ;
        RECT 36.885 64.840 37.175 64.885 ;
        RECT 37.790 64.840 38.110 64.900 ;
        RECT 36.885 64.700 38.110 64.840 ;
        RECT 36.885 64.655 37.175 64.700 ;
        RECT 37.790 64.640 38.110 64.700 ;
        RECT 39.185 64.840 39.475 64.885 ;
        RECT 42.390 64.840 42.710 64.900 ;
        RECT 39.185 64.700 42.710 64.840 ;
        RECT 39.185 64.655 39.475 64.700 ;
        RECT 42.390 64.640 42.710 64.700 ;
        RECT 53.430 64.640 53.750 64.900 ;
        RECT 53.890 64.640 54.210 64.900 ;
        RECT 63.090 64.840 63.410 64.900 ;
        RECT 66.785 64.840 67.075 64.885 ;
        RECT 75.970 64.840 76.290 64.900 ;
        RECT 63.090 64.700 70.220 64.840 ;
        RECT 63.090 64.640 63.410 64.700 ;
        RECT 66.785 64.655 67.075 64.700 ;
        RECT 13.870 64.500 14.190 64.560 ;
        RECT 14.805 64.500 15.095 64.545 ;
        RECT 17.550 64.500 17.870 64.560 ;
        RECT 13.870 64.360 17.870 64.500 ;
        RECT 13.870 64.300 14.190 64.360 ;
        RECT 14.805 64.315 15.095 64.360 ;
        RECT 17.550 64.300 17.870 64.360 ;
        RECT 18.010 64.500 18.330 64.560 ;
        RECT 19.405 64.500 19.695 64.545 ;
        RECT 26.840 64.500 26.980 64.640 ;
        RECT 18.010 64.360 26.980 64.500 ;
        RECT 34.110 64.500 34.430 64.560 ;
        RECT 36.410 64.500 36.730 64.560 ;
        RECT 38.725 64.500 39.015 64.545 ;
        RECT 34.110 64.360 39.015 64.500 ;
        RECT 18.010 64.300 18.330 64.360 ;
        RECT 19.405 64.315 19.695 64.360 ;
        RECT 34.110 64.300 34.430 64.360 ;
        RECT 36.410 64.300 36.730 64.360 ;
        RECT 38.725 64.315 39.015 64.360 ;
        RECT 12.965 63.975 13.255 64.205 ;
        RECT 13.410 64.160 13.730 64.220 ;
        RECT 18.470 64.160 18.790 64.220 ;
        RECT 13.410 64.020 18.790 64.160 ;
        RECT 13.040 63.480 13.180 63.975 ;
        RECT 13.410 63.960 13.730 64.020 ;
        RECT 18.470 63.960 18.790 64.020 ;
        RECT 18.945 64.160 19.235 64.205 ;
        RECT 22.150 64.160 22.470 64.220 ;
        RECT 23.545 64.160 23.835 64.205 ;
        RECT 31.825 64.160 32.115 64.205 ;
        RECT 38.250 64.160 38.570 64.220 ;
        RECT 18.945 64.020 23.835 64.160 ;
        RECT 18.945 63.975 19.235 64.020 ;
        RECT 16.630 63.820 16.950 63.880 ;
        RECT 19.020 63.820 19.160 63.975 ;
        RECT 22.150 63.960 22.470 64.020 ;
        RECT 23.545 63.975 23.835 64.020 ;
        RECT 25.000 64.020 38.570 64.160 ;
        RECT 16.630 63.680 19.160 63.820 ;
        RECT 20.325 63.820 20.615 63.865 ;
        RECT 24.450 63.820 24.770 63.880 ;
        RECT 20.325 63.680 24.770 63.820 ;
        RECT 16.630 63.620 16.950 63.680 ;
        RECT 20.325 63.635 20.615 63.680 ;
        RECT 24.450 63.620 24.770 63.680 ;
        RECT 17.105 63.480 17.395 63.525 ;
        RECT 13.040 63.340 17.395 63.480 ;
        RECT 17.105 63.295 17.395 63.340 ;
        RECT 17.550 63.480 17.870 63.540 ;
        RECT 25.000 63.480 25.140 64.020 ;
        RECT 31.825 63.975 32.115 64.020 ;
        RECT 38.250 63.960 38.570 64.020 ;
        RECT 51.145 64.160 51.435 64.205 ;
        RECT 64.010 64.160 64.330 64.220 ;
        RECT 64.930 64.160 65.250 64.220 ;
        RECT 65.865 64.160 66.155 64.205 ;
        RECT 51.145 64.020 51.820 64.160 ;
        RECT 51.145 63.975 51.435 64.020 ;
        RECT 25.370 63.820 25.690 63.880 ;
        RECT 29.065 63.820 29.355 63.865 ;
        RECT 39.170 63.820 39.490 63.880 ;
        RECT 39.645 63.820 39.935 63.865 ;
        RECT 25.370 63.680 39.935 63.820 ;
        RECT 25.370 63.620 25.690 63.680 ;
        RECT 29.065 63.635 29.355 63.680 ;
        RECT 39.170 63.620 39.490 63.680 ;
        RECT 39.645 63.635 39.935 63.680 ;
        RECT 17.550 63.340 25.140 63.480 ;
        RECT 30.430 63.480 30.750 63.540 ;
        RECT 34.570 63.480 34.890 63.540 ;
        RECT 42.850 63.480 43.170 63.540 ;
        RECT 51.680 63.525 51.820 64.020 ;
        RECT 64.010 64.020 66.155 64.160 ;
        RECT 64.010 63.960 64.330 64.020 ;
        RECT 64.930 63.960 65.250 64.020 ;
        RECT 65.865 63.975 66.155 64.020 ;
        RECT 67.705 63.975 67.995 64.205 ;
        RECT 52.050 63.820 52.370 63.880 ;
        RECT 53.430 63.820 53.750 63.880 ;
        RECT 54.365 63.820 54.655 63.865 ;
        RECT 52.050 63.680 54.655 63.820 ;
        RECT 52.050 63.620 52.370 63.680 ;
        RECT 53.430 63.620 53.750 63.680 ;
        RECT 54.365 63.635 54.655 63.680 ;
        RECT 65.390 63.820 65.710 63.880 ;
        RECT 67.780 63.820 67.920 63.975 ;
        RECT 65.390 63.680 67.920 63.820 ;
        RECT 70.080 63.820 70.220 64.700 ;
        RECT 70.540 64.700 76.290 64.840 ;
        RECT 70.540 64.205 70.680 64.700 ;
        RECT 75.970 64.640 76.290 64.700 ;
        RECT 78.270 64.840 78.590 64.900 ;
        RECT 79.205 64.840 79.495 64.885 ;
        RECT 78.270 64.700 79.495 64.840 ;
        RECT 78.270 64.640 78.590 64.700 ;
        RECT 79.205 64.655 79.495 64.700 ;
        RECT 92.530 64.840 92.850 64.900 ;
        RECT 93.925 64.840 94.215 64.885 ;
        RECT 92.530 64.700 94.215 64.840 ;
        RECT 92.530 64.640 92.850 64.700 ;
        RECT 93.925 64.655 94.215 64.700 ;
        RECT 96.670 64.840 96.990 64.900 ;
        RECT 102.665 64.840 102.955 64.885 ;
        RECT 103.110 64.840 103.430 64.900 ;
        RECT 96.670 64.700 103.430 64.840 ;
        RECT 96.670 64.640 96.990 64.700 ;
        RECT 102.665 64.655 102.955 64.700 ;
        RECT 103.110 64.640 103.430 64.700 ;
        RECT 113.230 64.840 113.550 64.900 ;
        RECT 120.605 64.840 120.895 64.885 ;
        RECT 113.230 64.700 120.895 64.840 ;
        RECT 113.230 64.640 113.550 64.700 ;
        RECT 120.605 64.655 120.895 64.700 ;
        RECT 71.845 64.500 72.135 64.545 ;
        RECT 72.290 64.500 72.610 64.560 ;
        RECT 71.845 64.360 72.610 64.500 ;
        RECT 71.845 64.315 72.135 64.360 ;
        RECT 72.290 64.300 72.610 64.360 ;
        RECT 74.125 64.500 74.775 64.545 ;
        RECT 77.725 64.500 78.015 64.545 ;
        RECT 80.125 64.500 80.415 64.545 ;
        RECT 74.125 64.360 80.415 64.500 ;
        RECT 74.125 64.315 74.775 64.360 ;
        RECT 77.425 64.315 78.015 64.360 ;
        RECT 80.125 64.315 80.415 64.360 ;
        RECT 93.450 64.500 93.770 64.560 ;
        RECT 102.205 64.500 102.495 64.545 ;
        RECT 104.950 64.500 105.270 64.560 ;
        RECT 93.450 64.360 105.270 64.500 ;
        RECT 70.465 63.975 70.755 64.205 ;
        RECT 70.930 64.160 71.220 64.205 ;
        RECT 72.765 64.160 73.055 64.205 ;
        RECT 76.345 64.160 76.635 64.205 ;
        RECT 70.930 64.020 76.635 64.160 ;
        RECT 70.930 63.975 71.220 64.020 ;
        RECT 72.765 63.975 73.055 64.020 ;
        RECT 76.345 63.975 76.635 64.020 ;
        RECT 77.425 64.000 77.715 64.315 ;
        RECT 93.450 64.300 93.770 64.360 ;
        RECT 102.205 64.315 102.495 64.360 ;
        RECT 104.950 64.300 105.270 64.360 ;
        RECT 115.525 64.500 116.175 64.545 ;
        RECT 119.125 64.500 119.415 64.545 ;
        RECT 115.525 64.360 119.415 64.500 ;
        RECT 115.525 64.315 116.175 64.360 ;
        RECT 118.825 64.315 119.415 64.360 ;
        RECT 118.825 64.220 119.115 64.315 ;
        RECT 80.585 64.160 80.875 64.205 ;
        RECT 81.950 64.160 82.270 64.220 ;
        RECT 80.585 64.020 82.270 64.160 ;
        RECT 80.585 63.975 80.875 64.020 ;
        RECT 81.950 63.960 82.270 64.020 ;
        RECT 87.930 63.960 88.250 64.220 ;
        RECT 88.850 63.960 89.170 64.220 ;
        RECT 94.830 64.160 95.150 64.220 ;
        RECT 96.225 64.160 96.515 64.205 ;
        RECT 89.400 64.020 95.150 64.160 ;
        RECT 89.400 63.820 89.540 64.020 ;
        RECT 94.830 63.960 95.150 64.020 ;
        RECT 95.840 64.020 96.515 64.160 ;
        RECT 70.080 63.680 89.540 63.820 ;
        RECT 90.245 63.820 90.535 63.865 ;
        RECT 92.990 63.820 93.310 63.880 ;
        RECT 90.245 63.680 93.310 63.820 ;
        RECT 65.390 63.620 65.710 63.680 ;
        RECT 90.245 63.635 90.535 63.680 ;
        RECT 92.990 63.620 93.310 63.680 ;
        RECT 95.840 63.525 95.980 64.020 ;
        RECT 96.225 63.975 96.515 64.020 ;
        RECT 110.930 64.160 111.250 64.220 ;
        RECT 111.865 64.160 112.155 64.205 ;
        RECT 110.930 64.020 112.155 64.160 ;
        RECT 110.930 63.960 111.250 64.020 ;
        RECT 111.865 63.975 112.155 64.020 ;
        RECT 112.330 64.160 112.620 64.205 ;
        RECT 114.165 64.160 114.455 64.205 ;
        RECT 117.745 64.160 118.035 64.205 ;
        RECT 112.330 64.020 118.035 64.160 ;
        RECT 112.330 63.975 112.620 64.020 ;
        RECT 114.165 63.975 114.455 64.020 ;
        RECT 117.745 63.975 118.035 64.020 ;
        RECT 118.750 64.000 119.115 64.220 ;
        RECT 118.750 63.960 119.070 64.000 ;
        RECT 103.585 63.820 103.875 63.865 ;
        RECT 105.410 63.820 105.730 63.880 ;
        RECT 103.585 63.680 105.730 63.820 ;
        RECT 103.585 63.635 103.875 63.680 ;
        RECT 105.410 63.620 105.730 63.680 ;
        RECT 113.245 63.820 113.535 63.865 ;
        RECT 118.290 63.820 118.610 63.880 ;
        RECT 113.245 63.680 118.610 63.820 ;
        RECT 113.245 63.635 113.535 63.680 ;
        RECT 118.290 63.620 118.610 63.680 ;
        RECT 30.430 63.340 32.960 63.480 ;
        RECT 17.550 63.280 17.870 63.340 ;
        RECT 30.430 63.280 30.750 63.340 ;
        RECT 12.045 63.140 12.335 63.185 ;
        RECT 12.490 63.140 12.810 63.200 ;
        RECT 12.045 63.000 12.810 63.140 ;
        RECT 12.045 62.955 12.335 63.000 ;
        RECT 12.490 62.940 12.810 63.000 ;
        RECT 21.230 62.940 21.550 63.200 ;
        RECT 21.690 63.140 22.010 63.200 ;
        RECT 25.845 63.140 26.135 63.185 ;
        RECT 21.690 63.000 26.135 63.140 ;
        RECT 21.690 62.940 22.010 63.000 ;
        RECT 25.845 62.955 26.135 63.000 ;
        RECT 31.810 63.140 32.130 63.200 ;
        RECT 32.285 63.140 32.575 63.185 ;
        RECT 31.810 63.000 32.575 63.140 ;
        RECT 32.820 63.140 32.960 63.340 ;
        RECT 34.570 63.340 43.170 63.480 ;
        RECT 34.570 63.280 34.890 63.340 ;
        RECT 42.850 63.280 43.170 63.340 ;
        RECT 43.400 63.340 50.900 63.480 ;
        RECT 43.400 63.140 43.540 63.340 ;
        RECT 32.820 63.000 43.540 63.140 ;
        RECT 31.810 62.940 32.130 63.000 ;
        RECT 32.285 62.955 32.575 63.000 ;
        RECT 50.210 62.940 50.530 63.200 ;
        RECT 50.760 63.140 50.900 63.340 ;
        RECT 51.605 63.295 51.895 63.525 ;
        RECT 71.335 63.480 71.625 63.525 ;
        RECT 73.225 63.480 73.515 63.525 ;
        RECT 76.345 63.480 76.635 63.525 ;
        RECT 62.030 63.340 68.840 63.480 ;
        RECT 62.030 63.140 62.170 63.340 ;
        RECT 68.700 63.185 68.840 63.340 ;
        RECT 71.335 63.340 76.635 63.480 ;
        RECT 71.335 63.295 71.625 63.340 ;
        RECT 73.225 63.295 73.515 63.340 ;
        RECT 76.345 63.295 76.635 63.340 ;
        RECT 81.580 63.340 87.700 63.480 ;
        RECT 50.760 63.000 62.170 63.140 ;
        RECT 68.625 63.140 68.915 63.185 ;
        RECT 81.580 63.140 81.720 63.340 ;
        RECT 68.625 63.000 81.720 63.140 ;
        RECT 86.550 63.140 86.870 63.200 ;
        RECT 87.025 63.140 87.315 63.185 ;
        RECT 86.550 63.000 87.315 63.140 ;
        RECT 87.560 63.140 87.700 63.340 ;
        RECT 95.765 63.295 96.055 63.525 ;
        RECT 112.735 63.480 113.025 63.525 ;
        RECT 114.625 63.480 114.915 63.525 ;
        RECT 117.745 63.480 118.035 63.525 ;
        RECT 112.735 63.340 118.035 63.480 ;
        RECT 112.735 63.295 113.025 63.340 ;
        RECT 114.625 63.295 114.915 63.340 ;
        RECT 117.745 63.295 118.035 63.340 ;
        RECT 96.670 63.140 96.990 63.200 ;
        RECT 87.560 63.000 96.990 63.140 ;
        RECT 68.625 62.955 68.915 63.000 ;
        RECT 86.550 62.940 86.870 63.000 ;
        RECT 87.025 62.955 87.315 63.000 ;
        RECT 96.670 62.940 96.990 63.000 ;
        RECT 97.145 63.140 97.435 63.185 ;
        RECT 97.590 63.140 97.910 63.200 ;
        RECT 97.145 63.000 97.910 63.140 ;
        RECT 97.145 62.955 97.435 63.000 ;
        RECT 97.590 62.940 97.910 63.000 ;
        RECT 98.970 63.140 99.290 63.200 ;
        RECT 100.365 63.140 100.655 63.185 ;
        RECT 98.970 63.000 100.655 63.140 ;
        RECT 98.970 62.940 99.290 63.000 ;
        RECT 100.365 62.955 100.655 63.000 ;
        RECT 5.520 62.320 123.740 62.800 ;
        RECT 16.630 61.920 16.950 62.180 ;
        RECT 18.470 62.120 18.790 62.180 ;
        RECT 36.410 62.165 36.730 62.180 ;
        RECT 18.470 61.980 34.570 62.120 ;
        RECT 18.470 61.920 18.790 61.980 ;
        RECT 8.775 61.780 9.065 61.825 ;
        RECT 10.665 61.780 10.955 61.825 ;
        RECT 13.785 61.780 14.075 61.825 ;
        RECT 8.775 61.640 14.075 61.780 ;
        RECT 8.775 61.595 9.065 61.640 ;
        RECT 10.665 61.595 10.955 61.640 ;
        RECT 13.785 61.595 14.075 61.640 ;
        RECT 19.865 61.595 20.155 61.825 ;
        RECT 27.690 61.780 27.980 61.825 ;
        RECT 29.550 61.780 29.840 61.825 ;
        RECT 32.330 61.780 32.620 61.825 ;
        RECT 27.690 61.640 32.620 61.780 ;
        RECT 34.430 61.780 34.570 61.980 ;
        RECT 36.195 61.935 36.730 62.165 ;
        RECT 64.025 62.120 64.315 62.165 ;
        RECT 88.850 62.120 89.170 62.180 ;
        RECT 36.410 61.920 36.730 61.935 ;
        RECT 48.920 61.980 61.020 62.120 ;
        RECT 48.920 61.780 49.060 61.980 ;
        RECT 34.430 61.640 49.060 61.780 ;
        RECT 49.310 61.780 49.600 61.825 ;
        RECT 51.170 61.780 51.460 61.825 ;
        RECT 53.950 61.780 54.240 61.825 ;
        RECT 49.310 61.640 54.240 61.780 ;
        RECT 27.690 61.595 27.980 61.640 ;
        RECT 29.550 61.595 29.840 61.640 ;
        RECT 32.330 61.595 32.620 61.640 ;
        RECT 49.310 61.595 49.600 61.640 ;
        RECT 51.170 61.595 51.460 61.640 ;
        RECT 53.950 61.595 54.240 61.640 ;
        RECT 7.905 60.915 8.195 61.145 ;
        RECT 8.370 61.100 8.660 61.145 ;
        RECT 10.205 61.100 10.495 61.145 ;
        RECT 13.785 61.100 14.075 61.145 ;
        RECT 8.370 60.960 14.075 61.100 ;
        RECT 8.370 60.915 8.660 60.960 ;
        RECT 10.205 60.915 10.495 60.960 ;
        RECT 13.785 60.915 14.075 60.960 ;
        RECT 14.790 61.120 15.110 61.160 ;
        RECT 7.980 60.760 8.120 60.915 ;
        RECT 14.790 60.900 15.155 61.120 ;
        RECT 18.025 61.100 18.315 61.145 ;
        RECT 19.940 61.100 20.080 61.595 ;
        RECT 23.085 61.440 23.375 61.485 ;
        RECT 24.450 61.440 24.770 61.500 ;
        RECT 23.085 61.300 24.770 61.440 ;
        RECT 23.085 61.255 23.375 61.300 ;
        RECT 24.450 61.240 24.770 61.300 ;
        RECT 28.130 61.440 28.450 61.500 ;
        RECT 29.065 61.440 29.355 61.485 ;
        RECT 28.130 61.300 29.355 61.440 ;
        RECT 28.130 61.240 28.450 61.300 ;
        RECT 29.065 61.255 29.355 61.300 ;
        RECT 42.850 61.440 43.170 61.500 ;
        RECT 48.845 61.440 49.135 61.485 ;
        RECT 42.850 61.300 49.135 61.440 ;
        RECT 42.850 61.240 43.170 61.300 ;
        RECT 48.845 61.255 49.135 61.300 ;
        RECT 50.210 61.440 50.530 61.500 ;
        RECT 50.685 61.440 50.975 61.485 ;
        RECT 50.210 61.300 50.975 61.440 ;
        RECT 50.210 61.240 50.530 61.300 ;
        RECT 50.685 61.255 50.975 61.300 ;
        RECT 18.025 60.960 20.080 61.100 ;
        RECT 22.150 61.100 22.470 61.160 ;
        RECT 27.225 61.100 27.515 61.145 ;
        RECT 32.330 61.100 32.620 61.145 ;
        RECT 22.150 60.960 27.515 61.100 ;
        RECT 18.025 60.915 18.315 60.960 ;
        RECT 22.150 60.900 22.470 60.960 ;
        RECT 27.225 60.915 27.515 60.960 ;
        RECT 30.085 60.960 32.620 61.100 ;
        RECT 8.810 60.760 9.130 60.820 ;
        RECT 7.980 60.620 9.130 60.760 ;
        RECT 8.810 60.560 9.130 60.620 ;
        RECT 9.270 60.560 9.590 60.820 ;
        RECT 14.865 60.805 15.155 60.900 ;
        RECT 11.565 60.760 12.215 60.805 ;
        RECT 14.865 60.760 15.455 60.805 ;
        RECT 21.230 60.760 21.550 60.820 ;
        RECT 30.085 60.805 30.300 60.960 ;
        RECT 32.330 60.915 32.620 60.960 ;
        RECT 38.250 61.100 38.570 61.160 ;
        RECT 46.085 61.100 46.375 61.145 ;
        RECT 47.465 61.100 47.755 61.145 ;
        RECT 53.950 61.100 54.240 61.145 ;
        RECT 38.250 60.960 47.755 61.100 ;
        RECT 38.250 60.900 38.570 60.960 ;
        RECT 46.085 60.915 46.375 60.960 ;
        RECT 47.465 60.915 47.755 60.960 ;
        RECT 51.705 60.960 54.240 61.100 ;
        RECT 11.565 60.620 15.455 60.760 ;
        RECT 11.565 60.575 12.215 60.620 ;
        RECT 15.165 60.575 15.455 60.620 ;
        RECT 15.800 60.620 21.550 60.760 ;
        RECT 11.110 60.420 11.430 60.480 ;
        RECT 15.800 60.420 15.940 60.620 ;
        RECT 21.230 60.560 21.550 60.620 ;
        RECT 21.705 60.760 21.995 60.805 ;
        RECT 28.150 60.760 28.440 60.805 ;
        RECT 30.010 60.760 30.300 60.805 ;
        RECT 21.705 60.620 27.900 60.760 ;
        RECT 21.705 60.575 21.995 60.620 ;
        RECT 11.110 60.280 15.940 60.420 ;
        RECT 17.105 60.420 17.395 60.465 ;
        RECT 17.550 60.420 17.870 60.480 ;
        RECT 17.105 60.280 17.870 60.420 ;
        RECT 11.110 60.220 11.430 60.280 ;
        RECT 17.105 60.235 17.395 60.280 ;
        RECT 17.550 60.220 17.870 60.280 ;
        RECT 22.165 60.420 22.455 60.465 ;
        RECT 22.610 60.420 22.930 60.480 ;
        RECT 22.165 60.280 22.930 60.420 ;
        RECT 27.760 60.420 27.900 60.620 ;
        RECT 28.150 60.620 30.300 60.760 ;
        RECT 28.150 60.575 28.440 60.620 ;
        RECT 30.010 60.575 30.300 60.620 ;
        RECT 30.930 60.760 31.220 60.805 ;
        RECT 31.810 60.760 32.130 60.820 ;
        RECT 51.705 60.805 51.920 60.960 ;
        RECT 53.950 60.915 54.240 60.960 ;
        RECT 34.190 60.760 34.480 60.805 ;
        RECT 30.930 60.620 34.480 60.760 ;
        RECT 30.930 60.575 31.220 60.620 ;
        RECT 31.810 60.560 32.130 60.620 ;
        RECT 34.190 60.575 34.480 60.620 ;
        RECT 49.770 60.760 50.060 60.805 ;
        RECT 51.630 60.760 51.920 60.805 ;
        RECT 52.550 60.760 52.840 60.805 ;
        RECT 55.810 60.760 56.100 60.805 ;
        RECT 49.770 60.620 51.920 60.760 ;
        RECT 49.770 60.575 50.060 60.620 ;
        RECT 51.630 60.575 51.920 60.620 ;
        RECT 52.140 60.620 56.100 60.760 ;
        RECT 60.880 60.760 61.020 61.980 ;
        RECT 62.030 61.980 89.170 62.120 ;
        RECT 62.030 61.440 62.170 61.980 ;
        RECT 64.025 61.935 64.315 61.980 ;
        RECT 88.850 61.920 89.170 61.980 ;
        RECT 92.530 62.120 92.850 62.180 ;
        RECT 93.925 62.120 94.215 62.165 ;
        RECT 92.530 61.980 94.215 62.120 ;
        RECT 92.530 61.920 92.850 61.980 ;
        RECT 93.925 61.935 94.215 61.980 ;
        RECT 103.110 62.120 103.430 62.180 ;
        RECT 114.165 62.120 114.455 62.165 ;
        RECT 118.290 62.120 118.610 62.180 ;
        RECT 118.765 62.120 119.055 62.165 ;
        RECT 103.110 61.980 114.455 62.120 ;
        RECT 103.110 61.920 103.430 61.980 ;
        RECT 86.055 61.780 86.345 61.825 ;
        RECT 87.945 61.780 88.235 61.825 ;
        RECT 91.065 61.780 91.355 61.825 ;
        RECT 86.055 61.640 91.355 61.780 ;
        RECT 86.055 61.595 86.345 61.640 ;
        RECT 87.945 61.595 88.235 61.640 ;
        RECT 91.065 61.595 91.355 61.640 ;
        RECT 97.095 61.780 97.385 61.825 ;
        RECT 98.985 61.780 99.275 61.825 ;
        RECT 102.105 61.780 102.395 61.825 ;
        RECT 97.095 61.640 102.395 61.780 ;
        RECT 97.095 61.595 97.385 61.640 ;
        RECT 98.985 61.595 99.275 61.640 ;
        RECT 102.105 61.595 102.395 61.640 ;
        RECT 104.950 61.580 105.270 61.840 ;
        RECT 106.295 61.780 106.585 61.825 ;
        RECT 108.185 61.780 108.475 61.825 ;
        RECT 111.305 61.780 111.595 61.825 ;
        RECT 106.295 61.640 111.595 61.780 ;
        RECT 106.295 61.595 106.585 61.640 ;
        RECT 108.185 61.595 108.475 61.640 ;
        RECT 111.305 61.595 111.595 61.640 ;
        RECT 61.340 61.300 62.170 61.440 ;
        RECT 63.105 61.440 63.395 61.485 ;
        RECT 63.105 61.300 65.620 61.440 ;
        RECT 61.340 61.145 61.480 61.300 ;
        RECT 63.105 61.255 63.395 61.300 ;
        RECT 65.480 61.160 65.620 61.300 ;
        RECT 86.550 61.240 86.870 61.500 ;
        RECT 96.225 61.440 96.515 61.485 ;
        RECT 105.425 61.440 105.715 61.485 ;
        RECT 110.470 61.440 110.790 61.500 ;
        RECT 96.225 61.300 110.790 61.440 ;
        RECT 111.940 61.440 112.080 61.980 ;
        RECT 114.165 61.935 114.455 61.980 ;
        RECT 116.080 61.980 117.140 62.120 ;
        RECT 112.310 61.780 112.630 61.840 ;
        RECT 116.080 61.780 116.220 61.980 ;
        RECT 112.310 61.640 116.220 61.780 ;
        RECT 117.000 61.780 117.140 61.980 ;
        RECT 118.290 61.980 119.055 62.120 ;
        RECT 118.290 61.920 118.610 61.980 ;
        RECT 118.765 61.935 119.055 61.980 ;
        RECT 117.000 61.640 117.600 61.780 ;
        RECT 112.310 61.580 112.630 61.640 ;
        RECT 111.940 61.300 116.680 61.440 ;
        RECT 96.225 61.255 96.515 61.300 ;
        RECT 105.425 61.255 105.715 61.300 ;
        RECT 110.470 61.240 110.790 61.300 ;
        RECT 61.265 60.915 61.555 61.145 ;
        RECT 63.550 60.900 63.870 61.160 ;
        RECT 64.470 60.900 64.790 61.160 ;
        RECT 64.930 60.900 65.250 61.160 ;
        RECT 65.390 60.900 65.710 61.160 ;
        RECT 70.465 61.100 70.755 61.145 ;
        RECT 70.080 60.960 70.755 61.100 ;
        RECT 70.080 60.820 70.220 60.960 ;
        RECT 70.465 60.915 70.755 60.960 ;
        RECT 82.410 61.100 82.730 61.160 ;
        RECT 116.540 61.145 116.680 61.300 ;
        RECT 116.910 61.240 117.230 61.500 ;
        RECT 117.460 61.485 117.600 61.640 ;
        RECT 117.385 61.255 117.675 61.485 ;
        RECT 85.185 61.100 85.475 61.145 ;
        RECT 82.410 60.960 85.475 61.100 ;
        RECT 82.410 60.900 82.730 60.960 ;
        RECT 85.185 60.915 85.475 60.960 ;
        RECT 85.650 61.100 85.940 61.145 ;
        RECT 87.485 61.100 87.775 61.145 ;
        RECT 91.065 61.100 91.355 61.145 ;
        RECT 85.650 60.960 91.355 61.100 ;
        RECT 85.650 60.915 85.940 60.960 ;
        RECT 87.485 60.915 87.775 60.960 ;
        RECT 91.065 60.915 91.355 60.960 ;
        RECT 69.990 60.760 70.310 60.820 ;
        RECT 60.880 60.620 70.310 60.760 ;
        RECT 31.350 60.420 31.670 60.480 ;
        RECT 27.760 60.280 31.670 60.420 ;
        RECT 22.165 60.235 22.455 60.280 ;
        RECT 22.610 60.220 22.930 60.280 ;
        RECT 31.350 60.220 31.670 60.280 ;
        RECT 46.530 60.220 46.850 60.480 ;
        RECT 47.925 60.420 48.215 60.465 ;
        RECT 52.140 60.420 52.280 60.620 ;
        RECT 52.550 60.575 52.840 60.620 ;
        RECT 55.810 60.575 56.100 60.620 ;
        RECT 69.990 60.560 70.310 60.620 ;
        RECT 71.830 60.760 72.150 60.820 ;
        RECT 75.510 60.760 75.830 60.820 ;
        RECT 71.830 60.620 75.830 60.760 ;
        RECT 71.830 60.560 72.150 60.620 ;
        RECT 75.510 60.560 75.830 60.620 ;
        RECT 88.845 60.760 89.495 60.805 ;
        RECT 90.230 60.760 90.550 60.820 ;
        RECT 92.145 60.805 92.435 61.120 ;
        RECT 96.690 61.100 96.980 61.145 ;
        RECT 98.525 61.100 98.815 61.145 ;
        RECT 102.105 61.100 102.395 61.145 ;
        RECT 96.690 60.960 102.395 61.100 ;
        RECT 96.690 60.915 96.980 60.960 ;
        RECT 98.525 60.915 98.815 60.960 ;
        RECT 102.105 60.915 102.395 60.960 ;
        RECT 92.145 60.760 92.735 60.805 ;
        RECT 88.845 60.620 92.735 60.760 ;
        RECT 88.845 60.575 89.495 60.620 ;
        RECT 90.230 60.560 90.550 60.620 ;
        RECT 92.445 60.575 92.735 60.620 ;
        RECT 97.590 60.560 97.910 60.820 ;
        RECT 99.885 60.760 100.535 60.805 ;
        RECT 101.270 60.760 101.590 60.820 ;
        RECT 103.185 60.805 103.475 61.120 ;
        RECT 105.890 61.100 106.180 61.145 ;
        RECT 107.725 61.100 108.015 61.145 ;
        RECT 111.305 61.100 111.595 61.145 ;
        RECT 105.890 60.960 111.595 61.100 ;
        RECT 105.890 60.915 106.180 60.960 ;
        RECT 107.725 60.915 108.015 60.960 ;
        RECT 111.305 60.915 111.595 60.960 ;
        RECT 109.090 60.805 109.410 60.820 ;
        RECT 112.385 60.805 112.675 61.120 ;
        RECT 116.465 60.915 116.755 61.145 ;
        RECT 119.670 60.900 119.990 61.160 ;
        RECT 103.185 60.760 103.775 60.805 ;
        RECT 99.885 60.620 103.775 60.760 ;
        RECT 99.885 60.575 100.535 60.620 ;
        RECT 101.270 60.560 101.590 60.620 ;
        RECT 103.485 60.575 103.775 60.620 ;
        RECT 106.805 60.575 107.095 60.805 ;
        RECT 109.085 60.760 109.735 60.805 ;
        RECT 112.385 60.760 112.975 60.805 ;
        RECT 109.085 60.620 112.975 60.760 ;
        RECT 109.085 60.575 109.735 60.620 ;
        RECT 112.685 60.575 112.975 60.620 ;
        RECT 113.320 60.620 114.840 60.760 ;
        RECT 47.925 60.280 52.280 60.420 ;
        RECT 53.890 60.420 54.210 60.480 ;
        RECT 57.815 60.420 58.105 60.465 ;
        RECT 53.890 60.280 58.105 60.420 ;
        RECT 47.925 60.235 48.215 60.280 ;
        RECT 53.890 60.220 54.210 60.280 ;
        RECT 57.815 60.235 58.105 60.280 ;
        RECT 59.870 60.220 60.190 60.480 ;
        RECT 66.325 60.420 66.615 60.465 ;
        RECT 69.070 60.420 69.390 60.480 ;
        RECT 72.290 60.420 72.610 60.480 ;
        RECT 66.325 60.280 72.610 60.420 ;
        RECT 66.325 60.235 66.615 60.280 ;
        RECT 69.070 60.220 69.390 60.280 ;
        RECT 72.290 60.220 72.610 60.280 ;
        RECT 100.810 60.420 101.130 60.480 ;
        RECT 106.880 60.420 107.020 60.575 ;
        RECT 109.090 60.560 109.410 60.575 ;
        RECT 100.810 60.280 107.020 60.420 ;
        RECT 107.250 60.420 107.570 60.480 ;
        RECT 113.320 60.420 113.460 60.620 ;
        RECT 114.700 60.465 114.840 60.620 ;
        RECT 107.250 60.280 113.460 60.420 ;
        RECT 100.810 60.220 101.130 60.280 ;
        RECT 107.250 60.220 107.570 60.280 ;
        RECT 114.625 60.235 114.915 60.465 ;
        RECT 5.520 59.600 123.740 60.080 ;
        RECT 9.270 59.400 9.590 59.460 ;
        RECT 10.205 59.400 10.495 59.445 ;
        RECT 17.550 59.400 17.870 59.460 ;
        RECT 9.270 59.260 10.495 59.400 ;
        RECT 9.270 59.200 9.590 59.260 ;
        RECT 10.205 59.215 10.495 59.260 ;
        RECT 14.420 59.260 17.870 59.400 ;
        RECT 13.870 59.060 14.190 59.120 ;
        RECT 14.420 59.105 14.560 59.260 ;
        RECT 17.550 59.200 17.870 59.260 ;
        RECT 21.705 59.400 21.995 59.445 ;
        RECT 22.610 59.400 22.930 59.460 ;
        RECT 21.705 59.260 22.930 59.400 ;
        RECT 21.705 59.215 21.995 59.260 ;
        RECT 22.610 59.200 22.930 59.260 ;
        RECT 28.590 59.400 28.910 59.460 ;
        RECT 30.905 59.400 31.195 59.445 ;
        RECT 53.430 59.400 53.750 59.460 ;
        RECT 28.590 59.260 31.195 59.400 ;
        RECT 28.590 59.200 28.910 59.260 ;
        RECT 30.905 59.215 31.195 59.260 ;
        RECT 43.400 59.260 53.750 59.400 ;
        RECT 12.580 58.920 14.190 59.060 ;
        RECT 11.110 58.520 11.430 58.780 ;
        RECT 12.580 58.765 12.720 58.920 ;
        RECT 13.870 58.860 14.190 58.920 ;
        RECT 14.345 58.875 14.635 59.105 ;
        RECT 16.625 59.060 17.275 59.105 ;
        RECT 19.390 59.060 19.710 59.120 ;
        RECT 20.225 59.060 20.515 59.105 ;
        RECT 16.625 58.920 20.515 59.060 ;
        RECT 16.625 58.875 17.275 58.920 ;
        RECT 19.390 58.860 19.710 58.920 ;
        RECT 19.925 58.875 20.515 58.920 ;
        RECT 25.825 59.060 26.475 59.105 ;
        RECT 29.425 59.060 29.715 59.105 ;
        RECT 29.970 59.060 30.290 59.120 ;
        RECT 40.105 59.060 40.395 59.105 ;
        RECT 42.390 59.060 42.710 59.120 ;
        RECT 25.825 58.920 30.290 59.060 ;
        RECT 25.825 58.875 26.475 58.920 ;
        RECT 29.125 58.875 29.715 58.920 ;
        RECT 12.505 58.535 12.795 58.765 ;
        RECT 13.430 58.720 13.720 58.765 ;
        RECT 15.265 58.720 15.555 58.765 ;
        RECT 18.845 58.720 19.135 58.765 ;
        RECT 13.430 58.580 19.135 58.720 ;
        RECT 13.430 58.535 13.720 58.580 ;
        RECT 15.265 58.535 15.555 58.580 ;
        RECT 18.845 58.535 19.135 58.580 ;
        RECT 19.925 58.560 20.215 58.875 ;
        RECT 22.630 58.720 22.920 58.765 ;
        RECT 24.465 58.720 24.755 58.765 ;
        RECT 28.045 58.720 28.335 58.765 ;
        RECT 22.630 58.580 28.335 58.720 ;
        RECT 22.630 58.535 22.920 58.580 ;
        RECT 24.465 58.535 24.755 58.580 ;
        RECT 28.045 58.535 28.335 58.580 ;
        RECT 29.125 58.560 29.415 58.875 ;
        RECT 29.970 58.860 30.290 58.920 ;
        RECT 34.430 58.920 42.710 59.060 ;
        RECT 8.810 58.380 9.130 58.440 ;
        RECT 12.965 58.380 13.255 58.425 ;
        RECT 22.150 58.380 22.470 58.440 ;
        RECT 8.810 58.240 22.470 58.380 ;
        RECT 8.810 58.180 9.130 58.240 ;
        RECT 12.965 58.195 13.255 58.240 ;
        RECT 22.150 58.180 22.470 58.240 ;
        RECT 23.530 58.180 23.850 58.440 ;
        RECT 31.350 58.380 31.670 58.440 ;
        RECT 34.430 58.380 34.570 58.920 ;
        RECT 40.105 58.875 40.395 58.920 ;
        RECT 42.390 58.860 42.710 58.920 ;
        RECT 37.345 58.720 37.635 58.765 ;
        RECT 39.645 58.720 39.935 58.765 ;
        RECT 37.345 58.580 38.020 58.720 ;
        RECT 37.345 58.535 37.635 58.580 ;
        RECT 31.350 58.240 34.570 58.380 ;
        RECT 31.350 58.180 31.670 58.240 ;
        RECT 37.880 58.085 38.020 58.580 ;
        RECT 38.800 58.580 39.935 58.720 ;
        RECT 13.835 58.040 14.125 58.085 ;
        RECT 15.725 58.040 16.015 58.085 ;
        RECT 18.845 58.040 19.135 58.085 ;
        RECT 13.835 57.900 19.135 58.040 ;
        RECT 13.835 57.855 14.125 57.900 ;
        RECT 15.725 57.855 16.015 57.900 ;
        RECT 18.845 57.855 19.135 57.900 ;
        RECT 23.035 58.040 23.325 58.085 ;
        RECT 24.925 58.040 25.215 58.085 ;
        RECT 28.045 58.040 28.335 58.085 ;
        RECT 23.035 57.900 28.335 58.040 ;
        RECT 23.035 57.855 23.325 57.900 ;
        RECT 24.925 57.855 25.215 57.900 ;
        RECT 28.045 57.855 28.335 57.900 ;
        RECT 37.805 57.855 38.095 58.085 ;
        RECT 12.030 57.500 12.350 57.760 ;
        RECT 35.030 57.700 35.350 57.760 ;
        RECT 36.425 57.700 36.715 57.745 ;
        RECT 35.030 57.560 36.715 57.700 ;
        RECT 38.800 57.700 38.940 58.580 ;
        RECT 39.645 58.535 39.935 58.580 ;
        RECT 42.850 58.520 43.170 58.780 ;
        RECT 39.170 58.380 39.490 58.440 ;
        RECT 41.025 58.380 41.315 58.425 ;
        RECT 43.400 58.380 43.540 59.260 ;
        RECT 53.430 59.200 53.750 59.260 ;
        RECT 53.890 59.400 54.210 59.460 ;
        RECT 54.365 59.400 54.655 59.445 ;
        RECT 53.890 59.260 54.655 59.400 ;
        RECT 53.890 59.200 54.210 59.260 ;
        RECT 54.365 59.215 54.655 59.260 ;
        RECT 90.230 59.200 90.550 59.460 ;
        RECT 100.365 59.400 100.655 59.445 ;
        RECT 100.810 59.400 101.130 59.460 ;
        RECT 100.365 59.260 101.130 59.400 ;
        RECT 100.365 59.215 100.655 59.260 ;
        RECT 100.810 59.200 101.130 59.260 ;
        RECT 101.270 59.200 101.590 59.460 ;
        RECT 106.345 59.400 106.635 59.445 ;
        RECT 109.090 59.400 109.410 59.460 ;
        RECT 106.345 59.260 109.410 59.400 ;
        RECT 106.345 59.215 106.635 59.260 ;
        RECT 109.090 59.200 109.410 59.260 ;
        RECT 116.910 59.400 117.230 59.460 ;
        RECT 117.845 59.400 118.135 59.445 ;
        RECT 116.910 59.260 118.135 59.400 ;
        RECT 116.910 59.200 117.230 59.260 ;
        RECT 117.845 59.215 118.135 59.260 ;
        RECT 118.750 59.200 119.070 59.460 ;
        RECT 46.530 59.105 46.850 59.120 ;
        RECT 43.790 59.060 44.080 59.105 ;
        RECT 45.650 59.060 45.940 59.105 ;
        RECT 43.790 58.920 45.940 59.060 ;
        RECT 43.790 58.875 44.080 58.920 ;
        RECT 45.650 58.875 45.940 58.920 ;
        RECT 45.725 58.720 45.940 58.875 ;
        RECT 46.530 59.060 46.860 59.105 ;
        RECT 49.830 59.060 50.120 59.105 ;
        RECT 51.835 59.060 52.125 59.105 ;
        RECT 52.510 59.060 52.830 59.120 ;
        RECT 54.825 59.060 55.115 59.105 ;
        RECT 46.530 58.920 50.120 59.060 ;
        RECT 46.530 58.875 46.860 58.920 ;
        RECT 49.830 58.875 50.120 58.920 ;
        RECT 50.300 58.920 55.115 59.060 ;
        RECT 46.530 58.860 46.850 58.875 ;
        RECT 47.970 58.720 48.260 58.765 ;
        RECT 45.725 58.580 48.260 58.720 ;
        RECT 47.970 58.535 48.260 58.580 ;
        RECT 39.170 58.240 43.540 58.380 ;
        RECT 44.705 58.380 44.995 58.425 ;
        RECT 46.530 58.380 46.850 58.440 ;
        RECT 44.705 58.240 46.850 58.380 ;
        RECT 39.170 58.180 39.490 58.240 ;
        RECT 41.025 58.195 41.315 58.240 ;
        RECT 44.705 58.195 44.995 58.240 ;
        RECT 46.530 58.180 46.850 58.240 ;
        RECT 43.330 58.040 43.620 58.085 ;
        RECT 45.190 58.040 45.480 58.085 ;
        RECT 47.970 58.040 48.260 58.085 ;
        RECT 43.330 57.900 48.260 58.040 ;
        RECT 43.330 57.855 43.620 57.900 ;
        RECT 45.190 57.855 45.480 57.900 ;
        RECT 47.970 57.855 48.260 57.900 ;
        RECT 50.300 57.700 50.440 58.920 ;
        RECT 51.835 58.875 52.125 58.920 ;
        RECT 52.510 58.860 52.830 58.920 ;
        RECT 54.825 58.875 55.115 58.920 ;
        RECT 76.905 59.060 77.195 59.105 ;
        RECT 77.350 59.060 77.670 59.120 ;
        RECT 80.110 59.060 80.430 59.120 ;
        RECT 110.930 59.060 111.250 59.120 ;
        RECT 76.905 58.920 80.430 59.060 ;
        RECT 76.905 58.875 77.195 58.920 ;
        RECT 77.350 58.860 77.670 58.920 ;
        RECT 80.110 58.860 80.430 58.920 ;
        RECT 109.180 58.920 111.250 59.060 ;
        RECT 53.430 58.720 53.750 58.780 ;
        RECT 69.990 58.720 70.310 58.780 ;
        RECT 75.525 58.720 75.815 58.765 ;
        RECT 83.330 58.720 83.650 58.780 ;
        RECT 53.430 58.580 55.960 58.720 ;
        RECT 53.430 58.520 53.750 58.580 ;
        RECT 55.820 58.425 55.960 58.580 ;
        RECT 69.990 58.580 83.650 58.720 ;
        RECT 69.990 58.520 70.310 58.580 ;
        RECT 75.525 58.535 75.815 58.580 ;
        RECT 83.330 58.520 83.650 58.580 ;
        RECT 84.725 58.720 85.015 58.765 ;
        RECT 89.785 58.720 90.075 58.765 ;
        RECT 84.725 58.580 90.075 58.720 ;
        RECT 84.725 58.535 85.015 58.580 ;
        RECT 89.785 58.535 90.075 58.580 ;
        RECT 98.970 58.720 99.290 58.780 ;
        RECT 99.445 58.720 99.735 58.765 ;
        RECT 98.970 58.580 99.735 58.720 ;
        RECT 55.745 58.380 56.035 58.425 ;
        RECT 59.870 58.380 60.190 58.440 ;
        RECT 55.745 58.240 60.190 58.380 ;
        RECT 89.860 58.380 90.000 58.535 ;
        RECT 98.970 58.520 99.290 58.580 ;
        RECT 99.445 58.535 99.735 58.580 ;
        RECT 100.825 58.720 101.115 58.765 ;
        RECT 105.870 58.720 106.190 58.780 ;
        RECT 100.825 58.580 106.190 58.720 ;
        RECT 100.825 58.535 101.115 58.580 ;
        RECT 100.900 58.380 101.040 58.535 ;
        RECT 105.870 58.520 106.190 58.580 ;
        RECT 107.250 58.520 107.570 58.780 ;
        RECT 109.180 58.765 109.320 58.920 ;
        RECT 110.930 58.860 111.250 58.920 ;
        RECT 112.765 59.060 113.415 59.105 ;
        RECT 113.690 59.060 114.010 59.120 ;
        RECT 116.365 59.060 116.655 59.105 ;
        RECT 112.765 58.920 116.655 59.060 ;
        RECT 112.765 58.875 113.415 58.920 ;
        RECT 113.690 58.860 114.010 58.920 ;
        RECT 116.065 58.875 116.655 58.920 ;
        RECT 109.105 58.535 109.395 58.765 ;
        RECT 109.570 58.720 109.860 58.765 ;
        RECT 111.405 58.720 111.695 58.765 ;
        RECT 114.985 58.720 115.275 58.765 ;
        RECT 109.570 58.580 115.275 58.720 ;
        RECT 109.570 58.535 109.860 58.580 ;
        RECT 111.405 58.535 111.695 58.580 ;
        RECT 114.985 58.535 115.275 58.580 ;
        RECT 116.065 58.560 116.355 58.875 ;
        RECT 118.290 58.520 118.610 58.780 ;
        RECT 110.485 58.380 110.775 58.425 ;
        RECT 89.860 58.240 101.040 58.380 ;
        RECT 108.260 58.240 110.775 58.380 ;
        RECT 55.745 58.195 56.035 58.240 ;
        RECT 59.870 58.180 60.190 58.240 ;
        RECT 108.260 58.085 108.400 58.240 ;
        RECT 110.485 58.195 110.775 58.240 ;
        RECT 108.185 57.855 108.475 58.085 ;
        RECT 109.975 58.040 110.265 58.085 ;
        RECT 111.865 58.040 112.155 58.085 ;
        RECT 114.985 58.040 115.275 58.085 ;
        RECT 109.975 57.900 115.275 58.040 ;
        RECT 109.975 57.855 110.265 57.900 ;
        RECT 111.865 57.855 112.155 57.900 ;
        RECT 114.985 57.855 115.275 57.900 ;
        RECT 38.800 57.560 50.440 57.700 ;
        RECT 35.030 57.500 35.350 57.560 ;
        RECT 36.425 57.515 36.715 57.560 ;
        RECT 52.510 57.500 52.830 57.760 ;
        RECT 5.520 56.880 123.740 57.360 ;
        RECT 18.010 56.480 18.330 56.740 ;
        RECT 19.390 56.480 19.710 56.740 ;
        RECT 21.705 56.680 21.995 56.725 ;
        RECT 23.530 56.680 23.850 56.740 ;
        RECT 21.705 56.540 23.850 56.680 ;
        RECT 21.705 56.495 21.995 56.540 ;
        RECT 23.530 56.480 23.850 56.540 ;
        RECT 42.390 56.480 42.710 56.740 ;
        RECT 46.530 56.480 46.850 56.740 ;
        RECT 64.930 56.680 65.250 56.740 ;
        RECT 65.865 56.680 66.155 56.725 ;
        RECT 64.930 56.540 66.155 56.680 ;
        RECT 64.930 56.480 65.250 56.540 ;
        RECT 65.865 56.495 66.155 56.540 ;
        RECT 94.845 56.680 95.135 56.725 ;
        RECT 98.050 56.680 98.370 56.740 ;
        RECT 94.845 56.540 98.370 56.680 ;
        RECT 94.845 56.495 95.135 56.540 ;
        RECT 98.050 56.480 98.370 56.540 ;
        RECT 113.690 56.480 114.010 56.740 ;
        RECT 10.155 56.340 10.445 56.385 ;
        RECT 12.045 56.340 12.335 56.385 ;
        RECT 15.165 56.340 15.455 56.385 ;
        RECT 10.155 56.200 15.455 56.340 ;
        RECT 10.155 56.155 10.445 56.200 ;
        RECT 12.045 56.155 12.335 56.200 ;
        RECT 15.165 56.155 15.455 56.200 ;
        RECT 34.535 56.340 34.825 56.385 ;
        RECT 36.425 56.340 36.715 56.385 ;
        RECT 39.545 56.340 39.835 56.385 ;
        RECT 34.535 56.200 39.835 56.340 ;
        RECT 34.535 56.155 34.825 56.200 ;
        RECT 36.425 56.155 36.715 56.200 ;
        RECT 39.545 56.155 39.835 56.200 ;
        RECT 75.050 56.340 75.370 56.400 ;
        RECT 77.825 56.340 78.115 56.385 ;
        RECT 75.050 56.200 78.115 56.340 ;
        RECT 75.050 56.140 75.370 56.200 ;
        RECT 77.825 56.155 78.115 56.200 ;
        RECT 10.665 56.000 10.955 56.045 ;
        RECT 12.490 56.000 12.810 56.060 ;
        RECT 10.665 55.860 12.810 56.000 ;
        RECT 10.665 55.815 10.955 55.860 ;
        RECT 12.490 55.800 12.810 55.860 ;
        RECT 35.030 55.800 35.350 56.060 ;
        RECT 62.170 56.000 62.490 56.060 ;
        RECT 64.945 56.000 65.235 56.045 ;
        RECT 68.625 56.000 68.915 56.045 ;
        RECT 62.170 55.860 65.235 56.000 ;
        RECT 62.170 55.800 62.490 55.860 ;
        RECT 64.945 55.815 65.235 55.860 ;
        RECT 67.780 55.860 68.915 56.000 ;
        RECT 8.810 55.660 9.130 55.720 ;
        RECT 9.285 55.660 9.575 55.705 ;
        RECT 8.810 55.520 9.575 55.660 ;
        RECT 8.810 55.460 9.130 55.520 ;
        RECT 9.285 55.475 9.575 55.520 ;
        RECT 9.750 55.660 10.040 55.705 ;
        RECT 11.585 55.660 11.875 55.705 ;
        RECT 15.165 55.660 15.455 55.705 ;
        RECT 9.750 55.520 15.455 55.660 ;
        RECT 9.750 55.475 10.040 55.520 ;
        RECT 11.585 55.475 11.875 55.520 ;
        RECT 15.165 55.475 15.455 55.520 ;
        RECT 12.030 55.320 12.350 55.380 ;
        RECT 16.245 55.365 16.535 55.680 ;
        RECT 19.850 55.460 20.170 55.720 ;
        RECT 20.785 55.660 21.075 55.705 ;
        RECT 21.690 55.660 22.010 55.720 ;
        RECT 20.785 55.520 22.010 55.660 ;
        RECT 20.785 55.475 21.075 55.520 ;
        RECT 21.690 55.460 22.010 55.520 ;
        RECT 22.150 55.660 22.470 55.720 ;
        RECT 23.545 55.660 23.835 55.705 ;
        RECT 22.150 55.520 23.835 55.660 ;
        RECT 22.150 55.460 22.470 55.520 ;
        RECT 23.545 55.475 23.835 55.520 ;
        RECT 33.665 55.475 33.955 55.705 ;
        RECT 34.130 55.660 34.420 55.705 ;
        RECT 35.965 55.660 36.255 55.705 ;
        RECT 39.545 55.660 39.835 55.705 ;
        RECT 34.130 55.520 39.835 55.660 ;
        RECT 34.130 55.475 34.420 55.520 ;
        RECT 35.965 55.475 36.255 55.520 ;
        RECT 39.545 55.475 39.835 55.520 ;
        RECT 12.945 55.320 13.595 55.365 ;
        RECT 16.245 55.320 16.835 55.365 ;
        RECT 12.030 55.180 16.835 55.320 ;
        RECT 12.030 55.120 12.350 55.180 ;
        RECT 12.945 55.135 13.595 55.180 ;
        RECT 16.545 55.135 16.835 55.180 ;
        RECT 32.270 55.120 32.590 55.380 ;
        RECT 33.740 55.320 33.880 55.475 ;
        RECT 34.570 55.320 34.890 55.380 ;
        RECT 40.625 55.365 40.915 55.680 ;
        RECT 43.785 55.660 44.075 55.705 ;
        RECT 45.610 55.660 45.930 55.720 ;
        RECT 43.785 55.520 45.930 55.660 ;
        RECT 43.785 55.475 44.075 55.520 ;
        RECT 45.610 55.460 45.930 55.520 ;
        RECT 47.465 55.660 47.755 55.705 ;
        RECT 52.510 55.660 52.830 55.720 ;
        RECT 47.465 55.520 52.830 55.660 ;
        RECT 47.465 55.475 47.755 55.520 ;
        RECT 52.510 55.460 52.830 55.520 ;
        RECT 63.090 55.660 63.410 55.720 ;
        RECT 63.565 55.660 63.855 55.705 ;
        RECT 63.090 55.520 63.855 55.660 ;
        RECT 63.090 55.460 63.410 55.520 ;
        RECT 63.565 55.475 63.855 55.520 ;
        RECT 64.025 55.475 64.315 55.705 ;
        RECT 64.485 55.475 64.775 55.705 ;
        RECT 65.390 55.660 65.710 55.720 ;
        RECT 67.780 55.705 67.920 55.860 ;
        RECT 68.625 55.815 68.915 55.860 ;
        RECT 72.290 56.000 72.610 56.060 ;
        RECT 98.050 56.000 98.370 56.060 ;
        RECT 110.930 56.000 111.250 56.060 ;
        RECT 72.290 55.860 91.840 56.000 ;
        RECT 72.290 55.800 72.610 55.860 ;
        RECT 67.705 55.660 67.995 55.705 ;
        RECT 65.390 55.520 67.995 55.660 ;
        RECT 33.740 55.180 34.890 55.320 ;
        RECT 34.570 55.120 34.890 55.180 ;
        RECT 37.325 55.320 37.975 55.365 ;
        RECT 40.625 55.320 41.215 55.365 ;
        RECT 43.325 55.320 43.615 55.365 ;
        RECT 64.100 55.320 64.240 55.475 ;
        RECT 37.325 55.180 43.615 55.320 ;
        RECT 37.325 55.135 37.975 55.180 ;
        RECT 40.925 55.135 41.215 55.180 ;
        RECT 43.325 55.135 43.615 55.180 ;
        RECT 61.800 55.180 64.240 55.320 ;
        RECT 64.560 55.320 64.700 55.475 ;
        RECT 65.390 55.460 65.710 55.520 ;
        RECT 67.705 55.475 67.995 55.520 ;
        RECT 68.150 55.460 68.470 55.720 ;
        RECT 69.070 55.660 69.390 55.720 ;
        RECT 70.465 55.660 70.755 55.705 ;
        RECT 69.070 55.520 70.755 55.660 ;
        RECT 69.070 55.460 69.390 55.520 ;
        RECT 70.465 55.475 70.755 55.520 ;
        RECT 78.730 55.460 79.050 55.720 ;
        RECT 80.110 55.460 80.430 55.720 ;
        RECT 91.700 55.705 91.840 55.860 ;
        RECT 92.620 55.860 98.370 56.000 ;
        RECT 92.620 55.705 92.760 55.860 ;
        RECT 98.050 55.800 98.370 55.860 ;
        RECT 108.720 55.860 111.250 56.000 ;
        RECT 80.585 55.475 80.875 55.705 ;
        RECT 91.625 55.475 91.915 55.705 ;
        RECT 92.545 55.475 92.835 55.705 ;
        RECT 76.430 55.320 76.750 55.380 ;
        RECT 80.660 55.320 80.800 55.475 ;
        RECT 92.990 55.460 93.310 55.720 ;
        RECT 93.465 55.475 93.755 55.705 ;
        RECT 99.445 55.660 99.735 55.705 ;
        RECT 102.190 55.660 102.510 55.720 ;
        RECT 108.720 55.705 108.860 55.860 ;
        RECT 110.930 55.800 111.250 55.860 ;
        RECT 108.645 55.660 108.935 55.705 ;
        RECT 113.245 55.660 113.535 55.705 ;
        RECT 118.290 55.660 118.610 55.720 ;
        RECT 99.445 55.520 108.935 55.660 ;
        RECT 99.445 55.475 99.735 55.520 ;
        RECT 82.410 55.320 82.730 55.380 ;
        RECT 93.540 55.320 93.680 55.475 ;
        RECT 102.190 55.460 102.510 55.520 ;
        RECT 108.645 55.475 108.935 55.520 ;
        RECT 110.330 55.520 118.610 55.660 ;
        RECT 110.330 55.380 110.470 55.520 ;
        RECT 113.245 55.475 113.535 55.520 ;
        RECT 118.290 55.460 118.610 55.520 ;
        RECT 100.825 55.320 101.115 55.365 ;
        RECT 64.560 55.180 65.160 55.320 ;
        RECT 60.790 54.980 61.110 55.040 ;
        RECT 61.800 54.980 61.940 55.180 ;
        RECT 65.020 55.040 65.160 55.180 ;
        RECT 76.430 55.180 82.730 55.320 ;
        RECT 76.430 55.120 76.750 55.180 ;
        RECT 82.410 55.120 82.730 55.180 ;
        RECT 92.620 55.180 93.680 55.320 ;
        RECT 96.760 55.180 101.115 55.320 ;
        RECT 92.620 55.040 92.760 55.180 ;
        RECT 60.790 54.840 61.940 54.980 ;
        RECT 60.790 54.780 61.110 54.840 ;
        RECT 64.930 54.780 65.250 55.040 ;
        RECT 66.770 54.780 67.090 55.040 ;
        RECT 67.230 54.980 67.550 55.040 ;
        RECT 71.385 54.980 71.675 55.025 ;
        RECT 75.510 54.980 75.830 55.040 ;
        RECT 67.230 54.840 75.830 54.980 ;
        RECT 67.230 54.780 67.550 54.840 ;
        RECT 71.385 54.795 71.675 54.840 ;
        RECT 75.510 54.780 75.830 54.840 ;
        RECT 79.665 54.980 79.955 55.025 ;
        RECT 80.110 54.980 80.430 55.040 ;
        RECT 79.665 54.840 80.430 54.980 ;
        RECT 79.665 54.795 79.955 54.840 ;
        RECT 80.110 54.780 80.430 54.840 ;
        RECT 92.530 54.780 92.850 55.040 ;
        RECT 95.290 54.980 95.610 55.040 ;
        RECT 96.760 54.980 96.900 55.180 ;
        RECT 100.825 55.135 101.115 55.180 ;
        RECT 105.870 55.320 106.190 55.380 ;
        RECT 110.010 55.320 110.470 55.380 ;
        RECT 105.870 55.180 110.470 55.320 ;
        RECT 105.870 55.120 106.190 55.180 ;
        RECT 110.010 55.120 110.330 55.180 ;
        RECT 95.290 54.840 96.900 54.980 ;
        RECT 95.290 54.780 95.610 54.840 ;
        RECT 5.520 54.160 123.740 54.640 ;
        RECT 14.790 53.760 15.110 54.020 ;
        RECT 29.970 53.760 30.290 54.020 ;
        RECT 34.570 53.960 34.890 54.020 ;
        RECT 37.805 53.960 38.095 54.005 ;
        RECT 34.570 53.820 39.400 53.960 ;
        RECT 34.570 53.760 34.890 53.820 ;
        RECT 37.805 53.775 38.095 53.820 ;
        RECT 11.585 53.620 11.875 53.665 ;
        RECT 13.410 53.620 13.730 53.680 ;
        RECT 39.260 53.665 39.400 53.820 ;
        RECT 48.830 53.760 49.150 54.020 ;
        RECT 51.130 53.960 51.450 54.020 ;
        RECT 52.065 53.960 52.355 54.005 ;
        RECT 51.130 53.820 52.355 53.960 ;
        RECT 51.130 53.760 51.450 53.820 ;
        RECT 52.065 53.775 52.355 53.820 ;
        RECT 63.090 53.960 63.410 54.020 ;
        RECT 64.485 53.960 64.775 54.005 ;
        RECT 63.090 53.820 64.775 53.960 ;
        RECT 63.090 53.760 63.410 53.820 ;
        RECT 64.485 53.775 64.775 53.820 ;
        RECT 65.405 53.960 65.695 54.005 ;
        RECT 65.850 53.960 66.170 54.020 ;
        RECT 65.405 53.820 66.170 53.960 ;
        RECT 65.405 53.775 65.695 53.820 ;
        RECT 65.850 53.760 66.170 53.820 ;
        RECT 71.830 53.760 72.150 54.020 ;
        RECT 74.590 53.960 74.910 54.020 ;
        RECT 98.985 53.960 99.275 54.005 ;
        RECT 101.730 53.960 102.050 54.020 ;
        RECT 74.590 53.820 96.900 53.960 ;
        RECT 74.590 53.760 74.910 53.820 ;
        RECT 11.585 53.480 13.730 53.620 ;
        RECT 11.585 53.435 11.875 53.480 ;
        RECT 13.410 53.420 13.730 53.480 ;
        RECT 39.185 53.435 39.475 53.665 ;
        RECT 47.910 53.420 48.230 53.680 ;
        RECT 48.920 53.620 49.060 53.760 ;
        RECT 48.920 53.480 61.480 53.620 ;
        RECT 1.910 53.280 2.230 53.340 ;
        RECT 10.665 53.280 10.955 53.325 ;
        RECT 1.910 53.140 10.955 53.280 ;
        RECT 1.910 53.080 2.230 53.140 ;
        RECT 10.665 53.095 10.955 53.140 ;
        RECT 13.870 53.280 14.190 53.340 ;
        RECT 15.265 53.280 15.555 53.325 ;
        RECT 19.850 53.280 20.170 53.340 ;
        RECT 30.445 53.280 30.735 53.325 ;
        RECT 45.610 53.280 45.930 53.340 ;
        RECT 13.870 53.140 45.930 53.280 ;
        RECT 13.870 53.080 14.190 53.140 ;
        RECT 15.265 53.095 15.555 53.140 ;
        RECT 19.850 53.080 20.170 53.140 ;
        RECT 30.445 53.095 30.735 53.140 ;
        RECT 45.610 53.080 45.930 53.140 ;
        RECT 48.845 53.280 49.135 53.325 ;
        RECT 49.290 53.280 49.610 53.340 ;
        RECT 48.845 53.140 49.610 53.280 ;
        RECT 48.845 53.095 49.135 53.140 ;
        RECT 49.290 53.080 49.610 53.140 ;
        RECT 49.765 53.095 50.055 53.325 ;
        RECT 44.230 52.940 44.550 53.000 ;
        RECT 49.840 52.940 49.980 53.095 ;
        RECT 50.210 53.080 50.530 53.340 ;
        RECT 50.685 53.280 50.975 53.325 ;
        RECT 51.130 53.280 51.450 53.340 ;
        RECT 50.685 53.140 51.450 53.280 ;
        RECT 61.340 53.280 61.480 53.480 ;
        RECT 61.710 53.420 62.030 53.680 ;
        RECT 71.920 53.620 72.060 53.760 ;
        RECT 76.430 53.620 76.750 53.680 ;
        RECT 63.180 53.480 72.060 53.620 ;
        RECT 73.760 53.480 76.750 53.620 ;
        RECT 63.180 53.280 63.320 53.480 ;
        RECT 61.340 53.140 63.320 53.280 ;
        RECT 63.550 53.280 63.870 53.340 ;
        RECT 66.785 53.280 67.075 53.325 ;
        RECT 63.550 53.140 67.075 53.280 ;
        RECT 50.685 53.095 50.975 53.140 ;
        RECT 51.130 53.080 51.450 53.140 ;
        RECT 63.550 53.080 63.870 53.140 ;
        RECT 66.785 53.095 67.075 53.140 ;
        RECT 68.625 53.280 68.915 53.325 ;
        RECT 69.070 53.280 69.390 53.340 ;
        RECT 68.625 53.140 69.390 53.280 ;
        RECT 68.625 53.095 68.915 53.140 ;
        RECT 69.070 53.080 69.390 53.140 ;
        RECT 70.005 53.280 70.295 53.325 ;
        RECT 70.465 53.280 70.755 53.325 ;
        RECT 71.830 53.280 72.150 53.340 ;
        RECT 73.760 53.325 73.900 53.480 ;
        RECT 76.430 53.420 76.750 53.480 ;
        RECT 77.345 53.620 77.995 53.665 ;
        RECT 80.110 53.620 80.430 53.680 ;
        RECT 80.945 53.620 81.235 53.665 ;
        RECT 77.345 53.480 81.235 53.620 ;
        RECT 77.345 53.435 77.995 53.480 ;
        RECT 80.110 53.420 80.430 53.480 ;
        RECT 80.645 53.435 81.235 53.480 ;
        RECT 82.410 53.620 82.730 53.680 ;
        RECT 83.345 53.620 83.635 53.665 ;
        RECT 82.410 53.480 83.635 53.620 ;
        RECT 70.005 53.140 72.150 53.280 ;
        RECT 70.005 53.095 70.295 53.140 ;
        RECT 70.465 53.095 70.755 53.140 ;
        RECT 71.830 53.080 72.150 53.140 ;
        RECT 73.685 53.095 73.975 53.325 ;
        RECT 74.150 53.280 74.440 53.325 ;
        RECT 75.985 53.280 76.275 53.325 ;
        RECT 79.565 53.280 79.855 53.325 ;
        RECT 74.150 53.140 79.855 53.280 ;
        RECT 74.150 53.095 74.440 53.140 ;
        RECT 75.985 53.095 76.275 53.140 ;
        RECT 79.565 53.095 79.855 53.140 ;
        RECT 80.645 53.120 80.935 53.435 ;
        RECT 82.410 53.420 82.730 53.480 ;
        RECT 83.345 53.435 83.635 53.480 ;
        RECT 92.070 53.620 92.390 53.680 ;
        RECT 95.290 53.620 95.610 53.680 ;
        RECT 92.070 53.480 95.610 53.620 ;
        RECT 92.070 53.420 92.390 53.480 ;
        RECT 95.290 53.420 95.610 53.480 ;
        RECT 96.760 53.280 96.900 53.820 ;
        RECT 98.985 53.820 102.050 53.960 ;
        RECT 98.985 53.775 99.275 53.820 ;
        RECT 101.730 53.760 102.050 53.820 ;
        RECT 97.130 53.620 97.450 53.680 ;
        RECT 97.130 53.480 102.420 53.620 ;
        RECT 97.130 53.420 97.450 53.480 ;
        RECT 98.970 53.280 99.290 53.340 ;
        RECT 100.365 53.280 100.655 53.325 ;
        RECT 96.760 53.140 100.655 53.280 ;
        RECT 98.970 53.080 99.290 53.140 ;
        RECT 100.365 53.095 100.655 53.140 ;
        RECT 100.825 53.095 101.115 53.325 ;
        RECT 101.285 53.280 101.575 53.325 ;
        RECT 101.730 53.280 102.050 53.340 ;
        RECT 102.280 53.325 102.420 53.480 ;
        RECT 101.285 53.140 102.050 53.280 ;
        RECT 101.285 53.095 101.575 53.140 ;
        RECT 44.230 52.800 49.980 52.940 ;
        RECT 55.270 52.940 55.590 53.000 ;
        RECT 64.025 52.940 64.315 52.985 ;
        RECT 64.930 52.940 65.250 53.000 ;
        RECT 55.270 52.800 63.780 52.940 ;
        RECT 44.230 52.740 44.550 52.800 ;
        RECT 55.270 52.740 55.590 52.800 ;
        RECT 60.790 52.600 61.110 52.660 ;
        RECT 61.725 52.600 62.015 52.645 ;
        RECT 60.790 52.460 62.015 52.600 ;
        RECT 63.640 52.600 63.780 52.800 ;
        RECT 64.025 52.800 65.250 52.940 ;
        RECT 64.025 52.755 64.315 52.800 ;
        RECT 64.930 52.740 65.250 52.800 ;
        RECT 65.390 52.940 65.710 53.000 ;
        RECT 65.865 52.940 66.155 52.985 ;
        RECT 85.630 52.940 85.950 53.000 ;
        RECT 65.390 52.800 66.155 52.940 ;
        RECT 65.390 52.740 65.710 52.800 ;
        RECT 65.865 52.755 66.155 52.800 ;
        RECT 70.540 52.800 85.950 52.940 ;
        RECT 70.540 52.600 70.680 52.800 ;
        RECT 85.630 52.740 85.950 52.800 ;
        RECT 97.590 52.940 97.910 53.000 ;
        RECT 100.900 52.940 101.040 53.095 ;
        RECT 101.730 53.080 102.050 53.140 ;
        RECT 102.205 53.280 102.495 53.325 ;
        RECT 103.110 53.280 103.430 53.340 ;
        RECT 102.205 53.140 103.430 53.280 ;
        RECT 102.205 53.095 102.495 53.140 ;
        RECT 103.110 53.080 103.430 53.140 ;
        RECT 97.590 52.800 101.040 52.940 ;
        RECT 97.590 52.740 97.910 52.800 ;
        RECT 63.640 52.460 70.680 52.600 ;
        RECT 60.790 52.400 61.110 52.460 ;
        RECT 61.725 52.415 62.015 52.460 ;
        RECT 61.250 52.260 61.570 52.320 ;
        RECT 66.310 52.260 66.630 52.320 ;
        RECT 61.250 52.120 66.630 52.260 ;
        RECT 70.540 52.260 70.680 52.460 ;
        RECT 74.555 52.600 74.845 52.645 ;
        RECT 76.445 52.600 76.735 52.645 ;
        RECT 79.565 52.600 79.855 52.645 ;
        RECT 74.555 52.460 79.855 52.600 ;
        RECT 74.555 52.415 74.845 52.460 ;
        RECT 76.445 52.415 76.735 52.460 ;
        RECT 79.565 52.415 79.855 52.460 ;
        RECT 75.050 52.305 75.370 52.320 ;
        RECT 71.385 52.260 71.675 52.305 ;
        RECT 70.540 52.120 71.675 52.260 ;
        RECT 61.250 52.060 61.570 52.120 ;
        RECT 66.310 52.060 66.630 52.120 ;
        RECT 71.385 52.075 71.675 52.120 ;
        RECT 75.000 52.075 75.370 52.305 ;
        RECT 82.425 52.260 82.715 52.305 ;
        RECT 82.870 52.260 83.190 52.320 ;
        RECT 82.425 52.120 83.190 52.260 ;
        RECT 82.425 52.075 82.715 52.120 ;
        RECT 75.050 52.060 75.370 52.075 ;
        RECT 82.870 52.060 83.190 52.120 ;
        RECT 5.520 51.440 123.740 51.920 ;
        RECT 23.070 51.040 23.390 51.300 ;
        RECT 23.990 51.240 24.310 51.300 ;
        RECT 26.765 51.240 27.055 51.285 ;
        RECT 23.990 51.100 27.055 51.240 ;
        RECT 23.990 51.040 24.310 51.100 ;
        RECT 26.765 51.055 27.055 51.100 ;
        RECT 33.190 51.240 33.510 51.300 ;
        RECT 51.130 51.240 51.450 51.300 ;
        RECT 55.270 51.240 55.590 51.300 ;
        RECT 33.190 51.100 34.570 51.240 ;
        RECT 33.190 51.040 33.510 51.100 ;
        RECT 28.130 50.900 28.450 50.960 ;
        RECT 24.540 50.760 28.450 50.900 ;
        RECT 34.430 50.900 34.570 51.100 ;
        RECT 51.130 51.100 55.590 51.240 ;
        RECT 51.130 51.040 51.450 51.100 ;
        RECT 55.270 51.040 55.590 51.100 ;
        RECT 56.665 51.240 56.955 51.285 ;
        RECT 57.110 51.240 57.430 51.300 ;
        RECT 56.665 51.100 57.430 51.240 ;
        RECT 56.665 51.055 56.955 51.100 ;
        RECT 57.110 51.040 57.430 51.100 ;
        RECT 67.690 51.040 68.010 51.300 ;
        RECT 69.070 51.240 69.390 51.300 ;
        RECT 70.465 51.240 70.755 51.285 ;
        RECT 69.070 51.100 70.755 51.240 ;
        RECT 69.070 51.040 69.390 51.100 ;
        RECT 70.465 51.055 70.755 51.100 ;
        RECT 78.730 51.240 79.050 51.300 ;
        RECT 79.665 51.240 79.955 51.285 ;
        RECT 87.025 51.240 87.315 51.285 ;
        RECT 87.470 51.240 87.790 51.300 ;
        RECT 78.730 51.100 79.955 51.240 ;
        RECT 78.730 51.040 79.050 51.100 ;
        RECT 79.665 51.055 79.955 51.100 ;
        RECT 81.120 51.100 85.400 51.240 ;
        RECT 68.610 50.900 68.930 50.960 ;
        RECT 75.510 50.900 75.830 50.960 ;
        RECT 81.120 50.900 81.260 51.100 ;
        RECT 83.330 50.900 83.650 50.960 ;
        RECT 85.260 50.900 85.400 51.100 ;
        RECT 87.025 51.100 87.790 51.240 ;
        RECT 87.025 51.055 87.315 51.100 ;
        RECT 87.470 51.040 87.790 51.100 ;
        RECT 90.690 51.240 91.010 51.300 ;
        RECT 91.165 51.240 91.455 51.285 ;
        RECT 90.690 51.100 91.455 51.240 ;
        RECT 90.690 51.040 91.010 51.100 ;
        RECT 91.165 51.055 91.455 51.100 ;
        RECT 98.510 51.240 98.830 51.300 ;
        RECT 99.905 51.240 100.195 51.285 ;
        RECT 98.510 51.100 100.195 51.240 ;
        RECT 98.510 51.040 98.830 51.100 ;
        RECT 99.905 51.055 100.195 51.100 ;
        RECT 103.585 51.240 103.875 51.285 ;
        RECT 104.490 51.240 104.810 51.300 ;
        RECT 103.585 51.100 104.810 51.240 ;
        RECT 103.585 51.055 103.875 51.100 ;
        RECT 104.490 51.040 104.810 51.100 ;
        RECT 89.770 50.900 90.090 50.960 ;
        RECT 34.430 50.760 68.930 50.900 ;
        RECT 24.540 50.265 24.680 50.760 ;
        RECT 28.130 50.700 28.450 50.760 ;
        RECT 68.610 50.700 68.930 50.760 ;
        RECT 69.160 50.760 72.980 50.900 ;
        RECT 33.190 50.560 33.510 50.620 ;
        RECT 52.985 50.560 53.275 50.605 ;
        RECT 58.030 50.560 58.350 50.620 ;
        RECT 25.000 50.420 33.510 50.560 ;
        RECT 25.000 50.265 25.140 50.420 ;
        RECT 24.465 50.035 24.755 50.265 ;
        RECT 24.925 50.035 25.215 50.265 ;
        RECT 25.385 50.035 25.675 50.265 ;
        RECT 26.305 50.220 26.595 50.265 ;
        RECT 26.750 50.220 27.070 50.280 ;
        RECT 26.305 50.080 27.070 50.220 ;
        RECT 26.305 50.035 26.595 50.080 ;
        RECT 21.230 49.880 21.550 49.940 ;
        RECT 25.460 49.880 25.600 50.035 ;
        RECT 26.750 50.020 27.070 50.080 ;
        RECT 28.130 50.020 28.450 50.280 ;
        RECT 28.680 50.265 28.820 50.420 ;
        RECT 33.190 50.360 33.510 50.420 ;
        RECT 49.840 50.420 52.280 50.560 ;
        RECT 28.605 50.035 28.895 50.265 ;
        RECT 29.065 50.035 29.355 50.265 ;
        RECT 29.985 50.220 30.275 50.265 ;
        RECT 30.430 50.220 30.750 50.280 ;
        RECT 29.985 50.080 30.750 50.220 ;
        RECT 29.985 50.035 30.275 50.080 ;
        RECT 21.230 49.740 25.600 49.880 ;
        RECT 21.230 49.680 21.550 49.740 ;
        RECT 18.010 49.540 18.330 49.600 ;
        RECT 29.140 49.540 29.280 50.035 ;
        RECT 30.430 50.020 30.750 50.080 ;
        RECT 47.465 50.220 47.755 50.265 ;
        RECT 48.830 50.220 49.150 50.280 ;
        RECT 47.465 50.080 49.150 50.220 ;
        RECT 47.465 50.035 47.755 50.080 ;
        RECT 48.830 50.020 49.150 50.080 ;
        RECT 49.290 50.220 49.610 50.280 ;
        RECT 49.840 50.265 49.980 50.420 ;
        RECT 49.765 50.220 50.055 50.265 ;
        RECT 49.290 50.080 50.055 50.220 ;
        RECT 49.290 50.020 49.610 50.080 ;
        RECT 49.765 50.035 50.055 50.080 ;
        RECT 50.670 50.020 50.990 50.280 ;
        RECT 51.145 50.035 51.435 50.265 ;
        RECT 45.610 49.880 45.930 49.940 ;
        RECT 46.085 49.880 46.375 49.925 ;
        RECT 45.610 49.740 46.375 49.880 ;
        RECT 51.220 49.880 51.360 50.035 ;
        RECT 51.590 50.020 51.910 50.280 ;
        RECT 52.140 50.220 52.280 50.420 ;
        RECT 52.985 50.420 58.350 50.560 ;
        RECT 52.985 50.375 53.275 50.420 ;
        RECT 58.030 50.360 58.350 50.420 ;
        RECT 63.090 50.560 63.410 50.620 ;
        RECT 65.850 50.560 66.170 50.620 ;
        RECT 63.090 50.420 66.170 50.560 ;
        RECT 63.090 50.360 63.410 50.420 ;
        RECT 65.850 50.360 66.170 50.420 ;
        RECT 66.785 50.560 67.075 50.605 ;
        RECT 68.150 50.560 68.470 50.620 ;
        RECT 66.785 50.420 68.470 50.560 ;
        RECT 66.785 50.375 67.075 50.420 ;
        RECT 68.150 50.360 68.470 50.420 ;
        RECT 53.430 50.220 53.750 50.280 ;
        RECT 52.140 50.080 53.750 50.220 ;
        RECT 53.430 50.020 53.750 50.080 ;
        RECT 54.365 50.035 54.655 50.265 ;
        RECT 54.825 50.035 55.115 50.265 ;
        RECT 52.050 49.880 52.370 49.940 ;
        RECT 54.440 49.880 54.580 50.035 ;
        RECT 51.220 49.740 51.820 49.880 ;
        RECT 45.610 49.680 45.930 49.740 ;
        RECT 46.085 49.695 46.375 49.740 ;
        RECT 51.680 49.600 51.820 49.740 ;
        RECT 52.050 49.740 54.580 49.880 ;
        RECT 52.050 49.680 52.370 49.740 ;
        RECT 18.010 49.400 29.280 49.540 ;
        RECT 50.210 49.540 50.530 49.600 ;
        RECT 51.590 49.540 51.910 49.600 ;
        RECT 54.900 49.540 55.040 50.035 ;
        RECT 55.270 50.020 55.590 50.280 ;
        RECT 65.390 50.020 65.710 50.280 ;
        RECT 66.310 50.220 66.630 50.280 ;
        RECT 69.160 50.220 69.300 50.760 ;
        RECT 72.840 50.605 72.980 50.760 ;
        RECT 75.510 50.760 81.260 50.900 ;
        RECT 81.580 50.760 84.940 50.900 ;
        RECT 75.510 50.700 75.830 50.760 ;
        RECT 71.845 50.560 72.135 50.605 ;
        RECT 70.080 50.420 72.135 50.560 ;
        RECT 66.310 50.080 69.300 50.220 ;
        RECT 66.310 50.020 66.630 50.080 ;
        RECT 69.530 50.020 69.850 50.280 ;
        RECT 67.230 49.880 67.550 49.940 ;
        RECT 62.030 49.740 67.550 49.880 ;
        RECT 62.030 49.540 62.170 49.740 ;
        RECT 67.230 49.680 67.550 49.740 ;
        RECT 69.070 49.880 69.390 49.940 ;
        RECT 70.080 49.880 70.220 50.420 ;
        RECT 71.845 50.375 72.135 50.420 ;
        RECT 72.765 50.375 73.055 50.605 ;
        RECT 70.450 50.220 70.770 50.280 ;
        RECT 71.385 50.220 71.675 50.265 ;
        RECT 72.305 50.220 72.595 50.265 ;
        RECT 70.450 50.080 71.675 50.220 ;
        RECT 70.450 50.020 70.770 50.080 ;
        RECT 71.385 50.035 71.675 50.080 ;
        RECT 71.920 50.080 72.595 50.220 ;
        RECT 71.920 49.880 72.060 50.080 ;
        RECT 72.305 50.035 72.595 50.080 ;
        RECT 73.685 50.035 73.975 50.265 ;
        RECT 69.070 49.740 70.220 49.880 ;
        RECT 71.460 49.740 72.060 49.880 ;
        RECT 69.070 49.680 69.390 49.740 ;
        RECT 50.210 49.400 62.170 49.540 ;
        RECT 65.850 49.540 66.170 49.600 ;
        RECT 71.460 49.540 71.600 49.740 ;
        RECT 65.850 49.400 71.600 49.540 ;
        RECT 71.830 49.540 72.150 49.600 ;
        RECT 73.760 49.540 73.900 50.035 ;
        RECT 77.350 50.020 77.670 50.280 ;
        RECT 81.580 50.265 81.720 50.760 ;
        RECT 83.330 50.700 83.650 50.760 ;
        RECT 82.425 50.560 82.715 50.605 ;
        RECT 82.040 50.420 82.715 50.560 ;
        RECT 81.505 50.035 81.795 50.265 ;
        RECT 79.205 49.880 79.495 49.925 ;
        RECT 82.040 49.880 82.180 50.420 ;
        RECT 82.425 50.375 82.715 50.420 ;
        RECT 83.790 50.020 84.110 50.280 ;
        RECT 84.800 50.265 84.940 50.760 ;
        RECT 85.260 50.760 90.090 50.900 ;
        RECT 85.260 50.265 85.400 50.760 ;
        RECT 87.485 50.560 87.775 50.605 ;
        RECT 88.390 50.560 88.710 50.620 ;
        RECT 87.485 50.420 88.710 50.560 ;
        RECT 88.940 50.560 89.080 50.760 ;
        RECT 89.770 50.700 90.090 50.760 ;
        RECT 96.670 50.900 96.990 50.960 ;
        RECT 99.445 50.900 99.735 50.945 ;
        RECT 96.670 50.760 99.735 50.900 ;
        RECT 96.670 50.700 96.990 50.760 ;
        RECT 99.445 50.715 99.735 50.760 ;
        RECT 103.110 50.900 103.430 50.960 ;
        RECT 103.110 50.760 107.020 50.900 ;
        RECT 103.110 50.700 103.430 50.760 ;
        RECT 88.940 50.420 89.540 50.560 ;
        RECT 87.485 50.375 87.775 50.420 ;
        RECT 88.390 50.360 88.710 50.420 ;
        RECT 84.725 50.035 85.015 50.265 ;
        RECT 85.185 50.035 85.475 50.265 ;
        RECT 85.630 50.220 85.950 50.280 ;
        RECT 88.850 50.220 89.170 50.280 ;
        RECT 89.400 50.265 89.540 50.420 ;
        RECT 90.780 50.420 94.600 50.560 ;
        RECT 90.780 50.280 90.920 50.420 ;
        RECT 85.630 50.080 89.170 50.220 ;
        RECT 85.630 50.020 85.950 50.080 ;
        RECT 88.850 50.020 89.170 50.080 ;
        RECT 89.325 50.035 89.615 50.265 ;
        RECT 89.785 50.035 90.075 50.265 ;
        RECT 82.410 49.880 82.730 49.940 ;
        RECT 89.860 49.880 90.000 50.035 ;
        RECT 90.690 50.020 91.010 50.280 ;
        RECT 92.070 50.220 92.390 50.280 ;
        RECT 92.545 50.220 92.835 50.265 ;
        RECT 92.070 50.080 92.835 50.220 ;
        RECT 92.070 50.020 92.390 50.080 ;
        RECT 92.545 50.035 92.835 50.080 ;
        RECT 92.990 50.020 93.310 50.280 ;
        RECT 94.460 50.265 94.600 50.420 ;
        RECT 97.680 50.420 105.640 50.560 ;
        RECT 97.680 50.280 97.820 50.420 ;
        RECT 93.465 50.035 93.755 50.265 ;
        RECT 94.385 50.220 94.675 50.265 ;
        RECT 96.225 50.220 96.515 50.265 ;
        RECT 94.385 50.080 96.515 50.220 ;
        RECT 94.385 50.035 94.675 50.080 ;
        RECT 96.225 50.035 96.515 50.080 ;
        RECT 97.145 50.035 97.435 50.265 ;
        RECT 79.205 49.740 82.730 49.880 ;
        RECT 79.205 49.695 79.495 49.740 ;
        RECT 82.410 49.680 82.730 49.740 ;
        RECT 82.960 49.740 90.000 49.880 ;
        RECT 82.960 49.600 83.100 49.740 ;
        RECT 71.830 49.400 73.900 49.540 ;
        RECT 18.010 49.340 18.330 49.400 ;
        RECT 50.210 49.340 50.530 49.400 ;
        RECT 51.590 49.340 51.910 49.400 ;
        RECT 65.850 49.340 66.170 49.400 ;
        RECT 71.830 49.340 72.150 49.400 ;
        RECT 74.590 49.340 74.910 49.600 ;
        RECT 81.965 49.540 82.255 49.585 ;
        RECT 82.870 49.540 83.190 49.600 ;
        RECT 81.965 49.400 83.190 49.540 ;
        RECT 81.965 49.355 82.255 49.400 ;
        RECT 82.870 49.340 83.190 49.400 ;
        RECT 86.550 49.540 86.870 49.600 ;
        RECT 93.540 49.540 93.680 50.035 ;
        RECT 97.220 49.880 97.360 50.035 ;
        RECT 97.590 50.020 97.910 50.280 ;
        RECT 98.065 50.220 98.355 50.265 ;
        RECT 98.510 50.220 98.830 50.280 ;
        RECT 101.820 50.265 101.960 50.420 ;
        RECT 101.285 50.220 101.575 50.265 ;
        RECT 98.065 50.080 101.575 50.220 ;
        RECT 98.065 50.035 98.355 50.080 ;
        RECT 98.510 50.020 98.830 50.080 ;
        RECT 101.285 50.035 101.575 50.080 ;
        RECT 101.745 50.035 102.035 50.265 ;
        RECT 102.205 50.220 102.495 50.265 ;
        RECT 102.650 50.220 102.970 50.280 ;
        RECT 102.205 50.080 102.970 50.220 ;
        RECT 102.205 50.035 102.495 50.080 ;
        RECT 98.970 49.880 99.290 49.940 ;
        RECT 97.220 49.740 99.290 49.880 ;
        RECT 98.970 49.680 99.290 49.740 ;
        RECT 86.550 49.400 93.680 49.540 ;
        RECT 101.360 49.540 101.500 50.035 ;
        RECT 102.650 50.020 102.970 50.080 ;
        RECT 103.110 50.020 103.430 50.280 ;
        RECT 105.500 50.265 105.640 50.420 ;
        RECT 104.965 50.035 105.255 50.265 ;
        RECT 105.425 50.035 105.715 50.265 ;
        RECT 105.040 49.540 105.180 50.035 ;
        RECT 105.870 50.020 106.190 50.280 ;
        RECT 106.880 50.265 107.020 50.760 ;
        RECT 106.805 50.035 107.095 50.265 ;
        RECT 101.360 49.400 105.180 49.540 ;
        RECT 86.550 49.340 86.870 49.400 ;
        RECT 5.520 48.720 123.740 49.200 ;
        RECT 28.130 48.520 28.450 48.580 ;
        RECT 24.540 48.380 28.450 48.520 ;
        RECT 18.930 48.180 19.250 48.240 ;
        RECT 15.800 48.040 19.250 48.180 ;
        RECT 12.965 47.655 13.255 47.885 ;
        RECT 13.040 47.500 13.180 47.655 ;
        RECT 14.330 47.640 14.650 47.900 ;
        RECT 15.800 47.885 15.940 48.040 ;
        RECT 18.930 47.980 19.250 48.040 ;
        RECT 20.770 48.180 21.090 48.240 ;
        RECT 23.085 48.180 23.375 48.225 ;
        RECT 20.770 48.040 23.375 48.180 ;
        RECT 20.770 47.980 21.090 48.040 ;
        RECT 23.085 47.995 23.375 48.040 ;
        RECT 15.725 47.655 16.015 47.885 ;
        RECT 18.010 47.840 18.330 47.900 ;
        RECT 18.485 47.840 18.775 47.885 ;
        RECT 21.230 47.840 21.550 47.900 ;
        RECT 24.540 47.885 24.680 48.380 ;
        RECT 28.130 48.320 28.450 48.380 ;
        RECT 47.910 48.520 48.230 48.580 ;
        RECT 52.050 48.520 52.370 48.580 ;
        RECT 47.910 48.380 52.370 48.520 ;
        RECT 47.910 48.320 48.230 48.380 ;
        RECT 52.050 48.320 52.370 48.380 ;
        RECT 53.430 48.520 53.750 48.580 ;
        RECT 66.770 48.520 67.090 48.580 ;
        RECT 83.790 48.520 84.110 48.580 ;
        RECT 88.850 48.520 89.170 48.580 ;
        RECT 92.070 48.520 92.390 48.580 ;
        RECT 100.825 48.520 101.115 48.565 ;
        RECT 101.730 48.520 102.050 48.580 ;
        RECT 53.430 48.380 87.700 48.520 ;
        RECT 53.430 48.320 53.750 48.380 ;
        RECT 66.770 48.320 67.090 48.380 ;
        RECT 83.790 48.320 84.110 48.380 ;
        RECT 27.210 48.180 27.530 48.240 ;
        RECT 29.510 48.180 29.830 48.240 ;
        RECT 29.985 48.180 30.275 48.225 ;
        RECT 35.045 48.180 35.335 48.225 ;
        RECT 35.950 48.180 36.270 48.240 ;
        RECT 25.000 48.040 28.360 48.180 ;
        RECT 25.000 47.885 25.140 48.040 ;
        RECT 27.210 47.980 27.530 48.040 ;
        RECT 18.010 47.700 18.775 47.840 ;
        RECT 18.010 47.640 18.330 47.700 ;
        RECT 18.485 47.655 18.775 47.700 ;
        RECT 19.020 47.700 21.550 47.840 ;
        RECT 19.020 47.545 19.160 47.700 ;
        RECT 21.230 47.640 21.550 47.700 ;
        RECT 24.465 47.655 24.755 47.885 ;
        RECT 24.925 47.655 25.215 47.885 ;
        RECT 25.385 47.655 25.675 47.885 ;
        RECT 26.305 47.840 26.595 47.885 ;
        RECT 26.750 47.840 27.070 47.900 ;
        RECT 26.305 47.700 27.070 47.840 ;
        RECT 26.305 47.655 26.595 47.700 ;
        RECT 13.040 47.360 16.860 47.500 ;
        RECT 16.720 47.205 16.860 47.360 ;
        RECT 18.945 47.315 19.235 47.545 ;
        RECT 19.865 47.500 20.155 47.545 ;
        RECT 21.690 47.500 22.010 47.560 ;
        RECT 19.865 47.360 22.010 47.500 ;
        RECT 19.865 47.315 20.155 47.360 ;
        RECT 21.690 47.300 22.010 47.360 ;
        RECT 23.990 47.500 24.310 47.560 ;
        RECT 25.460 47.500 25.600 47.655 ;
        RECT 26.750 47.640 27.070 47.700 ;
        RECT 27.670 47.640 27.990 47.900 ;
        RECT 28.220 47.885 28.360 48.040 ;
        RECT 29.510 48.040 30.275 48.180 ;
        RECT 29.510 47.980 29.830 48.040 ;
        RECT 29.985 47.995 30.275 48.040 ;
        RECT 30.520 48.040 33.880 48.180 ;
        RECT 28.145 47.655 28.435 47.885 ;
        RECT 28.590 47.840 28.910 47.900 ;
        RECT 30.520 47.840 30.660 48.040 ;
        RECT 28.590 47.700 30.660 47.840 ;
        RECT 30.890 47.840 31.210 47.900 ;
        RECT 31.825 47.840 32.115 47.885 ;
        RECT 30.890 47.700 32.115 47.840 ;
        RECT 23.990 47.360 25.600 47.500 ;
        RECT 23.990 47.300 24.310 47.360 ;
        RECT 16.645 46.975 16.935 47.205 ;
        RECT 25.830 47.160 26.150 47.220 ;
        RECT 26.840 47.160 26.980 47.640 ;
        RECT 28.220 47.500 28.360 47.655 ;
        RECT 28.590 47.640 28.910 47.700 ;
        RECT 30.890 47.640 31.210 47.700 ;
        RECT 31.825 47.655 32.115 47.700 ;
        RECT 32.730 47.640 33.050 47.900 ;
        RECT 33.190 47.640 33.510 47.900 ;
        RECT 33.740 47.885 33.880 48.040 ;
        RECT 35.045 48.040 36.270 48.180 ;
        RECT 35.045 47.995 35.335 48.040 ;
        RECT 35.950 47.980 36.270 48.040 ;
        RECT 48.385 48.180 48.675 48.225 ;
        RECT 52.525 48.180 52.815 48.225 ;
        RECT 52.970 48.180 53.290 48.240 ;
        RECT 61.250 48.180 61.570 48.240 ;
        RECT 48.385 48.040 52.280 48.180 ;
        RECT 48.385 47.995 48.675 48.040 ;
        RECT 33.665 47.840 33.955 47.885 ;
        RECT 33.665 47.700 34.570 47.840 ;
        RECT 33.665 47.655 33.955 47.700 ;
        RECT 33.280 47.500 33.420 47.640 ;
        RECT 28.220 47.360 33.420 47.500 ;
        RECT 30.430 47.160 30.750 47.220 ;
        RECT 25.830 47.020 30.750 47.160 ;
        RECT 34.430 47.160 34.570 47.700 ;
        RECT 37.790 47.640 38.110 47.900 ;
        RECT 49.290 47.640 49.610 47.900 ;
        RECT 50.225 47.655 50.515 47.885 ;
        RECT 50.685 47.655 50.975 47.885 ;
        RECT 43.770 47.500 44.090 47.560 ;
        RECT 50.300 47.500 50.440 47.655 ;
        RECT 43.770 47.360 50.440 47.500 ;
        RECT 50.760 47.500 50.900 47.655 ;
        RECT 51.130 47.640 51.450 47.900 ;
        RECT 52.140 47.840 52.280 48.040 ;
        RECT 52.525 48.040 53.290 48.180 ;
        RECT 52.525 47.995 52.815 48.040 ;
        RECT 52.970 47.980 53.290 48.040 ;
        RECT 55.360 48.040 61.570 48.180 ;
        RECT 55.360 47.840 55.500 48.040 ;
        RECT 61.250 47.980 61.570 48.040 ;
        RECT 68.165 48.180 68.455 48.225 ;
        RECT 71.830 48.180 72.150 48.240 ;
        RECT 68.165 48.040 72.150 48.180 ;
        RECT 68.165 47.995 68.455 48.040 ;
        RECT 71.830 47.980 72.150 48.040 ;
        RECT 82.870 48.180 83.190 48.240 ;
        RECT 85.185 48.180 85.475 48.225 ;
        RECT 82.870 48.040 85.475 48.180 ;
        RECT 82.870 47.980 83.190 48.040 ;
        RECT 85.185 47.995 85.475 48.040 ;
        RECT 85.645 48.180 85.935 48.225 ;
        RECT 86.550 48.180 86.870 48.240 ;
        RECT 85.645 48.040 86.870 48.180 ;
        RECT 85.645 47.995 85.935 48.040 ;
        RECT 86.550 47.980 86.870 48.040 ;
        RECT 52.140 47.700 55.500 47.840 ;
        RECT 55.730 47.840 56.050 47.900 ;
        RECT 57.585 47.840 57.875 47.885 ;
        RECT 65.865 47.840 66.155 47.885 ;
        RECT 68.610 47.840 68.930 47.900 ;
        RECT 87.560 47.885 87.700 48.380 ;
        RECT 88.850 48.380 93.220 48.520 ;
        RECT 88.850 48.320 89.170 48.380 ;
        RECT 55.730 47.700 57.875 47.840 ;
        RECT 55.730 47.640 56.050 47.700 ;
        RECT 57.585 47.655 57.875 47.700 ;
        RECT 62.030 47.700 68.930 47.840 ;
        RECT 51.590 47.500 51.910 47.560 ;
        RECT 50.760 47.360 51.910 47.500 ;
        RECT 43.770 47.300 44.090 47.360 ;
        RECT 51.590 47.300 51.910 47.360 ;
        RECT 60.790 47.500 61.110 47.560 ;
        RECT 62.030 47.500 62.170 47.700 ;
        RECT 65.865 47.655 66.155 47.700 ;
        RECT 68.610 47.640 68.930 47.700 ;
        RECT 87.485 47.655 87.775 47.885 ;
        RECT 60.790 47.360 62.170 47.500 ;
        RECT 60.790 47.300 61.110 47.360 ;
        RECT 66.310 47.300 66.630 47.560 ;
        RECT 66.785 47.315 67.075 47.545 ;
        RECT 62.630 47.160 62.950 47.220 ;
        RECT 65.390 47.160 65.710 47.220 ;
        RECT 66.860 47.160 67.000 47.315 ;
        RECT 67.230 47.300 67.550 47.560 ;
        RECT 82.870 47.500 83.190 47.560 ;
        RECT 86.105 47.500 86.395 47.545 ;
        RECT 87.010 47.500 87.330 47.560 ;
        RECT 82.870 47.360 87.330 47.500 ;
        RECT 82.870 47.300 83.190 47.360 ;
        RECT 86.105 47.315 86.395 47.360 ;
        RECT 87.010 47.300 87.330 47.360 ;
        RECT 70.450 47.160 70.770 47.220 ;
        RECT 34.430 47.020 62.170 47.160 ;
        RECT 25.830 46.960 26.150 47.020 ;
        RECT 30.430 46.960 30.750 47.020 ;
        RECT 11.570 46.820 11.890 46.880 ;
        RECT 12.045 46.820 12.335 46.865 ;
        RECT 11.570 46.680 12.335 46.820 ;
        RECT 11.570 46.620 11.890 46.680 ;
        RECT 12.045 46.635 12.335 46.680 ;
        RECT 13.410 46.620 13.730 46.880 ;
        RECT 15.250 46.620 15.570 46.880 ;
        RECT 36.410 46.820 36.730 46.880 ;
        RECT 36.885 46.820 37.175 46.865 ;
        RECT 36.410 46.680 37.175 46.820 ;
        RECT 36.410 46.620 36.730 46.680 ;
        RECT 36.885 46.635 37.175 46.680 ;
        RECT 46.990 46.620 47.310 46.880 ;
        RECT 58.030 46.620 58.350 46.880 ;
        RECT 62.030 46.820 62.170 47.020 ;
        RECT 62.630 47.020 70.770 47.160 ;
        RECT 62.630 46.960 62.950 47.020 ;
        RECT 65.390 46.960 65.710 47.020 ;
        RECT 70.450 46.960 70.770 47.020 ;
        RECT 74.590 46.820 74.910 46.880 ;
        RECT 62.030 46.680 74.910 46.820 ;
        RECT 74.590 46.620 74.910 46.680 ;
        RECT 79.650 46.820 79.970 46.880 ;
        RECT 83.345 46.820 83.635 46.865 ;
        RECT 79.650 46.680 83.635 46.820 ;
        RECT 87.560 46.820 87.700 47.655 ;
        RECT 88.390 47.640 88.710 47.900 ;
        RECT 88.865 47.655 89.155 47.885 ;
        RECT 89.325 47.840 89.615 47.885 ;
        RECT 90.320 47.840 90.460 48.380 ;
        RECT 92.070 48.320 92.390 48.380 ;
        RECT 90.705 48.180 90.995 48.225 ;
        RECT 91.610 48.180 91.930 48.240 ;
        RECT 90.705 48.040 91.930 48.180 ;
        RECT 90.705 47.995 90.995 48.040 ;
        RECT 91.610 47.980 91.930 48.040 ;
        RECT 89.325 47.700 90.460 47.840 ;
        RECT 89.325 47.655 89.615 47.700 ;
        RECT 88.940 47.500 89.080 47.655 ;
        RECT 91.150 47.640 91.470 47.900 ;
        RECT 92.070 47.640 92.390 47.900 ;
        RECT 92.530 47.640 92.850 47.900 ;
        RECT 93.080 47.885 93.220 48.380 ;
        RECT 100.825 48.380 102.050 48.520 ;
        RECT 100.825 48.335 101.115 48.380 ;
        RECT 101.730 48.320 102.050 48.380 ;
        RECT 94.370 47.980 94.690 48.240 ;
        RECT 104.950 48.180 105.270 48.240 ;
        RECT 102.740 48.040 105.270 48.180 ;
        RECT 93.005 47.655 93.295 47.885 ;
        RECT 98.970 47.840 99.290 47.900 ;
        RECT 101.285 47.840 101.575 47.885 ;
        RECT 98.970 47.700 101.575 47.840 ;
        RECT 98.970 47.640 99.290 47.700 ;
        RECT 101.285 47.655 101.575 47.700 ;
        RECT 89.770 47.500 90.090 47.560 ;
        RECT 92.620 47.500 92.760 47.640 ;
        RECT 88.940 47.360 92.760 47.500 ;
        RECT 93.450 47.500 93.770 47.560 ;
        RECT 99.905 47.500 100.195 47.545 ;
        RECT 102.740 47.500 102.880 48.040 ;
        RECT 104.950 47.980 105.270 48.040 ;
        RECT 104.505 47.840 104.795 47.885 ;
        RECT 93.450 47.360 102.880 47.500 ;
        RECT 103.200 47.700 104.795 47.840 ;
        RECT 89.770 47.300 90.090 47.360 ;
        RECT 93.450 47.300 93.770 47.360 ;
        RECT 99.905 47.315 100.195 47.360 ;
        RECT 103.200 47.205 103.340 47.700 ;
        RECT 104.505 47.655 104.795 47.700 ;
        RECT 105.885 47.840 106.175 47.885 ;
        RECT 108.170 47.840 108.490 47.900 ;
        RECT 105.885 47.700 108.490 47.840 ;
        RECT 105.885 47.655 106.175 47.700 ;
        RECT 108.170 47.640 108.490 47.700 ;
        RECT 110.010 47.640 110.330 47.900 ;
        RECT 103.125 46.975 103.415 47.205 ;
        RECT 90.690 46.820 91.010 46.880 ;
        RECT 87.560 46.680 91.010 46.820 ;
        RECT 79.650 46.620 79.970 46.680 ;
        RECT 83.345 46.635 83.635 46.680 ;
        RECT 90.690 46.620 91.010 46.680 ;
        RECT 103.570 46.620 103.890 46.880 ;
        RECT 106.790 46.620 107.110 46.880 ;
        RECT 109.090 46.820 109.410 46.880 ;
        RECT 109.565 46.820 109.855 46.865 ;
        RECT 109.090 46.680 109.855 46.820 ;
        RECT 109.090 46.620 109.410 46.680 ;
        RECT 109.565 46.635 109.855 46.680 ;
        RECT 5.520 46.000 123.740 46.480 ;
        RECT 14.330 45.800 14.650 45.860 ;
        RECT 18.945 45.800 19.235 45.845 ;
        RECT 14.330 45.660 19.235 45.800 ;
        RECT 14.330 45.600 14.650 45.660 ;
        RECT 18.945 45.615 19.235 45.660 ;
        RECT 29.050 45.600 29.370 45.860 ;
        RECT 43.785 45.800 44.075 45.845 ;
        RECT 44.230 45.800 44.550 45.860 ;
        RECT 43.785 45.660 44.550 45.800 ;
        RECT 43.785 45.615 44.075 45.660 ;
        RECT 44.230 45.600 44.550 45.660 ;
        RECT 64.010 45.800 64.330 45.860 ;
        RECT 66.325 45.800 66.615 45.845 ;
        RECT 64.010 45.660 66.615 45.800 ;
        RECT 64.010 45.600 64.330 45.660 ;
        RECT 66.325 45.615 66.615 45.660 ;
        RECT 67.705 45.800 67.995 45.845 ;
        RECT 68.610 45.800 68.930 45.860 ;
        RECT 67.705 45.660 68.930 45.800 ;
        RECT 67.705 45.615 67.995 45.660 ;
        RECT 68.610 45.600 68.930 45.660 ;
        RECT 101.730 45.800 102.050 45.860 ;
        RECT 110.945 45.800 111.235 45.845 ;
        RECT 101.730 45.660 111.235 45.800 ;
        RECT 101.730 45.600 102.050 45.660 ;
        RECT 110.945 45.615 111.235 45.660 ;
        RECT 10.155 45.460 10.445 45.505 ;
        RECT 12.045 45.460 12.335 45.505 ;
        RECT 15.165 45.460 15.455 45.505 ;
        RECT 10.155 45.320 15.455 45.460 ;
        RECT 10.155 45.275 10.445 45.320 ;
        RECT 12.045 45.275 12.335 45.320 ;
        RECT 15.165 45.275 15.455 45.320 ;
        RECT 35.915 45.460 36.205 45.505 ;
        RECT 37.805 45.460 38.095 45.505 ;
        RECT 40.925 45.460 41.215 45.505 ;
        RECT 35.915 45.320 41.215 45.460 ;
        RECT 35.915 45.275 36.205 45.320 ;
        RECT 37.805 45.275 38.095 45.320 ;
        RECT 40.925 45.275 41.215 45.320 ;
        RECT 53.855 45.460 54.145 45.505 ;
        RECT 55.745 45.460 56.035 45.505 ;
        RECT 58.865 45.460 59.155 45.505 ;
        RECT 53.855 45.320 59.155 45.460 ;
        RECT 53.855 45.275 54.145 45.320 ;
        RECT 55.745 45.275 56.035 45.320 ;
        RECT 58.865 45.275 59.155 45.320 ;
        RECT 62.630 45.260 62.950 45.520 ;
        RECT 90.705 45.275 90.995 45.505 ;
        RECT 103.075 45.460 103.365 45.505 ;
        RECT 104.965 45.460 105.255 45.505 ;
        RECT 108.085 45.460 108.375 45.505 ;
        RECT 103.075 45.320 108.375 45.460 ;
        RECT 103.075 45.275 103.365 45.320 ;
        RECT 104.965 45.275 105.255 45.320 ;
        RECT 108.085 45.275 108.375 45.320 ;
        RECT 10.665 45.120 10.955 45.165 ;
        RECT 13.410 45.120 13.730 45.180 ;
        RECT 10.665 44.980 13.730 45.120 ;
        RECT 10.665 44.935 10.955 44.980 ;
        RECT 13.410 44.920 13.730 44.980 ;
        RECT 18.025 45.120 18.315 45.165 ;
        RECT 21.245 45.120 21.535 45.165 ;
        RECT 18.025 44.980 21.535 45.120 ;
        RECT 18.025 44.935 18.315 44.980 ;
        RECT 21.245 44.935 21.535 44.980 ;
        RECT 8.810 44.780 9.130 44.840 ;
        RECT 9.285 44.780 9.575 44.825 ;
        RECT 8.810 44.640 9.575 44.780 ;
        RECT 8.810 44.580 9.130 44.640 ;
        RECT 9.285 44.595 9.575 44.640 ;
        RECT 9.750 44.780 10.040 44.825 ;
        RECT 11.585 44.780 11.875 44.825 ;
        RECT 15.165 44.780 15.455 44.825 ;
        RECT 9.750 44.640 15.455 44.780 ;
        RECT 9.750 44.595 10.040 44.640 ;
        RECT 11.585 44.595 11.875 44.640 ;
        RECT 15.165 44.595 15.455 44.640 ;
        RECT 16.245 44.485 16.535 44.800 ;
        RECT 12.945 44.440 13.595 44.485 ;
        RECT 16.245 44.440 16.835 44.485 ;
        RECT 18.470 44.440 18.790 44.500 ;
        RECT 12.945 44.300 18.790 44.440 ;
        RECT 21.320 44.440 21.460 44.935 ;
        RECT 21.690 44.920 22.010 45.180 ;
        RECT 34.570 45.120 34.890 45.180 ;
        RECT 35.045 45.120 35.335 45.165 ;
        RECT 36.870 45.120 37.190 45.180 ;
        RECT 51.590 45.120 51.910 45.180 ;
        RECT 52.985 45.120 53.275 45.165 ;
        RECT 34.570 44.980 53.275 45.120 ;
        RECT 34.570 44.920 34.890 44.980 ;
        RECT 35.045 44.935 35.335 44.980 ;
        RECT 36.870 44.920 37.190 44.980 ;
        RECT 51.590 44.920 51.910 44.980 ;
        RECT 52.985 44.935 53.275 44.980 ;
        RECT 54.365 45.120 54.655 45.165 ;
        RECT 57.570 45.120 57.890 45.180 ;
        RECT 54.365 44.980 57.890 45.120 ;
        RECT 54.365 44.935 54.655 44.980 ;
        RECT 57.570 44.920 57.890 44.980 ;
        RECT 61.725 45.120 62.015 45.165 ;
        RECT 63.090 45.120 63.410 45.180 ;
        RECT 65.405 45.120 65.695 45.165 ;
        RECT 61.725 44.980 67.000 45.120 ;
        RECT 61.725 44.935 62.015 44.980 ;
        RECT 63.090 44.920 63.410 44.980 ;
        RECT 65.405 44.935 65.695 44.980 ;
        RECT 25.830 44.580 26.150 44.840 ;
        RECT 26.765 44.595 27.055 44.825 ;
        RECT 26.840 44.440 26.980 44.595 ;
        RECT 27.210 44.580 27.530 44.840 ;
        RECT 27.685 44.780 27.975 44.825 ;
        RECT 28.590 44.780 28.910 44.840 ;
        RECT 27.685 44.640 28.910 44.780 ;
        RECT 27.685 44.595 27.975 44.640 ;
        RECT 28.590 44.580 28.910 44.640 ;
        RECT 35.510 44.780 35.800 44.825 ;
        RECT 37.345 44.780 37.635 44.825 ;
        RECT 40.925 44.780 41.215 44.825 ;
        RECT 35.510 44.640 41.215 44.780 ;
        RECT 35.510 44.595 35.800 44.640 ;
        RECT 37.345 44.595 37.635 44.640 ;
        RECT 40.925 44.595 41.215 44.640 ;
        RECT 28.130 44.440 28.450 44.500 ;
        RECT 21.320 44.300 28.450 44.440 ;
        RECT 12.945 44.255 13.595 44.300 ;
        RECT 16.545 44.255 16.835 44.300 ;
        RECT 18.470 44.240 18.790 44.300 ;
        RECT 28.130 44.240 28.450 44.300 ;
        RECT 36.410 44.240 36.730 44.500 ;
        RECT 42.005 44.485 42.295 44.800 ;
        RECT 45.610 44.580 45.930 44.840 ;
        RECT 48.830 44.780 49.150 44.840 ;
        RECT 66.860 44.825 67.000 44.980 ;
        RECT 49.765 44.780 50.055 44.825 ;
        RECT 48.830 44.640 50.055 44.780 ;
        RECT 48.830 44.580 49.150 44.640 ;
        RECT 49.765 44.595 50.055 44.640 ;
        RECT 53.450 44.780 53.740 44.825 ;
        RECT 55.285 44.780 55.575 44.825 ;
        RECT 58.865 44.780 59.155 44.825 ;
        RECT 53.450 44.640 59.155 44.780 ;
        RECT 53.450 44.595 53.740 44.640 ;
        RECT 55.285 44.595 55.575 44.640 ;
        RECT 58.865 44.595 59.155 44.640 ;
        RECT 38.705 44.440 39.355 44.485 ;
        RECT 42.005 44.440 42.595 44.485 ;
        RECT 45.165 44.440 45.455 44.485 ;
        RECT 38.705 44.300 45.455 44.440 ;
        RECT 38.705 44.255 39.355 44.300 ;
        RECT 42.305 44.255 42.595 44.300 ;
        RECT 45.165 44.255 45.455 44.300 ;
        RECT 48.385 44.440 48.675 44.485 ;
        RECT 55.730 44.440 56.050 44.500 ;
        RECT 48.385 44.300 56.050 44.440 ;
        RECT 48.385 44.255 48.675 44.300 ;
        RECT 55.730 44.240 56.050 44.300 ;
        RECT 56.645 44.440 57.295 44.485 ;
        RECT 58.030 44.440 58.350 44.500 ;
        RECT 59.945 44.485 60.235 44.800 ;
        RECT 66.785 44.595 67.075 44.825 ;
        RECT 79.650 44.580 79.970 44.840 ;
        RECT 80.570 44.780 80.890 44.840 ;
        RECT 81.505 44.780 81.795 44.825 ;
        RECT 82.870 44.780 83.190 44.840 ;
        RECT 80.570 44.640 83.190 44.780 ;
        RECT 80.570 44.580 80.890 44.640 ;
        RECT 81.505 44.595 81.795 44.640 ;
        RECT 82.870 44.580 83.190 44.640 ;
        RECT 89.325 44.780 89.615 44.825 ;
        RECT 90.780 44.780 90.920 45.275 ;
        RECT 93.450 44.920 93.770 45.180 ;
        RECT 103.570 44.920 103.890 45.180 ;
        RECT 89.325 44.640 90.920 44.780 ;
        RECT 92.070 44.780 92.390 44.840 ;
        RECT 92.545 44.780 92.835 44.825 ;
        RECT 92.070 44.640 92.835 44.780 ;
        RECT 89.325 44.595 89.615 44.640 ;
        RECT 92.070 44.580 92.390 44.640 ;
        RECT 92.545 44.595 92.835 44.640 ;
        RECT 59.945 44.440 60.535 44.485 ;
        RECT 56.645 44.300 60.535 44.440 ;
        RECT 56.645 44.255 57.295 44.300 ;
        RECT 58.030 44.240 58.350 44.300 ;
        RECT 60.245 44.255 60.535 44.300 ;
        RECT 62.170 44.440 62.490 44.500 ;
        RECT 62.645 44.440 62.935 44.485 ;
        RECT 67.230 44.440 67.550 44.500 ;
        RECT 62.170 44.300 67.550 44.440 ;
        RECT 62.170 44.240 62.490 44.300 ;
        RECT 62.645 44.255 62.935 44.300 ;
        RECT 67.230 44.240 67.550 44.300 ;
        RECT 87.010 44.440 87.330 44.500 ;
        RECT 93.540 44.440 93.680 44.920 ;
        RECT 102.190 44.580 102.510 44.840 ;
        RECT 102.670 44.780 102.960 44.825 ;
        RECT 104.505 44.780 104.795 44.825 ;
        RECT 108.085 44.780 108.375 44.825 ;
        RECT 102.670 44.640 108.375 44.780 ;
        RECT 102.670 44.595 102.960 44.640 ;
        RECT 104.505 44.595 104.795 44.640 ;
        RECT 108.085 44.595 108.375 44.640 ;
        RECT 109.090 44.800 109.410 44.840 ;
        RECT 109.090 44.580 109.455 44.800 ;
        RECT 109.165 44.485 109.455 44.580 ;
        RECT 87.010 44.300 93.680 44.440 ;
        RECT 105.865 44.440 106.515 44.485 ;
        RECT 109.165 44.440 109.755 44.485 ;
        RECT 105.865 44.300 109.755 44.440 ;
        RECT 87.010 44.240 87.330 44.300 ;
        RECT 105.865 44.255 106.515 44.300 ;
        RECT 109.465 44.255 109.755 44.300 ;
        RECT 20.785 44.100 21.075 44.145 ;
        RECT 21.230 44.100 21.550 44.160 ;
        RECT 20.785 43.960 21.550 44.100 ;
        RECT 20.785 43.915 21.075 43.960 ;
        RECT 21.230 43.900 21.550 43.960 ;
        RECT 63.550 44.100 63.870 44.160 ;
        RECT 64.945 44.100 65.235 44.145 ;
        RECT 63.550 43.960 65.235 44.100 ;
        RECT 63.550 43.900 63.870 43.960 ;
        RECT 64.945 43.915 65.235 43.960 ;
        RECT 75.050 44.100 75.370 44.160 ;
        RECT 78.745 44.100 79.035 44.145 ;
        RECT 75.050 43.960 79.035 44.100 ;
        RECT 75.050 43.900 75.370 43.960 ;
        RECT 78.745 43.915 79.035 43.960 ;
        RECT 80.570 44.100 80.890 44.160 ;
        RECT 81.045 44.100 81.335 44.145 ;
        RECT 80.570 43.960 81.335 44.100 ;
        RECT 80.570 43.900 80.890 43.960 ;
        RECT 81.045 43.915 81.335 43.960 ;
        RECT 90.245 44.100 90.535 44.145 ;
        RECT 92.070 44.100 92.390 44.160 ;
        RECT 90.245 43.960 92.390 44.100 ;
        RECT 90.245 43.915 90.535 43.960 ;
        RECT 92.070 43.900 92.390 43.960 ;
        RECT 93.005 44.100 93.295 44.145 ;
        RECT 99.430 44.100 99.750 44.160 ;
        RECT 93.005 43.960 99.750 44.100 ;
        RECT 93.005 43.915 93.295 43.960 ;
        RECT 99.430 43.900 99.750 43.960 ;
        RECT 5.520 43.280 123.740 43.760 ;
        RECT 18.470 42.880 18.790 43.140 ;
        RECT 28.130 42.880 28.450 43.140 ;
        RECT 36.425 43.080 36.715 43.125 ;
        RECT 37.790 43.080 38.110 43.140 ;
        RECT 36.425 42.940 38.110 43.080 ;
        RECT 36.425 42.895 36.715 42.940 ;
        RECT 37.790 42.880 38.110 42.940 ;
        RECT 43.770 42.880 44.090 43.140 ;
        RECT 57.570 43.080 57.890 43.140 ;
        RECT 58.965 43.080 59.255 43.125 ;
        RECT 57.570 42.940 59.255 43.080 ;
        RECT 57.570 42.880 57.890 42.940 ;
        RECT 58.965 42.895 59.255 42.940 ;
        RECT 63.090 42.880 63.410 43.140 ;
        RECT 64.470 42.880 64.790 43.140 ;
        RECT 65.850 42.880 66.170 43.140 ;
        RECT 82.425 43.080 82.715 43.125 ;
        RECT 86.105 43.080 86.395 43.125 ;
        RECT 86.550 43.080 86.870 43.140 ;
        RECT 96.670 43.080 96.990 43.140 ;
        RECT 82.425 42.940 86.870 43.080 ;
        RECT 82.425 42.895 82.715 42.940 ;
        RECT 86.105 42.895 86.395 42.940 ;
        RECT 86.550 42.880 86.870 42.940 ;
        RECT 90.780 42.940 96.990 43.080 ;
        RECT 10.205 42.740 10.495 42.785 ;
        RECT 11.570 42.740 11.890 42.800 ;
        RECT 10.205 42.600 11.890 42.740 ;
        RECT 10.205 42.555 10.495 42.600 ;
        RECT 11.570 42.540 11.890 42.600 ;
        RECT 12.485 42.740 13.135 42.785 ;
        RECT 15.250 42.740 15.570 42.800 ;
        RECT 16.085 42.740 16.375 42.785 ;
        RECT 12.485 42.600 16.375 42.740 ;
        RECT 12.485 42.555 13.135 42.600 ;
        RECT 15.250 42.540 15.570 42.600 ;
        RECT 15.785 42.555 16.375 42.600 ;
        RECT 21.690 42.740 22.010 42.800 ;
        RECT 28.605 42.740 28.895 42.785 ;
        RECT 32.730 42.740 33.050 42.800 ;
        RECT 34.110 42.740 34.430 42.800 ;
        RECT 38.265 42.740 38.555 42.785 ;
        RECT 21.690 42.600 26.980 42.740 ;
        RECT 9.290 42.400 9.580 42.445 ;
        RECT 11.125 42.400 11.415 42.445 ;
        RECT 14.705 42.400 14.995 42.445 ;
        RECT 9.290 42.260 14.995 42.400 ;
        RECT 9.290 42.215 9.580 42.260 ;
        RECT 11.125 42.215 11.415 42.260 ;
        RECT 14.705 42.215 14.995 42.260 ;
        RECT 15.785 42.240 16.075 42.555 ;
        RECT 21.690 42.540 22.010 42.600 ;
        RECT 18.930 42.200 19.250 42.460 ;
        RECT 24.925 42.400 25.215 42.445 ;
        RECT 24.925 42.260 26.520 42.400 ;
        RECT 24.925 42.215 25.215 42.260 ;
        RECT 8.810 41.860 9.130 42.120 ;
        RECT 17.565 42.060 17.855 42.105 ;
        RECT 21.230 42.060 21.550 42.120 ;
        RECT 17.565 41.920 21.550 42.060 ;
        RECT 17.565 41.875 17.855 41.920 ;
        RECT 21.230 41.860 21.550 41.920 ;
        RECT 26.380 41.765 26.520 42.260 ;
        RECT 26.840 42.060 26.980 42.600 ;
        RECT 28.605 42.600 38.555 42.740 ;
        RECT 28.605 42.555 28.895 42.600 ;
        RECT 32.730 42.540 33.050 42.600 ;
        RECT 34.110 42.540 34.430 42.600 ;
        RECT 38.265 42.555 38.555 42.600 ;
        RECT 38.725 42.740 39.015 42.785 ;
        RECT 43.325 42.740 43.615 42.785 ;
        RECT 44.230 42.740 44.550 42.800 ;
        RECT 76.430 42.740 76.750 42.800 ;
        RECT 38.725 42.600 44.550 42.740 ;
        RECT 38.725 42.555 39.015 42.600 ;
        RECT 43.325 42.555 43.615 42.600 ;
        RECT 44.230 42.540 44.550 42.600 ;
        RECT 73.760 42.600 76.750 42.740 ;
        RECT 59.425 42.400 59.715 42.445 ;
        RECT 60.790 42.400 61.110 42.460 ;
        RECT 73.760 42.445 73.900 42.600 ;
        RECT 76.430 42.540 76.750 42.600 ;
        RECT 77.345 42.740 77.995 42.785 ;
        RECT 80.945 42.740 81.235 42.785 ;
        RECT 77.345 42.600 81.235 42.740 ;
        RECT 77.345 42.555 77.995 42.600 ;
        RECT 80.645 42.555 81.235 42.600 ;
        RECT 80.645 42.460 80.935 42.555 ;
        RECT 59.425 42.260 61.110 42.400 ;
        RECT 59.425 42.215 59.715 42.260 ;
        RECT 60.790 42.200 61.110 42.260 ;
        RECT 65.405 42.215 65.695 42.445 ;
        RECT 73.685 42.215 73.975 42.445 ;
        RECT 74.150 42.400 74.440 42.445 ;
        RECT 75.985 42.400 76.275 42.445 ;
        RECT 79.565 42.400 79.855 42.445 ;
        RECT 74.150 42.260 79.855 42.400 ;
        RECT 74.150 42.215 74.440 42.260 ;
        RECT 75.985 42.215 76.275 42.260 ;
        RECT 79.565 42.215 79.855 42.260 ;
        RECT 80.570 42.240 80.935 42.460 ;
        RECT 86.565 42.400 86.855 42.445 ;
        RECT 89.770 42.400 90.090 42.460 ;
        RECT 90.780 42.445 90.920 42.940 ;
        RECT 96.670 42.880 96.990 42.940 ;
        RECT 99.430 42.880 99.750 43.140 ;
        RECT 105.870 42.880 106.190 43.140 ;
        RECT 106.790 43.080 107.110 43.140 ;
        RECT 106.790 42.940 110.700 43.080 ;
        RECT 106.790 42.880 107.110 42.940 ;
        RECT 92.070 42.540 92.390 42.800 ;
        RECT 94.365 42.740 95.015 42.785 ;
        RECT 97.130 42.740 97.450 42.800 ;
        RECT 97.965 42.740 98.255 42.785 ;
        RECT 94.365 42.600 98.255 42.740 ;
        RECT 94.365 42.555 95.015 42.600 ;
        RECT 97.130 42.540 97.450 42.600 ;
        RECT 97.665 42.555 98.255 42.600 ;
        RECT 102.190 42.740 102.510 42.800 ;
        RECT 110.560 42.785 110.700 42.940 ;
        RECT 102.190 42.600 109.320 42.740 ;
        RECT 86.565 42.260 90.090 42.400 ;
        RECT 27.210 42.060 27.530 42.120 ;
        RECT 29.065 42.060 29.355 42.105 ;
        RECT 39.645 42.060 39.935 42.105 ;
        RECT 44.705 42.060 44.995 42.105 ;
        RECT 46.990 42.060 47.310 42.120 ;
        RECT 26.840 41.920 47.310 42.060 ;
        RECT 27.210 41.860 27.530 41.920 ;
        RECT 29.065 41.875 29.355 41.920 ;
        RECT 39.645 41.875 39.935 41.920 ;
        RECT 44.705 41.875 44.995 41.920 ;
        RECT 46.990 41.860 47.310 41.920 ;
        RECT 61.265 42.060 61.555 42.105 ;
        RECT 62.170 42.060 62.490 42.120 ;
        RECT 61.265 41.920 62.490 42.060 ;
        RECT 61.265 41.875 61.555 41.920 ;
        RECT 62.170 41.860 62.490 41.920 ;
        RECT 62.630 41.860 62.950 42.120 ;
        RECT 63.550 42.105 63.870 42.120 ;
        RECT 63.550 42.060 63.980 42.105 ;
        RECT 65.480 42.060 65.620 42.215 ;
        RECT 80.570 42.200 80.890 42.240 ;
        RECT 86.565 42.215 86.855 42.260 ;
        RECT 89.770 42.200 90.090 42.260 ;
        RECT 90.705 42.215 90.995 42.445 ;
        RECT 91.170 42.400 91.460 42.445 ;
        RECT 93.005 42.400 93.295 42.445 ;
        RECT 96.585 42.400 96.875 42.445 ;
        RECT 91.170 42.260 96.875 42.400 ;
        RECT 91.170 42.215 91.460 42.260 ;
        RECT 93.005 42.215 93.295 42.260 ;
        RECT 96.585 42.215 96.875 42.260 ;
        RECT 97.665 42.240 97.955 42.555 ;
        RECT 102.190 42.540 102.510 42.600 ;
        RECT 101.730 42.400 102.050 42.460 ;
        RECT 109.180 42.445 109.320 42.600 ;
        RECT 110.485 42.555 110.775 42.785 ;
        RECT 111.850 42.740 112.170 42.800 ;
        RECT 112.765 42.740 113.415 42.785 ;
        RECT 116.365 42.740 116.655 42.785 ;
        RECT 111.850 42.600 116.655 42.740 ;
        RECT 111.850 42.540 112.170 42.600 ;
        RECT 112.765 42.555 113.415 42.600 ;
        RECT 116.065 42.555 116.655 42.600 ;
        RECT 106.345 42.400 106.635 42.445 ;
        RECT 101.730 42.260 106.635 42.400 ;
        RECT 101.730 42.200 102.050 42.260 ;
        RECT 106.345 42.215 106.635 42.260 ;
        RECT 109.105 42.215 109.395 42.445 ;
        RECT 109.570 42.400 109.860 42.445 ;
        RECT 111.405 42.400 111.695 42.445 ;
        RECT 114.985 42.400 115.275 42.445 ;
        RECT 109.570 42.260 115.275 42.400 ;
        RECT 109.570 42.215 109.860 42.260 ;
        RECT 111.405 42.215 111.695 42.260 ;
        RECT 114.985 42.215 115.275 42.260 ;
        RECT 116.065 42.240 116.355 42.555 ;
        RECT 63.550 41.920 65.620 42.060 ;
        RECT 63.550 41.875 63.980 41.920 ;
        RECT 63.550 41.860 63.870 41.875 ;
        RECT 75.050 41.860 75.370 42.120 ;
        RECT 87.010 41.860 87.330 42.120 ;
        RECT 104.950 41.860 105.270 42.120 ;
        RECT 105.870 42.060 106.190 42.120 ;
        RECT 117.845 42.060 118.135 42.105 ;
        RECT 105.870 41.920 118.135 42.060 ;
        RECT 105.870 41.860 106.190 41.920 ;
        RECT 117.845 41.875 118.135 41.920 ;
        RECT 9.695 41.720 9.985 41.765 ;
        RECT 11.585 41.720 11.875 41.765 ;
        RECT 14.705 41.720 14.995 41.765 ;
        RECT 9.695 41.580 14.995 41.720 ;
        RECT 9.695 41.535 9.985 41.580 ;
        RECT 11.585 41.535 11.875 41.580 ;
        RECT 14.705 41.535 14.995 41.580 ;
        RECT 26.305 41.535 26.595 41.765 ;
        RECT 74.555 41.720 74.845 41.765 ;
        RECT 76.445 41.720 76.735 41.765 ;
        RECT 79.565 41.720 79.855 41.765 ;
        RECT 74.555 41.580 79.855 41.720 ;
        RECT 74.555 41.535 74.845 41.580 ;
        RECT 76.445 41.535 76.735 41.580 ;
        RECT 79.565 41.535 79.855 41.580 ;
        RECT 91.575 41.720 91.865 41.765 ;
        RECT 93.465 41.720 93.755 41.765 ;
        RECT 96.585 41.720 96.875 41.765 ;
        RECT 91.575 41.580 96.875 41.720 ;
        RECT 91.575 41.535 91.865 41.580 ;
        RECT 93.465 41.535 93.755 41.580 ;
        RECT 96.585 41.535 96.875 41.580 ;
        RECT 108.170 41.520 108.490 41.780 ;
        RECT 109.975 41.720 110.265 41.765 ;
        RECT 111.865 41.720 112.155 41.765 ;
        RECT 114.985 41.720 115.275 41.765 ;
        RECT 109.975 41.580 115.275 41.720 ;
        RECT 109.975 41.535 110.265 41.580 ;
        RECT 111.865 41.535 112.155 41.580 ;
        RECT 114.985 41.535 115.275 41.580 ;
        RECT 25.845 41.380 26.135 41.425 ;
        RECT 26.750 41.380 27.070 41.440 ;
        RECT 25.845 41.240 27.070 41.380 ;
        RECT 25.845 41.195 26.135 41.240 ;
        RECT 26.750 41.180 27.070 41.240 ;
        RECT 41.485 41.380 41.775 41.425 ;
        RECT 41.930 41.380 42.250 41.440 ;
        RECT 41.485 41.240 42.250 41.380 ;
        RECT 41.485 41.195 41.775 41.240 ;
        RECT 41.930 41.180 42.250 41.240 ;
        RECT 83.790 41.380 84.110 41.440 ;
        RECT 84.265 41.380 84.555 41.425 ;
        RECT 83.790 41.240 84.555 41.380 ;
        RECT 83.790 41.180 84.110 41.240 ;
        RECT 84.265 41.195 84.555 41.240 ;
        RECT 5.520 40.560 123.740 41.040 ;
        RECT 34.110 40.160 34.430 40.420 ;
        RECT 60.345 40.360 60.635 40.405 ;
        RECT 63.550 40.360 63.870 40.420 ;
        RECT 60.345 40.220 63.870 40.360 ;
        RECT 60.345 40.175 60.635 40.220 ;
        RECT 63.550 40.160 63.870 40.220 ;
        RECT 89.770 40.360 90.090 40.420 ;
        RECT 91.610 40.360 91.930 40.420 ;
        RECT 89.770 40.220 91.930 40.360 ;
        RECT 89.770 40.160 90.090 40.220 ;
        RECT 91.610 40.160 91.930 40.220 ;
        RECT 96.685 40.360 96.975 40.405 ;
        RECT 97.130 40.360 97.450 40.420 ;
        RECT 96.685 40.220 97.450 40.360 ;
        RECT 96.685 40.175 96.975 40.220 ;
        RECT 97.130 40.160 97.450 40.220 ;
        RECT 111.850 40.160 112.170 40.420 ;
        RECT 26.255 40.020 26.545 40.065 ;
        RECT 28.145 40.020 28.435 40.065 ;
        RECT 31.265 40.020 31.555 40.065 ;
        RECT 26.255 39.880 31.555 40.020 ;
        RECT 26.255 39.835 26.545 39.880 ;
        RECT 28.145 39.835 28.435 39.880 ;
        RECT 31.265 39.835 31.555 39.880 ;
        RECT 52.475 40.020 52.765 40.065 ;
        RECT 54.365 40.020 54.655 40.065 ;
        RECT 57.485 40.020 57.775 40.065 ;
        RECT 52.475 39.880 57.775 40.020 ;
        RECT 52.475 39.835 52.765 39.880 ;
        RECT 54.365 39.835 54.655 39.880 ;
        RECT 57.485 39.835 57.775 39.880 ;
        RECT 81.915 40.020 82.205 40.065 ;
        RECT 83.805 40.020 84.095 40.065 ;
        RECT 86.925 40.020 87.215 40.065 ;
        RECT 81.915 39.880 87.215 40.020 ;
        RECT 81.915 39.835 82.205 39.880 ;
        RECT 83.805 39.835 84.095 39.880 ;
        RECT 86.925 39.835 87.215 39.880 ;
        RECT 103.075 40.020 103.365 40.065 ;
        RECT 104.965 40.020 105.255 40.065 ;
        RECT 108.085 40.020 108.375 40.065 ;
        RECT 103.075 39.880 108.375 40.020 ;
        RECT 103.075 39.835 103.365 39.880 ;
        RECT 104.965 39.835 105.255 39.880 ;
        RECT 108.085 39.835 108.375 39.880 ;
        RECT 26.750 39.480 27.070 39.740 ;
        RECT 45.610 39.680 45.930 39.740 ;
        RECT 35.580 39.540 45.930 39.680 ;
        RECT 23.530 39.340 23.850 39.400 ;
        RECT 35.580 39.385 35.720 39.540 ;
        RECT 45.610 39.480 45.930 39.540 ;
        RECT 48.370 39.680 48.690 39.740 ;
        RECT 51.590 39.680 51.910 39.740 ;
        RECT 48.370 39.540 51.910 39.680 ;
        RECT 48.370 39.480 48.690 39.540 ;
        RECT 51.590 39.480 51.910 39.540 ;
        RECT 76.890 39.680 77.210 39.740 ;
        RECT 81.045 39.680 81.335 39.725 ;
        RECT 76.890 39.540 81.335 39.680 ;
        RECT 76.890 39.480 77.210 39.540 ;
        RECT 81.045 39.495 81.335 39.540 ;
        RECT 96.670 39.680 96.990 39.740 ;
        RECT 102.190 39.680 102.510 39.740 ;
        RECT 96.670 39.540 102.510 39.680 ;
        RECT 96.670 39.480 96.990 39.540 ;
        RECT 102.190 39.480 102.510 39.540 ;
        RECT 25.385 39.340 25.675 39.385 ;
        RECT 23.530 39.200 25.675 39.340 ;
        RECT 23.530 39.140 23.850 39.200 ;
        RECT 25.385 39.155 25.675 39.200 ;
        RECT 25.850 39.340 26.140 39.385 ;
        RECT 27.685 39.340 27.975 39.385 ;
        RECT 31.265 39.340 31.555 39.385 ;
        RECT 25.850 39.200 31.555 39.340 ;
        RECT 25.850 39.155 26.140 39.200 ;
        RECT 27.685 39.155 27.975 39.200 ;
        RECT 31.265 39.155 31.555 39.200 ;
        RECT 32.345 39.045 32.635 39.360 ;
        RECT 35.505 39.155 35.795 39.385 ;
        RECT 40.565 39.340 40.855 39.385 ;
        RECT 41.930 39.340 42.250 39.400 ;
        RECT 40.565 39.200 42.250 39.340 ;
        RECT 40.565 39.155 40.855 39.200 ;
        RECT 41.930 39.140 42.250 39.200 ;
        RECT 52.070 39.340 52.360 39.385 ;
        RECT 53.905 39.340 54.195 39.385 ;
        RECT 57.485 39.340 57.775 39.385 ;
        RECT 52.070 39.200 57.775 39.340 ;
        RECT 52.070 39.155 52.360 39.200 ;
        RECT 53.905 39.155 54.195 39.200 ;
        RECT 57.485 39.155 57.775 39.200 ;
        RECT 29.045 39.000 29.695 39.045 ;
        RECT 32.345 39.000 32.935 39.045 ;
        RECT 35.045 39.000 35.335 39.045 ;
        RECT 29.045 38.860 35.335 39.000 ;
        RECT 29.045 38.815 29.695 38.860 ;
        RECT 32.645 38.815 32.935 38.860 ;
        RECT 35.045 38.815 35.335 38.860 ;
        RECT 52.985 38.815 53.275 39.045 ;
        RECT 55.265 39.000 55.915 39.045 ;
        RECT 56.650 39.000 56.970 39.060 ;
        RECT 58.565 39.045 58.855 39.360 ;
        RECT 81.510 39.340 81.800 39.385 ;
        RECT 83.345 39.340 83.635 39.385 ;
        RECT 86.925 39.340 87.215 39.385 ;
        RECT 81.510 39.200 87.215 39.340 ;
        RECT 81.510 39.155 81.800 39.200 ;
        RECT 83.345 39.155 83.635 39.200 ;
        RECT 86.925 39.155 87.215 39.200 ;
        RECT 58.565 39.000 59.155 39.045 ;
        RECT 55.265 38.860 59.155 39.000 ;
        RECT 55.265 38.815 55.915 38.860 ;
        RECT 39.170 38.660 39.490 38.720 ;
        RECT 39.645 38.660 39.935 38.705 ;
        RECT 39.170 38.520 39.935 38.660 ;
        RECT 53.060 38.660 53.200 38.815 ;
        RECT 56.650 38.800 56.970 38.860 ;
        RECT 58.865 38.815 59.155 38.860 ;
        RECT 82.410 38.800 82.730 39.060 ;
        RECT 84.705 39.000 85.355 39.045 ;
        RECT 87.470 39.000 87.790 39.060 ;
        RECT 88.005 39.045 88.295 39.360 ;
        RECT 97.145 39.155 97.435 39.385 ;
        RECT 102.670 39.340 102.960 39.385 ;
        RECT 104.505 39.340 104.795 39.385 ;
        RECT 108.085 39.340 108.375 39.385 ;
        RECT 102.670 39.200 108.375 39.340 ;
        RECT 102.670 39.155 102.960 39.200 ;
        RECT 104.505 39.155 104.795 39.200 ;
        RECT 108.085 39.155 108.375 39.200 ;
        RECT 109.090 39.360 109.410 39.400 ;
        RECT 88.005 39.000 88.595 39.045 ;
        RECT 84.705 38.860 88.595 39.000 ;
        RECT 84.705 38.815 85.355 38.860 ;
        RECT 87.470 38.800 87.790 38.860 ;
        RECT 88.305 38.815 88.595 38.860 ;
        RECT 57.570 38.660 57.890 38.720 ;
        RECT 53.060 38.520 57.890 38.660 ;
        RECT 97.220 38.660 97.360 39.155 ;
        RECT 109.090 39.140 109.455 39.360 ;
        RECT 110.010 39.340 110.330 39.400 ;
        RECT 111.405 39.340 111.695 39.385 ;
        RECT 110.010 39.200 111.695 39.340 ;
        RECT 110.010 39.140 110.330 39.200 ;
        RECT 111.405 39.155 111.695 39.200 ;
        RECT 103.110 39.000 103.430 39.060 ;
        RECT 109.165 39.045 109.455 39.140 ;
        RECT 103.585 39.000 103.875 39.045 ;
        RECT 103.110 38.860 103.875 39.000 ;
        RECT 103.110 38.800 103.430 38.860 ;
        RECT 103.585 38.815 103.875 38.860 ;
        RECT 105.865 39.000 106.515 39.045 ;
        RECT 109.165 39.000 109.755 39.045 ;
        RECT 105.865 38.860 109.755 39.000 ;
        RECT 105.865 38.815 106.515 38.860 ;
        RECT 109.465 38.815 109.755 38.860 ;
        RECT 97.590 38.660 97.910 38.720 ;
        RECT 110.100 38.660 110.240 39.140 ;
        RECT 97.220 38.520 110.240 38.660 ;
        RECT 39.170 38.460 39.490 38.520 ;
        RECT 39.645 38.475 39.935 38.520 ;
        RECT 57.570 38.460 57.890 38.520 ;
        RECT 97.590 38.460 97.910 38.520 ;
        RECT 110.930 38.460 111.250 38.720 ;
        RECT 5.520 37.840 123.740 38.320 ;
        RECT 43.770 37.640 44.090 37.700 ;
        RECT 46.545 37.640 46.835 37.685 ;
        RECT 43.770 37.500 46.835 37.640 ;
        RECT 43.770 37.440 44.090 37.500 ;
        RECT 46.545 37.455 46.835 37.500 ;
        RECT 48.830 37.640 49.150 37.700 ;
        RECT 49.305 37.640 49.595 37.685 ;
        RECT 50.670 37.640 50.990 37.700 ;
        RECT 48.830 37.500 50.990 37.640 ;
        RECT 39.170 37.100 39.490 37.360 ;
        RECT 41.465 37.300 42.115 37.345 ;
        RECT 42.850 37.300 43.170 37.360 ;
        RECT 45.065 37.300 45.355 37.345 ;
        RECT 41.465 37.160 45.355 37.300 ;
        RECT 41.465 37.115 42.115 37.160 ;
        RECT 42.850 37.100 43.170 37.160 ;
        RECT 44.765 37.115 45.355 37.160 ;
        RECT 36.870 36.960 37.190 37.020 ;
        RECT 37.790 36.960 38.110 37.020 ;
        RECT 36.870 36.820 38.110 36.960 ;
        RECT 36.870 36.760 37.190 36.820 ;
        RECT 37.790 36.760 38.110 36.820 ;
        RECT 38.270 36.960 38.560 37.005 ;
        RECT 40.105 36.960 40.395 37.005 ;
        RECT 43.685 36.960 43.975 37.005 ;
        RECT 38.270 36.820 43.975 36.960 ;
        RECT 38.270 36.775 38.560 36.820 ;
        RECT 40.105 36.775 40.395 36.820 ;
        RECT 43.685 36.775 43.975 36.820 ;
        RECT 44.765 36.800 45.055 37.115 ;
        RECT 46.620 36.960 46.760 37.455 ;
        RECT 48.830 37.440 49.150 37.500 ;
        RECT 49.305 37.455 49.595 37.500 ;
        RECT 50.670 37.440 50.990 37.500 ;
        RECT 56.205 37.640 56.495 37.685 ;
        RECT 56.650 37.640 56.970 37.700 ;
        RECT 56.205 37.500 56.970 37.640 ;
        RECT 56.205 37.455 56.495 37.500 ;
        RECT 56.650 37.440 56.970 37.500 ;
        RECT 57.570 37.440 57.890 37.700 ;
        RECT 62.170 37.640 62.490 37.700 ;
        RECT 65.390 37.640 65.710 37.700 ;
        RECT 82.410 37.640 82.730 37.700 ;
        RECT 83.345 37.640 83.635 37.685 ;
        RECT 62.170 37.500 72.520 37.640 ;
        RECT 62.170 37.440 62.490 37.500 ;
        RECT 65.390 37.440 65.710 37.500 ;
        RECT 64.010 37.300 64.330 37.360 ;
        RECT 64.485 37.300 64.775 37.345 ;
        RECT 68.610 37.300 68.930 37.360 ;
        RECT 64.010 37.160 68.930 37.300 ;
        RECT 64.010 37.100 64.330 37.160 ;
        RECT 64.485 37.115 64.775 37.160 ;
        RECT 68.610 37.100 68.930 37.160 ;
        RECT 48.845 36.960 49.135 37.005 ;
        RECT 46.620 36.820 49.135 36.960 ;
        RECT 48.845 36.775 49.135 36.820 ;
        RECT 55.745 36.960 56.035 37.005 ;
        RECT 57.110 36.960 57.430 37.020 ;
        RECT 55.745 36.820 57.430 36.960 ;
        RECT 55.745 36.775 56.035 36.820 ;
        RECT 57.110 36.760 57.430 36.820 ;
        RECT 58.490 36.760 58.810 37.020 ;
        RECT 63.565 36.960 63.855 37.005 ;
        RECT 64.930 36.960 65.250 37.020 ;
        RECT 65.850 36.960 66.170 37.020 ;
        RECT 67.705 36.960 67.995 37.005 ;
        RECT 63.565 36.820 67.995 36.960 ;
        RECT 68.700 36.960 68.840 37.100 ;
        RECT 69.545 36.960 69.835 37.005 ;
        RECT 71.385 36.960 71.675 37.005 ;
        RECT 68.700 36.820 71.675 36.960 ;
        RECT 63.565 36.775 63.855 36.820 ;
        RECT 64.930 36.760 65.250 36.820 ;
        RECT 65.850 36.760 66.170 36.820 ;
        RECT 67.705 36.775 67.995 36.820 ;
        RECT 69.545 36.775 69.835 36.820 ;
        RECT 71.385 36.775 71.675 36.820 ;
        RECT 46.990 36.620 47.310 36.680 ;
        RECT 49.765 36.620 50.055 36.665 ;
        RECT 46.990 36.480 50.055 36.620 ;
        RECT 46.990 36.420 47.310 36.480 ;
        RECT 49.765 36.435 50.055 36.480 ;
        RECT 38.675 36.280 38.965 36.325 ;
        RECT 40.565 36.280 40.855 36.325 ;
        RECT 43.685 36.280 43.975 36.325 ;
        RECT 38.675 36.140 43.975 36.280 ;
        RECT 67.780 36.280 67.920 36.775 ;
        RECT 68.610 36.620 68.930 36.680 ;
        RECT 72.380 36.665 72.520 37.500 ;
        RECT 82.410 37.500 83.635 37.640 ;
        RECT 82.410 37.440 82.730 37.500 ;
        RECT 83.345 37.455 83.635 37.500 ;
        RECT 85.185 37.640 85.475 37.685 ;
        RECT 87.470 37.640 87.790 37.700 ;
        RECT 85.185 37.500 87.790 37.640 ;
        RECT 85.185 37.455 85.475 37.500 ;
        RECT 87.470 37.440 87.790 37.500 ;
        RECT 103.110 37.440 103.430 37.700 ;
        RECT 103.585 37.455 103.875 37.685 ;
        RECT 105.425 37.640 105.715 37.685 ;
        RECT 105.870 37.640 106.190 37.700 ;
        RECT 105.425 37.500 106.190 37.640 ;
        RECT 105.425 37.455 105.715 37.500 ;
        RECT 82.870 37.300 83.190 37.360 ;
        RECT 82.870 37.160 84.940 37.300 ;
        RECT 82.870 37.100 83.190 37.160 ;
        RECT 83.790 36.960 84.110 37.020 ;
        RECT 84.800 37.005 84.940 37.160 ;
        RECT 84.265 36.960 84.555 37.005 ;
        RECT 83.790 36.820 84.555 36.960 ;
        RECT 83.790 36.760 84.110 36.820 ;
        RECT 84.265 36.775 84.555 36.820 ;
        RECT 84.725 36.775 85.015 37.005 ;
        RECT 97.590 36.760 97.910 37.020 ;
        RECT 102.205 36.960 102.495 37.005 ;
        RECT 103.660 36.960 103.800 37.455 ;
        RECT 105.870 37.440 106.190 37.500 ;
        RECT 109.090 37.640 109.410 37.700 ;
        RECT 109.565 37.640 109.855 37.685 ;
        RECT 109.090 37.500 109.855 37.640 ;
        RECT 109.090 37.440 109.410 37.500 ;
        RECT 109.565 37.455 109.855 37.500 ;
        RECT 110.930 37.300 111.250 37.360 ;
        RECT 102.205 36.820 103.800 36.960 ;
        RECT 105.960 37.160 111.250 37.300 ;
        RECT 102.205 36.775 102.495 36.820 ;
        RECT 70.925 36.620 71.215 36.665 ;
        RECT 68.610 36.480 71.215 36.620 ;
        RECT 68.610 36.420 68.930 36.480 ;
        RECT 70.925 36.435 71.215 36.480 ;
        RECT 71.845 36.435 72.135 36.665 ;
        RECT 72.305 36.620 72.595 36.665 ;
        RECT 75.050 36.620 75.370 36.680 ;
        RECT 72.305 36.480 75.370 36.620 ;
        RECT 72.305 36.435 72.595 36.480 ;
        RECT 71.920 36.280 72.060 36.435 ;
        RECT 75.050 36.420 75.370 36.480 ;
        RECT 98.510 36.620 98.830 36.680 ;
        RECT 105.960 36.665 106.100 37.160 ;
        RECT 110.930 37.100 111.250 37.160 ;
        RECT 110.010 36.760 110.330 37.020 ;
        RECT 105.885 36.620 106.175 36.665 ;
        RECT 98.510 36.480 106.175 36.620 ;
        RECT 98.510 36.420 98.830 36.480 ;
        RECT 105.885 36.435 106.175 36.480 ;
        RECT 106.345 36.435 106.635 36.665 ;
        RECT 67.780 36.140 72.060 36.280 ;
        RECT 104.950 36.280 105.270 36.340 ;
        RECT 106.420 36.280 106.560 36.435 ;
        RECT 104.950 36.140 106.560 36.280 ;
        RECT 38.675 36.095 38.965 36.140 ;
        RECT 40.565 36.095 40.855 36.140 ;
        RECT 43.685 36.095 43.975 36.140 ;
        RECT 104.950 36.080 105.270 36.140 ;
        RECT 46.990 35.740 47.310 36.000 ;
        RECT 61.710 35.940 62.030 36.000 ;
        RECT 62.645 35.940 62.935 35.985 ;
        RECT 61.710 35.800 62.935 35.940 ;
        RECT 61.710 35.740 62.030 35.800 ;
        RECT 62.645 35.755 62.935 35.800 ;
        RECT 66.770 35.740 67.090 36.000 ;
        RECT 68.150 35.740 68.470 36.000 ;
        RECT 70.005 35.940 70.295 35.985 ;
        RECT 71.830 35.940 72.150 36.000 ;
        RECT 70.005 35.800 72.150 35.940 ;
        RECT 70.005 35.755 70.295 35.800 ;
        RECT 71.830 35.740 72.150 35.800 ;
        RECT 98.050 35.740 98.370 36.000 ;
        RECT 5.520 35.120 123.740 35.600 ;
        RECT 58.490 34.920 58.810 34.980 ;
        RECT 60.805 34.920 61.095 34.965 ;
        RECT 58.490 34.780 61.095 34.920 ;
        RECT 58.490 34.720 58.810 34.780 ;
        RECT 60.805 34.735 61.095 34.780 ;
        RECT 61.710 34.720 62.030 34.980 ;
        RECT 63.550 34.920 63.870 34.980 ;
        RECT 65.865 34.920 66.155 34.965 ;
        RECT 68.610 34.920 68.930 34.980 ;
        RECT 63.550 34.780 68.930 34.920 ;
        RECT 63.550 34.720 63.870 34.780 ;
        RECT 65.865 34.735 66.155 34.780 ;
        RECT 68.610 34.720 68.930 34.780 ;
        RECT 71.385 34.735 71.675 34.965 ;
        RECT 64.010 34.580 64.330 34.640 ;
        RECT 22.240 34.440 26.520 34.580 ;
        RECT 18.010 34.240 18.330 34.300 ;
        RECT 22.240 34.285 22.380 34.440 ;
        RECT 26.380 34.285 26.520 34.440 ;
        RECT 59.960 34.440 64.330 34.580 ;
        RECT 21.245 34.240 21.535 34.285 ;
        RECT 18.010 34.100 21.535 34.240 ;
        RECT 18.010 34.040 18.330 34.100 ;
        RECT 21.245 34.055 21.535 34.100 ;
        RECT 22.165 34.240 22.455 34.285 ;
        RECT 26.305 34.240 26.595 34.285 ;
        RECT 27.210 34.240 27.530 34.300 ;
        RECT 22.165 34.100 22.565 34.240 ;
        RECT 26.195 34.100 27.530 34.240 ;
        RECT 22.165 34.055 22.455 34.100 ;
        RECT 26.305 34.055 26.595 34.100 ;
        RECT 27.210 34.040 27.530 34.100 ;
        RECT 42.850 34.040 43.170 34.300 ;
        RECT 59.960 34.240 60.100 34.440 ;
        RECT 64.010 34.380 64.330 34.440 ;
        RECT 64.485 34.395 64.775 34.625 ;
        RECT 70.465 34.395 70.755 34.625 ;
        RECT 64.560 34.240 64.700 34.395 ;
        RECT 59.500 34.100 60.100 34.240 ;
        RECT 60.420 34.100 64.240 34.240 ;
        RECT 64.560 34.100 66.540 34.240 ;
        RECT 16.185 33.900 16.475 33.945 ;
        RECT 24.925 33.900 25.215 33.945 ;
        RECT 27.670 33.900 27.990 33.960 ;
        RECT 16.185 33.760 19.160 33.900 ;
        RECT 16.185 33.715 16.475 33.760 ;
        RECT 10.650 33.220 10.970 33.280 ;
        RECT 19.020 33.265 19.160 33.760 ;
        RECT 24.925 33.760 27.990 33.900 ;
        RECT 24.925 33.715 25.215 33.760 ;
        RECT 27.670 33.700 27.990 33.760 ;
        RECT 41.945 33.715 42.235 33.945 ;
        RECT 42.390 33.900 42.710 33.960 ;
        RECT 45.610 33.900 45.930 33.960 ;
        RECT 59.500 33.945 59.640 34.100 ;
        RECT 60.420 33.945 60.560 34.100 ;
        RECT 42.390 33.760 45.930 33.900 ;
        RECT 20.785 33.560 21.075 33.605 ;
        RECT 23.990 33.560 24.310 33.620 ;
        RECT 42.020 33.560 42.160 33.715 ;
        RECT 42.390 33.700 42.710 33.760 ;
        RECT 45.610 33.700 45.930 33.760 ;
        RECT 59.425 33.715 59.715 33.945 ;
        RECT 60.345 33.715 60.635 33.945 ;
        RECT 62.170 33.900 62.490 33.960 ;
        RECT 63.105 33.900 63.395 33.945 ;
        RECT 62.170 33.760 63.395 33.900 ;
        RECT 64.100 33.900 64.240 34.100 ;
        RECT 64.930 33.900 65.250 33.960 ;
        RECT 64.100 33.760 65.250 33.900 ;
        RECT 62.170 33.700 62.490 33.760 ;
        RECT 63.105 33.715 63.395 33.760 ;
        RECT 64.930 33.700 65.250 33.760 ;
        RECT 65.390 33.700 65.710 33.960 ;
        RECT 66.400 33.900 66.540 34.100 ;
        RECT 66.770 34.040 67.090 34.300 ;
        RECT 67.230 34.240 67.550 34.300 ;
        RECT 70.540 34.240 70.680 34.395 ;
        RECT 67.230 34.100 70.680 34.240 ;
        RECT 67.230 34.040 67.550 34.100 ;
        RECT 69.070 33.900 69.390 33.960 ;
        RECT 71.460 33.900 71.600 34.735 ;
        RECT 95.305 34.395 95.595 34.625 ;
        RECT 96.690 34.580 96.980 34.625 ;
        RECT 98.550 34.580 98.840 34.625 ;
        RECT 101.330 34.580 101.620 34.625 ;
        RECT 96.690 34.440 101.620 34.580 ;
        RECT 96.690 34.395 96.980 34.440 ;
        RECT 98.550 34.395 98.840 34.440 ;
        RECT 101.330 34.395 101.620 34.440 ;
        RECT 88.390 34.240 88.710 34.300 ;
        RECT 92.545 34.240 92.835 34.285 ;
        RECT 88.390 34.100 92.835 34.240 ;
        RECT 88.390 34.040 88.710 34.100 ;
        RECT 92.545 34.055 92.835 34.100 ;
        RECT 93.450 34.040 93.770 34.300 ;
        RECT 95.380 34.240 95.520 34.395 ;
        RECT 98.065 34.240 98.355 34.285 ;
        RECT 95.380 34.100 98.355 34.240 ;
        RECT 98.065 34.055 98.355 34.100 ;
        RECT 102.650 34.240 102.970 34.300 ;
        RECT 105.195 34.240 105.485 34.285 ;
        RECT 102.650 34.100 105.485 34.240 ;
        RECT 102.650 34.040 102.970 34.100 ;
        RECT 105.195 34.055 105.485 34.100 ;
        RECT 66.400 33.760 71.600 33.900 ;
        RECT 94.385 33.900 94.675 33.945 ;
        RECT 94.830 33.900 95.150 33.960 ;
        RECT 94.385 33.760 95.150 33.900 ;
        RECT 69.070 33.700 69.390 33.760 ;
        RECT 94.385 33.715 94.675 33.760 ;
        RECT 94.830 33.700 95.150 33.760 ;
        RECT 96.225 33.900 96.515 33.945 ;
        RECT 96.670 33.900 96.990 33.960 ;
        RECT 101.330 33.900 101.620 33.945 ;
        RECT 96.225 33.760 96.990 33.900 ;
        RECT 96.225 33.715 96.515 33.760 ;
        RECT 96.670 33.700 96.990 33.760 ;
        RECT 99.085 33.760 101.620 33.900 ;
        RECT 46.990 33.560 47.310 33.620 ;
        RECT 20.785 33.420 25.600 33.560 ;
        RECT 42.020 33.420 47.310 33.560 ;
        RECT 20.785 33.375 21.075 33.420 ;
        RECT 23.990 33.360 24.310 33.420 ;
        RECT 15.265 33.220 15.555 33.265 ;
        RECT 10.650 33.080 15.555 33.220 ;
        RECT 10.650 33.020 10.970 33.080 ;
        RECT 15.265 33.035 15.555 33.080 ;
        RECT 18.945 33.035 19.235 33.265 ;
        RECT 23.070 33.020 23.390 33.280 ;
        RECT 25.460 33.265 25.600 33.420 ;
        RECT 46.990 33.360 47.310 33.420 ;
        RECT 59.870 33.560 60.190 33.620 ;
        RECT 62.645 33.560 62.935 33.605 ;
        RECT 71.305 33.560 71.595 33.605 ;
        RECT 71.830 33.560 72.150 33.620 ;
        RECT 99.085 33.605 99.300 33.760 ;
        RECT 101.330 33.715 101.620 33.760 ;
        RECT 59.870 33.420 62.935 33.560 ;
        RECT 59.870 33.360 60.190 33.420 ;
        RECT 62.645 33.375 62.935 33.420 ;
        RECT 63.180 33.420 65.620 33.560 ;
        RECT 25.385 33.220 25.675 33.265 ;
        RECT 27.210 33.220 27.530 33.280 ;
        RECT 25.385 33.080 27.530 33.220 ;
        RECT 25.385 33.035 25.675 33.080 ;
        RECT 27.210 33.020 27.530 33.080 ;
        RECT 41.010 33.020 41.330 33.280 ;
        RECT 45.150 33.020 45.470 33.280 ;
        RECT 61.645 33.220 61.935 33.265 ;
        RECT 63.180 33.220 63.320 33.420 ;
        RECT 61.645 33.080 63.320 33.220 ;
        RECT 61.645 33.035 61.935 33.080 ;
        RECT 63.550 33.020 63.870 33.280 ;
        RECT 64.010 33.020 64.330 33.280 ;
        RECT 65.480 33.220 65.620 33.420 ;
        RECT 71.305 33.420 72.150 33.560 ;
        RECT 71.305 33.375 71.595 33.420 ;
        RECT 71.830 33.360 72.150 33.420 ;
        RECT 72.305 33.375 72.595 33.605 ;
        RECT 97.150 33.560 97.440 33.605 ;
        RECT 99.010 33.560 99.300 33.605 ;
        RECT 99.930 33.560 100.220 33.605 ;
        RECT 103.190 33.560 103.480 33.605 ;
        RECT 97.150 33.420 99.300 33.560 ;
        RECT 97.150 33.375 97.440 33.420 ;
        RECT 99.010 33.375 99.300 33.420 ;
        RECT 99.520 33.420 103.480 33.560 ;
        RECT 68.165 33.220 68.455 33.265 ;
        RECT 72.380 33.220 72.520 33.375 ;
        RECT 65.480 33.080 72.520 33.220 ;
        RECT 88.850 33.220 89.170 33.280 ;
        RECT 90.245 33.220 90.535 33.265 ;
        RECT 88.850 33.080 90.535 33.220 ;
        RECT 68.165 33.035 68.455 33.080 ;
        RECT 88.850 33.020 89.170 33.080 ;
        RECT 90.245 33.035 90.535 33.080 ;
        RECT 92.085 33.220 92.375 33.265 ;
        RECT 97.590 33.220 97.910 33.280 ;
        RECT 92.085 33.080 97.910 33.220 ;
        RECT 92.085 33.035 92.375 33.080 ;
        RECT 97.590 33.020 97.910 33.080 ;
        RECT 98.050 33.220 98.370 33.280 ;
        RECT 99.520 33.220 99.660 33.420 ;
        RECT 99.930 33.375 100.220 33.420 ;
        RECT 103.190 33.375 103.480 33.420 ;
        RECT 98.050 33.080 99.660 33.220 ;
        RECT 98.050 33.020 98.370 33.080 ;
        RECT 5.520 32.400 123.740 32.880 ;
        RECT 18.010 32.000 18.330 32.260 ;
        RECT 27.210 32.000 27.530 32.260 ;
        RECT 31.825 32.015 32.115 32.245 ;
        RECT 46.990 32.200 47.310 32.260 ;
        RECT 34.430 32.060 47.310 32.200 ;
        RECT 10.650 31.660 10.970 31.920 ;
        RECT 12.945 31.860 13.595 31.905 ;
        RECT 16.545 31.860 16.835 31.905 ;
        RECT 17.090 31.860 17.410 31.920 ;
        RECT 12.945 31.720 17.410 31.860 ;
        RECT 12.945 31.675 13.595 31.720 ;
        RECT 16.245 31.675 16.835 31.720 ;
        RECT 9.750 31.520 10.040 31.565 ;
        RECT 11.585 31.520 11.875 31.565 ;
        RECT 15.165 31.520 15.455 31.565 ;
        RECT 9.750 31.380 15.455 31.520 ;
        RECT 9.750 31.335 10.040 31.380 ;
        RECT 11.585 31.335 11.875 31.380 ;
        RECT 15.165 31.335 15.455 31.380 ;
        RECT 16.245 31.360 16.535 31.675 ;
        RECT 17.090 31.660 17.410 31.720 ;
        RECT 22.145 31.860 22.795 31.905 ;
        RECT 24.910 31.860 25.230 31.920 ;
        RECT 25.745 31.860 26.035 31.905 ;
        RECT 22.145 31.720 26.035 31.860 ;
        RECT 22.145 31.675 22.795 31.720 ;
        RECT 24.910 31.660 25.230 31.720 ;
        RECT 25.445 31.675 26.035 31.720 ;
        RECT 18.950 31.520 19.240 31.565 ;
        RECT 20.785 31.520 21.075 31.565 ;
        RECT 24.365 31.520 24.655 31.565 ;
        RECT 18.950 31.380 24.655 31.520 ;
        RECT 18.950 31.335 19.240 31.380 ;
        RECT 20.785 31.335 21.075 31.380 ;
        RECT 24.365 31.335 24.655 31.380 ;
        RECT 25.445 31.360 25.735 31.675 ;
        RECT 29.065 31.520 29.355 31.565 ;
        RECT 31.900 31.520 32.040 32.015 ;
        RECT 33.665 31.860 33.955 31.905 ;
        RECT 34.430 31.860 34.570 32.060 ;
        RECT 46.990 32.000 47.310 32.060 ;
        RECT 47.695 32.200 47.985 32.245 ;
        RECT 48.830 32.200 49.150 32.260 ;
        RECT 47.695 32.060 49.150 32.200 ;
        RECT 47.695 32.015 47.985 32.060 ;
        RECT 48.830 32.000 49.150 32.060 ;
        RECT 61.265 32.200 61.555 32.245 ;
        RECT 63.550 32.200 63.870 32.260 ;
        RECT 61.265 32.060 63.870 32.200 ;
        RECT 61.265 32.015 61.555 32.060 ;
        RECT 33.665 31.720 34.570 31.860 ;
        RECT 39.650 31.860 39.940 31.905 ;
        RECT 41.510 31.860 41.800 31.905 ;
        RECT 39.650 31.720 41.800 31.860 ;
        RECT 33.665 31.675 33.955 31.720 ;
        RECT 39.650 31.675 39.940 31.720 ;
        RECT 41.510 31.675 41.800 31.720 ;
        RECT 42.430 31.860 42.720 31.905 ;
        RECT 43.310 31.860 43.630 31.920 ;
        RECT 45.690 31.860 45.980 31.905 ;
        RECT 42.430 31.720 45.980 31.860 ;
        RECT 42.430 31.675 42.720 31.720 ;
        RECT 29.065 31.380 32.040 31.520 ;
        RECT 37.790 31.520 38.110 31.580 ;
        RECT 38.725 31.520 39.015 31.565 ;
        RECT 37.790 31.380 39.015 31.520 ;
        RECT 29.065 31.335 29.355 31.380 ;
        RECT 37.790 31.320 38.110 31.380 ;
        RECT 38.725 31.335 39.015 31.380 ;
        RECT 40.565 31.520 40.855 31.565 ;
        RECT 41.010 31.520 41.330 31.580 ;
        RECT 40.565 31.380 41.330 31.520 ;
        RECT 41.585 31.520 41.800 31.675 ;
        RECT 43.310 31.660 43.630 31.720 ;
        RECT 45.690 31.675 45.980 31.720 ;
        RECT 43.830 31.520 44.120 31.565 ;
        RECT 41.585 31.380 44.120 31.520 ;
        RECT 40.565 31.335 40.855 31.380 ;
        RECT 41.010 31.320 41.330 31.380 ;
        RECT 43.830 31.335 44.120 31.380 ;
        RECT 46.990 31.520 47.310 31.580 ;
        RECT 47.910 31.520 48.230 31.580 ;
        RECT 46.990 31.380 48.230 31.520 ;
        RECT 46.990 31.320 47.310 31.380 ;
        RECT 47.910 31.320 48.230 31.380 ;
        RECT 59.425 31.520 59.715 31.565 ;
        RECT 61.340 31.520 61.480 32.015 ;
        RECT 63.550 32.000 63.870 32.060 ;
        RECT 66.785 32.200 67.075 32.245 ;
        RECT 83.330 32.200 83.650 32.260 ;
        RECT 85.630 32.200 85.950 32.260 ;
        RECT 66.785 32.060 68.840 32.200 ;
        RECT 66.785 32.015 67.075 32.060 ;
        RECT 67.230 31.660 67.550 31.920 ;
        RECT 68.700 31.905 68.840 32.060 ;
        RECT 83.330 32.060 85.950 32.200 ;
        RECT 83.330 32.000 83.650 32.060 ;
        RECT 85.630 32.000 85.950 32.060 ;
        RECT 94.830 32.000 95.150 32.260 ;
        RECT 97.145 32.200 97.435 32.245 ;
        RECT 97.590 32.200 97.910 32.260 ;
        RECT 102.650 32.200 102.970 32.260 ;
        RECT 97.145 32.060 102.970 32.200 ;
        RECT 97.145 32.015 97.435 32.060 ;
        RECT 97.590 32.000 97.910 32.060 ;
        RECT 102.650 32.000 102.970 32.060 ;
        RECT 68.625 31.675 68.915 31.905 ;
        RECT 70.905 31.860 71.555 31.905 ;
        RECT 71.830 31.860 72.150 31.920 ;
        RECT 74.505 31.860 74.795 31.905 ;
        RECT 70.905 31.720 74.795 31.860 ;
        RECT 70.905 31.675 71.555 31.720 ;
        RECT 71.830 31.660 72.150 31.720 ;
        RECT 74.205 31.675 74.795 31.720 ;
        RECT 75.050 31.860 75.370 31.920 ;
        RECT 77.365 31.860 77.655 31.905 ;
        RECT 75.050 31.720 77.655 31.860 ;
        RECT 59.425 31.380 61.480 31.520 ;
        RECT 62.185 31.520 62.475 31.565 ;
        RECT 62.630 31.520 62.950 31.580 ;
        RECT 62.185 31.380 62.950 31.520 ;
        RECT 59.425 31.335 59.715 31.380 ;
        RECT 62.185 31.335 62.475 31.380 ;
        RECT 62.630 31.320 62.950 31.380 ;
        RECT 65.865 31.520 66.155 31.565 ;
        RECT 67.320 31.520 67.460 31.660 ;
        RECT 65.865 31.380 67.460 31.520 ;
        RECT 67.710 31.520 68.000 31.565 ;
        RECT 69.545 31.520 69.835 31.565 ;
        RECT 73.125 31.520 73.415 31.565 ;
        RECT 67.710 31.380 73.415 31.520 ;
        RECT 65.865 31.335 66.155 31.380 ;
        RECT 67.710 31.335 68.000 31.380 ;
        RECT 69.545 31.335 69.835 31.380 ;
        RECT 73.125 31.335 73.415 31.380 ;
        RECT 74.205 31.360 74.495 31.675 ;
        RECT 75.050 31.660 75.370 31.720 ;
        RECT 77.365 31.675 77.655 31.720 ;
        RECT 85.185 31.860 85.475 31.905 ;
        RECT 86.090 31.860 86.410 31.920 ;
        RECT 88.390 31.860 88.710 31.920 ;
        RECT 85.185 31.720 88.710 31.860 ;
        RECT 85.185 31.675 85.475 31.720 ;
        RECT 86.090 31.660 86.410 31.720 ;
        RECT 88.390 31.660 88.710 31.720 ;
        RECT 96.685 31.860 96.975 31.905 ;
        RECT 98.510 31.860 98.830 31.920 ;
        RECT 96.685 31.720 98.830 31.860 ;
        RECT 96.685 31.675 96.975 31.720 ;
        RECT 98.510 31.660 98.830 31.720 ;
        RECT 80.585 31.335 80.875 31.565 ;
        RECT 81.505 31.520 81.795 31.565 ;
        RECT 82.870 31.520 83.190 31.580 ;
        RECT 87.485 31.520 87.775 31.565 ;
        RECT 81.505 31.380 87.775 31.520 ;
        RECT 81.505 31.335 81.795 31.380 ;
        RECT 8.810 31.180 9.130 31.240 ;
        RECT 9.285 31.180 9.575 31.225 ;
        RECT 8.810 31.040 9.960 31.180 ;
        RECT 8.810 30.980 9.130 31.040 ;
        RECT 9.285 30.995 9.575 31.040 ;
        RECT 9.820 30.500 9.960 31.040 ;
        RECT 18.485 30.995 18.775 31.225 ;
        RECT 10.155 30.840 10.445 30.885 ;
        RECT 12.045 30.840 12.335 30.885 ;
        RECT 15.165 30.840 15.455 30.885 ;
        RECT 18.560 30.840 18.700 30.995 ;
        RECT 19.850 30.980 20.170 31.240 ;
        RECT 27.670 31.180 27.990 31.240 ;
        RECT 34.110 31.180 34.430 31.240 ;
        RECT 27.670 31.040 34.430 31.180 ;
        RECT 27.670 30.980 27.990 31.040 ;
        RECT 34.110 30.980 34.430 31.040 ;
        RECT 35.045 31.180 35.335 31.225 ;
        RECT 47.450 31.180 47.770 31.240 ;
        RECT 35.045 31.040 47.770 31.180 ;
        RECT 35.045 30.995 35.335 31.040 ;
        RECT 47.450 30.980 47.770 31.040 ;
        RECT 59.870 30.980 60.190 31.240 ;
        RECT 67.245 30.995 67.535 31.225 ;
        RECT 80.660 31.180 80.800 31.335 ;
        RECT 82.870 31.320 83.190 31.380 ;
        RECT 87.485 31.335 87.775 31.380 ;
        RECT 88.850 31.320 89.170 31.580 ;
        RECT 86.565 31.180 86.855 31.225 ;
        RECT 93.450 31.180 93.770 31.240 ;
        RECT 97.605 31.180 97.895 31.225 ;
        RECT 80.660 31.040 83.560 31.180 ;
        RECT 10.155 30.700 15.455 30.840 ;
        RECT 10.155 30.655 10.445 30.700 ;
        RECT 12.045 30.655 12.335 30.700 ;
        RECT 15.165 30.655 15.455 30.700 ;
        RECT 15.800 30.700 18.700 30.840 ;
        RECT 15.800 30.500 15.940 30.700 ;
        RECT 9.820 30.360 15.940 30.500 ;
        RECT 18.560 30.500 18.700 30.700 ;
        RECT 19.355 30.840 19.645 30.885 ;
        RECT 21.245 30.840 21.535 30.885 ;
        RECT 24.365 30.840 24.655 30.885 ;
        RECT 19.355 30.700 24.655 30.840 ;
        RECT 19.355 30.655 19.645 30.700 ;
        RECT 21.245 30.655 21.535 30.700 ;
        RECT 24.365 30.655 24.655 30.700 ;
        RECT 26.750 30.840 27.070 30.900 ;
        RECT 28.145 30.840 28.435 30.885 ;
        RECT 26.750 30.700 28.435 30.840 ;
        RECT 26.750 30.640 27.070 30.700 ;
        RECT 28.145 30.655 28.435 30.700 ;
        RECT 39.190 30.840 39.480 30.885 ;
        RECT 41.050 30.840 41.340 30.885 ;
        RECT 43.830 30.840 44.120 30.885 ;
        RECT 39.190 30.700 44.120 30.840 ;
        RECT 39.190 30.655 39.480 30.700 ;
        RECT 41.050 30.655 41.340 30.700 ;
        RECT 43.830 30.655 44.120 30.700 ;
        RECT 23.530 30.500 23.850 30.560 ;
        RECT 25.370 30.500 25.690 30.560 ;
        RECT 18.560 30.360 25.690 30.500 ;
        RECT 23.530 30.300 23.850 30.360 ;
        RECT 25.370 30.300 25.690 30.360 ;
        RECT 52.970 30.500 53.290 30.560 ;
        RECT 58.045 30.500 58.335 30.545 ;
        RECT 52.970 30.360 58.335 30.500 ;
        RECT 67.320 30.500 67.460 30.995 ;
        RECT 83.420 30.885 83.560 31.040 ;
        RECT 86.565 31.040 97.895 31.180 ;
        RECT 86.565 30.995 86.855 31.040 ;
        RECT 93.450 30.980 93.770 31.040 ;
        RECT 97.605 30.995 97.895 31.040 ;
        RECT 68.115 30.840 68.405 30.885 ;
        RECT 70.005 30.840 70.295 30.885 ;
        RECT 73.125 30.840 73.415 30.885 ;
        RECT 68.115 30.700 73.415 30.840 ;
        RECT 68.115 30.655 68.405 30.700 ;
        RECT 70.005 30.655 70.295 30.700 ;
        RECT 73.125 30.655 73.415 30.700 ;
        RECT 83.345 30.655 83.635 30.885 ;
        RECT 76.890 30.500 77.210 30.560 ;
        RECT 67.320 30.360 77.210 30.500 ;
        RECT 52.970 30.300 53.290 30.360 ;
        RECT 58.045 30.315 58.335 30.360 ;
        RECT 76.890 30.300 77.210 30.360 ;
        RECT 78.270 30.500 78.590 30.560 ;
        RECT 79.665 30.500 79.955 30.545 ;
        RECT 78.270 30.360 79.955 30.500 ;
        RECT 78.270 30.300 78.590 30.360 ;
        RECT 79.665 30.315 79.955 30.360 ;
        RECT 81.950 30.300 82.270 30.560 ;
        RECT 87.930 30.300 88.250 30.560 ;
        RECT 89.785 30.500 90.075 30.545 ;
        RECT 93.450 30.500 93.770 30.560 ;
        RECT 89.785 30.360 93.770 30.500 ;
        RECT 89.785 30.315 90.075 30.360 ;
        RECT 93.450 30.300 93.770 30.360 ;
        RECT 5.520 29.680 123.740 30.160 ;
        RECT 17.090 29.280 17.410 29.540 ;
        RECT 19.850 29.480 20.170 29.540 ;
        RECT 21.245 29.480 21.535 29.525 ;
        RECT 19.850 29.340 21.535 29.480 ;
        RECT 19.850 29.280 20.170 29.340 ;
        RECT 21.245 29.295 21.535 29.340 ;
        RECT 24.005 29.480 24.295 29.525 ;
        RECT 24.910 29.480 25.230 29.540 ;
        RECT 24.005 29.340 25.230 29.480 ;
        RECT 24.005 29.295 24.295 29.340 ;
        RECT 24.910 29.280 25.230 29.340 ;
        RECT 34.110 29.280 34.430 29.540 ;
        RECT 43.310 29.280 43.630 29.540 ;
        RECT 60.345 29.480 60.635 29.525 ;
        RECT 62.630 29.480 62.950 29.540 ;
        RECT 60.345 29.340 62.950 29.480 ;
        RECT 60.345 29.295 60.635 29.340 ;
        RECT 62.630 29.280 62.950 29.340 ;
        RECT 71.385 29.480 71.675 29.525 ;
        RECT 71.830 29.480 72.150 29.540 ;
        RECT 71.385 29.340 72.150 29.480 ;
        RECT 71.385 29.295 71.675 29.340 ;
        RECT 71.830 29.280 72.150 29.340 ;
        RECT 85.630 29.280 85.950 29.540 ;
        RECT 86.090 29.280 86.410 29.540 ;
        RECT 26.255 29.140 26.545 29.185 ;
        RECT 28.145 29.140 28.435 29.185 ;
        RECT 31.265 29.140 31.555 29.185 ;
        RECT 26.255 29.000 31.555 29.140 ;
        RECT 26.255 28.955 26.545 29.000 ;
        RECT 28.145 28.955 28.435 29.000 ;
        RECT 31.265 28.955 31.555 29.000 ;
        RECT 44.705 28.955 44.995 29.185 ;
        RECT 52.475 29.140 52.765 29.185 ;
        RECT 54.365 29.140 54.655 29.185 ;
        RECT 57.485 29.140 57.775 29.185 ;
        RECT 52.475 29.000 57.775 29.140 ;
        RECT 52.475 28.955 52.765 29.000 ;
        RECT 54.365 28.955 54.655 29.000 ;
        RECT 57.485 28.955 57.775 29.000 ;
        RECT 77.775 29.140 78.065 29.185 ;
        RECT 79.665 29.140 79.955 29.185 ;
        RECT 82.785 29.140 83.075 29.185 ;
        RECT 77.775 29.000 83.075 29.140 ;
        RECT 77.775 28.955 78.065 29.000 ;
        RECT 79.665 28.955 79.955 29.000 ;
        RECT 82.785 28.955 83.075 29.000 ;
        RECT 88.965 29.140 89.255 29.185 ;
        RECT 92.085 29.140 92.375 29.185 ;
        RECT 93.975 29.140 94.265 29.185 ;
        RECT 88.965 29.000 94.265 29.140 ;
        RECT 88.965 28.955 89.255 29.000 ;
        RECT 92.085 28.955 92.375 29.000 ;
        RECT 93.975 28.955 94.265 29.000 ;
        RECT 25.370 28.600 25.690 28.860 ;
        RECT 26.750 28.600 27.070 28.860 ;
        RECT 44.780 28.800 44.920 28.955 ;
        RECT 41.560 28.660 44.920 28.800 ;
        RECT 17.565 28.275 17.855 28.505 ;
        RECT 22.165 28.460 22.455 28.505 ;
        RECT 23.070 28.460 23.390 28.520 ;
        RECT 41.560 28.505 41.700 28.660 ;
        RECT 46.990 28.600 47.310 28.860 ;
        RECT 47.450 28.600 47.770 28.860 ;
        RECT 48.370 28.800 48.690 28.860 ;
        RECT 51.605 28.800 51.895 28.845 ;
        RECT 48.370 28.660 51.895 28.800 ;
        RECT 48.370 28.600 48.690 28.660 ;
        RECT 51.605 28.615 51.895 28.660 ;
        RECT 52.970 28.600 53.290 28.860 ;
        RECT 75.510 28.800 75.830 28.860 ;
        RECT 76.890 28.800 77.210 28.860 ;
        RECT 75.510 28.660 77.210 28.800 ;
        RECT 75.510 28.600 75.830 28.660 ;
        RECT 76.890 28.600 77.210 28.660 ;
        RECT 78.270 28.600 78.590 28.860 ;
        RECT 93.450 28.600 93.770 28.860 ;
        RECT 94.845 28.800 95.135 28.845 ;
        RECT 96.670 28.800 96.990 28.860 ;
        RECT 94.845 28.660 96.990 28.800 ;
        RECT 94.845 28.615 95.135 28.660 ;
        RECT 96.670 28.600 96.990 28.660 ;
        RECT 22.165 28.320 23.390 28.460 ;
        RECT 22.165 28.275 22.455 28.320 ;
        RECT 17.640 28.120 17.780 28.275 ;
        RECT 23.070 28.260 23.390 28.320 ;
        RECT 23.545 28.275 23.835 28.505 ;
        RECT 25.850 28.460 26.140 28.505 ;
        RECT 27.685 28.460 27.975 28.505 ;
        RECT 31.265 28.460 31.555 28.505 ;
        RECT 25.850 28.320 31.555 28.460 ;
        RECT 25.850 28.275 26.140 28.320 ;
        RECT 27.685 28.275 27.975 28.320 ;
        RECT 31.265 28.275 31.555 28.320 ;
        RECT 18.930 28.120 19.250 28.180 ;
        RECT 23.620 28.120 23.760 28.275 ;
        RECT 32.345 28.165 32.635 28.480 ;
        RECT 35.505 28.460 35.795 28.505 ;
        RECT 35.505 28.320 41.240 28.460 ;
        RECT 35.505 28.275 35.795 28.320 ;
        RECT 17.640 27.980 23.760 28.120 ;
        RECT 18.930 27.920 19.250 27.980 ;
        RECT 23.620 27.780 23.760 27.980 ;
        RECT 29.045 28.120 29.695 28.165 ;
        RECT 32.345 28.120 32.935 28.165 ;
        RECT 35.045 28.120 35.335 28.165 ;
        RECT 29.045 27.980 35.335 28.120 ;
        RECT 29.045 27.935 29.695 27.980 ;
        RECT 32.645 27.935 32.935 27.980 ;
        RECT 35.045 27.935 35.335 27.980 ;
        RECT 35.580 27.780 35.720 28.275 ;
        RECT 23.620 27.640 35.720 27.780 ;
        RECT 40.550 27.580 40.870 27.840 ;
        RECT 41.100 27.780 41.240 28.320 ;
        RECT 41.485 28.275 41.775 28.505 ;
        RECT 42.390 28.460 42.710 28.520 ;
        RECT 42.865 28.460 43.155 28.505 ;
        RECT 42.390 28.320 43.155 28.460 ;
        RECT 42.390 28.260 42.710 28.320 ;
        RECT 42.865 28.275 43.155 28.320 ;
        RECT 46.545 28.460 46.835 28.505 ;
        RECT 48.830 28.460 49.150 28.520 ;
        RECT 46.545 28.320 49.150 28.460 ;
        RECT 46.545 28.275 46.835 28.320 ;
        RECT 48.830 28.260 49.150 28.320 ;
        RECT 52.070 28.460 52.360 28.505 ;
        RECT 53.905 28.460 54.195 28.505 ;
        RECT 57.485 28.460 57.775 28.505 ;
        RECT 52.070 28.320 57.775 28.460 ;
        RECT 52.070 28.275 52.360 28.320 ;
        RECT 53.905 28.275 54.195 28.320 ;
        RECT 57.485 28.275 57.775 28.320 ;
        RECT 55.265 28.120 55.915 28.165 ;
        RECT 56.650 28.120 56.970 28.180 ;
        RECT 58.565 28.165 58.855 28.480 ;
        RECT 59.410 28.460 59.730 28.520 ;
        RECT 69.070 28.460 69.390 28.520 ;
        RECT 70.925 28.460 71.215 28.505 ;
        RECT 59.410 28.320 71.215 28.460 ;
        RECT 59.410 28.260 59.730 28.320 ;
        RECT 69.070 28.260 69.390 28.320 ;
        RECT 70.925 28.275 71.215 28.320 ;
        RECT 77.370 28.460 77.660 28.505 ;
        RECT 79.205 28.460 79.495 28.505 ;
        RECT 82.785 28.460 83.075 28.505 ;
        RECT 87.930 28.480 88.250 28.520 ;
        RECT 77.370 28.320 83.075 28.460 ;
        RECT 77.370 28.275 77.660 28.320 ;
        RECT 79.205 28.275 79.495 28.320 ;
        RECT 82.785 28.275 83.075 28.320 ;
        RECT 58.565 28.120 59.155 28.165 ;
        RECT 55.265 27.980 59.155 28.120 ;
        RECT 55.265 27.935 55.915 27.980 ;
        RECT 56.650 27.920 56.970 27.980 ;
        RECT 58.865 27.935 59.155 27.980 ;
        RECT 80.565 28.120 81.215 28.165 ;
        RECT 81.950 28.120 82.270 28.180 ;
        RECT 83.865 28.165 84.155 28.480 ;
        RECT 87.885 28.260 88.250 28.480 ;
        RECT 88.965 28.460 89.255 28.505 ;
        RECT 92.545 28.460 92.835 28.505 ;
        RECT 94.380 28.460 94.670 28.505 ;
        RECT 88.965 28.320 94.670 28.460 ;
        RECT 88.965 28.275 89.255 28.320 ;
        RECT 92.545 28.275 92.835 28.320 ;
        RECT 94.380 28.275 94.670 28.320 ;
        RECT 87.885 28.165 88.175 28.260 ;
        RECT 83.865 28.120 84.455 28.165 ;
        RECT 80.565 27.980 84.455 28.120 ;
        RECT 80.565 27.935 81.215 27.980 ;
        RECT 81.950 27.920 82.270 27.980 ;
        RECT 84.165 27.935 84.455 27.980 ;
        RECT 87.585 28.120 88.175 28.165 ;
        RECT 90.825 28.120 91.475 28.165 ;
        RECT 87.585 27.980 91.475 28.120 ;
        RECT 87.585 27.935 87.875 27.980 ;
        RECT 90.825 27.935 91.475 27.980 ;
        RECT 57.110 27.780 57.430 27.840 ;
        RECT 41.100 27.640 57.430 27.780 ;
        RECT 57.110 27.580 57.430 27.640 ;
        RECT 5.520 26.960 123.740 27.440 ;
        RECT 46.990 26.805 47.310 26.820 ;
        RECT 46.990 26.575 47.525 26.805 ;
        RECT 56.205 26.760 56.495 26.805 ;
        RECT 56.650 26.760 56.970 26.820 ;
        RECT 69.530 26.760 69.850 26.820 ;
        RECT 56.205 26.620 56.970 26.760 ;
        RECT 56.205 26.575 56.495 26.620 ;
        RECT 46.990 26.560 47.310 26.575 ;
        RECT 56.650 26.560 56.970 26.620 ;
        RECT 64.560 26.620 69.850 26.760 ;
        RECT 45.150 26.465 45.470 26.480 ;
        RECT 39.190 26.420 39.480 26.465 ;
        RECT 41.050 26.420 41.340 26.465 ;
        RECT 39.190 26.280 41.340 26.420 ;
        RECT 39.190 26.235 39.480 26.280 ;
        RECT 41.050 26.235 41.340 26.280 ;
        RECT 41.970 26.420 42.260 26.465 ;
        RECT 45.150 26.420 45.520 26.465 ;
        RECT 41.970 26.280 45.520 26.420 ;
        RECT 41.970 26.235 42.260 26.280 ;
        RECT 45.150 26.235 45.520 26.280 ;
        RECT 37.790 26.080 38.110 26.140 ;
        RECT 38.265 26.080 38.555 26.125 ;
        RECT 37.790 25.940 38.555 26.080 ;
        RECT 37.790 25.880 38.110 25.940 ;
        RECT 38.265 25.895 38.555 25.940 ;
        RECT 40.105 26.080 40.395 26.125 ;
        RECT 40.550 26.080 40.870 26.140 ;
        RECT 40.105 25.940 40.870 26.080 ;
        RECT 41.125 26.080 41.340 26.235 ;
        RECT 45.150 26.220 45.470 26.235 ;
        RECT 43.370 26.080 43.660 26.125 ;
        RECT 41.125 25.940 43.660 26.080 ;
        RECT 40.105 25.895 40.395 25.940 ;
        RECT 40.550 25.880 40.870 25.940 ;
        RECT 43.370 25.895 43.660 25.940 ;
        RECT 55.745 26.080 56.035 26.125 ;
        RECT 57.110 26.080 57.430 26.140 ;
        RECT 59.410 26.080 59.730 26.140 ;
        RECT 55.745 25.940 59.730 26.080 ;
        RECT 55.745 25.895 56.035 25.940 ;
        RECT 57.110 25.880 57.430 25.940 ;
        RECT 59.410 25.880 59.730 25.940 ;
        RECT 64.025 25.895 64.315 26.125 ;
        RECT 38.730 25.400 39.020 25.445 ;
        RECT 40.590 25.400 40.880 25.445 ;
        RECT 43.370 25.400 43.660 25.445 ;
        RECT 38.730 25.260 43.660 25.400 ;
        RECT 38.730 25.215 39.020 25.260 ;
        RECT 40.590 25.215 40.880 25.260 ;
        RECT 43.370 25.215 43.660 25.260 ;
        RECT 64.100 25.060 64.240 25.895 ;
        RECT 64.560 25.785 64.700 26.620 ;
        RECT 69.530 26.560 69.850 26.620 ;
        RECT 71.830 26.465 72.150 26.480 ;
        RECT 68.265 26.420 68.555 26.465 ;
        RECT 71.505 26.420 72.155 26.465 ;
        RECT 68.265 26.280 72.155 26.420 ;
        RECT 68.265 26.235 68.855 26.280 ;
        RECT 71.505 26.235 72.155 26.280 ;
        RECT 68.565 25.920 68.855 26.235 ;
        RECT 71.830 26.220 72.150 26.235 ;
        RECT 69.645 26.080 69.935 26.125 ;
        RECT 73.225 26.080 73.515 26.125 ;
        RECT 75.060 26.080 75.350 26.125 ;
        RECT 69.645 25.940 75.350 26.080 ;
        RECT 69.645 25.895 69.935 25.940 ;
        RECT 73.225 25.895 73.515 25.940 ;
        RECT 75.060 25.895 75.350 25.940 ;
        RECT 75.510 25.880 75.830 26.140 ;
        RECT 64.485 25.555 64.775 25.785 ;
        RECT 74.145 25.740 74.435 25.785 ;
        RECT 65.940 25.600 74.435 25.740 ;
        RECT 65.940 25.445 66.080 25.600 ;
        RECT 74.145 25.555 74.435 25.600 ;
        RECT 65.865 25.215 66.155 25.445 ;
        RECT 66.785 25.400 67.075 25.445 ;
        RECT 68.150 25.400 68.470 25.460 ;
        RECT 66.785 25.260 68.470 25.400 ;
        RECT 66.785 25.215 67.075 25.260 ;
        RECT 66.860 25.060 67.000 25.215 ;
        RECT 68.150 25.200 68.470 25.260 ;
        RECT 69.645 25.400 69.935 25.445 ;
        RECT 72.765 25.400 73.055 25.445 ;
        RECT 74.655 25.400 74.945 25.445 ;
        RECT 69.645 25.260 74.945 25.400 ;
        RECT 69.645 25.215 69.935 25.260 ;
        RECT 72.765 25.215 73.055 25.260 ;
        RECT 74.655 25.215 74.945 25.260 ;
        RECT 64.100 24.920 67.000 25.060 ;
        RECT 5.520 24.240 123.740 24.720 ;
        RECT 70.925 24.040 71.215 24.085 ;
        RECT 71.830 24.040 72.150 24.100 ;
        RECT 70.925 23.900 72.150 24.040 ;
        RECT 70.925 23.855 71.215 23.900 ;
        RECT 71.830 23.840 72.150 23.900 ;
        RECT 69.070 23.020 69.390 23.080 ;
        RECT 70.465 23.020 70.755 23.065 ;
        RECT 69.070 22.880 70.755 23.020 ;
        RECT 69.070 22.820 69.390 22.880 ;
        RECT 70.465 22.835 70.755 22.880 ;
        RECT 5.520 21.520 123.740 22.000 ;
        RECT 5.520 18.800 123.740 19.280 ;
        RECT 5.520 16.080 123.740 16.560 ;
        RECT 5.520 13.360 123.740 13.840 ;
        RECT 5.520 10.640 123.740 11.120 ;
      LAYER met2 ;
        RECT 10.030 138.990 11.800 139.130 ;
        RECT 3.380 118.310 3.520 138.395 ;
        RECT 9.580 127.655 11.460 128.025 ;
        RECT 3.780 123.770 4.040 124.090 ;
        RECT 3.840 120.205 3.980 123.770 ;
        RECT 9.580 122.215 11.460 122.585 ;
        RECT 11.660 122.050 11.800 138.990 ;
        RECT 21.320 138.990 22.630 139.130 ;
        RECT 35.790 138.990 36.180 139.130 ;
        RECT 16.260 123.750 16.400 138.395 ;
        RECT 17.580 124.110 17.840 124.430 ;
        RECT 16.200 123.430 16.460 123.750 ;
        RECT 17.640 122.050 17.780 124.110 ;
        RECT 19.880 123.430 20.140 123.750 ;
        RECT 18.960 122.750 19.220 123.070 ;
        RECT 11.600 121.730 11.860 122.050 ;
        RECT 17.580 121.730 17.840 122.050 ;
        RECT 19.020 121.710 19.160 122.750 ;
        RECT 18.960 121.390 19.220 121.710 ;
        RECT 18.040 120.710 18.300 121.030 ;
        RECT 7.920 120.370 8.180 120.690 ;
        RECT 8.380 120.370 8.640 120.690 ;
        RECT 3.770 119.835 4.050 120.205 ;
        RECT 3.320 117.990 3.580 118.310 ;
        RECT 7.980 117.630 8.120 120.370 ;
        RECT 7.920 117.310 8.180 117.630 ;
        RECT 7.980 112.870 8.120 117.310 ;
        RECT 8.440 116.610 8.580 120.370 ;
        RECT 18.100 118.650 18.240 120.710 ;
        RECT 18.040 118.330 18.300 118.650 ;
        RECT 19.420 118.330 19.680 118.650 ;
        RECT 15.280 117.990 15.540 118.310 ;
        RECT 9.580 116.775 11.460 117.145 ;
        RECT 15.340 116.610 15.480 117.990 ;
        RECT 8.380 116.290 8.640 116.610 ;
        RECT 15.280 116.290 15.540 116.610 ;
        RECT 12.060 115.270 12.320 115.590 ;
        RECT 12.520 115.270 12.780 115.590 ;
        RECT 7.920 112.550 8.180 112.870 ;
        RECT 7.980 101.990 8.120 112.550 ;
        RECT 9.580 111.335 11.460 111.705 ;
        RECT 9.580 105.895 11.460 106.265 ;
        RECT 11.600 103.710 11.860 104.030 ;
        RECT 7.920 101.670 8.180 101.990 ;
        RECT 7.980 99.270 8.120 101.670 ;
        RECT 9.580 100.455 11.460 100.825 ;
        RECT 11.660 99.610 11.800 103.710 ;
        RECT 11.600 99.290 11.860 99.610 ;
        RECT 7.920 98.950 8.180 99.270 ;
        RECT 7.980 88.390 8.120 98.950 ;
        RECT 9.580 95.015 11.460 95.385 ;
        RECT 11.600 90.110 11.860 90.430 ;
        RECT 9.580 89.575 11.460 89.945 ;
        RECT 11.660 88.730 11.800 90.110 ;
        RECT 11.600 88.410 11.860 88.730 ;
        RECT 7.920 88.070 8.180 88.390 ;
        RECT 7.980 86.010 8.120 88.070 ;
        RECT 7.920 85.690 8.180 86.010 ;
        RECT 11.600 85.350 11.860 85.670 ;
        RECT 9.580 84.135 11.460 84.505 ;
        RECT 11.660 83.970 11.800 85.350 ;
        RECT 11.600 83.650 11.860 83.970 ;
        RECT 9.580 78.695 11.460 79.065 ;
        RECT 12.120 78.530 12.260 115.270 ;
        RECT 12.060 78.210 12.320 78.530 ;
        RECT 12.580 78.190 12.720 115.270 ;
        RECT 16.200 113.230 16.460 113.550 ;
        RECT 14.360 112.550 14.620 112.870 ;
        RECT 14.420 111.170 14.560 112.550 ;
        RECT 14.360 110.850 14.620 111.170 ;
        RECT 16.260 110.490 16.400 113.230 ;
        RECT 16.200 110.170 16.460 110.490 ;
        RECT 16.660 109.830 16.920 110.150 ;
        RECT 16.720 104.710 16.860 109.830 ;
        RECT 18.960 107.450 19.220 107.770 ;
        RECT 19.020 105.730 19.160 107.450 ;
        RECT 18.960 105.410 19.220 105.730 ;
        RECT 18.960 104.730 19.220 105.050 ;
        RECT 16.660 104.390 16.920 104.710 ;
        RECT 18.040 104.050 18.300 104.370 ;
        RECT 13.900 103.710 14.160 104.030 ;
        RECT 14.360 103.710 14.620 104.030 ;
        RECT 16.200 103.710 16.460 104.030 ;
        RECT 13.960 102.670 14.100 103.710 ;
        RECT 13.900 102.350 14.160 102.670 ;
        RECT 14.420 101.310 14.560 103.710 ;
        RECT 16.260 101.650 16.400 103.710 ;
        RECT 18.100 103.010 18.240 104.050 ;
        RECT 18.040 102.690 18.300 103.010 ;
        RECT 19.020 101.990 19.160 104.730 ;
        RECT 18.960 101.670 19.220 101.990 ;
        RECT 16.200 101.330 16.460 101.650 ;
        RECT 14.360 100.990 14.620 101.310 ;
        RECT 18.500 100.990 18.760 101.310 ;
        RECT 18.560 98.930 18.700 100.990 ;
        RECT 18.500 98.610 18.760 98.930 ;
        RECT 16.200 91.130 16.460 91.450 ;
        RECT 14.820 87.730 15.080 88.050 ;
        RECT 13.440 86.030 13.700 86.350 ;
        RECT 13.500 82.950 13.640 86.030 ;
        RECT 14.880 82.950 15.020 87.730 ;
        RECT 16.260 85.670 16.400 91.130 ;
        RECT 16.660 90.790 16.920 91.110 ;
        RECT 16.720 89.410 16.860 90.790 ;
        RECT 16.660 89.090 16.920 89.410 ;
        RECT 16.720 86.350 16.860 89.090 ;
        RECT 16.660 86.030 16.920 86.350 ;
        RECT 18.960 85.690 19.220 86.010 ;
        RECT 16.200 85.350 16.460 85.670 ;
        RECT 17.580 84.670 17.840 84.990 ;
        RECT 13.440 82.630 13.700 82.950 ;
        RECT 13.900 82.630 14.160 82.950 ;
        RECT 14.820 82.630 15.080 82.950 ;
        RECT 12.520 77.870 12.780 78.190 ;
        RECT 11.140 76.510 11.400 76.830 ;
        RECT 11.200 75.130 11.340 76.510 ;
        RECT 13.960 75.130 14.100 82.630 ;
        RECT 17.640 82.610 17.780 84.670 ;
        RECT 17.580 82.290 17.840 82.610 ;
        RECT 19.020 79.890 19.160 85.690 ;
        RECT 19.480 81.250 19.620 118.330 ;
        RECT 19.940 117.970 20.080 123.430 ;
        RECT 20.800 122.980 21.060 123.070 ;
        RECT 20.400 122.840 21.060 122.980 ;
        RECT 20.400 121.370 20.540 122.840 ;
        RECT 20.800 122.750 21.060 122.840 ;
        RECT 20.340 121.050 20.600 121.370 ;
        RECT 19.880 117.650 20.140 117.970 ;
        RECT 20.400 117.630 20.540 121.050 ;
        RECT 21.320 118.310 21.460 138.990 ;
        RECT 24.580 124.935 26.460 125.305 ;
        RECT 21.720 123.770 21.980 124.090 ;
        RECT 21.780 121.030 21.920 123.770 ;
        RECT 26.780 122.750 27.040 123.070 ;
        RECT 21.720 120.710 21.980 121.030 ;
        RECT 24.580 119.495 26.460 119.865 ;
        RECT 26.840 118.990 26.980 122.750 ;
        RECT 29.140 122.050 29.280 138.395 ;
        RECT 33.680 123.770 33.940 124.090 ;
        RECT 29.540 122.750 29.800 123.070 ;
        RECT 29.080 121.730 29.340 122.050 ;
        RECT 29.600 120.690 29.740 122.750 ;
        RECT 33.740 121.030 33.880 123.770 ;
        RECT 33.680 120.710 33.940 121.030 ;
        RECT 29.540 120.370 29.800 120.690 ;
        RECT 30.000 120.030 30.260 120.350 ;
        RECT 35.520 120.030 35.780 120.350 ;
        RECT 30.060 119.330 30.200 120.030 ;
        RECT 30.000 119.010 30.260 119.330 ;
        RECT 35.580 118.990 35.720 120.030 ;
        RECT 26.780 118.670 27.040 118.990 ;
        RECT 35.520 118.670 35.780 118.990 ;
        RECT 30.920 118.330 31.180 118.650 ;
        RECT 21.260 117.990 21.520 118.310 ;
        RECT 28.160 117.990 28.420 118.310 ;
        RECT 20.340 117.310 20.600 117.630 ;
        RECT 20.400 109.810 20.540 117.310 ;
        RECT 28.220 116.610 28.360 117.990 ;
        RECT 28.160 116.290 28.420 116.610 ;
        RECT 26.780 115.270 27.040 115.590 ;
        RECT 24.580 114.055 26.460 114.425 ;
        RECT 20.800 111.870 21.060 112.190 ;
        RECT 20.340 109.490 20.600 109.810 ;
        RECT 20.400 107.430 20.540 109.490 ;
        RECT 20.860 109.470 21.000 111.870 ;
        RECT 22.180 110.170 22.440 110.490 ;
        RECT 20.800 109.150 21.060 109.470 ;
        RECT 21.260 109.150 21.520 109.470 ;
        RECT 20.340 107.110 20.600 107.430 ;
        RECT 19.880 103.710 20.140 104.030 ;
        RECT 19.940 102.330 20.080 103.710 ;
        RECT 19.880 102.010 20.140 102.330 ;
        RECT 19.940 100.290 20.080 102.010 ;
        RECT 19.880 99.970 20.140 100.290 ;
        RECT 19.940 96.550 20.080 99.970 ;
        RECT 19.880 96.230 20.140 96.550 ;
        RECT 20.400 94.170 20.540 107.110 ;
        RECT 20.860 102.670 21.000 109.150 ;
        RECT 20.800 102.350 21.060 102.670 ;
        RECT 21.320 101.990 21.460 109.150 ;
        RECT 22.240 105.050 22.380 110.170 ;
        RECT 24.020 109.150 24.280 109.470 ;
        RECT 24.080 108.110 24.220 109.150 ;
        RECT 24.580 108.615 26.460 108.985 ;
        RECT 24.020 107.790 24.280 108.110 ;
        RECT 22.180 104.730 22.440 105.050 ;
        RECT 21.720 104.390 21.980 104.710 ;
        RECT 21.780 102.330 21.920 104.390 ;
        RECT 25.390 104.195 25.670 104.565 ;
        RECT 25.400 104.050 25.660 104.195 ;
        RECT 23.560 103.710 23.820 104.030 ;
        RECT 21.720 102.010 21.980 102.330 ;
        RECT 21.260 101.670 21.520 101.990 ;
        RECT 23.620 101.650 23.760 103.710 ;
        RECT 24.580 103.175 26.460 103.545 ;
        RECT 26.320 102.350 26.580 102.670 ;
        RECT 23.560 101.330 23.820 101.650 ;
        RECT 23.620 99.950 23.760 101.330 ;
        RECT 23.560 99.630 23.820 99.950 ;
        RECT 26.380 99.270 26.520 102.350 ;
        RECT 22.180 98.950 22.440 99.270 ;
        RECT 26.320 98.950 26.580 99.270 ;
        RECT 21.720 98.610 21.980 98.930 ;
        RECT 20.800 96.570 21.060 96.890 ;
        RECT 20.340 93.850 20.600 94.170 ;
        RECT 20.340 90.790 20.600 91.110 ;
        RECT 20.400 85.670 20.540 90.790 ;
        RECT 19.880 85.350 20.140 85.670 ;
        RECT 20.340 85.350 20.600 85.670 ;
        RECT 19.940 82.610 20.080 85.350 ;
        RECT 19.880 82.290 20.140 82.610 ;
        RECT 19.420 80.930 19.680 81.250 ;
        RECT 15.740 79.570 16.000 79.890 ;
        RECT 18.960 79.570 19.220 79.890 ;
        RECT 15.800 76.830 15.940 79.570 ;
        RECT 19.880 77.250 20.140 77.510 ;
        RECT 20.400 77.250 20.540 85.350 ;
        RECT 20.860 79.550 21.000 96.570 ;
        RECT 21.260 79.910 21.520 80.230 ;
        RECT 20.800 79.230 21.060 79.550 ;
        RECT 21.320 77.760 21.460 79.910 ;
        RECT 21.780 78.530 21.920 98.610 ;
        RECT 22.240 96.890 22.380 98.950 ;
        RECT 24.020 98.270 24.280 98.590 ;
        RECT 22.180 96.570 22.440 96.890 ;
        RECT 23.100 96.570 23.360 96.890 ;
        RECT 23.160 92.130 23.300 96.570 ;
        RECT 23.560 95.550 23.820 95.870 ;
        RECT 23.620 93.830 23.760 95.550 ;
        RECT 23.560 93.510 23.820 93.830 ;
        RECT 23.100 91.810 23.360 92.130 ;
        RECT 24.080 89.410 24.220 98.270 ;
        RECT 24.580 97.735 26.460 98.105 ;
        RECT 24.580 92.295 26.460 92.665 ;
        RECT 26.840 89.410 26.980 115.270 ;
        RECT 27.700 113.230 27.960 113.550 ;
        RECT 27.760 110.490 27.900 113.230 ;
        RECT 29.540 111.870 29.800 112.190 ;
        RECT 29.600 110.490 29.740 111.870 ;
        RECT 27.700 110.170 27.960 110.490 ;
        RECT 29.540 110.170 29.800 110.490 ;
        RECT 27.700 109.210 27.960 109.470 ;
        RECT 27.300 109.150 27.960 109.210 ;
        RECT 27.300 109.070 27.900 109.150 ;
        RECT 27.300 104.370 27.440 109.070 ;
        RECT 27.700 106.430 27.960 106.750 ;
        RECT 27.760 104.710 27.900 106.430 ;
        RECT 27.700 104.390 27.960 104.710 ;
        RECT 27.240 104.050 27.500 104.370 ;
        RECT 27.300 101.990 27.440 104.050 ;
        RECT 27.240 101.670 27.500 101.990 ;
        RECT 27.760 101.650 27.900 104.390 ;
        RECT 29.540 102.350 29.800 102.670 ;
        RECT 28.160 102.010 28.420 102.330 ;
        RECT 27.700 101.330 27.960 101.650 ;
        RECT 27.760 99.270 27.900 101.330 ;
        RECT 28.220 99.270 28.360 102.010 ;
        RECT 28.620 100.990 28.880 101.310 ;
        RECT 27.700 98.950 27.960 99.270 ;
        RECT 28.160 98.950 28.420 99.270 ;
        RECT 27.240 96.570 27.500 96.890 ;
        RECT 27.300 93.490 27.440 96.570 ;
        RECT 27.240 93.170 27.500 93.490 ;
        RECT 24.020 89.090 24.280 89.410 ;
        RECT 26.780 89.090 27.040 89.410 ;
        RECT 27.240 88.750 27.500 89.070 ;
        RECT 23.100 88.410 23.360 88.730 ;
        RECT 22.180 85.350 22.440 85.670 ;
        RECT 22.240 82.950 22.380 85.350 ;
        RECT 22.180 82.630 22.440 82.950 ;
        RECT 22.240 82.270 22.380 82.630 ;
        RECT 22.180 81.950 22.440 82.270 ;
        RECT 22.640 80.250 22.900 80.570 ;
        RECT 22.180 79.230 22.440 79.550 ;
        RECT 21.720 78.210 21.980 78.530 ;
        RECT 21.320 77.620 21.920 77.760 ;
        RECT 19.880 77.190 20.540 77.250 ;
        RECT 20.800 77.190 21.060 77.510 ;
        RECT 19.940 77.110 20.540 77.190 ;
        RECT 15.280 76.510 15.540 76.830 ;
        RECT 15.740 76.510 16.000 76.830 ;
        RECT 15.340 75.130 15.480 76.510 ;
        RECT 11.140 74.810 11.400 75.130 ;
        RECT 13.900 74.810 14.160 75.130 ;
        RECT 15.280 74.810 15.540 75.130 ;
        RECT 8.840 73.790 9.100 74.110 ;
        RECT 11.600 73.790 11.860 74.110 ;
        RECT 13.440 73.790 13.700 74.110 ;
        RECT 8.900 72.410 9.040 73.790 ;
        RECT 9.580 73.255 11.460 73.625 ;
        RECT 8.380 72.090 8.640 72.410 ;
        RECT 8.840 72.090 9.100 72.410 ;
        RECT 8.440 69.350 8.580 72.090 ;
        RECT 11.660 69.350 11.800 73.790 ;
        RECT 13.500 71.730 13.640 73.790 ;
        RECT 13.960 72.070 14.100 74.810 ;
        RECT 15.800 73.090 15.940 76.510 ;
        RECT 17.120 74.810 17.380 75.130 ;
        RECT 15.740 72.770 16.000 73.090 ;
        RECT 13.900 71.750 14.160 72.070 ;
        RECT 13.440 71.410 13.700 71.730 ;
        RECT 8.380 69.030 8.640 69.350 ;
        RECT 11.600 69.030 11.860 69.350 ;
        RECT 8.440 60.930 8.580 69.030 ;
        RECT 9.580 67.815 11.460 68.185 ;
        RECT 13.960 64.590 14.100 71.750 ;
        RECT 17.180 70.370 17.320 74.810 ;
        RECT 20.400 74.790 20.540 77.110 ;
        RECT 20.340 74.470 20.600 74.790 ;
        RECT 17.580 71.070 17.840 71.390 ;
        RECT 17.120 70.050 17.380 70.370 ;
        RECT 17.640 70.030 17.780 71.070 ;
        RECT 17.580 69.710 17.840 70.030 ;
        RECT 18.500 69.370 18.760 69.690 ;
        RECT 13.900 64.270 14.160 64.590 ;
        RECT 17.580 64.270 17.840 64.590 ;
        RECT 18.040 64.270 18.300 64.590 ;
        RECT 13.440 63.930 13.700 64.250 ;
        RECT 12.520 62.910 12.780 63.230 ;
        RECT 9.580 62.375 11.460 62.745 ;
        RECT 8.440 60.850 9.040 60.930 ;
        RECT 8.440 60.790 9.100 60.850 ;
        RECT 8.840 60.530 9.100 60.790 ;
        RECT 9.300 60.530 9.560 60.850 ;
        RECT 8.900 58.470 9.040 60.530 ;
        RECT 9.360 59.490 9.500 60.530 ;
        RECT 11.140 60.190 11.400 60.510 ;
        RECT 9.300 59.170 9.560 59.490 ;
        RECT 11.200 58.810 11.340 60.190 ;
        RECT 11.140 58.490 11.400 58.810 ;
        RECT 8.840 58.150 9.100 58.470 ;
        RECT 8.900 55.750 9.040 58.150 ;
        RECT 12.060 57.470 12.320 57.790 ;
        RECT 9.580 56.935 11.460 57.305 ;
        RECT 8.840 55.430 9.100 55.750 ;
        RECT 1.940 53.050 2.200 53.370 ;
        RECT 2.000 52.205 2.140 53.050 ;
        RECT 1.930 51.835 2.210 52.205 ;
        RECT 8.900 44.870 9.040 55.430 ;
        RECT 12.120 55.410 12.260 57.470 ;
        RECT 12.580 56.090 12.720 62.910 ;
        RECT 12.520 55.770 12.780 56.090 ;
        RECT 12.060 55.090 12.320 55.410 ;
        RECT 13.500 53.710 13.640 63.930 ;
        RECT 16.660 63.590 16.920 63.910 ;
        RECT 16.720 62.210 16.860 63.590 ;
        RECT 17.640 63.570 17.780 64.270 ;
        RECT 17.580 63.250 17.840 63.570 ;
        RECT 16.660 61.890 16.920 62.210 ;
        RECT 14.820 60.870 15.080 61.190 ;
        RECT 13.900 58.830 14.160 59.150 ;
        RECT 13.440 53.390 13.700 53.710 ;
        RECT 13.960 53.370 14.100 58.830 ;
        RECT 14.880 54.050 15.020 60.870 ;
        RECT 17.580 60.190 17.840 60.510 ;
        RECT 17.640 59.490 17.780 60.190 ;
        RECT 17.580 59.170 17.840 59.490 ;
        RECT 18.100 56.770 18.240 64.270 ;
        RECT 18.560 64.250 18.700 69.370 ;
        RECT 18.500 63.930 18.760 64.250 ;
        RECT 18.560 62.210 18.700 63.930 ;
        RECT 18.500 61.890 18.760 62.210 ;
        RECT 19.420 58.830 19.680 59.150 ;
        RECT 19.480 56.770 19.620 58.830 ;
        RECT 18.040 56.450 18.300 56.770 ;
        RECT 19.420 56.450 19.680 56.770 ;
        RECT 19.880 55.430 20.140 55.750 ;
        RECT 14.820 53.730 15.080 54.050 ;
        RECT 19.940 53.370 20.080 55.430 ;
        RECT 13.900 53.050 14.160 53.370 ;
        RECT 19.880 53.050 20.140 53.370 ;
        RECT 9.580 51.495 11.460 51.865 ;
        RECT 18.040 49.310 18.300 49.630 ;
        RECT 18.100 47.930 18.240 49.310 ;
        RECT 20.860 48.270 21.000 77.190 ;
        RECT 21.260 76.850 21.520 77.170 ;
        RECT 21.320 70.370 21.460 76.850 ;
        RECT 21.780 71.730 21.920 77.620 ;
        RECT 22.240 75.470 22.380 79.230 ;
        RECT 22.700 75.810 22.840 80.250 ;
        RECT 22.640 75.490 22.900 75.810 ;
        RECT 22.180 75.150 22.440 75.470 ;
        RECT 21.720 71.410 21.980 71.730 ;
        RECT 22.180 71.070 22.440 71.390 ;
        RECT 21.260 70.050 21.520 70.370 ;
        RECT 22.240 64.250 22.380 71.070 ;
        RECT 23.160 69.770 23.300 88.410 ;
        RECT 23.560 88.070 23.820 88.390 ;
        RECT 23.620 73.090 23.760 88.070 ;
        RECT 24.020 87.730 24.280 88.050 ;
        RECT 24.080 83.970 24.220 87.730 ;
        RECT 24.580 86.855 26.460 87.225 ;
        RECT 25.860 85.690 26.120 86.010 ;
        RECT 26.320 85.690 26.580 86.010 ;
        RECT 24.020 83.650 24.280 83.970 ;
        RECT 25.920 83.290 26.060 85.690 ;
        RECT 26.380 83.290 26.520 85.690 ;
        RECT 27.300 85.670 27.440 88.750 ;
        RECT 27.240 85.350 27.500 85.670 ;
        RECT 25.860 82.970 26.120 83.290 ;
        RECT 26.320 82.970 26.580 83.290 ;
        RECT 24.020 81.950 24.280 82.270 ;
        RECT 25.920 82.180 26.060 82.970 ;
        RECT 27.240 82.630 27.500 82.950 ;
        RECT 25.920 82.040 26.980 82.180 ;
        RECT 24.080 80.650 24.220 81.950 ;
        RECT 24.580 81.415 26.460 81.785 ;
        RECT 24.080 80.570 24.680 80.650 ;
        RECT 26.840 80.570 26.980 82.040 ;
        RECT 27.300 81.250 27.440 82.630 ;
        RECT 27.240 80.930 27.500 81.250 ;
        RECT 27.300 80.570 27.440 80.930 ;
        RECT 24.080 80.510 24.740 80.570 ;
        RECT 24.480 80.250 24.740 80.510 ;
        RECT 25.400 80.250 25.660 80.570 ;
        RECT 26.780 80.250 27.040 80.570 ;
        RECT 27.240 80.250 27.500 80.570 ;
        RECT 25.460 77.510 25.600 80.250 ;
        RECT 26.840 77.850 26.980 80.250 ;
        RECT 26.780 77.530 27.040 77.850 ;
        RECT 24.480 77.420 24.740 77.510 ;
        RECT 24.080 77.280 24.740 77.420 ;
        RECT 24.080 75.130 24.220 77.280 ;
        RECT 24.480 77.190 24.740 77.280 ;
        RECT 25.400 77.190 25.660 77.510 ;
        RECT 27.300 77.170 27.440 80.250 ;
        RECT 28.680 78.530 28.820 100.990 ;
        RECT 29.600 98.930 29.740 102.350 ;
        RECT 29.540 98.610 29.800 98.930 ;
        RECT 29.080 98.270 29.340 98.590 ;
        RECT 29.140 84.990 29.280 98.270 ;
        RECT 29.600 97.230 29.740 98.610 ;
        RECT 29.540 96.910 29.800 97.230 ;
        RECT 30.980 86.690 31.120 118.330 ;
        RECT 36.040 118.310 36.180 138.990 ;
        RECT 53.980 138.990 54.830 139.130 ;
        RECT 74.430 138.990 74.820 139.130 ;
        RECT 80.870 138.990 81.260 139.130 ;
        RECT 87.310 138.990 88.620 139.130 ;
        RECT 39.580 127.655 41.460 128.025 ;
        RECT 38.740 123.660 39.000 123.750 ;
        RECT 38.740 123.520 39.400 123.660 ;
        RECT 38.740 123.430 39.000 123.520 ;
        RECT 39.260 123.070 39.400 123.520 ;
        RECT 39.200 122.750 39.460 123.070 ;
        RECT 39.260 121.370 39.400 122.750 ;
        RECT 39.580 122.215 41.460 122.585 ;
        RECT 42.020 122.050 42.160 138.395 ;
        RECT 45.640 123.770 45.900 124.090 ;
        RECT 41.960 121.730 42.220 122.050 ;
        RECT 45.700 121.710 45.840 123.770 ;
        RECT 46.100 123.430 46.360 123.750 ;
        RECT 48.460 123.490 48.600 138.395 ;
        RECT 46.160 122.050 46.300 123.430 ;
        RECT 47.540 123.410 48.600 123.490 ;
        RECT 49.320 123.430 49.580 123.750 ;
        RECT 53.980 123.490 54.120 138.990 ;
        RECT 54.580 124.935 56.460 125.305 ;
        RECT 57.140 123.770 57.400 124.090 ;
        RECT 47.480 123.350 48.600 123.410 ;
        RECT 47.480 123.090 47.740 123.350 ;
        RECT 49.380 122.050 49.520 123.430 ;
        RECT 53.980 123.410 55.040 123.490 ;
        RECT 53.980 123.350 55.100 123.410 ;
        RECT 54.840 123.090 55.100 123.350 ;
        RECT 46.100 121.730 46.360 122.050 ;
        RECT 49.320 121.730 49.580 122.050 ;
        RECT 45.640 121.390 45.900 121.710 ;
        RECT 57.200 121.370 57.340 123.770 ;
        RECT 61.340 123.750 61.480 138.395 ;
        RECT 61.740 124.110 62.000 124.430 ;
        RECT 58.980 123.430 59.240 123.750 ;
        RECT 61.280 123.430 61.540 123.750 ;
        RECT 59.040 121.710 59.180 123.430 ;
        RECT 61.800 122.050 61.940 124.110 ;
        RECT 67.260 123.430 67.520 123.750 ;
        RECT 61.740 121.730 62.000 122.050 ;
        RECT 58.980 121.390 59.240 121.710 ;
        RECT 39.200 121.050 39.460 121.370 ;
        RECT 52.080 121.050 52.340 121.370 ;
        RECT 57.140 121.050 57.400 121.370 ;
        RECT 36.440 120.370 36.700 120.690 ;
        RECT 36.500 119.330 36.640 120.370 ;
        RECT 36.440 119.010 36.700 119.330 ;
        RECT 33.220 117.990 33.480 118.310 ;
        RECT 35.980 117.990 36.240 118.310 ;
        RECT 33.280 116.610 33.420 117.990 ;
        RECT 33.220 116.290 33.480 116.610 ;
        RECT 36.440 115.270 36.700 115.590 ;
        RECT 35.980 112.550 36.240 112.870 ;
        RECT 32.300 111.870 32.560 112.190 ;
        RECT 32.360 109.810 32.500 111.870 ;
        RECT 32.300 109.490 32.560 109.810 ;
        RECT 32.760 107.450 33.020 107.770 ;
        RECT 31.380 103.710 31.640 104.030 ;
        RECT 31.440 94.170 31.580 103.710 ;
        RECT 32.820 103.010 32.960 107.450 ;
        RECT 36.040 105.730 36.180 112.550 ;
        RECT 35.980 105.410 36.240 105.730 ;
        RECT 35.060 104.730 35.320 105.050 ;
        RECT 32.760 102.690 33.020 103.010 ;
        RECT 35.120 101.990 35.260 104.730 ;
        RECT 35.980 102.350 36.240 102.670 ;
        RECT 35.060 101.670 35.320 101.990 ;
        RECT 36.040 99.610 36.180 102.350 ;
        RECT 35.980 99.290 36.240 99.610 ;
        RECT 34.600 98.270 34.860 98.590 ;
        RECT 32.760 96.570 33.020 96.890 ;
        RECT 32.300 94.530 32.560 94.850 ;
        RECT 31.380 93.850 31.640 94.170 ;
        RECT 32.360 91.790 32.500 94.530 ;
        RECT 32.820 92.130 32.960 96.570 ;
        RECT 33.220 95.550 33.480 95.870 ;
        RECT 33.280 94.170 33.420 95.550 ;
        RECT 33.220 93.850 33.480 94.170 ;
        RECT 32.760 91.810 33.020 92.130 ;
        RECT 32.300 91.470 32.560 91.790 ;
        RECT 31.840 88.750 32.100 89.070 ;
        RECT 30.920 86.370 31.180 86.690 ;
        RECT 31.900 86.010 32.040 88.750 ;
        RECT 32.360 86.010 32.500 91.470 ;
        RECT 34.660 89.410 34.800 98.270 ;
        RECT 36.500 89.410 36.640 115.270 ;
        RECT 39.260 112.870 39.400 121.050 ;
        RECT 48.860 120.710 49.120 121.030 ;
        RECT 51.620 120.710 51.880 121.030 ;
        RECT 46.560 118.330 46.820 118.650 ;
        RECT 39.580 116.775 41.460 117.145 ;
        RECT 45.180 113.230 45.440 113.550 ;
        RECT 41.960 112.890 42.220 113.210 ;
        RECT 39.200 112.550 39.460 112.870 ;
        RECT 39.260 107.340 39.400 112.550 ;
        RECT 39.580 111.335 41.460 111.705 ;
        RECT 42.020 111.170 42.160 112.890 ;
        RECT 41.960 110.850 42.220 111.170 ;
        RECT 45.240 110.490 45.380 113.230 ;
        RECT 45.180 110.170 45.440 110.490 ;
        RECT 42.420 109.830 42.680 110.150 ;
        RECT 39.660 107.340 39.920 107.430 ;
        RECT 39.260 107.200 39.920 107.340 ;
        RECT 39.260 104.370 39.400 107.200 ;
        RECT 39.660 107.110 39.920 107.200 ;
        RECT 39.580 105.895 41.460 106.265 ;
        RECT 39.200 104.050 39.460 104.370 ;
        RECT 39.260 96.210 39.400 104.050 ;
        RECT 42.480 103.010 42.620 109.830 ;
        RECT 44.710 104.195 44.990 104.565 ;
        RECT 44.720 104.050 44.980 104.195 ;
        RECT 42.420 102.690 42.680 103.010 ;
        RECT 39.580 100.455 41.460 100.825 ;
        RECT 43.800 98.950 44.060 99.270 ;
        RECT 39.200 95.890 39.460 96.210 ;
        RECT 36.900 95.550 37.160 95.870 ;
        RECT 36.960 93.490 37.100 95.550 ;
        RECT 36.900 93.170 37.160 93.490 ;
        RECT 38.740 91.530 39.000 91.790 ;
        RECT 39.260 91.530 39.400 95.890 ;
        RECT 39.580 95.015 41.460 95.385 ;
        RECT 39.660 92.830 39.920 93.150 ;
        RECT 39.720 92.130 39.860 92.830 ;
        RECT 39.660 91.810 39.920 92.130 ;
        RECT 38.740 91.470 39.400 91.530 ;
        RECT 38.800 91.390 39.400 91.470 ;
        RECT 34.600 89.090 34.860 89.410 ;
        RECT 36.440 89.090 36.700 89.410 ;
        RECT 35.980 88.410 36.240 88.730 ;
        RECT 35.520 88.070 35.780 88.390 ;
        RECT 35.060 87.730 35.320 88.050 ;
        RECT 35.120 86.690 35.260 87.730 ;
        RECT 35.060 86.370 35.320 86.690 ;
        RECT 34.140 86.030 34.400 86.350 ;
        RECT 30.920 85.690 31.180 86.010 ;
        RECT 31.840 85.690 32.100 86.010 ;
        RECT 32.300 85.690 32.560 86.010 ;
        RECT 29.540 85.010 29.800 85.330 ;
        RECT 29.080 84.670 29.340 84.990 ;
        RECT 29.600 79.970 29.740 85.010 ;
        RECT 29.140 79.830 29.740 79.970 ;
        RECT 28.620 78.210 28.880 78.530 ;
        RECT 28.160 77.190 28.420 77.510 ;
        RECT 27.240 76.850 27.500 77.170 ;
        RECT 24.580 75.975 26.460 76.345 ;
        RECT 28.220 75.810 28.360 77.190 ;
        RECT 28.160 75.490 28.420 75.810 ;
        RECT 24.020 74.810 24.280 75.130 ;
        RECT 24.480 74.810 24.740 75.130 ;
        RECT 25.400 74.810 25.660 75.130 ;
        RECT 27.700 74.810 27.960 75.130 ;
        RECT 28.620 75.040 28.880 75.130 ;
        RECT 28.220 74.900 28.880 75.040 ;
        RECT 23.560 72.770 23.820 73.090 ;
        RECT 24.540 72.750 24.680 74.810 ;
        RECT 24.480 72.430 24.740 72.750 ;
        RECT 24.020 71.410 24.280 71.730 ;
        RECT 23.160 69.630 23.760 69.770 ;
        RECT 23.100 69.030 23.360 69.350 ;
        RECT 23.160 64.930 23.300 69.030 ;
        RECT 23.100 64.610 23.360 64.930 ;
        RECT 23.160 64.330 23.300 64.610 ;
        RECT 22.180 63.930 22.440 64.250 ;
        RECT 22.700 64.190 23.300 64.330 ;
        RECT 21.260 62.910 21.520 63.230 ;
        RECT 21.720 62.910 21.980 63.230 ;
        RECT 21.320 60.850 21.460 62.910 ;
        RECT 21.260 60.530 21.520 60.850 ;
        RECT 21.780 55.750 21.920 62.910 ;
        RECT 22.180 60.870 22.440 61.190 ;
        RECT 22.240 58.470 22.380 60.870 ;
        RECT 22.700 60.510 22.840 64.190 ;
        RECT 23.620 62.170 23.760 69.630 ;
        RECT 23.160 62.030 23.760 62.170 ;
        RECT 22.640 60.190 22.900 60.510 ;
        RECT 22.700 59.490 22.840 60.190 ;
        RECT 22.640 59.170 22.900 59.490 ;
        RECT 22.180 58.150 22.440 58.470 ;
        RECT 22.240 55.750 22.380 58.150 ;
        RECT 21.720 55.430 21.980 55.750 ;
        RECT 22.180 55.430 22.440 55.750 ;
        RECT 23.160 51.330 23.300 62.030 ;
        RECT 23.560 58.150 23.820 58.470 ;
        RECT 23.620 56.770 23.760 58.150 ;
        RECT 23.560 56.450 23.820 56.770 ;
        RECT 24.080 51.330 24.220 71.410 ;
        RECT 25.460 71.390 25.600 74.810 ;
        RECT 27.760 72.750 27.900 74.810 ;
        RECT 28.220 74.110 28.360 74.900 ;
        RECT 28.620 74.810 28.880 74.900 ;
        RECT 28.160 73.790 28.420 74.110 ;
        RECT 27.700 72.430 27.960 72.750 ;
        RECT 26.780 71.750 27.040 72.070 ;
        RECT 27.240 71.750 27.500 72.070 ;
        RECT 25.400 71.070 25.660 71.390 ;
        RECT 24.580 70.535 26.460 70.905 ;
        RECT 25.860 69.370 26.120 69.690 ;
        RECT 25.920 69.010 26.060 69.370 ;
        RECT 25.860 68.690 26.120 69.010 ;
        RECT 24.580 65.095 26.460 65.465 ;
        RECT 26.840 64.930 26.980 71.750 ;
        RECT 27.300 69.690 27.440 71.750 ;
        RECT 27.760 70.030 27.900 72.430 ;
        RECT 28.220 72.410 28.360 73.790 ;
        RECT 28.160 72.090 28.420 72.410 ;
        RECT 27.700 69.710 27.960 70.030 ;
        RECT 27.240 69.370 27.500 69.690 ;
        RECT 28.220 69.010 28.360 72.090 ;
        RECT 28.620 71.750 28.880 72.070 ;
        RECT 28.160 68.690 28.420 69.010 ;
        RECT 28.680 66.970 28.820 71.750 ;
        RECT 28.620 66.650 28.880 66.970 ;
        RECT 28.160 65.630 28.420 65.950 ;
        RECT 26.780 64.610 27.040 64.930 ;
        RECT 24.480 63.590 24.740 63.910 ;
        RECT 25.400 63.590 25.660 63.910 ;
        RECT 24.540 62.170 24.680 63.590 ;
        RECT 25.460 62.170 25.600 63.590 ;
        RECT 24.540 62.030 25.600 62.170 ;
        RECT 24.540 61.530 24.680 62.030 ;
        RECT 28.220 61.530 28.360 65.630 ;
        RECT 28.680 64.930 28.820 66.650 ;
        RECT 28.620 64.610 28.880 64.930 ;
        RECT 24.480 61.210 24.740 61.530 ;
        RECT 28.160 61.210 28.420 61.530 ;
        RECT 24.580 59.655 26.460 60.025 ;
        RECT 28.680 59.490 28.820 64.610 ;
        RECT 28.620 59.170 28.880 59.490 ;
        RECT 24.580 54.215 26.460 54.585 ;
        RECT 23.100 51.010 23.360 51.330 ;
        RECT 24.020 51.010 24.280 51.330 ;
        RECT 28.160 50.670 28.420 50.990 ;
        RECT 28.220 50.310 28.360 50.670 ;
        RECT 26.780 49.990 27.040 50.310 ;
        RECT 28.160 49.990 28.420 50.310 ;
        RECT 21.260 49.650 21.520 49.970 ;
        RECT 18.960 47.950 19.220 48.270 ;
        RECT 20.800 47.950 21.060 48.270 ;
        RECT 14.360 47.610 14.620 47.930 ;
        RECT 18.040 47.610 18.300 47.930 ;
        RECT 11.600 46.590 11.860 46.910 ;
        RECT 13.440 46.590 13.700 46.910 ;
        RECT 9.580 46.055 11.460 46.425 ;
        RECT 8.840 44.550 9.100 44.870 ;
        RECT 8.900 42.150 9.040 44.550 ;
        RECT 11.660 42.830 11.800 46.590 ;
        RECT 13.500 45.210 13.640 46.590 ;
        RECT 14.420 45.890 14.560 47.610 ;
        RECT 15.280 46.590 15.540 46.910 ;
        RECT 14.360 45.570 14.620 45.890 ;
        RECT 13.440 44.890 13.700 45.210 ;
        RECT 15.340 42.830 15.480 46.590 ;
        RECT 11.600 42.510 11.860 42.830 ;
        RECT 15.280 42.510 15.540 42.830 ;
        RECT 8.840 41.830 9.100 42.150 ;
        RECT 8.900 31.270 9.040 41.830 ;
        RECT 9.580 40.615 11.460 40.985 ;
        RECT 9.580 35.175 11.460 35.545 ;
        RECT 18.100 34.330 18.240 47.610 ;
        RECT 18.500 44.210 18.760 44.530 ;
        RECT 18.560 43.170 18.700 44.210 ;
        RECT 18.500 42.850 18.760 43.170 ;
        RECT 19.020 42.490 19.160 47.950 ;
        RECT 21.320 47.930 21.460 49.650 ;
        RECT 24.580 48.775 26.460 49.145 ;
        RECT 26.840 47.930 26.980 49.990 ;
        RECT 28.220 48.610 28.360 49.990 ;
        RECT 28.160 48.290 28.420 48.610 ;
        RECT 27.240 47.950 27.500 48.270 ;
        RECT 28.220 48.010 28.360 48.290 ;
        RECT 21.260 47.610 21.520 47.930 ;
        RECT 26.780 47.610 27.040 47.930 ;
        RECT 21.320 44.190 21.460 47.610 ;
        RECT 21.720 47.270 21.980 47.590 ;
        RECT 24.020 47.270 24.280 47.590 ;
        RECT 21.780 45.210 21.920 47.270 ;
        RECT 21.720 44.890 21.980 45.210 ;
        RECT 21.260 43.870 21.520 44.190 ;
        RECT 18.960 42.170 19.220 42.490 ;
        RECT 18.040 34.010 18.300 34.330 ;
        RECT 10.680 32.990 10.940 33.310 ;
        RECT 10.740 31.950 10.880 32.990 ;
        RECT 18.100 32.290 18.240 34.010 ;
        RECT 18.040 31.970 18.300 32.290 ;
        RECT 10.680 31.630 10.940 31.950 ;
        RECT 17.120 31.630 17.380 31.950 ;
        RECT 8.840 30.950 9.100 31.270 ;
        RECT 9.580 29.735 11.460 30.105 ;
        RECT 17.180 29.570 17.320 31.630 ;
        RECT 17.120 29.250 17.380 29.570 ;
        RECT 19.020 28.210 19.160 42.170 ;
        RECT 21.320 42.150 21.460 43.870 ;
        RECT 21.780 42.830 21.920 44.890 ;
        RECT 21.720 42.510 21.980 42.830 ;
        RECT 21.260 41.830 21.520 42.150 ;
        RECT 23.560 39.110 23.820 39.430 ;
        RECT 23.100 32.990 23.360 33.310 ;
        RECT 19.880 30.950 20.140 31.270 ;
        RECT 19.940 29.570 20.080 30.950 ;
        RECT 19.880 29.250 20.140 29.570 ;
        RECT 23.160 28.550 23.300 32.990 ;
        RECT 23.620 30.590 23.760 39.110 ;
        RECT 24.080 33.650 24.220 47.270 ;
        RECT 25.860 46.930 26.120 47.250 ;
        RECT 25.920 44.870 26.060 46.930 ;
        RECT 27.300 44.870 27.440 47.950 ;
        RECT 28.220 47.930 28.820 48.010 ;
        RECT 27.700 47.610 27.960 47.930 ;
        RECT 28.220 47.870 28.880 47.930 ;
        RECT 28.620 47.610 28.880 47.870 ;
        RECT 25.860 44.550 26.120 44.870 ;
        RECT 27.240 44.550 27.500 44.870 ;
        RECT 24.580 43.335 26.460 43.705 ;
        RECT 27.240 41.830 27.500 42.150 ;
        RECT 26.780 41.150 27.040 41.470 ;
        RECT 26.840 39.770 26.980 41.150 ;
        RECT 26.780 39.450 27.040 39.770 ;
        RECT 24.580 37.895 26.460 38.265 ;
        RECT 27.300 34.330 27.440 41.830 ;
        RECT 27.240 34.010 27.500 34.330 ;
        RECT 27.760 33.990 27.900 47.610 ;
        RECT 28.680 44.870 28.820 47.610 ;
        RECT 29.140 45.890 29.280 79.830 ;
        RECT 29.540 79.230 29.800 79.550 ;
        RECT 29.600 77.510 29.740 79.230 ;
        RECT 29.540 77.190 29.800 77.510 ;
        RECT 29.540 76.510 29.800 76.830 ;
        RECT 29.600 48.270 29.740 76.510 ;
        RECT 30.980 73.090 31.120 85.690 ;
        RECT 34.200 85.670 34.340 86.030 ;
        RECT 34.140 85.350 34.400 85.670 ;
        RECT 34.600 77.190 34.860 77.510 ;
        RECT 33.220 74.810 33.480 75.130 ;
        RECT 31.380 74.470 31.640 74.790 ;
        RECT 30.920 72.770 31.180 73.090 ;
        RECT 30.460 63.250 30.720 63.570 ;
        RECT 30.000 58.830 30.260 59.150 ;
        RECT 30.060 54.050 30.200 58.830 ;
        RECT 30.000 53.730 30.260 54.050 ;
        RECT 30.520 50.310 30.660 63.250 ;
        RECT 31.440 60.510 31.580 74.470 ;
        RECT 33.280 72.070 33.420 74.810 ;
        RECT 33.220 71.750 33.480 72.070 ;
        RECT 34.140 71.750 34.400 72.070 ;
        RECT 33.280 69.350 33.420 71.750 ;
        RECT 33.220 69.030 33.480 69.350 ;
        RECT 34.200 66.630 34.340 71.750 ;
        RECT 34.660 66.970 34.800 77.190 ;
        RECT 35.060 73.790 35.320 74.110 ;
        RECT 35.120 72.070 35.260 73.790 ;
        RECT 35.580 73.090 35.720 88.070 ;
        RECT 35.520 72.770 35.780 73.090 ;
        RECT 35.060 71.750 35.320 72.070 ;
        RECT 35.520 71.410 35.780 71.730 ;
        RECT 35.580 70.370 35.720 71.410 ;
        RECT 35.520 70.050 35.780 70.370 ;
        RECT 34.600 66.650 34.860 66.970 ;
        RECT 34.140 66.310 34.400 66.630 ;
        RECT 34.200 64.590 34.340 66.310 ;
        RECT 34.140 64.270 34.400 64.590 ;
        RECT 34.660 63.570 34.800 66.650 ;
        RECT 34.600 63.250 34.860 63.570 ;
        RECT 31.840 62.910 32.100 63.230 ;
        RECT 31.900 60.850 32.040 62.910 ;
        RECT 31.840 60.530 32.100 60.850 ;
        RECT 31.380 60.190 31.640 60.510 ;
        RECT 31.440 58.470 31.580 60.190 ;
        RECT 31.380 58.150 31.640 58.470 ;
        RECT 32.290 55.235 32.570 55.605 ;
        RECT 34.660 55.410 34.800 63.250 ;
        RECT 35.060 57.470 35.320 57.790 ;
        RECT 35.120 56.090 35.260 57.470 ;
        RECT 35.060 55.770 35.320 56.090 ;
        RECT 32.300 55.090 32.560 55.235 ;
        RECT 34.600 55.090 34.860 55.410 ;
        RECT 34.660 54.050 34.800 55.090 ;
        RECT 34.600 53.730 34.860 54.050 ;
        RECT 33.220 51.010 33.480 51.330 ;
        RECT 33.280 50.650 33.420 51.010 ;
        RECT 33.220 50.330 33.480 50.650 ;
        RECT 30.460 49.990 30.720 50.310 ;
        RECT 29.540 47.950 29.800 48.270 ;
        RECT 30.520 48.010 30.660 49.990 ;
        RECT 30.520 47.930 31.120 48.010 ;
        RECT 33.280 47.930 33.420 50.330 ;
        RECT 30.520 47.870 31.180 47.930 ;
        RECT 30.520 47.250 30.660 47.870 ;
        RECT 30.920 47.610 31.180 47.870 ;
        RECT 32.760 47.610 33.020 47.930 ;
        RECT 33.220 47.610 33.480 47.930 ;
        RECT 30.460 46.930 30.720 47.250 ;
        RECT 29.080 45.570 29.340 45.890 ;
        RECT 28.620 44.550 28.880 44.870 ;
        RECT 28.160 44.210 28.420 44.530 ;
        RECT 28.220 43.170 28.360 44.210 ;
        RECT 28.160 42.850 28.420 43.170 ;
        RECT 32.820 42.830 32.960 47.610 ;
        RECT 34.660 45.210 34.800 53.730 ;
        RECT 36.040 48.270 36.180 88.410 ;
        RECT 37.820 81.950 38.080 82.270 ;
        RECT 37.880 80.570 38.020 81.950 ;
        RECT 39.260 80.570 39.400 91.390 ;
        RECT 40.120 91.130 40.380 91.450 ;
        RECT 40.180 90.430 40.320 91.130 ;
        RECT 40.120 90.110 40.380 90.430 ;
        RECT 39.580 89.575 41.460 89.945 ;
        RECT 43.860 88.300 44.000 98.950 ;
        RECT 45.180 98.270 45.440 98.590 ;
        RECT 45.240 97.230 45.380 98.270 ;
        RECT 45.180 96.910 45.440 97.230 ;
        RECT 44.720 95.550 44.980 95.870 ;
        RECT 44.780 94.850 44.920 95.550 ;
        RECT 44.720 94.530 44.980 94.850 ;
        RECT 46.100 93.850 46.360 94.170 ;
        RECT 44.260 91.470 44.520 91.790 ;
        RECT 44.320 89.410 44.460 91.470 ;
        RECT 46.160 91.110 46.300 93.850 ;
        RECT 46.620 93.570 46.760 118.330 ;
        RECT 47.480 109.150 47.740 109.470 ;
        RECT 47.540 107.770 47.680 109.150 ;
        RECT 47.480 107.450 47.740 107.770 ;
        RECT 47.020 106.430 47.280 106.750 ;
        RECT 47.080 103.010 47.220 106.430 ;
        RECT 47.940 104.730 48.200 105.050 ;
        RECT 47.020 102.690 47.280 103.010 ;
        RECT 48.000 101.990 48.140 104.730 ;
        RECT 47.940 101.670 48.200 101.990 ;
        RECT 48.920 97.570 49.060 120.710 ;
        RECT 49.780 120.370 50.040 120.690 ;
        RECT 49.840 118.990 49.980 120.370 ;
        RECT 49.780 118.670 50.040 118.990 ;
        RECT 49.780 111.870 50.040 112.190 ;
        RECT 49.840 110.470 49.980 111.870 ;
        RECT 50.700 110.470 50.960 110.490 ;
        RECT 49.840 110.330 50.960 110.470 ;
        RECT 51.680 110.470 51.820 120.710 ;
        RECT 52.140 118.650 52.280 121.050 ;
        RECT 55.760 120.710 56.020 121.030 ;
        RECT 55.820 120.350 55.960 120.710 ;
        RECT 67.320 120.690 67.460 123.430 ;
        RECT 67.260 120.370 67.520 120.690 ;
        RECT 55.760 120.030 56.020 120.350 ;
        RECT 60.820 120.030 61.080 120.350 ;
        RECT 54.580 119.495 56.460 119.865 ;
        RECT 52.080 118.330 52.340 118.650 ;
        RECT 54.580 114.055 56.460 114.425 ;
        RECT 58.980 113.230 59.240 113.550 ;
        RECT 55.300 112.550 55.560 112.870 ;
        RECT 55.360 111.170 55.500 112.550 ;
        RECT 55.760 111.870 56.020 112.190 ;
        RECT 55.300 110.850 55.560 111.170 ;
        RECT 51.680 110.330 52.280 110.470 ;
        RECT 50.700 110.170 50.960 110.330 ;
        RECT 49.320 109.830 49.580 110.150 ;
        RECT 49.380 105.730 49.520 109.830 ;
        RECT 50.240 109.150 50.500 109.470 ;
        RECT 50.300 108.110 50.440 109.150 ;
        RECT 50.240 107.790 50.500 108.110 ;
        RECT 49.320 105.410 49.580 105.730 ;
        RECT 50.760 102.330 50.900 110.170 ;
        RECT 51.620 109.830 51.880 110.150 ;
        RECT 51.680 107.770 51.820 109.830 ;
        RECT 51.620 107.450 51.880 107.770 ;
        RECT 50.700 102.010 50.960 102.330 ;
        RECT 48.860 97.250 49.120 97.570 ;
        RECT 47.480 95.550 47.740 95.870 ;
        RECT 46.620 93.430 47.220 93.570 ;
        RECT 46.560 92.830 46.820 93.150 ;
        RECT 46.620 92.130 46.760 92.830 ;
        RECT 46.560 91.810 46.820 92.130 ;
        RECT 46.100 90.790 46.360 91.110 ;
        RECT 45.180 90.110 45.440 90.430 ;
        RECT 45.240 89.410 45.380 90.110 ;
        RECT 44.260 89.090 44.520 89.410 ;
        RECT 45.180 89.090 45.440 89.410 ;
        RECT 44.260 88.300 44.520 88.390 ;
        RECT 43.860 88.160 44.520 88.300 ;
        RECT 44.260 88.070 44.520 88.160 ;
        RECT 39.580 84.135 41.460 84.505 ;
        RECT 43.800 81.950 44.060 82.270 ;
        RECT 37.820 80.250 38.080 80.570 ;
        RECT 39.200 80.250 39.460 80.570 ;
        RECT 43.860 79.550 44.000 81.950 ;
        RECT 44.320 80.650 44.460 88.070 ;
        RECT 46.160 88.050 46.300 90.790 ;
        RECT 47.080 90.770 47.220 93.430 ;
        RECT 47.540 93.150 47.680 95.550 ;
        RECT 50.240 93.510 50.500 93.830 ;
        RECT 47.480 92.830 47.740 93.150 ;
        RECT 47.020 90.450 47.280 90.770 ;
        RECT 47.540 88.390 47.680 92.830 ;
        RECT 50.300 91.450 50.440 93.510 ;
        RECT 50.240 91.130 50.500 91.450 ;
        RECT 47.940 90.110 48.200 90.430 ;
        RECT 48.000 88.730 48.140 90.110 ;
        RECT 47.940 88.410 48.200 88.730 ;
        RECT 47.480 88.070 47.740 88.390 ;
        RECT 46.100 87.730 46.360 88.050 ;
        RECT 47.480 87.390 47.740 87.710 ;
        RECT 47.540 83.290 47.680 87.390 ;
        RECT 48.000 83.290 48.140 88.410 ;
        RECT 50.300 83.290 50.440 91.130 ;
        RECT 51.160 87.390 51.420 87.710 ;
        RECT 47.480 82.970 47.740 83.290 ;
        RECT 47.940 82.970 48.200 83.290 ;
        RECT 50.240 82.970 50.500 83.290 ;
        RECT 44.720 81.950 44.980 82.270 ;
        RECT 44.780 81.250 44.920 81.950 ;
        RECT 44.720 80.930 44.980 81.250 ;
        RECT 44.320 80.510 44.920 80.650 ;
        RECT 45.180 80.590 45.440 80.910 ;
        RECT 36.440 79.230 36.700 79.550 ;
        RECT 43.800 79.230 44.060 79.550 ;
        RECT 36.500 77.850 36.640 79.230 ;
        RECT 39.580 78.695 41.460 79.065 ;
        RECT 43.860 78.530 44.000 79.230 ;
        RECT 43.800 78.210 44.060 78.530 ;
        RECT 36.440 77.530 36.700 77.850 ;
        RECT 44.780 77.510 44.920 80.510 ;
        RECT 45.240 78.530 45.380 80.590 ;
        RECT 45.180 78.210 45.440 78.530 ;
        RECT 44.720 77.190 44.980 77.510 ;
        RECT 41.500 76.850 41.760 77.170 ;
        RECT 41.560 75.810 41.700 76.850 ;
        RECT 41.500 75.490 41.760 75.810 ;
        RECT 38.280 74.810 38.540 75.130 ;
        RECT 38.340 72.070 38.480 74.810 ;
        RECT 39.580 73.255 41.460 73.625 ;
        RECT 38.280 71.750 38.540 72.070 ;
        RECT 38.340 69.690 38.480 71.750 ;
        RECT 44.780 70.030 44.920 77.190 ;
        RECT 47.540 75.810 47.680 82.970 ;
        RECT 47.940 82.290 48.200 82.610 ;
        RECT 48.000 81.250 48.140 82.290 ;
        RECT 47.940 80.930 48.200 81.250 ;
        RECT 50.300 80.570 50.440 82.970 ;
        RECT 50.240 80.250 50.500 80.570 ;
        RECT 47.480 75.490 47.740 75.810 ;
        RECT 50.700 71.750 50.960 72.070 ;
        RECT 49.320 71.070 49.580 71.390 ;
        RECT 49.380 70.030 49.520 71.070 ;
        RECT 44.720 69.710 44.980 70.030 ;
        RECT 49.320 69.710 49.580 70.030 ;
        RECT 37.820 69.370 38.080 69.690 ;
        RECT 38.280 69.370 38.540 69.690 ;
        RECT 36.440 68.350 36.700 68.670 ;
        RECT 36.500 66.970 36.640 68.350 ;
        RECT 36.440 66.650 36.700 66.970 ;
        RECT 37.880 64.930 38.020 69.370 ;
        RECT 37.820 64.610 38.080 64.930 ;
        RECT 36.440 64.270 36.700 64.590 ;
        RECT 36.500 62.210 36.640 64.270 ;
        RECT 38.340 64.250 38.480 69.370 ;
        RECT 42.880 69.030 43.140 69.350 ;
        RECT 46.560 69.030 46.820 69.350 ;
        RECT 39.200 68.350 39.460 68.670 ;
        RECT 38.740 67.330 39.000 67.650 ;
        RECT 38.800 65.690 38.940 67.330 ;
        RECT 39.260 66.290 39.400 68.350 ;
        RECT 39.580 67.815 41.460 68.185 ;
        RECT 39.200 65.970 39.460 66.290 ;
        RECT 42.420 65.970 42.680 66.290 ;
        RECT 38.800 65.550 39.400 65.690 ;
        RECT 38.280 63.930 38.540 64.250 ;
        RECT 36.440 61.890 36.700 62.210 ;
        RECT 38.340 61.190 38.480 63.930 ;
        RECT 39.260 63.910 39.400 65.550 ;
        RECT 42.480 64.930 42.620 65.970 ;
        RECT 42.420 64.610 42.680 64.930 ;
        RECT 39.200 63.590 39.460 63.910 ;
        RECT 38.280 60.870 38.540 61.190 ;
        RECT 39.260 58.470 39.400 63.590 ;
        RECT 42.940 63.570 43.080 69.030 ;
        RECT 46.620 67.650 46.760 69.030 ;
        RECT 46.560 67.330 46.820 67.650 ;
        RECT 50.760 66.630 50.900 71.750 ;
        RECT 50.700 66.310 50.960 66.630 ;
        RECT 42.880 63.250 43.140 63.570 ;
        RECT 39.580 62.375 41.460 62.745 ;
        RECT 42.940 61.530 43.080 63.250 ;
        RECT 50.240 62.910 50.500 63.230 ;
        RECT 50.300 61.530 50.440 62.910 ;
        RECT 42.880 61.210 43.140 61.530 ;
        RECT 50.240 61.210 50.500 61.530 ;
        RECT 42.420 58.830 42.680 59.150 ;
        RECT 39.200 58.150 39.460 58.470 ;
        RECT 39.580 56.935 41.460 57.305 ;
        RECT 42.480 56.770 42.620 58.830 ;
        RECT 42.940 58.810 43.080 61.210 ;
        RECT 46.560 60.190 46.820 60.510 ;
        RECT 46.620 59.150 46.760 60.190 ;
        RECT 46.560 58.830 46.820 59.150 ;
        RECT 42.880 58.490 43.140 58.810 ;
        RECT 46.560 58.150 46.820 58.470 ;
        RECT 46.620 56.770 46.760 58.150 ;
        RECT 42.420 56.450 42.680 56.770 ;
        RECT 46.560 56.450 46.820 56.770 ;
        RECT 45.640 55.430 45.900 55.750 ;
        RECT 45.700 53.370 45.840 55.430 ;
        RECT 47.930 54.555 48.210 54.925 ;
        RECT 48.000 53.710 48.140 54.555 ;
        RECT 51.220 54.050 51.360 87.390 ;
        RECT 52.140 82.270 52.280 110.330 ;
        RECT 55.820 110.150 55.960 111.870 ;
        RECT 57.140 110.170 57.400 110.490 ;
        RECT 55.760 109.830 56.020 110.150 ;
        RECT 56.680 109.490 56.940 109.810 ;
        RECT 54.580 108.615 56.460 108.985 ;
        RECT 53.000 106.430 53.260 106.750 ;
        RECT 53.060 104.710 53.200 106.430 ;
        RECT 53.000 104.390 53.260 104.710 ;
        RECT 53.060 101.990 53.200 104.390 ;
        RECT 56.740 104.030 56.880 109.490 ;
        RECT 57.200 107.430 57.340 110.170 ;
        RECT 58.060 109.830 58.320 110.150 ;
        RECT 58.120 108.110 58.260 109.830 ;
        RECT 59.040 108.450 59.180 113.230 ;
        RECT 60.880 110.470 61.020 120.030 ;
        RECT 67.780 119.330 67.920 138.395 ;
        RECT 69.580 127.655 71.460 128.025 ;
        RECT 74.160 123.770 74.420 124.090 ;
        RECT 69.100 123.430 69.360 123.750 ;
        RECT 67.720 119.010 67.980 119.330 ;
        RECT 66.340 117.310 66.600 117.630 ;
        RECT 61.280 111.870 61.540 112.190 ;
        RECT 60.420 110.330 61.020 110.470 ;
        RECT 58.980 108.130 59.240 108.450 ;
        RECT 58.060 107.790 58.320 108.110 ;
        RECT 57.140 107.110 57.400 107.430 ;
        RECT 57.200 105.730 57.340 107.110 ;
        RECT 57.140 105.410 57.400 105.730 ;
        RECT 58.980 104.390 59.240 104.710 ;
        RECT 56.680 103.710 56.940 104.030 ;
        RECT 57.140 103.710 57.400 104.030 ;
        RECT 54.580 103.175 56.460 103.545 ;
        RECT 53.000 101.670 53.260 101.990 ;
        RECT 53.460 101.330 53.720 101.650 ;
        RECT 52.540 93.510 52.800 93.830 ;
        RECT 53.000 93.510 53.260 93.830 ;
        RECT 52.600 90.770 52.740 93.510 ;
        RECT 53.060 91.110 53.200 93.510 ;
        RECT 53.000 90.790 53.260 91.110 ;
        RECT 52.540 90.450 52.800 90.770 ;
        RECT 52.600 82.950 52.740 90.450 ;
        RECT 53.060 82.950 53.200 90.790 ;
        RECT 52.540 82.630 52.800 82.950 ;
        RECT 53.000 82.630 53.260 82.950 ;
        RECT 52.080 81.950 52.340 82.270 ;
        RECT 52.080 80.480 52.340 80.570 ;
        RECT 52.600 80.480 52.740 82.630 ;
        RECT 53.060 80.570 53.200 82.630 ;
        RECT 52.080 80.340 52.740 80.480 ;
        RECT 52.080 80.250 52.340 80.340 ;
        RECT 52.600 76.830 52.740 80.340 ;
        RECT 53.000 80.250 53.260 80.570 ;
        RECT 53.520 79.550 53.660 101.330 ;
        RECT 53.920 100.990 54.180 101.310 ;
        RECT 53.980 90.430 54.120 100.990 ;
        RECT 54.580 97.735 56.460 98.105 ;
        RECT 56.740 96.890 56.880 103.710 ;
        RECT 54.840 96.570 55.100 96.890 ;
        RECT 55.760 96.570 56.020 96.890 ;
        RECT 56.680 96.570 56.940 96.890 ;
        RECT 54.900 93.685 55.040 96.570 ;
        RECT 55.820 94.850 55.960 96.570 ;
        RECT 55.760 94.530 56.020 94.850 ;
        RECT 56.740 94.170 56.880 96.570 ;
        RECT 56.680 93.850 56.940 94.170 ;
        RECT 54.830 93.315 55.110 93.685 ;
        RECT 54.580 92.295 56.460 92.665 ;
        RECT 54.380 91.130 54.640 91.450 ;
        RECT 53.920 90.110 54.180 90.430 ;
        RECT 54.440 87.620 54.580 91.130 ;
        RECT 54.840 90.790 55.100 91.110 ;
        RECT 54.900 87.710 55.040 90.790 ;
        RECT 53.980 87.480 54.580 87.620 ;
        RECT 53.460 79.230 53.720 79.550 ;
        RECT 52.540 76.510 52.800 76.830 ;
        RECT 52.080 74.810 52.340 75.130 ;
        RECT 52.140 72.750 52.280 74.810 ;
        RECT 52.540 74.470 52.800 74.790 ;
        RECT 52.080 72.430 52.340 72.750 ;
        RECT 52.080 66.650 52.340 66.970 ;
        RECT 52.140 63.910 52.280 66.650 ;
        RECT 52.080 63.590 52.340 63.910 ;
        RECT 52.600 59.150 52.740 74.470 ;
        RECT 53.460 73.000 53.720 73.090 ;
        RECT 53.980 73.000 54.120 87.480 ;
        RECT 54.840 87.390 55.100 87.710 ;
        RECT 54.580 86.855 56.460 87.225 ;
        RECT 56.740 86.010 56.880 93.850 ;
        RECT 56.680 85.690 56.940 86.010 ;
        RECT 57.200 83.970 57.340 103.710 ;
        RECT 59.040 102.330 59.180 104.390 ;
        RECT 58.980 102.010 59.240 102.330 ;
        RECT 57.600 100.990 57.860 101.310 ;
        RECT 57.660 95.870 57.800 100.990 ;
        RECT 58.520 96.910 58.780 97.230 ;
        RECT 57.600 95.550 57.860 95.870 ;
        RECT 57.140 83.650 57.400 83.970 ;
        RECT 58.060 82.970 58.320 83.290 ;
        RECT 55.760 82.860 56.020 82.950 ;
        RECT 55.760 82.720 57.340 82.860 ;
        RECT 55.760 82.630 56.020 82.720 ;
        RECT 54.580 81.415 56.460 81.785 ;
        RECT 56.680 80.250 56.940 80.570 ;
        RECT 54.580 75.975 56.460 76.345 ;
        RECT 56.740 75.810 56.880 80.250 ;
        RECT 55.300 75.490 55.560 75.810 ;
        RECT 56.680 75.490 56.940 75.810 ;
        RECT 54.380 74.810 54.640 75.130 ;
        RECT 53.460 72.860 54.120 73.000 ;
        RECT 53.460 72.770 53.720 72.860 ;
        RECT 54.440 72.750 54.580 74.810 ;
        RECT 55.360 74.790 55.500 75.490 ;
        RECT 55.760 74.810 56.020 75.130 ;
        RECT 55.300 74.470 55.560 74.790 ;
        RECT 52.990 72.235 53.270 72.605 ;
        RECT 54.380 72.430 54.640 72.750 ;
        RECT 52.540 58.830 52.800 59.150 ;
        RECT 52.540 57.470 52.800 57.790 ;
        RECT 52.600 55.750 52.740 57.470 ;
        RECT 52.540 55.430 52.800 55.750 ;
        RECT 48.860 53.730 49.120 54.050 ;
        RECT 51.160 53.730 51.420 54.050 ;
        RECT 47.940 53.390 48.200 53.710 ;
        RECT 45.640 53.050 45.900 53.370 ;
        RECT 44.260 52.710 44.520 53.030 ;
        RECT 39.580 51.495 41.460 51.865 ;
        RECT 35.980 47.950 36.240 48.270 ;
        RECT 37.820 47.610 38.080 47.930 ;
        RECT 36.440 46.590 36.700 46.910 ;
        RECT 34.600 44.890 34.860 45.210 ;
        RECT 36.500 44.530 36.640 46.590 ;
        RECT 36.900 44.890 37.160 45.210 ;
        RECT 36.440 44.210 36.700 44.530 ;
        RECT 32.760 42.510 33.020 42.830 ;
        RECT 34.140 42.510 34.400 42.830 ;
        RECT 34.200 40.450 34.340 42.510 ;
        RECT 34.140 40.130 34.400 40.450 ;
        RECT 36.960 37.050 37.100 44.890 ;
        RECT 37.880 43.170 38.020 47.610 ;
        RECT 43.800 47.270 44.060 47.590 ;
        RECT 39.580 46.055 41.460 46.425 ;
        RECT 43.860 43.170 44.000 47.270 ;
        RECT 44.320 45.890 44.460 52.710 ;
        RECT 45.700 49.970 45.840 53.050 ;
        RECT 48.920 50.310 49.060 53.730 ;
        RECT 49.320 53.050 49.580 53.370 ;
        RECT 50.240 53.050 50.500 53.370 ;
        RECT 51.160 53.050 51.420 53.370 ;
        RECT 49.380 50.310 49.520 53.050 ;
        RECT 48.860 49.990 49.120 50.310 ;
        RECT 49.320 49.990 49.580 50.310 ;
        RECT 45.640 49.650 45.900 49.970 ;
        RECT 44.260 45.570 44.520 45.890 ;
        RECT 37.820 42.850 38.080 43.170 ;
        RECT 43.800 42.850 44.060 43.170 ;
        RECT 41.960 41.150 42.220 41.470 ;
        RECT 39.580 40.615 41.460 40.985 ;
        RECT 42.020 39.430 42.160 41.150 ;
        RECT 41.960 39.110 42.220 39.430 ;
        RECT 39.200 38.430 39.460 38.750 ;
        RECT 39.260 37.390 39.400 38.430 ;
        RECT 43.860 37.730 44.000 42.850 ;
        RECT 44.320 42.830 44.460 45.570 ;
        RECT 45.700 44.870 45.840 49.650 ;
        RECT 47.940 48.290 48.200 48.610 ;
        RECT 47.020 46.590 47.280 46.910 ;
        RECT 45.640 44.550 45.900 44.870 ;
        RECT 44.260 42.510 44.520 42.830 ;
        RECT 45.700 39.770 45.840 44.550 ;
        RECT 47.080 42.150 47.220 46.590 ;
        RECT 47.020 41.830 47.280 42.150 ;
        RECT 45.640 39.450 45.900 39.770 ;
        RECT 43.800 37.410 44.060 37.730 ;
        RECT 39.200 37.070 39.460 37.390 ;
        RECT 42.880 37.070 43.140 37.390 ;
        RECT 36.900 36.730 37.160 37.050 ;
        RECT 37.820 36.730 38.080 37.050 ;
        RECT 27.700 33.670 27.960 33.990 ;
        RECT 24.020 33.330 24.280 33.650 ;
        RECT 27.240 32.990 27.500 33.310 ;
        RECT 24.580 32.455 26.460 32.825 ;
        RECT 27.300 32.290 27.440 32.990 ;
        RECT 27.240 31.970 27.500 32.290 ;
        RECT 24.940 31.630 25.200 31.950 ;
        RECT 23.560 30.270 23.820 30.590 ;
        RECT 25.000 29.570 25.140 31.630 ;
        RECT 27.760 31.270 27.900 33.670 ;
        RECT 37.880 31.610 38.020 36.730 ;
        RECT 39.580 35.175 41.460 35.545 ;
        RECT 42.940 34.330 43.080 37.070 ;
        RECT 42.880 34.010 43.140 34.330 ;
        RECT 45.700 33.990 45.840 39.450 ;
        RECT 47.080 36.710 47.220 41.830 ;
        RECT 47.020 36.620 47.280 36.710 ;
        RECT 47.020 36.480 47.680 36.620 ;
        RECT 47.020 36.390 47.280 36.480 ;
        RECT 47.020 35.710 47.280 36.030 ;
        RECT 42.420 33.670 42.680 33.990 ;
        RECT 45.640 33.670 45.900 33.990 ;
        RECT 41.040 32.990 41.300 33.310 ;
        RECT 41.100 31.610 41.240 32.990 ;
        RECT 37.820 31.290 38.080 31.610 ;
        RECT 41.040 31.290 41.300 31.610 ;
        RECT 27.700 30.950 27.960 31.270 ;
        RECT 34.140 30.950 34.400 31.270 ;
        RECT 26.780 30.610 27.040 30.930 ;
        RECT 25.400 30.270 25.660 30.590 ;
        RECT 24.940 29.250 25.200 29.570 ;
        RECT 25.460 28.890 25.600 30.270 ;
        RECT 26.840 28.890 26.980 30.610 ;
        RECT 34.200 29.570 34.340 30.950 ;
        RECT 34.140 29.250 34.400 29.570 ;
        RECT 25.400 28.570 25.660 28.890 ;
        RECT 26.780 28.570 27.040 28.890 ;
        RECT 23.100 28.230 23.360 28.550 ;
        RECT 18.960 27.890 19.220 28.210 ;
        RECT 24.580 27.015 26.460 27.385 ;
        RECT 37.880 26.170 38.020 31.290 ;
        RECT 39.580 29.735 41.460 30.105 ;
        RECT 42.480 28.550 42.620 33.670 ;
        RECT 47.080 33.650 47.220 35.710 ;
        RECT 47.020 33.330 47.280 33.650 ;
        RECT 45.180 32.990 45.440 33.310 ;
        RECT 43.340 31.630 43.600 31.950 ;
        RECT 43.400 29.570 43.540 31.630 ;
        RECT 43.340 29.250 43.600 29.570 ;
        RECT 42.420 28.230 42.680 28.550 ;
        RECT 40.580 27.550 40.840 27.870 ;
        RECT 40.640 26.170 40.780 27.550 ;
        RECT 45.240 26.510 45.380 32.990 ;
        RECT 47.020 31.970 47.280 32.290 ;
        RECT 47.080 31.610 47.220 31.970 ;
        RECT 47.020 31.290 47.280 31.610 ;
        RECT 47.080 28.890 47.220 31.290 ;
        RECT 47.540 31.270 47.680 36.480 ;
        RECT 48.000 31.610 48.140 48.290 ;
        RECT 48.920 44.870 49.060 49.990 ;
        RECT 49.380 47.930 49.520 49.990 ;
        RECT 50.300 49.630 50.440 53.050 ;
        RECT 51.220 51.330 51.360 53.050 ;
        RECT 51.160 51.010 51.420 51.330 ;
        RECT 50.700 49.990 50.960 50.310 ;
        RECT 51.220 50.220 51.360 51.010 ;
        RECT 51.620 50.220 51.880 50.310 ;
        RECT 51.220 50.080 51.880 50.220 ;
        RECT 50.240 49.310 50.500 49.630 ;
        RECT 49.320 47.610 49.580 47.930 ;
        RECT 48.860 44.550 49.120 44.870 ;
        RECT 48.400 39.450 48.660 39.770 ;
        RECT 47.940 31.290 48.200 31.610 ;
        RECT 47.480 30.950 47.740 31.270 ;
        RECT 47.540 28.890 47.680 30.950 ;
        RECT 48.460 28.890 48.600 39.450 ;
        RECT 50.760 37.730 50.900 49.990 ;
        RECT 51.220 47.930 51.360 50.080 ;
        RECT 51.620 49.990 51.880 50.080 ;
        RECT 52.080 49.650 52.340 49.970 ;
        RECT 51.620 49.310 51.880 49.630 ;
        RECT 51.160 47.610 51.420 47.930 ;
        RECT 51.680 47.590 51.820 49.310 ;
        RECT 52.140 48.610 52.280 49.650 ;
        RECT 52.080 48.290 52.340 48.610 ;
        RECT 53.060 48.270 53.200 72.235 ;
        RECT 55.820 72.070 55.960 74.810 ;
        RECT 57.200 73.090 57.340 82.720 ;
        RECT 57.600 79.910 57.860 80.230 ;
        RECT 57.140 72.770 57.400 73.090 ;
        RECT 54.380 71.980 54.640 72.070 ;
        RECT 53.980 71.840 54.640 71.980 ;
        RECT 53.460 69.370 53.720 69.690 ;
        RECT 53.520 66.630 53.660 69.370 ;
        RECT 53.460 66.310 53.720 66.630 ;
        RECT 53.520 64.930 53.660 66.310 ;
        RECT 53.980 64.930 54.120 71.840 ;
        RECT 54.380 71.750 54.640 71.840 ;
        RECT 55.760 71.750 56.020 72.070 ;
        RECT 54.580 70.535 56.460 70.905 ;
        RECT 54.580 65.095 56.460 65.465 ;
        RECT 53.460 64.610 53.720 64.930 ;
        RECT 53.920 64.610 54.180 64.930 ;
        RECT 53.460 63.590 53.720 63.910 ;
        RECT 53.520 59.490 53.660 63.590 ;
        RECT 53.980 60.510 54.120 64.610 ;
        RECT 57.660 62.170 57.800 79.910 ;
        RECT 57.200 62.030 57.800 62.170 ;
        RECT 53.920 60.190 54.180 60.510 ;
        RECT 53.980 59.490 54.120 60.190 ;
        RECT 54.580 59.655 56.460 60.025 ;
        RECT 53.460 59.170 53.720 59.490 ;
        RECT 53.920 59.170 54.180 59.490 ;
        RECT 53.520 58.810 53.660 59.170 ;
        RECT 53.460 58.490 53.720 58.810 ;
        RECT 54.580 54.215 56.460 54.585 ;
        RECT 55.300 52.710 55.560 53.030 ;
        RECT 55.360 51.330 55.500 52.710 ;
        RECT 57.200 51.330 57.340 62.030 ;
        RECT 55.300 51.010 55.560 51.330 ;
        RECT 57.140 51.010 57.400 51.330 ;
        RECT 55.360 50.310 55.500 51.010 ;
        RECT 58.120 50.650 58.260 82.970 ;
        RECT 58.580 73.090 58.720 96.910 ;
        RECT 59.440 87.390 59.700 87.710 ;
        RECT 59.500 86.010 59.640 87.390 ;
        RECT 59.440 85.690 59.700 86.010 ;
        RECT 60.420 81.250 60.560 110.330 ;
        RECT 61.340 108.530 61.480 111.870 ;
        RECT 64.960 109.490 65.220 109.810 ;
        RECT 61.740 109.150 62.000 109.470 ;
        RECT 60.880 108.390 61.480 108.530 ;
        RECT 61.800 108.450 61.940 109.150 ;
        RECT 65.020 108.450 65.160 109.490 ;
        RECT 60.880 108.110 61.020 108.390 ;
        RECT 61.740 108.130 62.000 108.450 ;
        RECT 64.960 108.130 65.220 108.450 ;
        RECT 60.820 107.790 61.080 108.110 ;
        RECT 60.880 102.330 61.020 107.790 ;
        RECT 61.800 105.050 61.940 108.130 ;
        RECT 62.660 107.110 62.920 107.430 ;
        RECT 62.720 105.730 62.860 107.110 ;
        RECT 62.660 105.410 62.920 105.730 ;
        RECT 61.740 104.730 62.000 105.050 ;
        RECT 60.820 102.010 61.080 102.330 ;
        RECT 66.400 101.990 66.540 117.310 ;
        RECT 69.160 116.270 69.300 123.430 ;
        RECT 69.580 122.215 71.460 122.585 ;
        RECT 74.220 122.050 74.360 123.770 ;
        RECT 74.680 123.750 74.820 138.990 ;
        RECT 74.620 123.430 74.880 123.750 ;
        RECT 81.120 122.050 81.260 138.990 ;
        RECT 84.580 124.935 86.460 125.305 ;
        RECT 88.480 123.750 88.620 138.990 ;
        RECT 92.620 138.990 93.470 139.130 ;
        RECT 100.190 138.990 101.960 139.130 ;
        RECT 113.070 138.990 114.380 139.130 ;
        RECT 89.800 123.770 90.060 124.090 ;
        RECT 83.360 123.430 83.620 123.750 ;
        RECT 87.960 123.430 88.220 123.750 ;
        RECT 88.420 123.430 88.680 123.750 ;
        RECT 74.160 121.730 74.420 122.050 ;
        RECT 81.060 121.730 81.320 122.050 ;
        RECT 74.160 120.940 74.420 121.030 ;
        RECT 74.160 120.800 75.280 120.940 ;
        RECT 74.160 120.710 74.420 120.800 ;
        RECT 75.140 120.350 75.280 120.800 ;
        RECT 75.540 120.370 75.800 120.690 ;
        RECT 76.000 120.370 76.260 120.690 ;
        RECT 71.860 120.030 72.120 120.350 ;
        RECT 75.080 120.030 75.340 120.350 ;
        RECT 71.920 118.990 72.060 120.030 ;
        RECT 75.140 118.990 75.280 120.030 ;
        RECT 71.860 118.670 72.120 118.990 ;
        RECT 75.080 118.670 75.340 118.990 ;
        RECT 73.700 118.330 73.960 118.650 ;
        RECT 71.860 117.990 72.120 118.310 ;
        RECT 69.580 116.775 71.460 117.145 ;
        RECT 71.920 116.610 72.060 117.990 ;
        RECT 73.760 117.630 73.900 118.330 ;
        RECT 75.600 118.310 75.740 120.370 ;
        RECT 76.060 119.330 76.200 120.370 ;
        RECT 76.000 119.010 76.260 119.330 ;
        RECT 75.540 117.990 75.800 118.310 ;
        RECT 73.700 117.310 73.960 117.630 ;
        RECT 71.860 116.290 72.120 116.610 ;
        RECT 69.100 115.950 69.360 116.270 ;
        RECT 72.320 115.270 72.580 115.590 ;
        RECT 69.580 111.335 71.460 111.705 ;
        RECT 69.580 105.895 71.460 106.265 ;
        RECT 68.180 104.050 68.440 104.370 ;
        RECT 68.240 103.010 68.380 104.050 ;
        RECT 68.180 102.690 68.440 103.010 ;
        RECT 67.260 102.010 67.520 102.330 ;
        RECT 66.340 101.670 66.600 101.990 ;
        RECT 62.200 96.230 62.460 96.550 ;
        RECT 62.260 94.850 62.400 96.230 ;
        RECT 64.960 95.550 65.220 95.870 ;
        RECT 62.200 94.530 62.460 94.850 ;
        RECT 61.280 93.170 61.540 93.490 ;
        RECT 61.340 92.130 61.480 93.170 ;
        RECT 64.500 92.890 64.760 93.150 ;
        RECT 64.100 92.830 64.760 92.890 ;
        RECT 64.100 92.750 64.700 92.830 ;
        RECT 61.280 91.810 61.540 92.130 ;
        RECT 61.280 91.130 61.540 91.450 ;
        RECT 61.340 83.290 61.480 91.130 ;
        RECT 64.100 91.110 64.240 92.750 ;
        RECT 65.020 92.130 65.160 95.550 ;
        RECT 64.960 91.810 65.220 92.130 ;
        RECT 64.040 90.790 64.300 91.110 ;
        RECT 62.660 88.070 62.920 88.390 ;
        RECT 62.200 86.030 62.460 86.350 ;
        RECT 61.280 82.970 61.540 83.290 ;
        RECT 62.260 82.950 62.400 86.030 ;
        RECT 62.720 83.970 62.860 88.070 ;
        RECT 64.100 88.050 64.240 90.790 ;
        RECT 64.040 87.730 64.300 88.050 ;
        RECT 62.660 83.650 62.920 83.970 ;
        RECT 64.100 82.950 64.240 87.730 ;
        RECT 65.020 85.670 65.160 91.810 ;
        RECT 64.960 85.350 65.220 85.670 ;
        RECT 64.960 82.970 65.220 83.290 ;
        RECT 62.200 82.630 62.460 82.950 ;
        RECT 64.040 82.630 64.300 82.950 ;
        RECT 60.360 80.930 60.620 81.250 ;
        RECT 62.200 80.930 62.460 81.250 ;
        RECT 59.440 74.810 59.700 75.130 ;
        RECT 58.520 72.770 58.780 73.090 ;
        RECT 58.980 71.925 59.240 72.070 ;
        RECT 58.970 71.555 59.250 71.925 ;
        RECT 59.040 67.650 59.180 71.555 ;
        RECT 59.500 71.390 59.640 74.810 ;
        RECT 61.280 72.430 61.540 72.750 ;
        RECT 61.340 72.070 61.480 72.430 ;
        RECT 59.900 71.750 60.160 72.070 ;
        RECT 61.280 71.750 61.540 72.070 ;
        RECT 59.440 71.070 59.700 71.390 ;
        RECT 59.500 70.370 59.640 71.070 ;
        RECT 59.440 70.050 59.700 70.370 ;
        RECT 59.960 69.690 60.100 71.750 ;
        RECT 61.340 70.370 61.480 71.750 ;
        RECT 61.280 70.050 61.540 70.370 ;
        RECT 62.260 69.690 62.400 80.930 ;
        RECT 62.660 77.530 62.920 77.850 ;
        RECT 62.720 75.810 62.860 77.530 ;
        RECT 62.660 75.490 62.920 75.810 ;
        RECT 64.040 75.325 64.300 75.470 ;
        RECT 64.030 74.955 64.310 75.325 ;
        RECT 63.120 73.790 63.380 74.110 ;
        RECT 59.900 69.370 60.160 69.690 ;
        RECT 62.200 69.600 62.460 69.690 ;
        RECT 62.200 69.460 62.860 69.600 ;
        RECT 62.200 69.370 62.460 69.460 ;
        RECT 60.360 69.090 60.620 69.350 ;
        RECT 60.360 69.030 62.400 69.090 ;
        RECT 60.420 68.950 62.400 69.030 ;
        RECT 62.260 68.670 62.400 68.950 ;
        RECT 62.200 68.350 62.460 68.670 ;
        RECT 58.980 67.330 59.240 67.650 ;
        RECT 62.260 67.310 62.400 68.350 ;
        RECT 62.200 66.990 62.460 67.310 ;
        RECT 62.720 62.170 62.860 69.460 ;
        RECT 63.180 64.930 63.320 73.790 ;
        RECT 64.040 71.750 64.300 72.070 ;
        RECT 64.100 69.690 64.240 71.750 ;
        RECT 64.040 69.370 64.300 69.690 ;
        RECT 64.100 67.050 64.240 69.370 ;
        RECT 65.020 68.670 65.160 82.970 ;
        RECT 66.400 81.250 66.540 101.670 ;
        RECT 67.320 98.930 67.460 102.010 ;
        RECT 69.580 100.455 71.460 100.825 ;
        RECT 67.260 98.610 67.520 98.930 ;
        RECT 67.320 98.445 67.460 98.610 ;
        RECT 67.250 98.075 67.530 98.445 ;
        RECT 68.180 98.270 68.440 98.590 ;
        RECT 71.860 98.270 72.120 98.590 ;
        RECT 68.240 97.230 68.380 98.270 ;
        RECT 68.180 96.910 68.440 97.230 ;
        RECT 71.920 96.890 72.060 98.270 ;
        RECT 71.860 96.570 72.120 96.890 ;
        RECT 69.580 95.015 71.460 95.385 ;
        RECT 66.800 93.510 67.060 93.830 ;
        RECT 71.860 93.510 72.120 93.830 ;
        RECT 66.860 92.130 67.000 93.510 ;
        RECT 66.800 91.810 67.060 92.130 ;
        RECT 71.920 90.770 72.060 93.510 ;
        RECT 71.860 90.450 72.120 90.770 ;
        RECT 69.580 89.575 71.460 89.945 ;
        RECT 69.100 88.410 69.360 88.730 ;
        RECT 68.180 88.070 68.440 88.390 ;
        RECT 68.240 86.350 68.380 88.070 ;
        RECT 68.640 87.730 68.900 88.050 ;
        RECT 68.180 86.030 68.440 86.350 ;
        RECT 67.720 85.690 67.980 86.010 ;
        RECT 67.780 84.990 67.920 85.690 ;
        RECT 67.260 84.670 67.520 84.990 ;
        RECT 67.720 84.670 67.980 84.990 ;
        RECT 67.320 82.950 67.460 84.670 ;
        RECT 68.240 82.950 68.380 86.030 ;
        RECT 68.700 85.330 68.840 87.730 ;
        RECT 68.640 85.010 68.900 85.330 ;
        RECT 68.700 83.290 68.840 85.010 ;
        RECT 69.160 84.990 69.300 88.410 ;
        RECT 69.100 84.670 69.360 84.990 ;
        RECT 68.640 82.970 68.900 83.290 ;
        RECT 67.260 82.630 67.520 82.950 ;
        RECT 68.180 82.630 68.440 82.950 ;
        RECT 67.720 81.950 67.980 82.270 ;
        RECT 66.340 80.930 66.600 81.250 ;
        RECT 65.420 80.590 65.680 80.910 ;
        RECT 65.480 74.450 65.620 80.590 ;
        RECT 67.780 80.230 67.920 81.950 ;
        RECT 67.720 79.910 67.980 80.230 ;
        RECT 67.720 79.230 67.980 79.550 ;
        RECT 66.800 77.190 67.060 77.510 ;
        RECT 66.340 76.510 66.600 76.830 ;
        RECT 66.400 75.470 66.540 76.510 ;
        RECT 66.340 75.150 66.600 75.470 ;
        RECT 65.880 74.810 66.140 75.130 ;
        RECT 65.420 74.130 65.680 74.450 ;
        RECT 65.480 71.390 65.620 74.130 ;
        RECT 65.420 71.070 65.680 71.390 ;
        RECT 65.940 69.690 66.080 74.810 ;
        RECT 65.420 69.370 65.680 69.690 ;
        RECT 65.880 69.370 66.140 69.690 ;
        RECT 64.960 68.350 65.220 68.670 ;
        RECT 63.640 66.910 64.240 67.050 ;
        RECT 63.120 64.610 63.380 64.930 ;
        RECT 63.640 63.650 63.780 66.910 ;
        RECT 65.480 66.630 65.620 69.370 ;
        RECT 64.040 66.310 64.300 66.630 ;
        RECT 65.420 66.310 65.680 66.630 ;
        RECT 64.100 64.250 64.240 66.310 ;
        RECT 64.500 65.970 64.760 66.290 ;
        RECT 64.040 63.930 64.300 64.250 ;
        RECT 63.640 63.510 64.240 63.650 ;
        RECT 62.720 62.030 63.780 62.170 ;
        RECT 63.640 61.190 63.780 62.030 ;
        RECT 63.580 60.870 63.840 61.190 ;
        RECT 59.900 60.190 60.160 60.510 ;
        RECT 59.960 58.470 60.100 60.190 ;
        RECT 59.900 58.150 60.160 58.470 ;
        RECT 62.200 55.770 62.460 56.090 ;
        RECT 60.820 54.750 61.080 55.070 ;
        RECT 60.880 52.690 61.020 54.750 ;
        RECT 61.740 53.450 62.000 53.710 ;
        RECT 62.260 53.450 62.400 55.770 ;
        RECT 63.120 55.430 63.380 55.750 ;
        RECT 63.180 54.050 63.320 55.430 ;
        RECT 63.120 53.730 63.380 54.050 ;
        RECT 61.740 53.390 62.400 53.450 ;
        RECT 61.800 53.310 62.400 53.390 ;
        RECT 60.820 52.370 61.080 52.690 ;
        RECT 58.060 50.330 58.320 50.650 ;
        RECT 53.460 49.990 53.720 50.310 ;
        RECT 55.300 49.990 55.560 50.310 ;
        RECT 53.520 48.610 53.660 49.990 ;
        RECT 54.580 48.775 56.460 49.145 ;
        RECT 53.460 48.290 53.720 48.610 ;
        RECT 53.000 47.950 53.260 48.270 ;
        RECT 55.760 47.610 56.020 47.930 ;
        RECT 51.620 47.270 51.880 47.590 ;
        RECT 51.620 44.890 51.880 45.210 ;
        RECT 51.680 39.770 51.820 44.890 ;
        RECT 55.820 44.610 55.960 47.610 ;
        RECT 60.880 47.590 61.020 52.370 ;
        RECT 61.280 52.030 61.540 52.350 ;
        RECT 61.340 48.270 61.480 52.030 ;
        RECT 61.280 47.950 61.540 48.270 ;
        RECT 60.820 47.270 61.080 47.590 ;
        RECT 58.060 46.590 58.320 46.910 ;
        RECT 57.600 44.890 57.860 45.210 ;
        RECT 55.820 44.530 57.340 44.610 ;
        RECT 55.760 44.470 57.340 44.530 ;
        RECT 55.760 44.210 56.020 44.470 ;
        RECT 54.580 43.335 56.460 43.705 ;
        RECT 51.620 39.450 51.880 39.770 ;
        RECT 56.680 38.770 56.940 39.090 ;
        RECT 54.580 37.895 56.460 38.265 ;
        RECT 56.740 37.730 56.880 38.770 ;
        RECT 48.860 37.410 49.120 37.730 ;
        RECT 50.700 37.410 50.960 37.730 ;
        RECT 56.680 37.410 56.940 37.730 ;
        RECT 48.920 32.290 49.060 37.410 ;
        RECT 57.200 37.050 57.340 44.470 ;
        RECT 57.660 43.170 57.800 44.890 ;
        RECT 58.120 44.530 58.260 46.590 ;
        RECT 58.060 44.210 58.320 44.530 ;
        RECT 57.600 42.850 57.860 43.170 ;
        RECT 60.880 42.490 61.020 47.270 ;
        RECT 62.260 44.530 62.400 53.310 ;
        RECT 63.180 50.650 63.320 53.730 ;
        RECT 63.640 53.370 63.780 60.870 ;
        RECT 63.580 53.050 63.840 53.370 ;
        RECT 63.120 50.330 63.380 50.650 ;
        RECT 62.660 46.930 62.920 47.250 ;
        RECT 62.720 45.550 62.860 46.930 ;
        RECT 64.100 45.890 64.240 63.510 ;
        RECT 64.560 61.190 64.700 65.970 ;
        RECT 64.960 63.930 65.220 64.250 ;
        RECT 65.020 61.190 65.160 63.930 ;
        RECT 65.480 63.910 65.620 66.310 ;
        RECT 65.420 63.590 65.680 63.910 ;
        RECT 65.480 61.190 65.620 63.590 ;
        RECT 64.500 60.870 64.760 61.190 ;
        RECT 64.960 60.870 65.220 61.190 ;
        RECT 65.420 60.870 65.680 61.190 ;
        RECT 64.040 45.570 64.300 45.890 ;
        RECT 62.660 45.230 62.920 45.550 ;
        RECT 62.200 44.210 62.460 44.530 ;
        RECT 60.820 42.170 61.080 42.490 ;
        RECT 62.260 42.150 62.400 44.210 ;
        RECT 62.720 42.570 62.860 45.230 ;
        RECT 63.120 44.890 63.380 45.210 ;
        RECT 63.180 43.170 63.320 44.890 ;
        RECT 63.580 43.870 63.840 44.190 ;
        RECT 63.120 42.850 63.380 43.170 ;
        RECT 62.720 42.430 63.320 42.570 ;
        RECT 62.200 41.830 62.460 42.150 ;
        RECT 62.660 41.830 62.920 42.150 ;
        RECT 57.600 38.430 57.860 38.750 ;
        RECT 57.660 37.730 57.800 38.430 ;
        RECT 62.260 37.730 62.400 41.830 ;
        RECT 57.600 37.410 57.860 37.730 ;
        RECT 62.200 37.410 62.460 37.730 ;
        RECT 57.140 36.730 57.400 37.050 ;
        RECT 58.520 36.730 58.780 37.050 ;
        RECT 54.580 32.455 56.460 32.825 ;
        RECT 48.860 31.970 49.120 32.290 ;
        RECT 47.020 28.570 47.280 28.890 ;
        RECT 47.480 28.570 47.740 28.890 ;
        RECT 48.400 28.570 48.660 28.890 ;
        RECT 47.080 26.850 47.220 28.570 ;
        RECT 48.920 28.550 49.060 31.970 ;
        RECT 53.000 30.270 53.260 30.590 ;
        RECT 53.060 28.890 53.200 30.270 ;
        RECT 53.000 28.570 53.260 28.890 ;
        RECT 48.860 28.230 49.120 28.550 ;
        RECT 56.680 27.890 56.940 28.210 ;
        RECT 54.580 27.015 56.460 27.385 ;
        RECT 56.740 26.850 56.880 27.890 ;
        RECT 57.200 27.870 57.340 36.730 ;
        RECT 58.580 35.010 58.720 36.730 ;
        RECT 61.740 35.710 62.000 36.030 ;
        RECT 61.800 35.010 61.940 35.710 ;
        RECT 58.520 34.690 58.780 35.010 ;
        RECT 61.740 34.690 62.000 35.010 ;
        RECT 62.260 33.990 62.400 37.410 ;
        RECT 62.200 33.670 62.460 33.990 ;
        RECT 59.900 33.330 60.160 33.650 ;
        RECT 59.960 31.270 60.100 33.330 ;
        RECT 62.720 31.610 62.860 41.830 ;
        RECT 63.180 34.920 63.320 42.430 ;
        RECT 63.640 42.150 63.780 43.870 ;
        RECT 64.560 43.170 64.700 60.870 ;
        RECT 65.020 56.770 65.160 60.870 ;
        RECT 64.960 56.450 65.220 56.770 ;
        RECT 65.480 55.750 65.620 60.870 ;
        RECT 65.420 55.430 65.680 55.750 ;
        RECT 64.960 54.750 65.220 55.070 ;
        RECT 65.020 53.030 65.160 54.750 ;
        RECT 65.480 53.030 65.620 55.430 ;
        RECT 65.940 54.050 66.080 69.370 ;
        RECT 66.400 68.670 66.540 75.150 ;
        RECT 66.860 72.070 67.000 77.190 ;
        RECT 67.780 75.130 67.920 79.230 ;
        RECT 68.240 78.190 68.380 82.630 ;
        RECT 68.180 77.870 68.440 78.190 ;
        RECT 68.700 77.850 68.840 82.970 ;
        RECT 68.640 77.530 68.900 77.850 ;
        RECT 69.160 77.510 69.300 84.670 ;
        RECT 69.580 84.135 71.460 84.505 ;
        RECT 71.920 83.630 72.060 90.450 ;
        RECT 71.860 83.310 72.120 83.630 ;
        RECT 71.860 82.290 72.120 82.610 ;
        RECT 71.920 81.250 72.060 82.290 ;
        RECT 71.860 80.930 72.120 81.250 ;
        RECT 69.580 78.695 71.460 79.065 ;
        RECT 69.100 77.190 69.360 77.510 ;
        RECT 67.720 74.810 67.980 75.130 ;
        RECT 66.800 71.750 67.060 72.070 ;
        RECT 67.780 69.010 67.920 74.810 ;
        RECT 68.180 72.090 68.440 72.410 ;
        RECT 67.720 68.690 67.980 69.010 ;
        RECT 66.340 68.350 66.600 68.670 ;
        RECT 68.240 67.650 68.380 72.090 ;
        RECT 68.640 69.370 68.900 69.690 ;
        RECT 68.180 67.330 68.440 67.650 ;
        RECT 68.700 66.290 68.840 69.370 ;
        RECT 68.640 65.970 68.900 66.290 ;
        RECT 69.160 60.510 69.300 77.190 ;
        RECT 72.380 74.645 72.520 115.270 ;
        RECT 73.760 110.470 73.900 117.310 ;
        RECT 75.600 115.590 75.740 117.990 ;
        RECT 75.540 115.270 75.800 115.590 ;
        RECT 77.840 115.270 78.100 115.590 ;
        RECT 75.600 112.870 75.740 115.270 ;
        RECT 77.900 113.890 78.040 115.270 ;
        RECT 80.600 114.930 80.860 115.250 ;
        RECT 80.660 113.890 80.800 114.930 ;
        RECT 77.840 113.570 78.100 113.890 ;
        RECT 80.600 113.570 80.860 113.890 ;
        RECT 75.540 112.550 75.800 112.870 ;
        RECT 75.600 110.490 75.740 112.550 ;
        RECT 82.900 111.870 83.160 112.190 ;
        RECT 73.760 110.330 74.360 110.470 ;
        RECT 72.780 109.830 73.040 110.150 ;
        RECT 72.840 108.450 72.980 109.830 ;
        RECT 72.780 108.130 73.040 108.450 ;
        RECT 74.220 107.770 74.360 110.330 ;
        RECT 75.540 110.170 75.800 110.490 ;
        RECT 79.680 110.170 79.940 110.490 ;
        RECT 74.160 107.450 74.420 107.770 ;
        RECT 75.080 107.450 75.340 107.770 ;
        RECT 75.140 98.930 75.280 107.450 ;
        RECT 75.600 105.050 75.740 110.170 ;
        RECT 76.460 109.490 76.720 109.810 ;
        RECT 76.520 105.730 76.660 109.490 ;
        RECT 79.740 108.450 79.880 110.170 ;
        RECT 79.680 108.360 79.940 108.450 ;
        RECT 78.820 108.220 79.940 108.360 ;
        RECT 77.380 107.790 77.640 108.110 ;
        RECT 76.920 107.110 77.180 107.430 ;
        RECT 76.460 105.410 76.720 105.730 ;
        RECT 75.540 104.730 75.800 105.050 ;
        RECT 75.080 98.610 75.340 98.930 ;
        RECT 74.620 96.910 74.880 97.230 ;
        RECT 72.780 95.550 73.040 95.870 ;
        RECT 72.840 94.170 72.980 95.550 ;
        RECT 74.680 94.850 74.820 96.910 ;
        RECT 74.620 94.530 74.880 94.850 ;
        RECT 72.780 93.850 73.040 94.170 ;
        RECT 75.140 93.830 75.280 98.610 ;
        RECT 75.600 97.570 75.740 104.730 ;
        RECT 76.980 104.710 77.120 107.110 ;
        RECT 76.920 104.390 77.180 104.710 ;
        RECT 76.920 98.950 77.180 99.270 ;
        RECT 75.540 97.250 75.800 97.570 ;
        RECT 75.080 93.510 75.340 93.830 ;
        RECT 75.140 91.790 75.280 93.510 ;
        RECT 75.080 91.470 75.340 91.790 ;
        RECT 74.160 83.310 74.420 83.630 ;
        RECT 74.220 82.950 74.360 83.310 ;
        RECT 73.240 82.630 73.500 82.950 ;
        RECT 74.160 82.630 74.420 82.950 ;
        RECT 73.300 79.550 73.440 82.630 ;
        RECT 74.220 82.270 74.360 82.630 ;
        RECT 74.160 81.950 74.420 82.270 ;
        RECT 73.240 79.230 73.500 79.550 ;
        RECT 73.300 77.170 73.440 79.230 ;
        RECT 73.240 76.850 73.500 77.170 ;
        RECT 72.310 74.275 72.590 74.645 ;
        RECT 71.860 73.965 72.120 74.110 ;
        RECT 69.580 73.255 71.460 73.625 ;
        RECT 71.850 73.595 72.130 73.965 ;
        RECT 73.300 72.070 73.440 76.850 ;
        RECT 74.220 73.090 74.360 81.950 ;
        RECT 75.140 80.480 75.280 91.470 ;
        RECT 75.600 88.390 75.740 97.250 ;
        RECT 76.980 94.850 77.120 98.950 ;
        RECT 76.920 94.530 77.180 94.850 ;
        RECT 75.540 88.070 75.800 88.390 ;
        RECT 75.540 80.480 75.800 80.570 ;
        RECT 75.140 80.340 75.800 80.480 ;
        RECT 75.540 80.250 75.800 80.340 ;
        RECT 74.160 72.770 74.420 73.090 ;
        RECT 74.220 72.410 74.360 72.770 ;
        RECT 74.160 72.090 74.420 72.410 ;
        RECT 73.240 71.750 73.500 72.070 ;
        RECT 71.400 71.070 71.660 71.390 ;
        RECT 71.460 69.690 71.600 71.070 ;
        RECT 71.400 69.370 71.660 69.690 ;
        RECT 74.220 69.010 74.360 72.090 ;
        RECT 74.160 68.690 74.420 69.010 ;
        RECT 72.320 68.350 72.580 68.670 ;
        RECT 69.580 67.815 71.460 68.185 ;
        RECT 72.380 64.590 72.520 68.350 ;
        RECT 72.320 64.270 72.580 64.590 ;
        RECT 69.580 62.375 71.460 62.745 ;
        RECT 75.600 60.850 75.740 80.250 ;
        RECT 76.000 79.910 76.260 80.230 ;
        RECT 76.060 77.850 76.200 79.910 ;
        RECT 76.000 77.530 76.260 77.850 ;
        RECT 76.060 66.630 76.200 77.530 ;
        RECT 76.460 71.750 76.720 72.070 ;
        RECT 76.520 70.370 76.660 71.750 ;
        RECT 76.460 70.050 76.720 70.370 ;
        RECT 76.460 68.350 76.720 68.670 ;
        RECT 76.520 67.650 76.660 68.350 ;
        RECT 76.460 67.330 76.720 67.650 ;
        RECT 76.000 66.310 76.260 66.630 ;
        RECT 76.060 64.930 76.200 66.310 ;
        RECT 76.000 64.610 76.260 64.930 ;
        RECT 76.060 62.170 76.200 64.610 ;
        RECT 76.060 62.030 76.660 62.170 ;
        RECT 70.020 60.530 70.280 60.850 ;
        RECT 71.860 60.530 72.120 60.850 ;
        RECT 75.540 60.530 75.800 60.850 ;
        RECT 69.100 60.190 69.360 60.510 ;
        RECT 70.080 58.810 70.220 60.530 ;
        RECT 70.020 58.490 70.280 58.810 ;
        RECT 69.580 56.935 71.460 57.305 ;
        RECT 68.180 55.430 68.440 55.750 ;
        RECT 69.100 55.430 69.360 55.750 ;
        RECT 66.800 54.750 67.060 55.070 ;
        RECT 67.260 54.750 67.520 55.070 ;
        RECT 65.880 53.730 66.140 54.050 ;
        RECT 64.960 52.710 65.220 53.030 ;
        RECT 65.420 52.710 65.680 53.030 ;
        RECT 65.020 52.260 65.160 52.710 ;
        RECT 66.330 52.515 66.610 52.885 ;
        RECT 66.400 52.350 66.540 52.515 ;
        RECT 65.020 52.120 65.620 52.260 ;
        RECT 65.480 50.310 65.620 52.120 ;
        RECT 66.340 52.030 66.600 52.350 ;
        RECT 65.880 50.330 66.140 50.650 ;
        RECT 65.420 49.990 65.680 50.310 ;
        RECT 65.480 47.250 65.620 49.990 ;
        RECT 65.940 49.630 66.080 50.330 ;
        RECT 66.340 49.990 66.600 50.310 ;
        RECT 65.880 49.310 66.140 49.630 ;
        RECT 65.940 47.500 66.080 49.310 ;
        RECT 66.400 48.010 66.540 49.990 ;
        RECT 66.860 48.610 67.000 54.750 ;
        RECT 67.320 49.970 67.460 54.750 ;
        RECT 67.710 51.155 67.990 51.525 ;
        RECT 67.720 51.010 67.980 51.155 ;
        RECT 68.240 50.650 68.380 55.430 ;
        RECT 69.160 53.370 69.300 55.430 ;
        RECT 71.920 54.050 72.060 60.530 ;
        RECT 72.320 60.190 72.580 60.510 ;
        RECT 72.380 56.090 72.520 60.190 ;
        RECT 75.080 56.110 75.340 56.430 ;
        RECT 72.320 55.770 72.580 56.090 ;
        RECT 71.860 53.730 72.120 54.050 ;
        RECT 74.620 53.730 74.880 54.050 ;
        RECT 69.100 53.050 69.360 53.370 ;
        RECT 71.860 53.050 72.120 53.370 ;
        RECT 69.160 51.330 69.300 53.050 ;
        RECT 69.580 51.495 71.460 51.865 ;
        RECT 69.100 51.010 69.360 51.330 ;
        RECT 68.640 50.845 68.900 50.990 ;
        RECT 68.180 50.330 68.440 50.650 ;
        RECT 68.630 50.475 68.910 50.845 ;
        RECT 69.160 50.730 69.300 51.010 ;
        RECT 69.160 50.590 69.760 50.730 ;
        RECT 67.260 49.650 67.520 49.970 ;
        RECT 66.800 48.290 67.060 48.610 ;
        RECT 66.400 47.870 67.460 48.010 ;
        RECT 67.320 47.590 67.460 47.870 ;
        RECT 66.340 47.500 66.600 47.590 ;
        RECT 65.940 47.360 66.600 47.500 ;
        RECT 65.420 46.930 65.680 47.250 ;
        RECT 65.940 43.170 66.080 47.360 ;
        RECT 66.340 47.270 66.600 47.360 ;
        RECT 67.260 47.270 67.520 47.590 ;
        RECT 67.320 44.530 67.460 47.270 ;
        RECT 67.260 44.210 67.520 44.530 ;
        RECT 64.500 42.850 64.760 43.170 ;
        RECT 65.880 42.850 66.140 43.170 ;
        RECT 63.580 41.830 63.840 42.150 ;
        RECT 63.640 40.450 63.780 41.830 ;
        RECT 63.580 40.130 63.840 40.450 ;
        RECT 65.420 37.410 65.680 37.730 ;
        RECT 64.040 37.070 64.300 37.390 ;
        RECT 63.580 34.920 63.840 35.010 ;
        RECT 63.180 34.780 63.840 34.920 ;
        RECT 63.580 34.690 63.840 34.780 ;
        RECT 63.640 33.310 63.780 34.690 ;
        RECT 64.100 34.670 64.240 37.070 ;
        RECT 64.960 36.730 65.220 37.050 ;
        RECT 64.040 34.350 64.300 34.670 ;
        RECT 64.100 33.310 64.240 34.350 ;
        RECT 65.020 33.990 65.160 36.730 ;
        RECT 65.480 33.990 65.620 37.410 ;
        RECT 65.940 37.050 66.080 42.850 ;
        RECT 65.880 36.730 66.140 37.050 ;
        RECT 68.240 36.030 68.380 50.330 ;
        RECT 69.620 50.310 69.760 50.590 ;
        RECT 69.560 49.990 69.820 50.310 ;
        RECT 70.480 49.990 70.740 50.310 ;
        RECT 69.100 49.650 69.360 49.970 ;
        RECT 69.160 48.010 69.300 49.650 ;
        RECT 68.700 47.930 69.300 48.010 ;
        RECT 68.640 47.870 69.300 47.930 ;
        RECT 68.640 47.610 68.900 47.870 ;
        RECT 68.700 45.890 68.840 47.610 ;
        RECT 70.540 47.250 70.680 49.990 ;
        RECT 71.920 49.630 72.060 53.050 ;
        RECT 74.680 49.630 74.820 53.730 ;
        RECT 75.140 52.350 75.280 56.110 ;
        RECT 76.520 55.410 76.660 62.030 ;
        RECT 77.440 59.150 77.580 107.790 ;
        RECT 78.820 104.710 78.960 108.220 ;
        RECT 79.680 108.130 79.940 108.220 ;
        RECT 80.600 107.110 80.860 107.430 ;
        RECT 80.660 105.390 80.800 107.110 ;
        RECT 80.600 105.070 80.860 105.390 ;
        RECT 82.960 104.710 83.100 111.870 ;
        RECT 83.420 111.170 83.560 123.430 ;
        RECT 88.020 122.050 88.160 123.430 ;
        RECT 89.860 122.050 90.000 123.770 ;
        RECT 92.620 123.750 92.760 138.990 ;
        RECT 99.580 127.655 101.460 128.025 ;
        RECT 93.020 123.770 93.280 124.090 ;
        RECT 92.560 123.430 92.820 123.750 ;
        RECT 93.080 122.050 93.220 123.770 ;
        RECT 93.480 123.430 93.740 123.750 ;
        RECT 87.960 121.730 88.220 122.050 ;
        RECT 89.800 121.730 90.060 122.050 ;
        RECT 93.020 121.730 93.280 122.050 ;
        RECT 89.800 120.710 90.060 121.030 ;
        RECT 92.560 120.710 92.820 121.030 ;
        RECT 84.580 119.495 86.460 119.865 ;
        RECT 83.820 114.590 84.080 114.910 ;
        RECT 83.880 113.890 84.020 114.590 ;
        RECT 84.580 114.055 86.460 114.425 ;
        RECT 83.820 113.570 84.080 113.890 ;
        RECT 86.580 113.230 86.840 113.550 ;
        RECT 85.660 112.550 85.920 112.870 ;
        RECT 83.360 110.850 83.620 111.170 ;
        RECT 83.420 107.680 83.560 110.850 ;
        RECT 85.720 110.490 85.860 112.550 ;
        RECT 85.660 110.170 85.920 110.490 ;
        RECT 84.580 108.615 86.460 108.985 ;
        RECT 83.820 107.680 84.080 107.770 ;
        RECT 83.420 107.540 84.080 107.680 ;
        RECT 83.820 107.450 84.080 107.540 ;
        RECT 83.360 106.770 83.620 107.090 ;
        RECT 78.760 104.390 79.020 104.710 ;
        RECT 79.680 104.390 79.940 104.710 ;
        RECT 82.900 104.390 83.160 104.710 ;
        RECT 79.740 101.990 79.880 104.390 ;
        RECT 80.600 103.710 80.860 104.030 ;
        RECT 79.680 101.670 79.940 101.990 ;
        RECT 79.220 95.550 79.480 95.870 ;
        RECT 78.760 93.510 79.020 93.830 ;
        RECT 78.300 88.070 78.560 88.390 ;
        RECT 78.360 86.350 78.500 88.070 ;
        RECT 78.300 86.030 78.560 86.350 ;
        RECT 77.840 79.230 78.100 79.550 ;
        RECT 77.900 77.850 78.040 79.230 ;
        RECT 77.840 77.530 78.100 77.850 ;
        RECT 78.820 75.325 78.960 93.510 ;
        RECT 79.280 93.490 79.420 95.550 ;
        RECT 79.220 93.170 79.480 93.490 ;
        RECT 80.140 90.110 80.400 90.430 ;
        RECT 80.200 88.730 80.340 90.110 ;
        RECT 80.140 88.410 80.400 88.730 ;
        RECT 79.220 80.250 79.480 80.570 ;
        RECT 79.280 78.530 79.420 80.250 ;
        RECT 79.220 78.210 79.480 78.530 ;
        RECT 78.750 74.955 79.030 75.325 ;
        RECT 78.760 74.810 79.020 74.955 ;
        RECT 78.300 74.470 78.560 74.790 ;
        RECT 78.360 71.390 78.500 74.470 ;
        RECT 80.660 74.110 80.800 103.710 ;
        RECT 83.420 102.330 83.560 106.770 ;
        RECT 83.880 105.050 84.020 107.450 ;
        RECT 86.640 105.730 86.780 113.230 ;
        RECT 87.040 112.890 87.300 113.210 ;
        RECT 86.580 105.410 86.840 105.730 ;
        RECT 83.820 104.730 84.080 105.050 ;
        RECT 86.640 104.030 86.780 105.410 ;
        RECT 86.580 103.710 86.840 104.030 ;
        RECT 84.580 103.175 86.460 103.545 ;
        RECT 87.100 103.010 87.240 112.890 ;
        RECT 87.960 112.550 88.220 112.870 ;
        RECT 88.020 110.830 88.160 112.550 ;
        RECT 89.340 111.870 89.600 112.190 ;
        RECT 87.960 110.510 88.220 110.830 ;
        RECT 88.020 107.430 88.160 110.510 ;
        RECT 87.960 107.110 88.220 107.430 ;
        RECT 87.040 102.690 87.300 103.010 ;
        RECT 87.500 102.690 87.760 103.010 ;
        RECT 83.360 102.010 83.620 102.330 ;
        RECT 87.560 101.990 87.700 102.690 ;
        RECT 87.500 101.670 87.760 101.990 ;
        RECT 88.020 101.900 88.160 107.110 ;
        RECT 89.400 104.370 89.540 111.870 ;
        RECT 89.860 105.730 90.000 120.710 ;
        RECT 92.620 118.990 92.760 120.710 ;
        RECT 93.540 119.330 93.680 123.430 ;
        RECT 96.240 122.750 96.500 123.070 ;
        RECT 96.300 121.030 96.440 122.750 ;
        RECT 99.580 122.215 101.460 122.585 ;
        RECT 96.240 120.710 96.500 121.030 ;
        RECT 93.480 119.010 93.740 119.330 ;
        RECT 92.560 118.670 92.820 118.990 ;
        RECT 90.720 118.330 90.980 118.650 ;
        RECT 91.180 118.330 91.440 118.650 ;
        RECT 90.260 109.490 90.520 109.810 ;
        RECT 89.800 105.410 90.060 105.730 ;
        RECT 89.800 104.730 90.060 105.050 ;
        RECT 89.340 104.050 89.600 104.370 ;
        RECT 88.880 103.710 89.140 104.030 ;
        RECT 88.940 102.670 89.080 103.710 ;
        RECT 88.880 102.350 89.140 102.670 ;
        RECT 89.340 101.900 89.600 101.990 ;
        RECT 88.020 101.760 89.600 101.900 ;
        RECT 89.340 101.670 89.600 101.760 ;
        RECT 84.580 97.735 86.460 98.105 ;
        RECT 84.280 94.190 84.540 94.510 ;
        RECT 84.340 93.830 84.480 94.190 ;
        RECT 86.180 94.110 87.240 94.250 ;
        RECT 84.280 93.570 84.540 93.830 ;
        RECT 82.960 93.510 84.540 93.570 ;
        RECT 82.960 93.430 84.480 93.510 ;
        RECT 86.180 93.490 86.320 94.110 ;
        RECT 86.580 93.510 86.840 93.830 ;
        RECT 82.960 90.770 83.100 93.430 ;
        RECT 86.120 93.170 86.380 93.490 ;
        RECT 83.820 92.830 84.080 93.150 ;
        RECT 83.880 92.130 84.020 92.830 ;
        RECT 84.580 92.295 86.460 92.665 ;
        RECT 83.820 91.810 84.080 92.130 ;
        RECT 85.660 91.810 85.920 92.130 ;
        RECT 83.820 91.130 84.080 91.450 ;
        RECT 82.900 90.450 83.160 90.770 ;
        RECT 81.980 88.410 82.240 88.730 ;
        RECT 82.040 80.570 82.180 88.410 ;
        RECT 81.980 80.250 82.240 80.570 ;
        RECT 81.520 79.230 81.780 79.550 ;
        RECT 81.580 77.170 81.720 79.230 ;
        RECT 81.520 76.850 81.780 77.170 ;
        RECT 81.060 74.810 81.320 75.130 ;
        RECT 81.120 74.450 81.260 74.810 ;
        RECT 81.060 74.130 81.320 74.450 ;
        RECT 80.600 73.790 80.860 74.110 ;
        RECT 78.300 71.070 78.560 71.390 ;
        RECT 78.360 69.690 78.500 71.070 ;
        RECT 82.040 69.690 82.180 80.250 ;
        RECT 82.960 80.230 83.100 90.450 ;
        RECT 83.360 85.690 83.620 86.010 ;
        RECT 83.420 83.970 83.560 85.690 ;
        RECT 83.880 84.990 84.020 91.130 ;
        RECT 85.720 89.070 85.860 91.810 ;
        RECT 86.640 91.530 86.780 93.510 ;
        RECT 87.100 92.130 87.240 94.110 ;
        RECT 88.420 93.510 88.680 93.830 ;
        RECT 88.480 92.130 88.620 93.510 ;
        RECT 87.040 91.810 87.300 92.130 ;
        RECT 88.420 91.810 88.680 92.130 ;
        RECT 86.180 91.450 86.780 91.530 ;
        RECT 86.120 91.390 86.780 91.450 ;
        RECT 86.120 91.130 86.380 91.390 ;
        RECT 86.580 90.790 86.840 91.110 ;
        RECT 85.660 88.750 85.920 89.070 ;
        RECT 84.580 86.855 86.460 87.225 ;
        RECT 83.820 84.670 84.080 84.990 ;
        RECT 83.360 83.650 83.620 83.970 ;
        RECT 83.880 83.290 84.020 84.670 ;
        RECT 83.820 82.970 84.080 83.290 ;
        RECT 86.640 82.950 86.780 90.790 ;
        RECT 86.580 82.630 86.840 82.950 ;
        RECT 83.820 81.950 84.080 82.270 ;
        RECT 83.880 81.250 84.020 81.950 ;
        RECT 84.580 81.415 86.460 81.785 ;
        RECT 83.820 80.930 84.080 81.250 ;
        RECT 83.360 80.250 83.620 80.570 ;
        RECT 82.900 79.910 83.160 80.230 ;
        RECT 82.960 75.470 83.100 79.910 ;
        RECT 82.900 75.150 83.160 75.470 ;
        RECT 83.420 75.325 83.560 80.250 ;
        RECT 83.880 78.190 84.020 80.930 ;
        RECT 86.580 80.480 86.840 80.570 ;
        RECT 87.100 80.480 87.240 91.810 ;
        RECT 88.880 82.630 89.140 82.950 ;
        RECT 86.580 80.340 87.240 80.480 ;
        RECT 86.580 80.250 86.840 80.340 ;
        RECT 83.820 77.870 84.080 78.190 ;
        RECT 83.820 76.510 84.080 76.830 ;
        RECT 83.350 74.955 83.630 75.325 ;
        RECT 83.880 75.130 84.020 76.510 ;
        RECT 84.580 75.975 86.460 76.345 ;
        RECT 83.360 74.810 83.620 74.955 ;
        RECT 83.820 74.810 84.080 75.130 ;
        RECT 83.880 70.370 84.020 74.810 ;
        RECT 86.640 74.790 86.780 80.250 ;
        RECT 88.420 79.910 88.680 80.230 ;
        RECT 86.580 74.470 86.840 74.790 ;
        RECT 87.500 74.470 87.760 74.790 ;
        RECT 84.580 70.535 86.460 70.905 ;
        RECT 82.440 70.050 82.700 70.370 ;
        RECT 83.820 70.050 84.080 70.370 ;
        RECT 78.300 69.370 78.560 69.690 ;
        RECT 81.980 69.370 82.240 69.690 ;
        RECT 78.360 64.930 78.500 69.370 ;
        RECT 80.600 68.350 80.860 68.670 ;
        RECT 80.660 66.290 80.800 68.350 ;
        RECT 82.040 66.970 82.180 69.370 ;
        RECT 82.500 67.650 82.640 70.050 ;
        RECT 82.440 67.330 82.700 67.650 ;
        RECT 81.980 66.650 82.240 66.970 ;
        RECT 80.600 65.970 80.860 66.290 ;
        RECT 78.300 64.610 78.560 64.930 ;
        RECT 82.040 64.250 82.180 66.650 ;
        RECT 83.360 66.310 83.620 66.630 ;
        RECT 81.980 63.930 82.240 64.250 ;
        RECT 82.440 60.870 82.700 61.190 ;
        RECT 77.380 58.830 77.640 59.150 ;
        RECT 80.140 58.830 80.400 59.150 ;
        RECT 80.200 55.750 80.340 58.830 ;
        RECT 78.760 55.430 79.020 55.750 ;
        RECT 80.140 55.490 80.400 55.750 ;
        RECT 80.140 55.430 80.800 55.490 ;
        RECT 76.460 55.090 76.720 55.410 ;
        RECT 75.540 54.750 75.800 55.070 ;
        RECT 75.080 52.030 75.340 52.350 ;
        RECT 75.600 50.990 75.740 54.750 ;
        RECT 76.520 53.710 76.660 55.090 ;
        RECT 76.460 53.390 76.720 53.710 ;
        RECT 75.540 50.670 75.800 50.990 ;
        RECT 71.860 49.310 72.120 49.630 ;
        RECT 74.620 49.310 74.880 49.630 ;
        RECT 71.920 48.270 72.060 49.310 ;
        RECT 71.860 47.950 72.120 48.270 ;
        RECT 70.480 46.930 70.740 47.250 ;
        RECT 74.680 46.910 74.820 49.310 ;
        RECT 74.620 46.590 74.880 46.910 ;
        RECT 69.580 46.055 71.460 46.425 ;
        RECT 68.640 45.570 68.900 45.890 ;
        RECT 68.700 37.390 68.840 45.570 ;
        RECT 75.080 43.870 75.340 44.190 ;
        RECT 75.140 42.150 75.280 43.870 ;
        RECT 76.520 42.830 76.660 53.390 ;
        RECT 77.370 52.515 77.650 52.885 ;
        RECT 77.440 50.310 77.580 52.515 ;
        RECT 78.820 51.330 78.960 55.430 ;
        RECT 80.200 55.350 80.800 55.430 ;
        RECT 82.500 55.410 82.640 60.870 ;
        RECT 83.420 58.810 83.560 66.310 ;
        RECT 84.580 65.095 86.460 65.465 ;
        RECT 86.580 62.910 86.840 63.230 ;
        RECT 86.640 61.530 86.780 62.910 ;
        RECT 86.580 61.210 86.840 61.530 ;
        RECT 84.580 59.655 86.460 60.025 ;
        RECT 83.360 58.490 83.620 58.810 ;
        RECT 80.140 54.750 80.400 55.070 ;
        RECT 80.200 53.710 80.340 54.750 ;
        RECT 80.140 53.390 80.400 53.710 ;
        RECT 78.760 51.010 79.020 51.330 ;
        RECT 77.380 49.990 77.640 50.310 ;
        RECT 79.680 46.590 79.940 46.910 ;
        RECT 79.740 44.870 79.880 46.590 ;
        RECT 80.660 44.870 80.800 55.350 ;
        RECT 82.440 55.090 82.700 55.410 ;
        RECT 82.500 53.710 82.640 55.090 ;
        RECT 84.580 54.215 86.460 54.585 ;
        RECT 82.440 53.390 82.700 53.710 ;
        RECT 85.660 52.710 85.920 53.030 ;
        RECT 82.900 52.030 83.160 52.350 ;
        RECT 82.440 49.650 82.700 49.970 ;
        RECT 82.500 47.500 82.640 49.650 ;
        RECT 82.960 49.630 83.100 52.030 ;
        RECT 83.360 50.670 83.620 50.990 ;
        RECT 82.900 49.310 83.160 49.630 ;
        RECT 82.960 48.270 83.100 49.310 ;
        RECT 82.900 47.950 83.160 48.270 ;
        RECT 82.900 47.500 83.160 47.590 ;
        RECT 82.500 47.360 83.160 47.500 ;
        RECT 82.900 47.270 83.160 47.360 ;
        RECT 79.680 44.550 79.940 44.870 ;
        RECT 80.600 44.550 80.860 44.870 ;
        RECT 82.900 44.550 83.160 44.870 ;
        RECT 80.600 43.870 80.860 44.190 ;
        RECT 76.460 42.740 76.720 42.830 ;
        RECT 76.460 42.600 77.120 42.740 ;
        RECT 76.460 42.510 76.720 42.600 ;
        RECT 75.080 41.830 75.340 42.150 ;
        RECT 69.580 40.615 71.460 40.985 ;
        RECT 76.980 39.770 77.120 42.600 ;
        RECT 80.660 42.490 80.800 43.870 ;
        RECT 80.600 42.170 80.860 42.490 ;
        RECT 76.920 39.450 77.180 39.770 ;
        RECT 68.640 37.070 68.900 37.390 ;
        RECT 68.640 36.390 68.900 36.710 ;
        RECT 75.080 36.390 75.340 36.710 ;
        RECT 66.800 35.710 67.060 36.030 ;
        RECT 68.180 35.710 68.440 36.030 ;
        RECT 66.860 34.330 67.000 35.710 ;
        RECT 66.800 34.010 67.060 34.330 ;
        RECT 67.260 34.010 67.520 34.330 ;
        RECT 64.960 33.670 65.220 33.990 ;
        RECT 65.420 33.670 65.680 33.990 ;
        RECT 63.580 32.990 63.840 33.310 ;
        RECT 64.040 32.990 64.300 33.310 ;
        RECT 63.640 32.290 63.780 32.990 ;
        RECT 63.580 31.970 63.840 32.290 ;
        RECT 67.320 31.950 67.460 34.010 ;
        RECT 67.260 31.630 67.520 31.950 ;
        RECT 62.660 31.290 62.920 31.610 ;
        RECT 59.900 30.950 60.160 31.270 ;
        RECT 62.720 29.570 62.860 31.290 ;
        RECT 62.660 29.250 62.920 29.570 ;
        RECT 59.440 28.230 59.700 28.550 ;
        RECT 57.140 27.550 57.400 27.870 ;
        RECT 47.020 26.530 47.280 26.850 ;
        RECT 56.680 26.530 56.940 26.850 ;
        RECT 45.180 26.190 45.440 26.510 ;
        RECT 57.200 26.170 57.340 27.550 ;
        RECT 59.500 26.170 59.640 28.230 ;
        RECT 37.820 25.850 38.080 26.170 ;
        RECT 40.580 25.850 40.840 26.170 ;
        RECT 57.140 25.850 57.400 26.170 ;
        RECT 59.440 25.850 59.700 26.170 ;
        RECT 68.240 25.490 68.380 35.710 ;
        RECT 68.700 35.010 68.840 36.390 ;
        RECT 71.860 35.710 72.120 36.030 ;
        RECT 69.580 35.175 71.460 35.545 ;
        RECT 68.640 34.690 68.900 35.010 ;
        RECT 69.100 33.670 69.360 33.990 ;
        RECT 69.160 28.970 69.300 33.670 ;
        RECT 71.920 33.650 72.060 35.710 ;
        RECT 71.860 33.330 72.120 33.650 ;
        RECT 75.140 31.950 75.280 36.390 ;
        RECT 71.860 31.630 72.120 31.950 ;
        RECT 75.080 31.630 75.340 31.950 ;
        RECT 69.580 29.735 71.460 30.105 ;
        RECT 71.920 29.570 72.060 31.630 ;
        RECT 76.980 30.590 77.120 39.450 ;
        RECT 82.440 38.770 82.700 39.090 ;
        RECT 82.500 37.730 82.640 38.770 ;
        RECT 82.440 37.410 82.700 37.730 ;
        RECT 82.960 37.390 83.100 44.550 ;
        RECT 82.900 37.070 83.160 37.390 ;
        RECT 82.960 31.610 83.100 37.070 ;
        RECT 83.420 32.290 83.560 50.670 ;
        RECT 85.720 50.310 85.860 52.710 ;
        RECT 87.560 51.330 87.700 74.470 ;
        RECT 87.960 65.630 88.220 65.950 ;
        RECT 88.020 64.250 88.160 65.630 ;
        RECT 87.960 63.930 88.220 64.250 ;
        RECT 87.500 51.010 87.760 51.330 ;
        RECT 88.480 50.650 88.620 79.910 ;
        RECT 88.940 77.850 89.080 82.630 ;
        RECT 89.860 79.550 90.000 104.730 ;
        RECT 90.320 104.710 90.460 109.490 ;
        RECT 90.260 104.565 90.520 104.710 ;
        RECT 90.250 104.195 90.530 104.565 ;
        RECT 90.780 91.530 90.920 118.330 ;
        RECT 91.240 94.850 91.380 118.330 ;
        RECT 93.020 114.930 93.280 115.250 ;
        RECT 92.100 113.570 92.360 113.890 ;
        RECT 92.160 109.470 92.300 113.570 ;
        RECT 92.560 112.890 92.820 113.210 ;
        RECT 92.620 111.170 92.760 112.890 ;
        RECT 92.560 110.850 92.820 111.170 ;
        RECT 92.100 109.150 92.360 109.470 ;
        RECT 92.160 104.710 92.300 109.150 ;
        RECT 92.560 105.410 92.820 105.730 ;
        RECT 91.640 104.390 91.900 104.710 ;
        RECT 92.100 104.390 92.360 104.710 ;
        RECT 91.700 102.670 91.840 104.390 ;
        RECT 91.640 102.350 91.900 102.670 ;
        RECT 92.100 102.010 92.360 102.330 ;
        RECT 91.640 100.990 91.900 101.310 ;
        RECT 91.180 94.530 91.440 94.850 ;
        RECT 90.320 91.390 90.920 91.530 ;
        RECT 90.320 81.250 90.460 91.390 ;
        RECT 90.720 90.790 90.980 91.110 ;
        RECT 90.260 80.930 90.520 81.250 ;
        RECT 89.800 79.230 90.060 79.550 ;
        RECT 88.880 77.530 89.140 77.850 ;
        RECT 90.260 75.150 90.520 75.470 ;
        RECT 89.340 74.810 89.600 75.130 ;
        RECT 88.870 74.275 89.150 74.645 ;
        RECT 88.880 74.130 89.140 74.275 ;
        RECT 88.880 71.750 89.140 72.070 ;
        RECT 88.940 69.010 89.080 71.750 ;
        RECT 89.400 70.370 89.540 74.810 ;
        RECT 89.800 71.750 90.060 72.070 ;
        RECT 89.340 70.050 89.600 70.370 ;
        RECT 88.880 68.690 89.140 69.010 ;
        RECT 89.860 66.970 90.000 71.750 ;
        RECT 90.320 70.030 90.460 75.150 ;
        RECT 90.260 69.710 90.520 70.030 ;
        RECT 89.800 66.650 90.060 66.970 ;
        RECT 88.880 63.930 89.140 64.250 ;
        RECT 88.940 62.210 89.080 63.930 ;
        RECT 88.880 61.890 89.140 62.210 ;
        RECT 90.260 60.530 90.520 60.850 ;
        RECT 90.320 59.490 90.460 60.530 ;
        RECT 90.260 59.170 90.520 59.490 ;
        RECT 90.780 51.330 90.920 90.790 ;
        RECT 91.700 90.430 91.840 100.990 ;
        RECT 91.640 90.110 91.900 90.430 ;
        RECT 92.160 87.450 92.300 102.010 ;
        RECT 92.620 92.130 92.760 105.410 ;
        RECT 92.560 91.810 92.820 92.130 ;
        RECT 91.240 87.310 92.300 87.450 ;
        RECT 91.240 74.110 91.380 87.310 ;
        RECT 93.080 75.810 93.220 114.930 ;
        RECT 96.300 112.870 96.440 120.710 ;
        RECT 97.620 120.370 97.880 120.690 ;
        RECT 99.920 120.370 100.180 120.690 ;
        RECT 97.680 119.330 97.820 120.370 ;
        RECT 99.980 119.330 100.120 120.370 ;
        RECT 101.820 120.350 101.960 138.990 ;
        RECT 105.900 123.770 106.160 124.090 ;
        RECT 103.140 123.090 103.400 123.410 ;
        RECT 101.760 120.030 102.020 120.350 ;
        RECT 103.200 119.330 103.340 123.090 ;
        RECT 105.960 122.050 106.100 123.770 ;
        RECT 106.420 123.750 106.560 138.395 ;
        RECT 111.880 126.150 112.140 126.470 ;
        RECT 111.940 124.770 112.080 126.150 ;
        RECT 113.720 125.810 113.980 126.130 ;
        RECT 111.880 124.450 112.140 124.770 ;
        RECT 106.360 123.430 106.620 123.750 ;
        RECT 105.900 121.730 106.160 122.050 ;
        RECT 111.940 121.370 112.080 124.450 ;
        RECT 108.660 121.050 108.920 121.370 ;
        RECT 111.880 121.050 112.140 121.370 ;
        RECT 108.720 120.770 108.860 121.050 ;
        RECT 106.820 120.370 107.080 120.690 ;
        RECT 108.720 120.630 109.320 120.770 ;
        RECT 106.880 119.330 107.020 120.370 ;
        RECT 97.620 119.010 97.880 119.330 ;
        RECT 99.920 119.010 100.180 119.330 ;
        RECT 103.140 119.010 103.400 119.330 ;
        RECT 106.820 119.010 107.080 119.330 ;
        RECT 98.540 118.330 98.800 118.650 ;
        RECT 103.140 118.330 103.400 118.650 ;
        RECT 105.900 118.330 106.160 118.650 ;
        RECT 96.240 112.550 96.500 112.870 ;
        RECT 97.160 112.550 97.420 112.870 ;
        RECT 93.480 109.150 93.740 109.470 ;
        RECT 93.540 107.090 93.680 109.150 ;
        RECT 93.480 106.770 93.740 107.090 ;
        RECT 93.540 102.330 93.680 106.770 ;
        RECT 96.300 102.670 96.440 112.550 ;
        RECT 96.700 111.870 96.960 112.190 ;
        RECT 96.760 108.110 96.900 111.870 ;
        RECT 97.220 111.170 97.360 112.550 ;
        RECT 97.160 110.850 97.420 111.170 ;
        RECT 98.080 110.170 98.340 110.490 ;
        RECT 98.140 109.470 98.280 110.170 ;
        RECT 98.080 109.150 98.340 109.470 ;
        RECT 96.700 107.790 96.960 108.110 ;
        RECT 96.240 102.350 96.500 102.670 ;
        RECT 93.480 102.010 93.740 102.330 ;
        RECT 95.320 102.010 95.580 102.330 ;
        RECT 94.400 100.990 94.660 101.310 ;
        RECT 94.460 94.850 94.600 100.990 ;
        RECT 95.380 99.270 95.520 102.010 ;
        RECT 98.140 101.990 98.280 109.150 ;
        RECT 98.080 101.670 98.340 101.990 ;
        RECT 97.160 101.330 97.420 101.650 ;
        RECT 95.320 98.950 95.580 99.270 ;
        RECT 97.220 98.590 97.360 101.330 ;
        RECT 97.620 99.290 97.880 99.610 ;
        RECT 96.700 98.270 96.960 98.590 ;
        RECT 97.160 98.270 97.420 98.590 ;
        RECT 96.760 94.850 96.900 98.270 ;
        RECT 97.220 96.890 97.360 98.270 ;
        RECT 97.680 97.230 97.820 99.290 ;
        RECT 97.620 96.910 97.880 97.230 ;
        RECT 97.160 96.570 97.420 96.890 ;
        RECT 98.600 94.850 98.740 118.330 ;
        RECT 99.580 116.775 101.460 117.145 ;
        RECT 101.760 113.570 102.020 113.890 ;
        RECT 99.580 111.335 101.460 111.705 ;
        RECT 101.820 107.770 101.960 113.570 ;
        RECT 102.220 113.230 102.480 113.550 ;
        RECT 102.280 110.490 102.420 113.230 ;
        RECT 102.220 110.170 102.480 110.490 ;
        RECT 102.680 109.830 102.940 110.150 ;
        RECT 101.760 107.450 102.020 107.770 ;
        RECT 99.580 105.895 101.460 106.265 ;
        RECT 102.740 104.710 102.880 109.830 ;
        RECT 102.680 104.390 102.940 104.710 ;
        RECT 100.840 103.710 101.100 104.030 ;
        RECT 100.900 102.670 101.040 103.710 ;
        RECT 102.680 102.690 102.940 103.010 ;
        RECT 100.840 102.350 101.100 102.670 ;
        RECT 99.000 101.670 99.260 101.990 ;
        RECT 99.060 100.290 99.200 101.670 ;
        RECT 99.580 100.455 101.460 100.825 ;
        RECT 99.000 99.970 99.260 100.290 ;
        RECT 102.740 98.590 102.880 102.690 ;
        RECT 102.680 98.270 102.940 98.590 ;
        RECT 102.220 96.910 102.480 97.230 ;
        RECT 101.760 96.570 102.020 96.890 ;
        RECT 99.580 95.015 101.460 95.385 ;
        RECT 94.400 94.530 94.660 94.850 ;
        RECT 96.700 94.530 96.960 94.850 ;
        RECT 98.540 94.530 98.800 94.850 ;
        RECT 99.000 93.850 99.260 94.170 ;
        RECT 93.480 93.510 93.740 93.830 ;
        RECT 94.400 93.510 94.660 93.830 ;
        RECT 93.540 75.810 93.680 93.510 ;
        RECT 93.940 80.250 94.200 80.570 ;
        RECT 93.020 75.490 93.280 75.810 ;
        RECT 93.480 75.490 93.740 75.810 ;
        RECT 92.100 74.810 92.360 75.130 ;
        RECT 91.640 74.470 91.900 74.790 ;
        RECT 91.180 73.790 91.440 74.110 ;
        RECT 91.180 71.925 91.440 72.070 ;
        RECT 91.170 71.555 91.450 71.925 ;
        RECT 91.240 69.690 91.380 71.555 ;
        RECT 91.180 69.370 91.440 69.690 ;
        RECT 90.720 51.010 90.980 51.330 ;
        RECT 89.800 50.670 90.060 50.990 ;
        RECT 88.420 50.330 88.680 50.650 ;
        RECT 83.820 49.990 84.080 50.310 ;
        RECT 85.660 49.990 85.920 50.310 ;
        RECT 88.880 49.990 89.140 50.310 ;
        RECT 83.880 48.610 84.020 49.990 ;
        RECT 86.580 49.310 86.840 49.630 ;
        RECT 84.580 48.775 86.460 49.145 ;
        RECT 83.820 48.290 84.080 48.610 ;
        RECT 86.640 48.270 86.780 49.310 ;
        RECT 88.940 48.610 89.080 49.990 ;
        RECT 88.880 48.290 89.140 48.610 ;
        RECT 86.580 47.950 86.840 48.270 ;
        RECT 84.580 43.335 86.460 43.705 ;
        RECT 86.640 43.170 86.780 47.950 ;
        RECT 88.420 47.610 88.680 47.930 ;
        RECT 87.040 47.270 87.300 47.590 ;
        RECT 87.100 44.530 87.240 47.270 ;
        RECT 87.040 44.210 87.300 44.530 ;
        RECT 86.580 42.850 86.840 43.170 ;
        RECT 87.100 42.150 87.240 44.210 ;
        RECT 87.040 41.830 87.300 42.150 ;
        RECT 83.820 41.150 84.080 41.470 ;
        RECT 83.880 37.050 84.020 41.150 ;
        RECT 87.500 38.770 87.760 39.090 ;
        RECT 84.580 37.895 86.460 38.265 ;
        RECT 87.560 37.730 87.700 38.770 ;
        RECT 87.500 37.410 87.760 37.730 ;
        RECT 83.820 36.730 84.080 37.050 ;
        RECT 88.480 34.330 88.620 47.610 ;
        RECT 89.860 47.590 90.000 50.670 ;
        RECT 90.720 49.990 90.980 50.310 ;
        RECT 90.780 48.010 90.920 49.990 ;
        RECT 91.700 48.270 91.840 74.470 ;
        RECT 92.160 73.090 92.300 74.810 ;
        RECT 92.560 74.470 92.820 74.790 ;
        RECT 92.100 72.770 92.360 73.090 ;
        RECT 92.620 71.730 92.760 74.470 ;
        RECT 92.560 71.410 92.820 71.730 ;
        RECT 92.620 69.690 92.760 71.410 ;
        RECT 94.000 70.370 94.140 80.250 ;
        RECT 93.940 70.050 94.200 70.370 ;
        RECT 92.560 69.370 92.820 69.690 ;
        RECT 93.480 69.370 93.740 69.690 ;
        RECT 93.940 69.370 94.200 69.690 ;
        RECT 92.560 66.650 92.820 66.970 ;
        RECT 93.020 66.650 93.280 66.970 ;
        RECT 92.620 64.930 92.760 66.650 ;
        RECT 92.560 64.610 92.820 64.930 ;
        RECT 92.620 62.210 92.760 64.610 ;
        RECT 93.080 63.910 93.220 66.650 ;
        RECT 93.540 64.590 93.680 69.370 ;
        RECT 94.000 69.010 94.140 69.370 ;
        RECT 93.940 68.690 94.200 69.010 ;
        RECT 93.480 64.270 93.740 64.590 ;
        RECT 93.020 63.590 93.280 63.910 ;
        RECT 92.560 61.890 92.820 62.210 ;
        RECT 92.090 55.235 92.370 55.605 ;
        RECT 93.020 55.430 93.280 55.750 ;
        RECT 92.160 53.710 92.300 55.235 ;
        RECT 92.560 54.750 92.820 55.070 ;
        RECT 92.100 53.390 92.360 53.710 ;
        RECT 92.620 52.940 92.760 54.750 ;
        RECT 92.160 52.800 92.760 52.940 ;
        RECT 92.160 50.310 92.300 52.800 ;
        RECT 93.080 50.310 93.220 55.430 ;
        RECT 92.100 49.990 92.360 50.310 ;
        RECT 93.020 50.050 93.280 50.310 ;
        RECT 92.620 49.990 93.280 50.050 ;
        RECT 92.160 48.610 92.300 49.990 ;
        RECT 92.620 49.910 93.220 49.990 ;
        RECT 92.100 48.290 92.360 48.610 ;
        RECT 90.780 47.930 91.380 48.010 ;
        RECT 91.640 47.950 91.900 48.270 ;
        RECT 92.620 47.930 92.760 49.910 ;
        RECT 94.460 48.270 94.600 93.510 ;
        RECT 95.780 93.170 96.040 93.490 ;
        RECT 95.320 88.070 95.580 88.390 ;
        RECT 95.380 86.010 95.520 88.070 ;
        RECT 95.320 85.690 95.580 86.010 ;
        RECT 95.840 81.250 95.980 93.170 ;
        RECT 97.620 91.130 97.880 91.450 ;
        RECT 96.700 85.690 96.960 86.010 ;
        RECT 95.780 80.930 96.040 81.250 ;
        RECT 96.240 80.590 96.500 80.910 ;
        RECT 94.860 80.250 95.120 80.570 ;
        RECT 94.920 64.250 95.060 80.250 ;
        RECT 96.300 76.570 96.440 80.590 ;
        RECT 96.760 77.170 96.900 85.690 ;
        RECT 97.160 79.570 97.420 79.890 ;
        RECT 96.700 76.850 96.960 77.170 ;
        RECT 96.300 76.430 96.900 76.570 ;
        RECT 96.760 75.810 96.900 76.430 ;
        RECT 96.700 75.490 96.960 75.810 ;
        RECT 97.220 75.210 97.360 79.570 ;
        RECT 97.680 75.810 97.820 91.130 ;
        RECT 98.080 86.030 98.340 86.350 ;
        RECT 97.620 75.490 97.880 75.810 ;
        RECT 97.220 75.130 97.820 75.210 ;
        RECT 95.320 74.810 95.580 75.130 ;
        RECT 97.220 75.070 97.880 75.130 ;
        RECT 97.620 74.810 97.880 75.070 ;
        RECT 95.380 74.530 95.520 74.810 ;
        RECT 96.700 74.530 96.960 74.790 ;
        RECT 95.380 74.470 96.960 74.530 ;
        RECT 95.380 74.390 96.900 74.470 ;
        RECT 95.380 72.070 95.520 74.390 ;
        RECT 97.680 74.110 97.820 74.810 ;
        RECT 97.620 73.790 97.880 74.110 ;
        RECT 95.320 71.750 95.580 72.070 ;
        RECT 95.380 69.690 95.520 71.750 ;
        RECT 97.680 69.690 97.820 73.790 ;
        RECT 95.320 69.370 95.580 69.690 ;
        RECT 96.700 69.370 96.960 69.690 ;
        RECT 97.620 69.370 97.880 69.690 ;
        RECT 96.760 64.930 96.900 69.370 ;
        RECT 97.160 69.030 97.420 69.350 ;
        RECT 96.700 64.610 96.960 64.930 ;
        RECT 94.860 63.930 95.120 64.250 ;
        RECT 96.700 62.970 96.960 63.230 ;
        RECT 97.220 62.970 97.360 69.030 ;
        RECT 97.680 69.010 97.820 69.370 ;
        RECT 97.620 68.690 97.880 69.010 ;
        RECT 96.700 62.910 97.360 62.970 ;
        RECT 97.620 62.910 97.880 63.230 ;
        RECT 96.760 62.830 97.360 62.910 ;
        RECT 96.690 62.035 96.970 62.405 ;
        RECT 95.320 54.750 95.580 55.070 ;
        RECT 95.380 53.710 95.520 54.750 ;
        RECT 95.320 53.390 95.580 53.710 ;
        RECT 96.760 50.990 96.900 62.035 ;
        RECT 97.220 53.710 97.360 62.830 ;
        RECT 97.680 60.850 97.820 62.910 ;
        RECT 97.620 60.530 97.880 60.850 ;
        RECT 98.140 56.770 98.280 86.030 ;
        RECT 98.540 85.350 98.800 85.670 ;
        RECT 98.080 56.450 98.340 56.770 ;
        RECT 98.080 55.770 98.340 56.090 ;
        RECT 97.160 53.390 97.420 53.710 ;
        RECT 97.620 52.710 97.880 53.030 ;
        RECT 96.700 50.670 96.960 50.990 ;
        RECT 97.680 50.845 97.820 52.710 ;
        RECT 97.610 50.475 97.890 50.845 ;
        RECT 97.680 50.310 97.820 50.475 ;
        RECT 97.620 49.990 97.880 50.310 ;
        RECT 94.400 47.950 94.660 48.270 ;
        RECT 90.780 47.870 91.440 47.930 ;
        RECT 89.800 47.270 90.060 47.590 ;
        RECT 90.780 46.910 90.920 47.870 ;
        RECT 91.180 47.610 91.440 47.870 ;
        RECT 92.100 47.610 92.360 47.930 ;
        RECT 92.560 47.610 92.820 47.930 ;
        RECT 90.720 46.590 90.980 46.910 ;
        RECT 92.160 44.870 92.300 47.610 ;
        RECT 93.480 47.270 93.740 47.590 ;
        RECT 93.540 45.210 93.680 47.270 ;
        RECT 93.480 44.890 93.740 45.210 ;
        RECT 92.100 44.610 92.360 44.870 ;
        RECT 91.700 44.550 92.360 44.610 ;
        RECT 91.700 44.470 92.300 44.550 ;
        RECT 89.800 42.170 90.060 42.490 ;
        RECT 89.860 40.450 90.000 42.170 ;
        RECT 91.700 40.450 91.840 44.470 ;
        RECT 92.100 43.870 92.360 44.190 ;
        RECT 92.160 42.830 92.300 43.870 ;
        RECT 92.100 42.510 92.360 42.830 ;
        RECT 89.800 40.130 90.060 40.450 ;
        RECT 91.640 40.130 91.900 40.450 ;
        RECT 93.540 34.330 93.680 44.890 ;
        RECT 96.700 42.850 96.960 43.170 ;
        RECT 96.760 39.770 96.900 42.850 ;
        RECT 97.160 42.510 97.420 42.830 ;
        RECT 97.220 40.450 97.360 42.510 ;
        RECT 97.160 40.130 97.420 40.450 ;
        RECT 96.700 39.450 96.960 39.770 ;
        RECT 88.420 34.010 88.680 34.330 ;
        RECT 93.480 34.010 93.740 34.330 ;
        RECT 84.580 32.455 86.460 32.825 ;
        RECT 83.360 31.970 83.620 32.290 ;
        RECT 85.660 31.970 85.920 32.290 ;
        RECT 82.900 31.290 83.160 31.610 ;
        RECT 76.920 30.270 77.180 30.590 ;
        RECT 78.300 30.270 78.560 30.590 ;
        RECT 81.980 30.270 82.240 30.590 ;
        RECT 71.860 29.250 72.120 29.570 ;
        RECT 69.160 28.830 69.760 28.970 ;
        RECT 76.980 28.890 77.120 30.270 ;
        RECT 78.360 28.890 78.500 30.270 ;
        RECT 69.100 28.230 69.360 28.550 ;
        RECT 68.180 25.170 68.440 25.490 ;
        RECT 9.580 24.295 11.460 24.665 ;
        RECT 39.580 24.295 41.460 24.665 ;
        RECT 69.160 23.110 69.300 28.230 ;
        RECT 69.620 26.850 69.760 28.830 ;
        RECT 75.540 28.570 75.800 28.890 ;
        RECT 76.920 28.570 77.180 28.890 ;
        RECT 78.300 28.570 78.560 28.890 ;
        RECT 69.560 26.530 69.820 26.850 ;
        RECT 71.860 26.190 72.120 26.510 ;
        RECT 69.580 24.295 71.460 24.665 ;
        RECT 71.920 24.130 72.060 26.190 ;
        RECT 75.600 26.170 75.740 28.570 ;
        RECT 82.040 28.210 82.180 30.270 ;
        RECT 85.720 29.570 85.860 31.970 ;
        RECT 88.480 31.950 88.620 34.010 ;
        RECT 88.880 32.990 89.140 33.310 ;
        RECT 86.120 31.630 86.380 31.950 ;
        RECT 88.420 31.630 88.680 31.950 ;
        RECT 86.180 29.570 86.320 31.630 ;
        RECT 88.940 31.610 89.080 32.990 ;
        RECT 88.880 31.290 89.140 31.610 ;
        RECT 93.540 31.270 93.680 34.010 ;
        RECT 96.760 33.990 96.900 39.450 ;
        RECT 97.620 38.430 97.880 38.750 ;
        RECT 97.680 37.050 97.820 38.430 ;
        RECT 97.620 36.730 97.880 37.050 ;
        RECT 98.140 36.450 98.280 55.770 ;
        RECT 98.600 51.330 98.740 85.350 ;
        RECT 99.060 63.765 99.200 93.850 ;
        RECT 99.580 89.575 101.460 89.945 ;
        RECT 101.820 88.810 101.960 96.570 ;
        RECT 102.280 93.830 102.420 96.910 ;
        RECT 102.740 94.170 102.880 98.270 ;
        RECT 102.680 93.850 102.940 94.170 ;
        RECT 102.220 93.510 102.480 93.830 ;
        RECT 102.680 92.830 102.940 93.150 ;
        RECT 101.360 88.670 101.960 88.810 ;
        RECT 100.380 87.730 100.640 88.050 ;
        RECT 100.440 86.690 100.580 87.730 ;
        RECT 100.380 86.370 100.640 86.690 ;
        RECT 101.360 84.990 101.500 88.670 ;
        RECT 101.760 88.070 102.020 88.390 ;
        RECT 101.300 84.670 101.560 84.990 ;
        RECT 99.580 84.135 101.460 84.505 ;
        RECT 101.820 83.970 101.960 88.070 ;
        RECT 102.220 85.690 102.480 86.010 ;
        RECT 101.760 83.650 102.020 83.970 ;
        RECT 99.460 82.630 99.720 82.950 ;
        RECT 100.380 82.630 100.640 82.950 ;
        RECT 100.840 82.805 101.100 82.950 ;
        RECT 99.520 80.570 99.660 82.630 ;
        RECT 99.460 80.250 99.720 80.570 ;
        RECT 100.440 79.890 100.580 82.630 ;
        RECT 100.830 82.435 101.110 82.805 ;
        RECT 101.300 82.630 101.560 82.950 ;
        RECT 100.900 81.250 101.040 82.435 ;
        RECT 100.840 80.930 101.100 81.250 ;
        RECT 100.900 80.570 101.040 80.930 ;
        RECT 101.360 80.570 101.500 82.630 ;
        RECT 102.280 81.250 102.420 85.690 ;
        RECT 102.740 84.990 102.880 92.830 ;
        RECT 103.200 89.410 103.340 118.330 ;
        RECT 104.520 117.990 104.780 118.310 ;
        RECT 104.060 111.870 104.320 112.190 ;
        RECT 104.120 109.810 104.260 111.870 ;
        RECT 104.060 109.490 104.320 109.810 ;
        RECT 103.600 92.830 103.860 93.150 ;
        RECT 104.060 92.830 104.320 93.150 ;
        RECT 103.660 89.410 103.800 92.830 ;
        RECT 103.140 89.090 103.400 89.410 ;
        RECT 103.600 89.090 103.860 89.410 ;
        RECT 104.120 89.070 104.260 92.830 ;
        RECT 104.580 89.070 104.720 117.990 ;
        RECT 104.980 112.890 105.240 113.210 ;
        RECT 104.060 88.750 104.320 89.070 ;
        RECT 104.520 88.750 104.780 89.070 ;
        RECT 103.600 88.410 103.860 88.730 ;
        RECT 103.140 87.390 103.400 87.710 ;
        RECT 102.680 84.670 102.940 84.990 ;
        RECT 102.220 80.930 102.480 81.250 ;
        RECT 100.840 80.250 101.100 80.570 ;
        RECT 101.300 80.250 101.560 80.570 ;
        RECT 100.380 79.570 100.640 79.890 ;
        RECT 101.360 79.550 101.500 80.250 ;
        RECT 102.680 79.910 102.940 80.230 ;
        RECT 101.300 79.230 101.560 79.550 ;
        RECT 99.580 78.695 101.460 79.065 ;
        RECT 100.840 74.810 101.100 75.130 ;
        RECT 102.220 74.810 102.480 75.130 ;
        RECT 100.900 74.110 101.040 74.810 ;
        RECT 100.840 73.790 101.100 74.110 ;
        RECT 101.760 73.790 102.020 74.110 ;
        RECT 99.580 73.255 101.460 73.625 ;
        RECT 101.820 72.070 101.960 73.790 ;
        RECT 101.760 71.750 102.020 72.070 ;
        RECT 102.280 70.370 102.420 74.810 ;
        RECT 102.740 71.390 102.880 79.910 ;
        RECT 102.680 71.070 102.940 71.390 ;
        RECT 99.920 70.050 100.180 70.370 ;
        RECT 102.220 70.050 102.480 70.370 ;
        RECT 99.980 69.690 100.120 70.050 ;
        RECT 103.200 69.770 103.340 87.390 ;
        RECT 99.920 69.370 100.180 69.690 ;
        RECT 101.820 69.630 103.340 69.770 ;
        RECT 99.580 67.815 101.460 68.185 ;
        RECT 98.990 63.395 99.270 63.765 ;
        RECT 99.000 62.910 99.260 63.230 ;
        RECT 99.060 58.810 99.200 62.910 ;
        RECT 99.580 62.375 101.460 62.745 ;
        RECT 101.300 60.530 101.560 60.850 ;
        RECT 100.840 60.190 101.100 60.510 ;
        RECT 100.900 59.490 101.040 60.190 ;
        RECT 101.360 59.490 101.500 60.530 ;
        RECT 100.840 59.170 101.100 59.490 ;
        RECT 101.300 59.170 101.560 59.490 ;
        RECT 99.000 58.490 99.260 58.810 ;
        RECT 99.580 56.935 101.460 57.305 ;
        RECT 101.820 54.050 101.960 69.630 ;
        RECT 103.140 69.030 103.400 69.350 ;
        RECT 103.200 66.630 103.340 69.030 ;
        RECT 103.140 66.310 103.400 66.630 ;
        RECT 103.140 64.610 103.400 64.930 ;
        RECT 103.200 62.210 103.340 64.610 ;
        RECT 103.140 61.890 103.400 62.210 ;
        RECT 103.660 62.170 103.800 88.410 ;
        RECT 104.060 88.070 104.320 88.390 ;
        RECT 104.520 88.070 104.780 88.390 ;
        RECT 104.120 86.690 104.260 88.070 ;
        RECT 104.060 86.370 104.320 86.690 ;
        RECT 104.060 85.010 104.320 85.330 ;
        RECT 104.120 70.030 104.260 85.010 ;
        RECT 104.580 82.270 104.720 88.070 ;
        RECT 105.040 86.690 105.180 112.890 ;
        RECT 105.440 109.150 105.700 109.470 ;
        RECT 105.500 104.030 105.640 109.150 ;
        RECT 105.440 103.710 105.700 104.030 ;
        RECT 105.500 100.290 105.640 103.710 ;
        RECT 105.440 99.970 105.700 100.290 ;
        RECT 105.960 89.410 106.100 118.330 ;
        RECT 109.180 118.310 109.320 120.630 ;
        RECT 113.260 120.030 113.520 120.350 ;
        RECT 109.120 117.990 109.380 118.310 ;
        RECT 110.500 117.990 110.760 118.310 ;
        RECT 109.180 110.150 109.320 117.990 ;
        RECT 110.560 113.890 110.700 117.990 ;
        RECT 113.320 115.590 113.460 120.030 ;
        RECT 113.780 119.330 113.920 125.810 ;
        RECT 114.240 122.050 114.380 138.990 ;
        RECT 117.920 138.990 119.230 139.130 ;
        RECT 117.400 125.810 117.660 126.130 ;
        RECT 114.580 124.935 116.460 125.305 ;
        RECT 117.460 122.050 117.600 125.810 ;
        RECT 114.180 121.730 114.440 122.050 ;
        RECT 117.400 121.730 117.660 122.050 ;
        RECT 114.580 119.495 116.460 119.865 ;
        RECT 117.920 119.330 118.060 138.990 ;
        RECT 125.740 127.490 125.880 138.395 ;
        RECT 125.680 127.170 125.940 127.490 ;
        RECT 113.720 119.010 113.980 119.330 ;
        RECT 117.860 119.010 118.120 119.330 ;
        RECT 114.180 118.670 114.440 118.990 ;
        RECT 114.240 116.610 114.380 118.670 ;
        RECT 114.180 116.290 114.440 116.610 ;
        RECT 113.260 115.270 113.520 115.590 ;
        RECT 114.580 114.055 116.460 114.425 ;
        RECT 110.500 113.570 110.760 113.890 ;
        RECT 113.260 110.170 113.520 110.490 ;
        RECT 109.120 109.830 109.380 110.150 ;
        RECT 109.580 109.830 109.840 110.150 ;
        RECT 107.280 109.150 107.540 109.470 ;
        RECT 107.340 107.770 107.480 109.150 ;
        RECT 107.280 107.450 107.540 107.770 ;
        RECT 109.180 107.430 109.320 109.830 ;
        RECT 109.640 108.450 109.780 109.830 ;
        RECT 109.580 108.130 109.840 108.450 ;
        RECT 110.500 107.450 110.760 107.770 ;
        RECT 109.120 107.110 109.380 107.430 ;
        RECT 109.180 104.370 109.320 107.110 ;
        RECT 110.560 105.730 110.700 107.450 ;
        RECT 110.500 105.410 110.760 105.730 ;
        RECT 113.320 105.050 113.460 110.170 ;
        RECT 117.400 109.830 117.660 110.150 ;
        RECT 114.580 108.615 116.460 108.985 ;
        RECT 116.480 107.790 116.740 108.110 ;
        RECT 114.640 106.430 114.900 106.750 ;
        RECT 113.260 104.730 113.520 105.050 ;
        RECT 109.120 104.050 109.380 104.370 ;
        RECT 109.180 101.990 109.320 104.050 ;
        RECT 113.320 101.990 113.460 104.730 ;
        RECT 114.700 104.710 114.840 106.430 ;
        RECT 116.540 105.730 116.680 107.790 ;
        RECT 116.480 105.410 116.740 105.730 ;
        RECT 117.460 104.710 117.600 109.830 ;
        RECT 113.720 104.390 113.980 104.710 ;
        RECT 114.640 104.390 114.900 104.710 ;
        RECT 117.400 104.390 117.660 104.710 ;
        RECT 109.120 101.670 109.380 101.990 ;
        RECT 111.880 101.670 112.140 101.990 ;
        RECT 113.260 101.670 113.520 101.990 ;
        RECT 109.180 99.270 109.320 101.670 ;
        RECT 110.040 100.990 110.300 101.310 ;
        RECT 109.120 98.950 109.380 99.270 ;
        RECT 109.580 98.950 109.840 99.270 ;
        RECT 109.180 97.230 109.320 98.950 ;
        RECT 109.120 96.910 109.380 97.230 ;
        RECT 105.900 89.090 106.160 89.410 ;
        RECT 105.440 87.390 105.700 87.710 ;
        RECT 104.980 86.370 105.240 86.690 ;
        RECT 105.500 86.350 105.640 87.390 ;
        RECT 105.440 86.030 105.700 86.350 ;
        RECT 104.980 85.690 105.240 86.010 ;
        RECT 105.040 83.630 105.180 85.690 ;
        RECT 109.180 85.670 109.320 96.910 ;
        RECT 109.640 96.890 109.780 98.950 ;
        RECT 110.100 96.890 110.240 100.990 ;
        RECT 109.580 96.570 109.840 96.890 ;
        RECT 110.040 96.570 110.300 96.890 ;
        RECT 110.500 96.570 110.760 96.890 ;
        RECT 110.560 94.850 110.700 96.570 ;
        RECT 111.940 96.210 112.080 101.670 ;
        RECT 113.320 99.610 113.460 101.670 ;
        RECT 113.260 99.290 113.520 99.610 ;
        RECT 111.880 95.890 112.140 96.210 ;
        RECT 110.500 94.530 110.760 94.850 ;
        RECT 111.940 94.170 112.080 95.890 ;
        RECT 113.320 94.510 113.460 99.290 ;
        RECT 113.260 94.190 113.520 94.510 ;
        RECT 111.880 93.850 112.140 94.170 ;
        RECT 113.780 93.490 113.920 104.390 ;
        RECT 114.580 103.175 116.460 103.545 ;
        RECT 117.460 102.330 117.600 104.390 ;
        RECT 117.400 102.010 117.660 102.330 ;
        RECT 114.180 100.990 114.440 101.310 ;
        RECT 114.240 98.930 114.380 100.990 ;
        RECT 117.460 99.270 117.600 102.010 ;
        RECT 117.400 98.950 117.660 99.270 ;
        RECT 114.180 98.610 114.440 98.930 ;
        RECT 117.860 98.270 118.120 98.590 ;
        RECT 114.580 97.735 116.460 98.105 ;
        RECT 117.920 97.230 118.060 98.270 ;
        RECT 117.860 96.910 118.120 97.230 ;
        RECT 113.720 93.170 113.980 93.490 ;
        RECT 114.580 92.295 116.460 92.665 ;
        RECT 112.340 88.070 112.600 88.390 ;
        RECT 116.940 88.070 117.200 88.390 ;
        RECT 109.120 85.350 109.380 85.670 ;
        RECT 110.960 85.350 111.220 85.670 ;
        RECT 104.980 83.310 105.240 83.630 ;
        RECT 109.180 83.290 109.320 85.350 ;
        RECT 109.120 82.970 109.380 83.290 ;
        RECT 104.980 82.805 105.240 82.950 ;
        RECT 104.970 82.435 105.250 82.805 ;
        RECT 106.820 82.630 107.080 82.950 ;
        RECT 104.520 81.950 104.780 82.270 ;
        RECT 106.880 79.890 107.020 82.630 ;
        RECT 110.500 81.950 110.760 82.270 ;
        RECT 110.560 80.910 110.700 81.950 ;
        RECT 111.020 81.250 111.160 85.350 ;
        RECT 111.420 81.950 111.680 82.270 ;
        RECT 110.960 80.930 111.220 81.250 ;
        RECT 110.500 80.590 110.760 80.910 ;
        RECT 111.480 80.570 111.620 81.950 ;
        RECT 112.400 81.250 112.540 88.070 ;
        RECT 113.720 87.390 113.980 87.710 ;
        RECT 114.180 87.390 114.440 87.710 ;
        RECT 113.260 83.650 113.520 83.970 ;
        RECT 113.320 82.870 113.460 83.650 ;
        RECT 113.780 83.290 113.920 87.390 ;
        RECT 114.240 86.090 114.380 87.390 ;
        RECT 114.580 86.855 116.460 87.225 ;
        RECT 114.640 86.090 114.900 86.350 ;
        RECT 114.240 86.030 114.900 86.090 ;
        RECT 114.240 85.950 114.840 86.030 ;
        RECT 117.000 86.010 117.140 88.070 ;
        RECT 116.940 85.690 117.200 86.010 ;
        RECT 117.000 85.410 117.140 85.690 ;
        RECT 117.000 85.270 117.600 85.410 ;
        RECT 116.940 84.670 117.200 84.990 ;
        RECT 113.720 82.970 113.980 83.290 ;
        RECT 112.860 82.730 113.460 82.870 ;
        RECT 112.340 80.930 112.600 81.250 ;
        RECT 112.860 80.650 113.000 82.730 ;
        RECT 114.180 82.630 114.440 82.950 ;
        RECT 111.420 80.250 111.680 80.570 ;
        RECT 112.400 80.510 113.000 80.650 ;
        RECT 113.260 80.590 113.520 80.910 ;
        RECT 112.400 79.890 112.540 80.510 ;
        RECT 106.820 79.570 107.080 79.890 ;
        RECT 112.340 79.570 112.600 79.890 ;
        RECT 110.500 77.190 110.760 77.510 ;
        RECT 110.960 77.190 111.220 77.510 ;
        RECT 110.560 75.810 110.700 77.190 ;
        RECT 110.500 75.490 110.760 75.810 ;
        RECT 111.020 72.410 111.160 77.190 ;
        RECT 112.400 72.410 112.540 79.570 ;
        RECT 113.320 76.830 113.460 80.590 ;
        RECT 113.720 80.250 113.980 80.570 ;
        RECT 113.260 76.510 113.520 76.830 ;
        RECT 113.320 75.810 113.460 76.510 ;
        RECT 113.260 75.490 113.520 75.810 ;
        RECT 112.800 74.470 113.060 74.790 ;
        RECT 110.960 72.090 111.220 72.410 ;
        RECT 112.340 72.090 112.600 72.410 ;
        RECT 110.500 71.750 110.760 72.070 ;
        RECT 104.520 71.070 104.780 71.390 ;
        RECT 104.060 69.710 104.320 70.030 ;
        RECT 104.580 69.350 104.720 71.070 ;
        RECT 104.520 69.030 104.780 69.350 ;
        RECT 105.440 68.690 105.700 69.010 ;
        RECT 105.500 66.970 105.640 68.690 ;
        RECT 105.440 66.650 105.700 66.970 ;
        RECT 104.980 64.270 105.240 64.590 ;
        RECT 103.660 62.030 104.720 62.170 ;
        RECT 102.220 55.430 102.480 55.750 ;
        RECT 101.760 53.730 102.020 54.050 ;
        RECT 99.000 53.050 99.260 53.370 ;
        RECT 101.760 53.050 102.020 53.370 ;
        RECT 98.540 51.010 98.800 51.330 ;
        RECT 99.060 50.730 99.200 53.050 ;
        RECT 99.580 51.495 101.460 51.865 ;
        RECT 98.600 50.590 99.200 50.730 ;
        RECT 98.600 50.310 98.740 50.590 ;
        RECT 98.540 49.990 98.800 50.310 ;
        RECT 99.000 49.650 99.260 49.970 ;
        RECT 99.060 47.930 99.200 49.650 ;
        RECT 101.820 48.610 101.960 53.050 ;
        RECT 101.760 48.290 102.020 48.610 ;
        RECT 99.000 47.610 99.260 47.930 ;
        RECT 99.060 45.290 99.200 47.610 ;
        RECT 99.580 46.055 101.460 46.425 ;
        RECT 101.820 45.890 101.960 48.290 ;
        RECT 101.760 45.570 102.020 45.890 ;
        RECT 99.060 45.150 99.660 45.290 ;
        RECT 99.520 44.190 99.660 45.150 ;
        RECT 99.460 43.870 99.720 44.190 ;
        RECT 99.520 43.170 99.660 43.870 ;
        RECT 99.460 42.850 99.720 43.170 ;
        RECT 101.820 42.490 101.960 45.570 ;
        RECT 102.280 44.870 102.420 55.430 ;
        RECT 103.140 53.050 103.400 53.370 ;
        RECT 103.200 50.990 103.340 53.050 ;
        RECT 104.580 51.330 104.720 62.030 ;
        RECT 105.040 61.870 105.180 64.270 ;
        RECT 105.500 63.910 105.640 66.650 ;
        RECT 110.560 66.630 110.700 71.750 ;
        RECT 111.020 69.690 111.160 72.090 ;
        RECT 110.960 69.370 111.220 69.690 ;
        RECT 110.500 66.310 110.760 66.630 ;
        RECT 111.020 64.250 111.160 69.370 ;
        RECT 112.400 66.970 112.540 72.090 ;
        RECT 112.340 66.650 112.600 66.970 ;
        RECT 110.960 63.930 111.220 64.250 ;
        RECT 105.440 63.590 105.700 63.910 ;
        RECT 104.980 61.550 105.240 61.870 ;
        RECT 111.020 61.610 111.160 63.930 ;
        RECT 112.400 61.870 112.540 66.650 ;
        RECT 112.860 65.950 113.000 74.470 ;
        RECT 113.260 74.130 113.520 74.450 ;
        RECT 113.320 66.290 113.460 74.130 ;
        RECT 113.780 72.070 113.920 80.250 ;
        RECT 114.240 80.230 114.380 82.630 ;
        RECT 117.000 82.270 117.140 84.670 ;
        RECT 116.940 81.950 117.200 82.270 ;
        RECT 114.580 81.415 116.460 81.785 ;
        RECT 117.000 81.250 117.140 81.950 ;
        RECT 116.940 80.930 117.200 81.250 ;
        RECT 117.460 80.650 117.600 85.270 ;
        RECT 118.780 84.670 119.040 84.990 ;
        RECT 118.840 82.610 118.980 84.670 ;
        RECT 118.780 82.290 119.040 82.610 ;
        RECT 117.000 80.570 117.600 80.650 ;
        RECT 116.940 80.510 117.600 80.570 ;
        RECT 116.940 80.250 117.200 80.510 ;
        RECT 114.180 79.910 114.440 80.230 ;
        RECT 114.240 72.070 114.380 79.910 ;
        RECT 116.480 79.230 116.740 79.550 ;
        RECT 116.540 77.170 116.680 79.230 ;
        RECT 116.480 76.850 116.740 77.170 ;
        RECT 114.580 75.975 116.460 76.345 ;
        RECT 115.100 74.470 115.360 74.790 ;
        RECT 115.160 72.410 115.300 74.470 ;
        RECT 115.100 72.090 115.360 72.410 ;
        RECT 113.720 71.750 113.980 72.070 ;
        RECT 114.180 71.750 114.440 72.070 ;
        RECT 113.720 71.070 113.980 71.390 ;
        RECT 116.940 71.070 117.200 71.390 ;
        RECT 113.780 70.370 113.920 71.070 ;
        RECT 114.580 70.535 116.460 70.905 ;
        RECT 113.720 70.050 113.980 70.370 ;
        RECT 117.000 69.350 117.140 71.070 ;
        RECT 117.400 69.710 117.660 70.030 ;
        RECT 116.940 69.030 117.200 69.350 ;
        RECT 117.460 67.650 117.600 69.710 ;
        RECT 117.400 67.330 117.660 67.650 ;
        RECT 113.260 65.970 113.520 66.290 ;
        RECT 116.940 65.970 117.200 66.290 ;
        RECT 112.800 65.630 113.060 65.950 ;
        RECT 113.320 64.930 113.460 65.970 ;
        RECT 114.580 65.095 116.460 65.465 ;
        RECT 113.260 64.610 113.520 64.930 ;
        RECT 110.560 61.530 111.160 61.610 ;
        RECT 112.340 61.550 112.600 61.870 ;
        RECT 117.000 61.530 117.140 65.970 ;
        RECT 119.700 65.630 119.960 65.950 ;
        RECT 118.780 63.930 119.040 64.250 ;
        RECT 118.320 63.590 118.580 63.910 ;
        RECT 118.380 62.210 118.520 63.590 ;
        RECT 118.320 61.890 118.580 62.210 ;
        RECT 110.500 61.470 111.160 61.530 ;
        RECT 110.500 61.210 110.760 61.470 ;
        RECT 109.120 60.530 109.380 60.850 ;
        RECT 107.280 60.190 107.540 60.510 ;
        RECT 107.340 58.810 107.480 60.190 ;
        RECT 109.180 59.490 109.320 60.530 ;
        RECT 109.120 59.170 109.380 59.490 ;
        RECT 111.020 59.150 111.160 61.470 ;
        RECT 116.940 61.210 117.200 61.530 ;
        RECT 114.580 59.655 116.460 60.025 ;
        RECT 117.000 59.490 117.140 61.210 ;
        RECT 118.840 59.490 118.980 63.930 ;
        RECT 119.760 61.190 119.900 65.630 ;
        RECT 119.700 60.870 119.960 61.190 ;
        RECT 116.940 59.170 117.200 59.490 ;
        RECT 118.780 59.170 119.040 59.490 ;
        RECT 110.960 58.830 111.220 59.150 ;
        RECT 113.720 58.830 113.980 59.150 ;
        RECT 105.900 58.490 106.160 58.810 ;
        RECT 107.280 58.490 107.540 58.810 ;
        RECT 105.960 55.410 106.100 58.490 ;
        RECT 111.020 56.090 111.160 58.830 ;
        RECT 113.780 56.770 113.920 58.830 ;
        RECT 118.320 58.490 118.580 58.810 ;
        RECT 113.720 56.450 113.980 56.770 ;
        RECT 110.960 55.770 111.220 56.090 ;
        RECT 118.380 55.750 118.520 58.490 ;
        RECT 118.320 55.430 118.580 55.750 ;
        RECT 105.900 55.090 106.160 55.410 ;
        RECT 110.040 55.090 110.300 55.410 ;
        RECT 104.520 51.010 104.780 51.330 ;
        RECT 103.140 50.670 103.400 50.990 ;
        RECT 103.200 50.310 103.340 50.670 ;
        RECT 102.680 49.990 102.940 50.310 ;
        RECT 103.140 49.990 103.400 50.310 ;
        RECT 105.900 49.990 106.160 50.310 ;
        RECT 102.220 44.550 102.480 44.870 ;
        RECT 102.280 42.830 102.420 44.550 ;
        RECT 102.220 42.510 102.480 42.830 ;
        RECT 101.760 42.170 102.020 42.490 ;
        RECT 99.580 40.615 101.460 40.985 ;
        RECT 102.280 39.770 102.420 42.510 ;
        RECT 102.220 39.450 102.480 39.770 ;
        RECT 98.540 36.450 98.800 36.710 ;
        RECT 98.140 36.390 98.800 36.450 ;
        RECT 98.140 36.310 98.740 36.390 ;
        RECT 98.080 35.710 98.340 36.030 ;
        RECT 94.860 33.670 95.120 33.990 ;
        RECT 96.700 33.670 96.960 33.990 ;
        RECT 94.920 32.290 95.060 33.670 ;
        RECT 94.860 31.970 95.120 32.290 ;
        RECT 93.480 30.950 93.740 31.270 ;
        RECT 87.960 30.270 88.220 30.590 ;
        RECT 93.480 30.270 93.740 30.590 ;
        RECT 85.660 29.250 85.920 29.570 ;
        RECT 86.120 29.250 86.380 29.570 ;
        RECT 88.020 28.550 88.160 30.270 ;
        RECT 93.540 28.890 93.680 30.270 ;
        RECT 96.760 28.890 96.900 33.670 ;
        RECT 98.140 33.310 98.280 35.710 ;
        RECT 97.620 32.990 97.880 33.310 ;
        RECT 98.080 32.990 98.340 33.310 ;
        RECT 97.680 32.290 97.820 32.990 ;
        RECT 97.620 31.970 97.880 32.290 ;
        RECT 98.600 31.950 98.740 36.310 ;
        RECT 99.580 35.175 101.460 35.545 ;
        RECT 102.740 34.330 102.880 49.990 ;
        RECT 104.980 47.950 105.240 48.270 ;
        RECT 103.600 46.590 103.860 46.910 ;
        RECT 103.660 45.210 103.800 46.590 ;
        RECT 103.600 44.890 103.860 45.210 ;
        RECT 105.040 42.150 105.180 47.950 ;
        RECT 105.960 43.170 106.100 49.990 ;
        RECT 110.100 47.930 110.240 55.090 ;
        RECT 114.580 54.215 116.460 54.585 ;
        RECT 114.580 48.775 116.460 49.145 ;
        RECT 108.200 47.610 108.460 47.930 ;
        RECT 110.040 47.610 110.300 47.930 ;
        RECT 106.820 46.590 107.080 46.910 ;
        RECT 106.880 43.170 107.020 46.590 ;
        RECT 105.900 42.850 106.160 43.170 ;
        RECT 106.820 42.850 107.080 43.170 ;
        RECT 105.960 42.150 106.100 42.850 ;
        RECT 104.980 41.830 105.240 42.150 ;
        RECT 105.900 41.830 106.160 42.150 ;
        RECT 103.140 38.770 103.400 39.090 ;
        RECT 103.200 37.730 103.340 38.770 ;
        RECT 103.140 37.410 103.400 37.730 ;
        RECT 105.040 36.370 105.180 41.830 ;
        RECT 105.960 37.730 106.100 41.830 ;
        RECT 108.260 41.810 108.400 47.610 ;
        RECT 109.120 46.590 109.380 46.910 ;
        RECT 109.180 44.870 109.320 46.590 ;
        RECT 109.120 44.550 109.380 44.870 ;
        RECT 108.200 41.490 108.460 41.810 ;
        RECT 110.100 39.430 110.240 47.610 ;
        RECT 114.580 43.335 116.460 43.705 ;
        RECT 111.880 42.510 112.140 42.830 ;
        RECT 111.940 40.450 112.080 42.510 ;
        RECT 111.880 40.130 112.140 40.450 ;
        RECT 109.120 39.110 109.380 39.430 ;
        RECT 110.040 39.110 110.300 39.430 ;
        RECT 109.180 37.730 109.320 39.110 ;
        RECT 105.900 37.410 106.160 37.730 ;
        RECT 109.120 37.410 109.380 37.730 ;
        RECT 110.100 37.050 110.240 39.110 ;
        RECT 110.960 38.430 111.220 38.750 ;
        RECT 111.020 37.390 111.160 38.430 ;
        RECT 114.580 37.895 116.460 38.265 ;
        RECT 110.960 37.070 111.220 37.390 ;
        RECT 110.040 36.730 110.300 37.050 ;
        RECT 104.980 36.050 105.240 36.370 ;
        RECT 102.680 34.010 102.940 34.330 ;
        RECT 102.740 32.290 102.880 34.010 ;
        RECT 114.580 32.455 116.460 32.825 ;
        RECT 102.680 31.970 102.940 32.290 ;
        RECT 98.540 31.630 98.800 31.950 ;
        RECT 99.580 29.735 101.460 30.105 ;
        RECT 93.480 28.570 93.740 28.890 ;
        RECT 96.700 28.570 96.960 28.890 ;
        RECT 87.960 28.230 88.220 28.550 ;
        RECT 81.980 27.890 82.240 28.210 ;
        RECT 84.580 27.015 86.460 27.385 ;
        RECT 114.580 27.015 116.460 27.385 ;
        RECT 75.540 25.850 75.800 26.170 ;
        RECT 99.580 24.295 101.460 24.665 ;
        RECT 71.860 23.810 72.120 24.130 ;
        RECT 69.100 22.790 69.360 23.110 ;
        RECT 24.580 21.575 26.460 21.945 ;
        RECT 54.580 21.575 56.460 21.945 ;
        RECT 84.580 21.575 86.460 21.945 ;
        RECT 114.580 21.575 116.460 21.945 ;
        RECT 9.580 18.855 11.460 19.225 ;
        RECT 39.580 18.855 41.460 19.225 ;
        RECT 69.580 18.855 71.460 19.225 ;
        RECT 99.580 18.855 101.460 19.225 ;
        RECT 24.580 16.135 26.460 16.505 ;
        RECT 54.580 16.135 56.460 16.505 ;
        RECT 84.580 16.135 86.460 16.505 ;
        RECT 114.580 16.135 116.460 16.505 ;
        RECT 9.580 13.415 11.460 13.785 ;
        RECT 39.580 13.415 41.460 13.785 ;
        RECT 69.580 13.415 71.460 13.785 ;
        RECT 99.580 13.415 101.460 13.785 ;
        RECT 24.580 10.695 26.460 11.065 ;
        RECT 54.580 10.695 56.460 11.065 ;
        RECT 84.580 10.695 86.460 11.065 ;
        RECT 114.580 10.695 116.460 11.065 ;
      LAYER met3 ;
        RECT 9.530 127.675 11.510 128.005 ;
        RECT 39.530 127.675 41.510 128.005 ;
        RECT 69.530 127.675 71.510 128.005 ;
        RECT 99.530 127.675 101.510 128.005 ;
        RECT 24.530 124.955 26.510 125.285 ;
        RECT 54.530 124.955 56.510 125.285 ;
        RECT 84.530 124.955 86.510 125.285 ;
        RECT 114.530 124.955 116.510 125.285 ;
        RECT 9.530 122.235 11.510 122.565 ;
        RECT 39.530 122.235 41.510 122.565 ;
        RECT 69.530 122.235 71.510 122.565 ;
        RECT 99.530 122.235 101.510 122.565 ;
        RECT 3.745 120.170 4.075 120.185 ;
        RECT 2.000 119.870 4.075 120.170 ;
        RECT 3.745 119.855 4.075 119.870 ;
        RECT 24.530 119.515 26.510 119.845 ;
        RECT 54.530 119.515 56.510 119.845 ;
        RECT 84.530 119.515 86.510 119.845 ;
        RECT 114.530 119.515 116.510 119.845 ;
        RECT 9.530 116.795 11.510 117.125 ;
        RECT 39.530 116.795 41.510 117.125 ;
        RECT 69.530 116.795 71.510 117.125 ;
        RECT 99.530 116.795 101.510 117.125 ;
        RECT 24.530 114.075 26.510 114.405 ;
        RECT 54.530 114.075 56.510 114.405 ;
        RECT 84.530 114.075 86.510 114.405 ;
        RECT 114.530 114.075 116.510 114.405 ;
        RECT 9.530 111.355 11.510 111.685 ;
        RECT 39.530 111.355 41.510 111.685 ;
        RECT 69.530 111.355 71.510 111.685 ;
        RECT 99.530 111.355 101.510 111.685 ;
        RECT 24.530 108.635 26.510 108.965 ;
        RECT 54.530 108.635 56.510 108.965 ;
        RECT 84.530 108.635 86.510 108.965 ;
        RECT 114.530 108.635 116.510 108.965 ;
        RECT 9.530 105.915 11.510 106.245 ;
        RECT 39.530 105.915 41.510 106.245 ;
        RECT 69.530 105.915 71.510 106.245 ;
        RECT 99.530 105.915 101.510 106.245 ;
        RECT 25.365 104.530 25.695 104.545 ;
        RECT 44.685 104.530 45.015 104.545 ;
        RECT 72.030 104.530 72.410 104.540 ;
        RECT 90.225 104.530 90.555 104.545 ;
        RECT 25.365 104.230 90.555 104.530 ;
        RECT 25.365 104.215 25.695 104.230 ;
        RECT 44.685 104.215 45.015 104.230 ;
        RECT 72.030 104.220 72.410 104.230 ;
        RECT 90.225 104.215 90.555 104.230 ;
        RECT 24.530 103.195 26.510 103.525 ;
        RECT 54.530 103.195 56.510 103.525 ;
        RECT 84.530 103.195 86.510 103.525 ;
        RECT 114.530 103.195 116.510 103.525 ;
        RECT 9.530 100.475 11.510 100.805 ;
        RECT 39.530 100.475 41.510 100.805 ;
        RECT 69.530 100.475 71.510 100.805 ;
        RECT 99.530 100.475 101.510 100.805 ;
        RECT 67.225 98.410 67.555 98.425 ;
        RECT 68.350 98.410 68.730 98.420 ;
        RECT 67.225 98.110 68.730 98.410 ;
        RECT 67.225 98.095 67.555 98.110 ;
        RECT 68.350 98.100 68.730 98.110 ;
        RECT 24.530 97.755 26.510 98.085 ;
        RECT 54.530 97.755 56.510 98.085 ;
        RECT 84.530 97.755 86.510 98.085 ;
        RECT 114.530 97.755 116.510 98.085 ;
        RECT 9.530 95.035 11.510 95.365 ;
        RECT 39.530 95.035 41.510 95.365 ;
        RECT 69.530 95.035 71.510 95.365 ;
        RECT 99.530 95.035 101.510 95.365 ;
        RECT 53.630 93.650 54.010 93.660 ;
        RECT 54.805 93.650 55.135 93.665 ;
        RECT 53.630 93.350 55.135 93.650 ;
        RECT 53.630 93.340 54.010 93.350 ;
        RECT 54.805 93.335 55.135 93.350 ;
        RECT 24.530 92.315 26.510 92.645 ;
        RECT 54.530 92.315 56.510 92.645 ;
        RECT 84.530 92.315 86.510 92.645 ;
        RECT 114.530 92.315 116.510 92.645 ;
        RECT 9.530 89.595 11.510 89.925 ;
        RECT 39.530 89.595 41.510 89.925 ;
        RECT 69.530 89.595 71.510 89.925 ;
        RECT 99.530 89.595 101.510 89.925 ;
        RECT 24.530 86.875 26.510 87.205 ;
        RECT 54.530 86.875 56.510 87.205 ;
        RECT 84.530 86.875 86.510 87.205 ;
        RECT 114.530 86.875 116.510 87.205 ;
        RECT 20.510 86.170 20.890 86.180 ;
        RECT 2.000 85.870 20.890 86.170 ;
        RECT 20.510 85.860 20.890 85.870 ;
        RECT 9.530 84.155 11.510 84.485 ;
        RECT 39.530 84.155 41.510 84.485 ;
        RECT 69.530 84.155 71.510 84.485 ;
        RECT 99.530 84.155 101.510 84.485 ;
        RECT 100.805 82.770 101.135 82.785 ;
        RECT 104.945 82.770 105.275 82.785 ;
        RECT 100.805 82.470 105.275 82.770 ;
        RECT 100.805 82.455 101.135 82.470 ;
        RECT 104.945 82.455 105.275 82.470 ;
        RECT 24.530 81.435 26.510 81.765 ;
        RECT 54.530 81.435 56.510 81.765 ;
        RECT 84.530 81.435 86.510 81.765 ;
        RECT 114.530 81.435 116.510 81.765 ;
        RECT 9.530 78.715 11.510 79.045 ;
        RECT 39.530 78.715 41.510 79.045 ;
        RECT 69.530 78.715 71.510 79.045 ;
        RECT 99.530 78.715 101.510 79.045 ;
        RECT 24.530 75.995 26.510 76.325 ;
        RECT 54.530 75.995 56.510 76.325 ;
        RECT 84.530 75.995 86.510 76.325 ;
        RECT 114.530 75.995 116.510 76.325 ;
        RECT 20.510 75.290 20.890 75.300 ;
        RECT 64.005 75.290 64.335 75.305 ;
        RECT 20.510 74.990 64.335 75.290 ;
        RECT 20.510 74.980 20.890 74.990 ;
        RECT 64.005 74.975 64.335 74.990 ;
        RECT 78.725 75.290 79.055 75.305 ;
        RECT 83.325 75.290 83.655 75.305 ;
        RECT 78.725 74.990 83.655 75.290 ;
        RECT 78.725 74.975 79.055 74.990 ;
        RECT 83.325 74.975 83.655 74.990 ;
        RECT 72.285 74.610 72.615 74.625 ;
        RECT 88.845 74.610 89.175 74.625 ;
        RECT 72.285 74.310 89.175 74.610 ;
        RECT 72.285 74.295 72.615 74.310 ;
        RECT 88.845 74.295 89.175 74.310 ;
        RECT 71.825 73.940 72.155 73.945 ;
        RECT 71.825 73.930 72.410 73.940 ;
        RECT 71.825 73.630 72.610 73.930 ;
        RECT 71.825 73.620 72.410 73.630 ;
        RECT 71.825 73.615 72.155 73.620 ;
        RECT 9.530 73.275 11.510 73.605 ;
        RECT 39.530 73.275 41.510 73.605 ;
        RECT 69.530 73.275 71.510 73.605 ;
        RECT 99.530 73.275 101.510 73.605 ;
        RECT 52.965 72.570 53.295 72.585 ;
        RECT 53.630 72.570 54.010 72.580 ;
        RECT 52.965 72.270 54.010 72.570 ;
        RECT 52.965 72.255 53.295 72.270 ;
        RECT 53.630 72.260 54.010 72.270 ;
        RECT 58.945 71.890 59.275 71.905 ;
        RECT 91.145 71.890 91.475 71.905 ;
        RECT 58.945 71.590 91.475 71.890 ;
        RECT 58.945 71.575 59.275 71.590 ;
        RECT 91.145 71.575 91.475 71.590 ;
        RECT 24.530 70.555 26.510 70.885 ;
        RECT 54.530 70.555 56.510 70.885 ;
        RECT 84.530 70.555 86.510 70.885 ;
        RECT 114.530 70.555 116.510 70.885 ;
        RECT 9.530 67.835 11.510 68.165 ;
        RECT 39.530 67.835 41.510 68.165 ;
        RECT 69.530 67.835 71.510 68.165 ;
        RECT 99.530 67.835 101.510 68.165 ;
        RECT 24.530 65.115 26.510 65.445 ;
        RECT 54.530 65.115 56.510 65.445 ;
        RECT 84.530 65.115 86.510 65.445 ;
        RECT 114.530 65.115 116.510 65.445 ;
        RECT 98.965 63.730 99.295 63.745 ;
        RECT 96.910 63.430 99.295 63.730 ;
        RECT 9.530 62.395 11.510 62.725 ;
        RECT 39.530 62.395 41.510 62.725 ;
        RECT 69.530 62.395 71.510 62.725 ;
        RECT 96.910 62.385 97.210 63.430 ;
        RECT 98.965 63.415 99.295 63.430 ;
        RECT 99.530 62.395 101.510 62.725 ;
        RECT 96.665 62.070 97.210 62.385 ;
        RECT 96.665 62.055 96.995 62.070 ;
        RECT 24.530 59.675 26.510 60.005 ;
        RECT 54.530 59.675 56.510 60.005 ;
        RECT 84.530 59.675 86.510 60.005 ;
        RECT 114.530 59.675 116.510 60.005 ;
        RECT 9.530 56.955 11.510 57.285 ;
        RECT 39.530 56.955 41.510 57.285 ;
        RECT 69.530 56.955 71.510 57.285 ;
        RECT 99.530 56.955 101.510 57.285 ;
        RECT 32.265 55.570 32.595 55.585 ;
        RECT 72.030 55.570 72.410 55.580 ;
        RECT 92.065 55.570 92.395 55.585 ;
        RECT 32.265 55.270 92.395 55.570 ;
        RECT 32.265 55.255 32.595 55.270 ;
        RECT 47.230 54.890 47.530 55.270 ;
        RECT 72.030 55.260 72.410 55.270 ;
        RECT 92.065 55.255 92.395 55.270 ;
        RECT 47.905 54.890 48.235 54.905 ;
        RECT 47.230 54.590 48.235 54.890 ;
        RECT 47.905 54.575 48.235 54.590 ;
        RECT 24.530 54.235 26.510 54.565 ;
        RECT 54.530 54.235 56.510 54.565 ;
        RECT 84.530 54.235 86.510 54.565 ;
        RECT 114.530 54.235 116.510 54.565 ;
        RECT 66.305 52.850 66.635 52.865 ;
        RECT 77.345 52.850 77.675 52.865 ;
        RECT 66.305 52.550 77.675 52.850 ;
        RECT 66.305 52.535 66.635 52.550 ;
        RECT 77.345 52.535 77.675 52.550 ;
        RECT 2.000 51.855 2.235 52.185 ;
        RECT 9.530 51.515 11.510 51.845 ;
        RECT 39.530 51.515 41.510 51.845 ;
        RECT 69.530 51.515 71.510 51.845 ;
        RECT 99.530 51.515 101.510 51.845 ;
        RECT 67.685 51.490 68.015 51.505 ;
        RECT 68.350 51.490 68.730 51.500 ;
        RECT 67.685 51.190 68.730 51.490 ;
        RECT 67.685 51.175 68.015 51.190 ;
        RECT 68.350 51.180 68.730 51.190 ;
        RECT 68.605 50.810 68.935 50.825 ;
        RECT 97.585 50.810 97.915 50.825 ;
        RECT 68.605 50.510 97.915 50.810 ;
        RECT 68.605 50.495 68.935 50.510 ;
        RECT 97.585 50.495 97.915 50.510 ;
        RECT 24.530 48.795 26.510 49.125 ;
        RECT 54.530 48.795 56.510 49.125 ;
        RECT 84.530 48.795 86.510 49.125 ;
        RECT 114.530 48.795 116.510 49.125 ;
        RECT 9.530 46.075 11.510 46.405 ;
        RECT 39.530 46.075 41.510 46.405 ;
        RECT 69.530 46.075 71.510 46.405 ;
        RECT 99.530 46.075 101.510 46.405 ;
        RECT 24.530 43.355 26.510 43.685 ;
        RECT 54.530 43.355 56.510 43.685 ;
        RECT 84.530 43.355 86.510 43.685 ;
        RECT 114.530 43.355 116.510 43.685 ;
        RECT 9.530 40.635 11.510 40.965 ;
        RECT 39.530 40.635 41.510 40.965 ;
        RECT 69.530 40.635 71.510 40.965 ;
        RECT 99.530 40.635 101.510 40.965 ;
        RECT 24.530 37.915 26.510 38.245 ;
        RECT 54.530 37.915 56.510 38.245 ;
        RECT 84.530 37.915 86.510 38.245 ;
        RECT 114.530 37.915 116.510 38.245 ;
        RECT 9.530 35.195 11.510 35.525 ;
        RECT 39.530 35.195 41.510 35.525 ;
        RECT 69.530 35.195 71.510 35.525 ;
        RECT 99.530 35.195 101.510 35.525 ;
        RECT 24.530 32.475 26.510 32.805 ;
        RECT 54.530 32.475 56.510 32.805 ;
        RECT 84.530 32.475 86.510 32.805 ;
        RECT 114.530 32.475 116.510 32.805 ;
        RECT 9.530 29.755 11.510 30.085 ;
        RECT 39.530 29.755 41.510 30.085 ;
        RECT 69.530 29.755 71.510 30.085 ;
        RECT 99.530 29.755 101.510 30.085 ;
        RECT 24.530 27.035 26.510 27.365 ;
        RECT 54.530 27.035 56.510 27.365 ;
        RECT 84.530 27.035 86.510 27.365 ;
        RECT 114.530 27.035 116.510 27.365 ;
        RECT 9.530 24.315 11.510 24.645 ;
        RECT 39.530 24.315 41.510 24.645 ;
        RECT 69.530 24.315 71.510 24.645 ;
        RECT 99.530 24.315 101.510 24.645 ;
        RECT 24.530 21.595 26.510 21.925 ;
        RECT 54.530 21.595 56.510 21.925 ;
        RECT 84.530 21.595 86.510 21.925 ;
        RECT 114.530 21.595 116.510 21.925 ;
        RECT 9.530 18.875 11.510 19.205 ;
        RECT 39.530 18.875 41.510 19.205 ;
        RECT 69.530 18.875 71.510 19.205 ;
        RECT 99.530 18.875 101.510 19.205 ;
        RECT 24.530 16.155 26.510 16.485 ;
        RECT 54.530 16.155 56.510 16.485 ;
        RECT 84.530 16.155 86.510 16.485 ;
        RECT 114.530 16.155 116.510 16.485 ;
        RECT 9.530 13.435 11.510 13.765 ;
        RECT 39.530 13.435 41.510 13.765 ;
        RECT 69.530 13.435 71.510 13.765 ;
        RECT 99.530 13.435 101.510 13.765 ;
        RECT 24.530 10.715 26.510 11.045 ;
        RECT 54.530 10.715 56.510 11.045 ;
        RECT 84.530 10.715 86.510 11.045 ;
        RECT 114.530 10.715 116.510 11.045 ;
      LAYER met4 ;
        RECT 72.055 104.215 72.385 104.545 ;
        RECT 68.375 98.095 68.705 98.425 ;
        RECT 53.655 93.335 53.985 93.665 ;
        RECT 20.535 85.855 20.865 86.185 ;
        RECT 20.550 75.305 20.850 85.855 ;
        RECT 20.535 74.975 20.865 75.305 ;
        RECT 53.670 72.585 53.970 93.335 ;
        RECT 53.655 72.255 53.985 72.585 ;
        RECT 68.390 51.505 68.690 98.095 ;
        RECT 72.070 73.945 72.370 104.215 ;
        RECT 72.055 73.615 72.385 73.945 ;
        RECT 72.070 55.585 72.370 73.615 ;
        RECT 72.055 55.255 72.385 55.585 ;
        RECT 68.375 51.175 68.705 51.505 ;
  END
END digital_top
END LIBRARY

