VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 853.044495 ;
    ANTENNADIFFAREA 1113.359375 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.805 211.185 14.975 211.375 ;
        RECT 18.485 211.185 18.655 211.375 ;
        RECT 24.005 211.185 24.175 211.375 ;
        RECT 25.845 211.185 26.015 211.375 ;
        RECT 31.365 211.185 31.535 211.375 ;
        RECT 36.885 211.185 37.055 211.375 ;
        RECT 38.725 211.185 38.895 211.375 ;
        RECT 44.245 211.185 44.415 211.375 ;
        RECT 49.765 211.185 49.935 211.375 ;
        RECT 51.605 211.185 51.775 211.375 ;
        RECT 57.125 211.185 57.295 211.375 ;
        RECT 62.645 211.185 62.815 211.375 ;
        RECT 64.485 211.185 64.655 211.375 ;
        RECT 70.005 211.185 70.175 211.375 ;
        RECT 75.525 211.185 75.695 211.375 ;
        RECT 77.365 211.185 77.535 211.375 ;
        RECT 82.885 211.185 83.055 211.375 ;
        RECT 88.405 211.185 88.575 211.375 ;
        RECT 90.245 211.185 90.415 211.375 ;
        RECT 95.765 211.185 95.935 211.375 ;
        RECT 101.285 211.185 101.455 211.375 ;
        RECT 103.125 211.185 103.295 211.375 ;
        RECT 108.645 211.185 108.815 211.375 ;
        RECT 114.165 211.185 114.335 211.375 ;
        RECT 115.140 211.235 115.260 211.345 ;
        RECT 120.605 211.185 120.775 211.375 ;
        RECT 126.125 211.185 126.295 211.375 ;
        RECT 127.505 211.185 127.675 211.375 ;
        RECT 14.665 210.375 16.035 211.185 ;
        RECT 16.045 210.375 18.795 211.185 ;
        RECT 18.805 210.375 24.315 211.185 ;
        RECT 24.335 210.315 24.765 211.100 ;
        RECT 24.785 210.375 26.155 211.185 ;
        RECT 26.165 210.375 31.675 211.185 ;
        RECT 31.685 210.375 37.195 211.185 ;
        RECT 37.215 210.315 37.645 211.100 ;
        RECT 37.665 210.375 39.035 211.185 ;
        RECT 39.045 210.375 44.555 211.185 ;
        RECT 44.565 210.375 50.075 211.185 ;
        RECT 50.095 210.315 50.525 211.100 ;
        RECT 50.545 210.375 51.915 211.185 ;
        RECT 51.925 210.375 57.435 211.185 ;
        RECT 57.445 210.375 62.955 211.185 ;
        RECT 62.975 210.315 63.405 211.100 ;
        RECT 63.425 210.375 64.795 211.185 ;
        RECT 64.805 210.375 70.315 211.185 ;
        RECT 70.325 210.375 75.835 211.185 ;
        RECT 75.855 210.315 76.285 211.100 ;
        RECT 76.305 210.375 77.675 211.185 ;
        RECT 77.685 210.375 83.195 211.185 ;
        RECT 83.205 210.375 88.715 211.185 ;
        RECT 88.735 210.315 89.165 211.100 ;
        RECT 89.185 210.375 90.555 211.185 ;
        RECT 90.565 210.375 96.075 211.185 ;
        RECT 96.085 210.375 101.595 211.185 ;
        RECT 101.615 210.315 102.045 211.100 ;
        RECT 102.065 210.375 103.435 211.185 ;
        RECT 103.445 210.375 108.955 211.185 ;
        RECT 108.965 210.375 114.475 211.185 ;
        RECT 114.495 210.315 114.925 211.100 ;
        RECT 115.405 210.375 120.915 211.185 ;
        RECT 120.925 210.375 126.435 211.185 ;
        RECT 126.445 210.375 127.815 211.185 ;
      LAYER nwell ;
        RECT 14.470 207.155 128.010 209.985 ;
      LAYER pwell ;
        RECT 14.665 205.955 16.035 206.765 ;
        RECT 16.045 205.955 18.795 206.765 ;
        RECT 18.805 205.955 24.315 206.765 ;
        RECT 24.335 206.040 24.765 206.825 ;
        RECT 25.245 205.955 27.995 206.765 ;
        RECT 28.005 205.955 33.515 206.765 ;
        RECT 33.525 205.955 39.035 206.765 ;
        RECT 39.045 205.955 44.555 206.765 ;
        RECT 44.565 205.955 50.075 206.765 ;
        RECT 50.095 206.040 50.525 206.825 ;
        RECT 50.545 205.955 56.055 206.765 ;
        RECT 56.065 205.955 61.575 206.765 ;
        RECT 61.585 205.955 67.095 206.765 ;
        RECT 67.105 205.955 72.615 206.765 ;
        RECT 72.635 205.955 73.985 206.865 ;
        RECT 74.490 206.635 75.835 206.865 ;
        RECT 74.005 205.955 75.835 206.635 ;
        RECT 75.855 206.040 76.285 206.825 ;
        RECT 77.225 205.955 80.335 206.865 ;
        RECT 81.365 205.955 85.035 206.765 ;
        RECT 85.045 205.955 90.555 206.765 ;
        RECT 90.565 205.955 96.075 206.765 ;
        RECT 96.085 205.955 101.595 206.765 ;
        RECT 101.615 206.040 102.045 206.825 ;
        RECT 102.525 205.955 104.355 206.765 ;
        RECT 104.365 205.955 109.875 206.765 ;
        RECT 109.885 205.955 115.395 206.765 ;
        RECT 115.405 205.955 120.915 206.765 ;
        RECT 120.925 205.955 126.435 206.765 ;
        RECT 126.445 205.955 127.815 206.765 ;
        RECT 14.805 205.745 14.975 205.955 ;
        RECT 16.645 205.790 16.805 205.900 ;
        RECT 18.485 205.765 18.655 205.955 ;
        RECT 20.325 205.745 20.495 205.935 ;
        RECT 24.005 205.765 24.175 205.955 ;
        RECT 24.980 205.795 25.100 205.905 ;
        RECT 25.845 205.745 26.015 205.935 ;
        RECT 27.685 205.765 27.855 205.955 ;
        RECT 31.365 205.745 31.535 205.935 ;
        RECT 33.205 205.765 33.375 205.955 ;
        RECT 36.885 205.745 37.055 205.935 ;
        RECT 37.860 205.795 37.980 205.905 ;
        RECT 38.725 205.765 38.895 205.955 ;
        RECT 40.565 205.745 40.735 205.935 ;
        RECT 44.245 205.765 44.415 205.955 ;
        RECT 46.085 205.745 46.255 205.935 ;
        RECT 49.765 205.765 49.935 205.955 ;
        RECT 51.605 205.745 51.775 205.935 ;
        RECT 55.745 205.765 55.915 205.955 ;
        RECT 57.125 205.745 57.295 205.935 ;
        RECT 61.265 205.765 61.435 205.955 ;
        RECT 62.645 205.745 62.815 205.935 ;
        RECT 64.485 205.745 64.655 205.935 ;
        RECT 65.865 205.745 66.035 205.935 ;
        RECT 66.785 205.765 66.955 205.955 ;
        RECT 67.245 205.745 67.415 205.935 ;
        RECT 72.305 205.765 72.475 205.955 ;
        RECT 72.765 205.765 72.935 205.955 ;
        RECT 74.145 205.765 74.315 205.955 ;
        RECT 76.905 205.800 77.065 205.910 ;
        RECT 77.365 205.745 77.535 205.935 ;
        RECT 80.125 205.765 80.295 205.955 ;
        RECT 81.045 205.800 81.205 205.910 ;
        RECT 84.725 205.765 84.895 205.955 ;
        RECT 86.565 205.745 86.735 205.935 ;
        RECT 88.405 205.745 88.575 205.935 ;
        RECT 89.380 205.795 89.500 205.905 ;
        RECT 90.245 205.765 90.415 205.955 ;
        RECT 92.085 205.745 92.255 205.935 ;
        RECT 95.765 205.765 95.935 205.955 ;
        RECT 97.605 205.745 97.775 205.935 ;
        RECT 101.285 205.765 101.455 205.955 ;
        RECT 102.260 205.795 102.380 205.905 ;
        RECT 103.125 205.745 103.295 205.935 ;
        RECT 104.045 205.765 104.215 205.955 ;
        RECT 108.645 205.745 108.815 205.935 ;
        RECT 109.565 205.765 109.735 205.955 ;
        RECT 114.165 205.745 114.335 205.935 ;
        RECT 115.085 205.905 115.255 205.955 ;
        RECT 115.085 205.795 115.260 205.905 ;
        RECT 115.085 205.765 115.255 205.795 ;
        RECT 120.605 205.745 120.775 205.955 ;
        RECT 126.125 205.745 126.295 205.955 ;
        RECT 127.505 205.745 127.675 205.955 ;
        RECT 14.665 204.935 16.035 205.745 ;
        RECT 16.965 204.935 20.635 205.745 ;
        RECT 20.645 204.935 26.155 205.745 ;
        RECT 26.165 204.935 31.675 205.745 ;
        RECT 31.685 204.935 37.195 205.745 ;
        RECT 37.215 204.875 37.645 205.660 ;
        RECT 38.125 204.935 40.875 205.745 ;
        RECT 40.885 204.935 46.395 205.745 ;
        RECT 46.405 204.935 51.915 205.745 ;
        RECT 51.925 204.935 57.435 205.745 ;
        RECT 57.445 204.935 62.955 205.745 ;
        RECT 62.975 204.875 63.405 205.660 ;
        RECT 63.425 204.935 64.795 205.745 ;
        RECT 64.815 204.835 66.165 205.745 ;
        RECT 67.115 204.835 68.465 205.745 ;
        RECT 68.485 205.065 77.675 205.745 ;
        RECT 77.685 205.065 86.875 205.745 ;
        RECT 68.485 204.835 69.405 205.065 ;
        RECT 72.235 204.845 73.165 205.065 ;
        RECT 77.685 204.835 78.605 205.065 ;
        RECT 81.435 204.845 82.365 205.065 ;
        RECT 86.885 204.935 88.715 205.745 ;
        RECT 88.735 204.875 89.165 205.660 ;
        RECT 89.645 204.935 92.395 205.745 ;
        RECT 92.405 204.935 97.915 205.745 ;
        RECT 97.925 204.935 103.435 205.745 ;
        RECT 103.445 204.935 108.955 205.745 ;
        RECT 108.965 204.935 114.475 205.745 ;
        RECT 114.495 204.875 114.925 205.660 ;
        RECT 115.405 204.935 120.915 205.745 ;
        RECT 120.925 204.935 126.435 205.745 ;
        RECT 126.445 204.935 127.815 205.745 ;
      LAYER nwell ;
        RECT 14.470 201.715 128.010 204.545 ;
      LAYER pwell ;
        RECT 14.665 200.515 16.035 201.325 ;
        RECT 16.045 200.515 18.795 201.325 ;
        RECT 18.805 200.515 24.315 201.325 ;
        RECT 24.335 200.600 24.765 201.385 ;
        RECT 25.245 200.515 27.995 201.325 ;
        RECT 28.005 200.515 33.515 201.325 ;
        RECT 33.525 200.515 39.035 201.325 ;
        RECT 39.045 200.515 44.555 201.325 ;
        RECT 44.565 200.515 50.075 201.325 ;
        RECT 50.095 200.600 50.525 201.385 ;
        RECT 50.545 200.515 54.215 201.325 ;
        RECT 54.225 200.515 59.735 201.325 ;
        RECT 64.255 201.195 65.185 201.415 ;
        RECT 67.905 201.195 70.115 201.425 ;
        RECT 59.745 200.515 70.115 201.195 ;
        RECT 70.325 201.195 71.255 201.425 ;
        RECT 70.325 200.515 73.995 201.195 ;
        RECT 74.005 200.515 75.835 201.195 ;
        RECT 75.855 200.600 76.285 201.385 ;
        RECT 76.765 201.195 77.685 201.425 ;
        RECT 79.525 201.195 80.445 201.425 ;
        RECT 83.275 201.195 84.205 201.415 ;
        RECT 76.765 200.515 79.055 201.195 ;
        RECT 79.525 200.515 88.715 201.195 ;
        RECT 88.725 200.515 90.555 201.325 ;
        RECT 90.565 200.515 96.075 201.325 ;
        RECT 96.085 200.515 101.595 201.325 ;
        RECT 101.615 200.600 102.045 201.385 ;
        RECT 102.525 200.515 104.355 201.325 ;
        RECT 104.365 200.515 109.875 201.325 ;
        RECT 109.885 200.515 115.395 201.325 ;
        RECT 115.405 200.515 120.915 201.325 ;
        RECT 120.925 200.515 126.435 201.325 ;
        RECT 126.445 200.515 127.815 201.325 ;
        RECT 14.805 200.305 14.975 200.515 ;
        RECT 16.645 200.350 16.805 200.460 ;
        RECT 18.485 200.325 18.655 200.515 ;
        RECT 20.325 200.305 20.495 200.495 ;
        RECT 24.005 200.325 24.175 200.515 ;
        RECT 24.980 200.355 25.100 200.465 ;
        RECT 25.845 200.305 26.015 200.495 ;
        RECT 27.685 200.325 27.855 200.515 ;
        RECT 31.365 200.305 31.535 200.495 ;
        RECT 33.205 200.325 33.375 200.515 ;
        RECT 36.885 200.305 37.055 200.495 ;
        RECT 37.860 200.355 37.980 200.465 ;
        RECT 38.725 200.325 38.895 200.515 ;
        RECT 40.565 200.305 40.735 200.495 ;
        RECT 44.245 200.325 44.415 200.515 ;
        RECT 46.085 200.305 46.255 200.495 ;
        RECT 49.765 200.325 49.935 200.515 ;
        RECT 51.605 200.305 51.775 200.495 ;
        RECT 53.905 200.325 54.075 200.515 ;
        RECT 57.125 200.305 57.295 200.495 ;
        RECT 59.425 200.325 59.595 200.515 ;
        RECT 59.885 200.325 60.055 200.515 ;
        RECT 62.645 200.305 62.815 200.495 ;
        RECT 63.620 200.355 63.740 200.465 ;
        RECT 67.245 200.305 67.415 200.495 ;
        RECT 68.625 200.305 68.795 200.495 ;
        RECT 70.465 200.305 70.635 200.495 ;
        RECT 73.685 200.325 73.855 200.515 ;
        RECT 75.065 200.305 75.235 200.495 ;
        RECT 75.525 200.325 75.695 200.515 ;
        RECT 76.500 200.355 76.620 200.465 ;
        RECT 78.745 200.305 78.915 200.515 ;
        RECT 79.260 200.355 79.380 200.465 ;
        RECT 81.045 200.325 81.215 200.495 ;
        RECT 81.045 200.305 81.210 200.325 ;
        RECT 82.430 200.305 82.600 200.495 ;
        RECT 82.885 200.305 83.055 200.495 ;
        RECT 84.265 200.305 84.435 200.495 ;
        RECT 86.565 200.305 86.735 200.495 ;
        RECT 88.405 200.305 88.575 200.515 ;
        RECT 89.380 200.355 89.500 200.465 ;
        RECT 90.245 200.325 90.415 200.515 ;
        RECT 91.165 200.305 91.335 200.495 ;
        RECT 95.765 200.325 95.935 200.515 ;
        RECT 96.685 200.305 96.855 200.495 ;
        RECT 101.285 200.325 101.455 200.515 ;
        RECT 102.260 200.355 102.380 200.465 ;
        RECT 104.045 200.325 104.215 200.515 ;
        RECT 105.885 200.305 106.055 200.495 ;
        RECT 108.645 200.305 108.815 200.495 ;
        RECT 109.565 200.325 109.735 200.515 ;
        RECT 114.165 200.305 114.335 200.495 ;
        RECT 115.085 200.465 115.255 200.515 ;
        RECT 115.085 200.355 115.260 200.465 ;
        RECT 115.085 200.325 115.255 200.355 ;
        RECT 120.605 200.305 120.775 200.515 ;
        RECT 126.125 200.305 126.295 200.515 ;
        RECT 127.505 200.305 127.675 200.515 ;
        RECT 14.665 199.495 16.035 200.305 ;
        RECT 16.965 199.495 20.635 200.305 ;
        RECT 20.645 199.495 26.155 200.305 ;
        RECT 26.165 199.495 31.675 200.305 ;
        RECT 31.685 199.495 37.195 200.305 ;
        RECT 37.215 199.435 37.645 200.220 ;
        RECT 38.125 199.495 40.875 200.305 ;
        RECT 40.885 199.495 46.395 200.305 ;
        RECT 46.405 199.495 51.915 200.305 ;
        RECT 51.925 199.495 57.435 200.305 ;
        RECT 57.445 199.495 62.955 200.305 ;
        RECT 62.975 199.435 63.405 200.220 ;
        RECT 63.885 199.495 67.555 200.305 ;
        RECT 67.565 199.525 68.935 200.305 ;
        RECT 68.945 199.625 70.775 200.305 ;
        RECT 70.795 200.265 71.715 200.305 ;
        RECT 70.785 200.075 71.715 200.265 ;
        RECT 73.805 200.075 75.375 200.305 ;
        RECT 70.785 199.715 75.375 200.075 ;
        RECT 70.795 199.625 75.375 199.715 ;
        RECT 75.480 199.625 78.945 200.305 ;
        RECT 79.375 199.625 81.210 200.305 ;
        RECT 70.795 199.395 73.795 199.625 ;
        RECT 75.480 199.395 76.400 199.625 ;
        RECT 79.375 199.395 80.305 199.625 ;
        RECT 81.365 199.395 82.715 200.305 ;
        RECT 82.745 199.525 84.115 200.305 ;
        RECT 84.135 199.395 85.485 200.305 ;
        RECT 85.515 199.395 86.865 200.305 ;
        RECT 86.885 199.495 88.715 200.305 ;
        RECT 88.735 199.435 89.165 200.220 ;
        RECT 89.645 199.495 91.475 200.305 ;
        RECT 91.485 199.495 96.995 200.305 ;
        RECT 97.005 199.625 106.195 200.305 ;
        RECT 97.005 199.395 97.925 199.625 ;
        RECT 100.755 199.405 101.685 199.625 ;
        RECT 106.205 199.495 108.955 200.305 ;
        RECT 108.965 199.495 114.475 200.305 ;
        RECT 114.495 199.435 114.925 200.220 ;
        RECT 115.405 199.495 120.915 200.305 ;
        RECT 120.925 199.495 126.435 200.305 ;
        RECT 126.445 199.495 127.815 200.305 ;
      LAYER nwell ;
        RECT 14.470 196.275 128.010 199.105 ;
      LAYER pwell ;
        RECT 14.665 195.075 16.035 195.885 ;
        RECT 16.045 195.075 18.795 195.885 ;
        RECT 18.805 195.075 24.315 195.885 ;
        RECT 24.335 195.160 24.765 195.945 ;
        RECT 25.245 195.075 27.995 195.885 ;
        RECT 28.005 195.075 33.515 195.885 ;
        RECT 33.525 195.075 39.035 195.885 ;
        RECT 39.045 195.075 44.555 195.885 ;
        RECT 44.565 195.075 50.075 195.885 ;
        RECT 50.095 195.160 50.525 195.945 ;
        RECT 51.005 195.075 52.835 195.885 ;
        RECT 52.855 195.075 54.205 195.985 ;
        RECT 56.880 195.755 57.800 195.985 ;
        RECT 54.335 195.075 57.800 195.755 ;
        RECT 57.905 195.075 63.415 195.885 ;
        RECT 63.425 195.075 68.935 195.885 ;
        RECT 68.945 195.755 69.865 195.985 ;
        RECT 68.945 195.075 71.235 195.755 ;
        RECT 71.245 195.075 74.165 195.985 ;
        RECT 74.465 195.075 75.835 195.885 ;
        RECT 75.855 195.160 76.285 195.945 ;
        RECT 76.305 195.075 79.975 195.885 ;
        RECT 79.985 195.075 85.495 195.885 ;
        RECT 85.875 195.875 86.795 195.985 ;
        RECT 85.875 195.755 88.210 195.875 ;
        RECT 92.875 195.755 93.795 195.975 ;
        RECT 85.875 195.075 95.155 195.755 ;
        RECT 95.165 195.075 97.915 195.885 ;
        RECT 100.580 195.755 101.500 195.985 ;
        RECT 98.035 195.075 101.500 195.755 ;
        RECT 101.615 195.160 102.045 195.945 ;
        RECT 102.065 195.075 104.815 195.885 ;
        RECT 104.825 195.075 110.335 195.885 ;
        RECT 110.345 195.755 111.265 195.985 ;
        RECT 114.095 195.755 115.025 195.975 ;
        RECT 110.345 195.075 119.535 195.755 ;
        RECT 119.545 195.075 120.915 195.885 ;
        RECT 120.925 195.075 126.435 195.885 ;
        RECT 126.445 195.075 127.815 195.885 ;
        RECT 14.805 194.865 14.975 195.075 ;
        RECT 16.645 194.910 16.805 195.020 ;
        RECT 18.485 194.885 18.655 195.075 ;
        RECT 20.325 194.865 20.495 195.055 ;
        RECT 24.005 194.885 24.175 195.075 ;
        RECT 24.980 194.915 25.100 195.025 ;
        RECT 25.845 194.865 26.015 195.055 ;
        RECT 27.685 194.885 27.855 195.075 ;
        RECT 31.365 194.865 31.535 195.055 ;
        RECT 33.205 194.885 33.375 195.075 ;
        RECT 36.885 194.865 37.055 195.055 ;
        RECT 38.265 194.910 38.425 195.020 ;
        RECT 38.725 194.885 38.895 195.075 ;
        RECT 41.945 194.865 42.115 195.055 ;
        RECT 44.245 194.885 44.415 195.075 ;
        RECT 47.465 194.865 47.635 195.055 ;
        RECT 48.845 194.865 49.015 195.055 ;
        RECT 49.305 194.865 49.475 195.055 ;
        RECT 49.765 194.885 49.935 195.075 ;
        RECT 50.740 194.915 50.860 195.025 ;
        RECT 52.525 194.885 52.695 195.075 ;
        RECT 53.905 194.885 54.075 195.075 ;
        RECT 54.365 194.885 54.535 195.075 ;
        RECT 58.965 194.910 59.125 195.020 ;
        RECT 62.645 194.865 62.815 195.055 ;
        RECT 63.105 194.885 63.275 195.075 ;
        RECT 64.945 194.865 65.115 195.055 ;
        RECT 66.325 194.865 66.495 195.055 ;
        RECT 66.840 194.915 66.960 195.025 ;
        RECT 68.625 194.865 68.795 195.075 ;
        RECT 14.665 194.055 16.035 194.865 ;
        RECT 16.965 194.055 20.635 194.865 ;
        RECT 20.645 194.055 26.155 194.865 ;
        RECT 26.165 194.055 31.675 194.865 ;
        RECT 31.685 194.055 37.195 194.865 ;
        RECT 37.215 193.995 37.645 194.780 ;
        RECT 38.585 194.055 42.255 194.865 ;
        RECT 42.265 194.055 47.775 194.865 ;
        RECT 47.795 193.955 49.145 194.865 ;
        RECT 49.165 194.185 58.355 194.865 ;
        RECT 53.675 193.965 54.605 194.185 ;
        RECT 57.435 193.955 58.355 194.185 ;
        RECT 59.285 194.055 62.955 194.865 ;
        RECT 62.975 193.995 63.405 194.780 ;
        RECT 63.425 194.055 65.255 194.865 ;
        RECT 65.275 193.955 66.625 194.865 ;
        RECT 67.105 194.055 68.935 194.865 ;
        RECT 69.085 194.835 69.255 195.055 ;
        RECT 70.925 194.885 71.095 195.075 ;
        RECT 71.390 194.885 71.560 195.075 ;
        RECT 71.210 194.835 72.155 194.865 ;
        RECT 69.085 194.635 72.155 194.835 ;
        RECT 68.945 194.155 72.155 194.635 ;
        RECT 68.945 193.955 69.875 194.155 ;
        RECT 71.210 193.955 72.155 194.155 ;
        RECT 72.165 194.835 73.110 194.865 ;
        RECT 75.065 194.835 75.235 195.055 ;
        RECT 75.525 194.885 75.695 195.075 ;
        RECT 78.745 194.865 78.915 195.055 ;
        RECT 79.665 194.885 79.835 195.075 ;
        RECT 84.265 194.865 84.435 195.055 ;
        RECT 85.185 194.885 85.355 195.075 ;
        RECT 88.130 194.865 88.300 195.055 ;
        RECT 90.245 194.865 90.415 195.055 ;
        RECT 93.005 194.865 93.175 195.055 ;
        RECT 93.465 194.865 93.635 195.055 ;
        RECT 94.845 194.865 95.015 195.075 ;
        RECT 97.605 194.885 97.775 195.075 ;
        RECT 98.065 194.885 98.235 195.075 ;
        RECT 104.505 194.885 104.675 195.075 ;
        RECT 104.965 194.865 105.135 195.055 ;
        RECT 108.645 194.865 108.815 195.055 ;
        RECT 109.105 194.865 109.275 195.055 ;
        RECT 110.025 194.885 110.195 195.075 ;
        RECT 113.890 194.865 114.060 195.055 ;
        RECT 116.005 194.865 116.175 195.055 ;
        RECT 116.925 194.910 117.085 195.020 ;
        RECT 119.225 194.885 119.395 195.075 ;
        RECT 120.605 194.865 120.775 195.075 ;
        RECT 126.125 194.865 126.295 195.075 ;
        RECT 127.505 194.865 127.675 195.075 ;
        RECT 72.165 194.635 75.235 194.835 ;
        RECT 72.165 194.155 75.375 194.635 ;
        RECT 72.165 193.955 73.110 194.155 ;
        RECT 74.445 193.955 75.375 194.155 ;
        RECT 75.385 194.055 79.055 194.865 ;
        RECT 79.065 194.055 84.575 194.865 ;
        RECT 84.815 194.185 88.715 194.865 ;
        RECT 87.785 193.955 88.715 194.185 ;
        RECT 88.735 193.995 89.165 194.780 ;
        RECT 89.195 193.955 90.545 194.865 ;
        RECT 90.565 194.055 93.315 194.865 ;
        RECT 93.335 193.955 94.685 194.865 ;
        RECT 94.705 194.185 103.810 194.865 ;
        RECT 103.905 194.055 105.275 194.865 ;
        RECT 105.285 194.055 108.955 194.865 ;
        RECT 108.975 193.955 110.325 194.865 ;
        RECT 110.575 194.185 114.475 194.865 ;
        RECT 113.545 193.955 114.475 194.185 ;
        RECT 114.495 193.995 114.925 194.780 ;
        RECT 114.955 193.955 116.305 194.865 ;
        RECT 117.245 194.055 120.915 194.865 ;
        RECT 120.925 194.055 126.435 194.865 ;
        RECT 126.445 194.055 127.815 194.865 ;
      LAYER nwell ;
        RECT 14.470 190.835 128.010 193.665 ;
      LAYER pwell ;
        RECT 14.665 189.635 16.035 190.445 ;
        RECT 16.045 189.635 18.795 190.445 ;
        RECT 18.805 189.635 24.315 190.445 ;
        RECT 24.335 189.720 24.765 190.505 ;
        RECT 25.245 189.635 30.755 190.445 ;
        RECT 30.765 189.635 36.275 190.445 ;
        RECT 36.655 190.435 37.575 190.545 ;
        RECT 36.655 190.315 38.990 190.435 ;
        RECT 43.655 190.315 44.575 190.535 ;
        RECT 49.145 190.315 50.075 190.545 ;
        RECT 36.655 189.635 45.935 190.315 ;
        RECT 46.175 189.635 50.075 190.315 ;
        RECT 50.095 189.720 50.525 190.505 ;
        RECT 51.005 189.635 52.375 190.415 ;
        RECT 52.385 190.315 53.305 190.545 ;
        RECT 56.135 190.315 57.065 190.535 ;
        RECT 61.625 190.315 62.965 190.545 ;
        RECT 65.795 190.315 66.725 190.535 ;
        RECT 52.385 189.635 61.575 190.315 ;
        RECT 61.625 189.635 71.235 190.315 ;
        RECT 71.245 189.635 74.355 190.545 ;
        RECT 74.465 189.635 75.835 190.445 ;
        RECT 75.855 189.720 76.285 190.505 ;
        RECT 76.305 189.635 78.595 190.545 ;
        RECT 79.525 189.635 83.195 190.445 ;
        RECT 83.575 190.435 84.495 190.545 ;
        RECT 83.575 190.315 85.910 190.435 ;
        RECT 90.575 190.315 91.495 190.535 ;
        RECT 83.575 189.635 92.855 190.315 ;
        RECT 92.865 189.635 94.235 190.415 ;
        RECT 100.665 190.315 101.595 190.545 ;
        RECT 94.625 189.635 97.050 190.315 ;
        RECT 97.695 189.635 101.595 190.315 ;
        RECT 101.615 189.720 102.045 190.505 ;
        RECT 102.065 189.635 103.435 190.415 ;
        RECT 103.445 189.635 104.815 190.445 ;
        RECT 108.025 190.315 108.955 190.545 ;
        RECT 105.055 189.635 108.955 190.315 ;
        RECT 108.965 190.315 109.885 190.545 ;
        RECT 112.715 190.315 113.645 190.535 ;
        RECT 108.965 189.635 118.155 190.315 ;
        RECT 118.165 189.635 119.535 190.415 ;
        RECT 119.545 189.635 120.915 190.445 ;
        RECT 120.925 189.635 126.435 190.445 ;
        RECT 126.445 189.635 127.815 190.445 ;
        RECT 14.805 189.425 14.975 189.635 ;
        RECT 16.240 189.475 16.360 189.585 ;
        RECT 18.025 189.425 18.195 189.615 ;
        RECT 18.485 189.445 18.655 189.635 ;
        RECT 23.545 189.425 23.715 189.615 ;
        RECT 24.005 189.445 24.175 189.635 ;
        RECT 24.980 189.475 25.100 189.585 ;
        RECT 29.065 189.425 29.235 189.615 ;
        RECT 30.445 189.425 30.615 189.635 ;
        RECT 31.825 189.425 31.995 189.615 ;
        RECT 35.505 189.425 35.675 189.615 ;
        RECT 35.965 189.425 36.135 189.635 ;
        RECT 45.625 189.445 45.795 189.635 ;
        RECT 46.545 189.425 46.715 189.615 ;
        RECT 49.490 189.445 49.660 189.635 ;
        RECT 50.740 189.475 50.860 189.585 ;
        RECT 52.065 189.445 52.235 189.635 ;
        RECT 55.745 189.425 55.915 189.615 ;
        RECT 59.610 189.425 59.780 189.615 ;
        RECT 61.265 189.425 61.435 189.635 ;
        RECT 62.645 189.425 62.815 189.615 ;
        RECT 63.620 189.475 63.740 189.585 ;
        RECT 64.025 189.425 64.195 189.615 ;
        RECT 70.005 189.425 70.175 189.615 ;
        RECT 70.925 189.445 71.095 189.635 ;
        RECT 74.145 189.445 74.315 189.635 ;
        RECT 75.525 189.425 75.695 189.635 ;
        RECT 76.450 189.445 76.620 189.635 ;
        RECT 79.205 189.480 79.365 189.590 ;
        RECT 81.045 189.425 81.215 189.615 ;
        RECT 82.885 189.445 83.055 189.635 ;
        RECT 86.565 189.425 86.735 189.615 ;
        RECT 87.945 189.425 88.115 189.615 ;
        RECT 88.460 189.475 88.580 189.585 ;
        RECT 89.325 189.425 89.495 189.615 ;
        RECT 92.085 189.425 92.255 189.615 ;
        RECT 92.545 189.445 92.715 189.635 ;
        RECT 93.005 189.445 93.175 189.635 ;
        RECT 97.145 189.445 97.315 189.615 ;
        RECT 97.605 189.425 97.775 189.615 ;
        RECT 101.010 189.445 101.180 189.635 ;
        RECT 102.205 189.445 102.375 189.635 ;
        RECT 104.505 189.445 104.675 189.635 ;
        RECT 106.805 189.425 106.975 189.615 ;
        RECT 108.370 189.445 108.540 189.635 ;
        RECT 110.485 189.425 110.655 189.615 ;
        RECT 111.000 189.475 111.120 189.585 ;
        RECT 112.785 189.425 112.955 189.615 ;
        RECT 113.245 189.425 113.415 189.615 ;
        RECT 115.140 189.475 115.260 189.585 ;
        RECT 117.845 189.445 118.015 189.635 ;
        RECT 119.225 189.445 119.395 189.635 ;
        RECT 120.605 189.425 120.775 189.635 ;
        RECT 126.125 189.425 126.295 189.635 ;
        RECT 127.505 189.425 127.675 189.635 ;
        RECT 14.665 188.615 16.035 189.425 ;
        RECT 16.505 188.615 18.335 189.425 ;
        RECT 18.345 188.615 23.855 189.425 ;
        RECT 23.865 188.615 29.375 189.425 ;
        RECT 29.395 188.515 30.745 189.425 ;
        RECT 30.765 188.615 32.135 189.425 ;
        RECT 32.145 188.615 35.815 189.425 ;
        RECT 35.835 188.515 37.185 189.425 ;
        RECT 37.215 188.555 37.645 189.340 ;
        RECT 37.665 188.745 46.855 189.425 ;
        RECT 46.950 188.745 56.055 189.425 ;
        RECT 56.295 188.745 60.195 189.425 ;
        RECT 37.665 188.515 38.585 188.745 ;
        RECT 41.415 188.525 42.345 188.745 ;
        RECT 59.265 188.515 60.195 188.745 ;
        RECT 60.205 188.645 61.575 189.425 ;
        RECT 61.585 188.615 62.955 189.425 ;
        RECT 62.975 188.555 63.405 189.340 ;
        RECT 63.995 188.745 67.460 189.425 ;
        RECT 66.540 188.515 67.460 188.745 ;
        RECT 67.565 188.615 70.315 189.425 ;
        RECT 70.325 188.615 75.835 189.425 ;
        RECT 75.845 188.615 81.355 189.425 ;
        RECT 81.365 188.615 86.875 189.425 ;
        RECT 86.895 188.515 88.245 189.425 ;
        RECT 88.735 188.555 89.165 189.340 ;
        RECT 89.185 188.645 90.555 189.425 ;
        RECT 90.565 188.615 92.395 189.425 ;
        RECT 92.405 188.615 97.915 189.425 ;
        RECT 97.925 188.745 107.115 189.425 ;
        RECT 107.220 188.745 110.685 189.425 ;
        RECT 97.925 188.515 98.845 188.745 ;
        RECT 101.675 188.525 102.605 188.745 ;
        RECT 107.220 188.515 108.140 188.745 ;
        RECT 111.265 188.615 113.095 189.425 ;
        RECT 113.105 188.645 114.475 189.425 ;
        RECT 114.495 188.555 114.925 189.340 ;
        RECT 115.405 188.615 120.915 189.425 ;
        RECT 120.925 188.615 126.435 189.425 ;
        RECT 126.445 188.615 127.815 189.425 ;
      LAYER nwell ;
        RECT 14.470 185.395 128.010 188.225 ;
      LAYER pwell ;
        RECT 14.665 184.195 16.035 185.005 ;
        RECT 16.045 184.195 18.795 185.005 ;
        RECT 18.805 184.195 24.315 185.005 ;
        RECT 24.335 184.280 24.765 185.065 ;
        RECT 24.785 184.195 26.155 185.005 ;
        RECT 26.165 184.875 27.085 185.105 ;
        RECT 29.915 184.875 30.845 185.095 ;
        RECT 26.165 184.195 35.355 184.875 ;
        RECT 35.825 184.195 38.575 185.005 ;
        RECT 38.595 184.195 39.945 185.105 ;
        RECT 43.165 184.875 44.095 185.105 ;
        RECT 40.195 184.195 44.095 184.875 ;
        RECT 44.105 184.875 45.035 185.105 ;
        RECT 44.105 184.195 48.005 184.875 ;
        RECT 48.715 184.195 50.065 185.105 ;
        RECT 50.095 184.280 50.525 185.065 ;
        RECT 50.545 184.875 51.465 185.105 ;
        RECT 54.295 184.875 55.225 185.095 ;
        RECT 50.545 184.195 59.735 184.875 ;
        RECT 60.205 184.195 65.715 185.005 ;
        RECT 65.725 184.195 71.235 185.005 ;
        RECT 71.255 184.875 74.255 185.105 ;
        RECT 71.255 184.785 75.835 184.875 ;
        RECT 71.245 184.425 75.835 184.785 ;
        RECT 71.245 184.235 72.175 184.425 ;
        RECT 71.255 184.195 72.175 184.235 ;
        RECT 74.265 184.195 75.835 184.425 ;
        RECT 75.855 184.280 76.285 185.065 ;
        RECT 76.305 184.195 79.055 185.005 ;
        RECT 79.065 184.195 84.575 185.005 ;
        RECT 87.785 184.875 88.715 185.105 ;
        RECT 84.815 184.195 88.715 184.875 ;
        RECT 88.725 184.195 94.235 185.005 ;
        RECT 96.900 184.875 97.820 185.105 ;
        RECT 94.355 184.195 97.820 184.875 ;
        RECT 98.845 184.195 100.215 184.975 ;
        RECT 100.235 184.195 101.585 185.105 ;
        RECT 101.615 184.280 102.045 185.065 ;
        RECT 102.620 184.875 103.540 185.105 ;
        RECT 109.320 184.875 110.240 185.105 ;
        RECT 113.000 184.875 113.920 185.105 ;
        RECT 102.620 184.195 106.085 184.875 ;
        RECT 106.775 184.195 110.240 184.875 ;
        RECT 110.455 184.195 113.920 184.875 ;
        RECT 114.025 184.195 115.395 185.005 ;
        RECT 115.405 184.195 120.915 185.005 ;
        RECT 120.925 184.195 126.435 185.005 ;
        RECT 126.445 184.195 127.815 185.005 ;
        RECT 14.805 183.985 14.975 184.195 ;
        RECT 16.240 184.035 16.360 184.145 ;
        RECT 18.485 184.005 18.655 184.195 ;
        RECT 21.705 183.985 21.875 184.175 ;
        RECT 22.165 183.985 22.335 184.175 ;
        RECT 24.005 184.005 24.175 184.195 ;
        RECT 25.845 184.005 26.015 184.195 ;
        RECT 26.765 183.985 26.935 184.175 ;
        RECT 27.225 183.985 27.395 184.175 ;
        RECT 31.180 183.985 31.350 184.175 ;
        RECT 35.045 184.145 35.215 184.195 ;
        RECT 35.045 184.035 35.220 184.145 ;
        RECT 35.560 184.035 35.680 184.145 ;
        RECT 35.045 184.005 35.215 184.035 ;
        RECT 36.885 183.985 37.055 184.175 ;
        RECT 37.805 183.985 37.975 184.175 ;
        RECT 38.265 184.005 38.435 184.195 ;
        RECT 38.725 184.005 38.895 184.195 ;
        RECT 41.485 183.985 41.655 184.175 ;
        RECT 43.510 184.005 43.680 184.195 ;
        RECT 44.520 184.005 44.690 184.195 ;
        RECT 45.165 183.985 45.335 184.175 ;
        RECT 48.440 184.035 48.560 184.145 ;
        RECT 48.845 184.005 49.015 184.195 ;
        RECT 49.765 183.985 49.935 184.175 ;
        RECT 51.145 183.985 51.315 184.175 ;
        RECT 51.605 183.985 51.775 184.175 ;
        RECT 55.745 183.985 55.915 184.175 ;
        RECT 56.260 184.035 56.380 184.145 ;
        RECT 58.965 183.985 59.135 184.175 ;
        RECT 59.425 184.005 59.595 184.195 ;
        RECT 59.940 184.035 60.060 184.145 ;
        RECT 60.345 183.985 60.515 184.175 ;
        RECT 60.860 184.035 60.980 184.145 ;
        RECT 62.645 183.985 62.815 184.175 ;
        RECT 63.620 184.035 63.740 184.145 ;
        RECT 65.405 184.005 65.575 184.195 ;
        RECT 66.325 183.985 66.495 184.175 ;
        RECT 66.785 184.005 66.955 184.175 ;
        RECT 66.885 183.985 66.955 184.005 ;
        RECT 70.005 183.985 70.175 184.175 ;
        RECT 70.925 184.005 71.095 184.195 ;
        RECT 75.525 184.005 75.695 184.195 ;
        RECT 78.285 184.005 78.455 184.175 ;
        RECT 78.745 184.005 78.915 184.195 ;
        RECT 79.205 184.030 79.365 184.140 ;
        RECT 84.265 184.005 84.435 184.195 ;
        RECT 88.130 184.005 88.300 184.195 ;
        RECT 78.285 183.985 78.355 184.005 ;
        RECT 88.405 183.985 88.575 184.175 ;
        RECT 90.245 183.985 90.415 184.175 ;
        RECT 91.625 183.985 91.795 184.175 ;
        RECT 93.925 184.005 94.095 184.195 ;
        RECT 94.385 184.005 94.555 184.195 ;
        RECT 95.305 183.985 95.475 184.175 ;
        RECT 98.525 184.040 98.685 184.150 ;
        RECT 98.985 184.005 99.155 184.195 ;
        RECT 99.170 183.985 99.340 184.175 ;
        RECT 100.365 184.005 100.535 184.195 ;
        RECT 102.205 184.145 102.375 184.175 ;
        RECT 102.205 184.035 102.380 184.145 ;
        RECT 102.205 183.985 102.375 184.035 ;
        RECT 105.885 184.005 106.055 184.195 ;
        RECT 106.805 184.175 106.975 184.195 ;
        RECT 106.070 183.985 106.240 184.175 ;
        RECT 106.400 184.035 106.520 184.145 ;
        RECT 106.805 184.005 106.980 184.175 ;
        RECT 110.485 184.005 110.655 184.195 ;
        RECT 106.810 183.985 106.980 184.005 ;
        RECT 113.890 183.985 114.060 184.175 ;
        RECT 115.085 184.005 115.255 184.195 ;
        RECT 115.545 184.030 115.705 184.140 ;
        RECT 120.605 184.005 120.775 184.195 ;
        RECT 124.745 183.985 124.915 184.175 ;
        RECT 126.125 183.985 126.295 184.195 ;
        RECT 127.505 183.985 127.675 184.195 ;
        RECT 14.665 183.175 16.035 183.985 ;
        RECT 16.505 183.175 22.015 183.985 ;
        RECT 22.025 183.205 23.395 183.985 ;
        RECT 23.500 183.305 26.965 183.985 ;
        RECT 27.195 183.305 30.660 183.985 ;
        RECT 23.500 183.075 24.420 183.305 ;
        RECT 29.740 183.075 30.660 183.305 ;
        RECT 30.765 183.305 34.665 183.985 ;
        RECT 30.765 183.075 31.695 183.305 ;
        RECT 35.365 183.175 37.195 183.985 ;
        RECT 37.215 183.115 37.645 183.900 ;
        RECT 37.775 183.305 41.240 183.985 ;
        RECT 41.455 183.305 44.920 183.985 ;
        RECT 45.135 183.305 48.600 183.985 ;
        RECT 40.320 183.075 41.240 183.305 ;
        RECT 44.000 183.075 44.920 183.305 ;
        RECT 47.680 183.075 48.600 183.305 ;
        RECT 48.705 183.205 50.075 183.985 ;
        RECT 50.085 183.205 51.455 183.985 ;
        RECT 51.465 183.205 52.835 183.985 ;
        RECT 52.845 183.075 56.005 183.985 ;
        RECT 56.525 183.175 59.275 183.985 ;
        RECT 59.295 183.075 60.645 183.985 ;
        RECT 61.125 183.175 62.955 183.985 ;
        RECT 62.975 183.115 63.405 183.900 ;
        RECT 63.885 183.175 66.635 183.985 ;
        RECT 66.885 183.755 69.155 183.985 ;
        RECT 69.865 183.755 74.290 183.985 ;
        RECT 76.085 183.755 78.355 183.985 ;
        RECT 66.885 183.075 69.640 183.755 ;
        RECT 69.865 183.075 75.230 183.755 ;
        RECT 75.600 183.075 78.355 183.755 ;
        RECT 79.525 183.305 88.715 183.985 ;
        RECT 79.525 183.075 80.445 183.305 ;
        RECT 83.275 183.085 84.205 183.305 ;
        RECT 88.735 183.115 89.165 183.900 ;
        RECT 89.195 183.075 90.545 183.985 ;
        RECT 90.565 183.175 91.935 183.985 ;
        RECT 91.945 183.175 95.615 183.985 ;
        RECT 95.855 183.305 99.755 183.985 ;
        RECT 98.825 183.075 99.755 183.305 ;
        RECT 99.765 183.175 102.515 183.985 ;
        RECT 102.755 183.305 106.655 183.985 ;
        RECT 105.725 183.075 106.655 183.305 ;
        RECT 106.665 183.075 110.140 183.985 ;
        RECT 110.575 183.305 114.475 183.985 ;
        RECT 113.545 183.075 114.475 183.305 ;
        RECT 114.495 183.115 114.925 183.900 ;
        RECT 115.865 183.305 125.055 183.985 ;
        RECT 115.865 183.075 116.785 183.305 ;
        RECT 119.615 183.085 120.545 183.305 ;
        RECT 125.065 183.175 126.435 183.985 ;
        RECT 126.445 183.175 127.815 183.985 ;
      LAYER nwell ;
        RECT 14.470 179.955 128.010 182.785 ;
      LAYER pwell ;
        RECT 14.665 178.755 16.035 179.565 ;
        RECT 16.045 178.755 18.795 179.565 ;
        RECT 18.805 178.755 24.315 179.565 ;
        RECT 24.335 178.840 24.765 179.625 ;
        RECT 29.295 179.435 30.225 179.655 ;
        RECT 33.055 179.435 33.975 179.665 ;
        RECT 24.785 178.755 33.975 179.435 ;
        RECT 34.080 179.435 35.000 179.665 ;
        RECT 34.080 178.755 37.545 179.435 ;
        RECT 38.125 178.755 41.600 179.665 ;
        RECT 42.265 178.755 45.740 179.665 ;
        RECT 49.145 179.435 50.075 179.665 ;
        RECT 46.175 178.755 50.075 179.435 ;
        RECT 50.095 178.840 50.525 179.625 ;
        RECT 53.200 179.435 54.120 179.665 ;
        RECT 50.655 178.755 54.120 179.435 ;
        RECT 54.225 178.755 56.055 179.565 ;
        RECT 56.065 179.435 56.995 179.665 ;
        RECT 56.065 178.755 59.965 179.435 ;
        RECT 60.215 178.755 62.955 179.435 ;
        RECT 62.965 178.755 65.715 179.565 ;
        RECT 65.735 178.755 67.085 179.665 ;
        RECT 67.105 179.435 68.450 179.665 ;
        RECT 67.105 178.755 68.935 179.435 ;
        RECT 68.945 178.755 71.685 179.435 ;
        RECT 71.945 178.985 74.700 179.665 ;
        RECT 71.945 178.755 74.215 178.985 ;
        RECT 75.855 178.840 76.285 179.625 ;
        RECT 78.960 179.435 79.880 179.665 ;
        RECT 76.415 178.755 79.880 179.435 ;
        RECT 80.180 178.755 83.655 179.665 ;
        RECT 83.665 178.755 85.495 179.565 ;
        RECT 88.705 179.435 89.635 179.665 ;
        RECT 85.735 178.755 89.635 179.435 ;
        RECT 89.645 178.755 91.015 179.535 ;
        RECT 91.035 178.755 92.385 179.665 ;
        RECT 92.405 179.435 93.325 179.665 ;
        RECT 96.155 179.435 97.085 179.655 ;
        RECT 92.405 178.755 101.595 179.435 ;
        RECT 101.615 178.840 102.045 179.625 ;
        RECT 102.160 179.435 103.080 179.665 ;
        RECT 105.840 179.435 106.760 179.665 ;
        RECT 102.160 178.755 105.625 179.435 ;
        RECT 105.840 178.755 109.305 179.435 ;
        RECT 109.895 178.755 111.245 179.665 ;
        RECT 111.265 179.435 112.185 179.665 ;
        RECT 115.015 179.435 115.945 179.655 ;
        RECT 111.265 178.755 120.455 179.435 ;
        RECT 120.475 178.755 121.825 179.665 ;
        RECT 121.845 178.755 123.215 179.535 ;
        RECT 123.685 178.755 126.435 179.565 ;
        RECT 126.445 178.755 127.815 179.565 ;
        RECT 14.805 178.545 14.975 178.755 ;
        RECT 18.485 178.565 18.655 178.755 ;
        RECT 19.405 178.545 19.575 178.735 ;
        RECT 24.005 178.565 24.175 178.755 ;
        RECT 24.925 178.545 25.095 178.755 ;
        RECT 26.305 178.545 26.475 178.735 ;
        RECT 26.765 178.545 26.935 178.735 ;
        RECT 36.885 178.545 37.055 178.735 ;
        RECT 37.345 178.565 37.515 178.755 ;
        RECT 37.860 178.595 37.980 178.705 ;
        RECT 38.270 178.565 38.440 178.755 ;
        RECT 41.210 178.545 41.380 178.735 ;
        RECT 42.000 178.595 42.120 178.705 ;
        RECT 42.410 178.700 42.580 178.755 ;
        RECT 42.405 178.590 42.580 178.700 ;
        RECT 42.410 178.565 42.580 178.590 ;
        RECT 42.865 178.545 43.035 178.735 ;
        RECT 49.490 178.565 49.660 178.755 ;
        RECT 49.760 178.545 49.930 178.735 ;
        RECT 50.225 178.545 50.395 178.735 ;
        RECT 50.685 178.565 50.855 178.755 ;
        RECT 55.745 178.565 55.915 178.755 ;
        RECT 56.480 178.565 56.650 178.755 ;
        RECT 62.645 178.545 62.815 178.755 ;
        RECT 64.485 178.545 64.655 178.735 ;
        RECT 65.405 178.565 65.575 178.755 ;
        RECT 65.865 178.565 66.035 178.755 ;
        RECT 67.245 178.545 67.415 178.735 ;
        RECT 68.625 178.565 68.795 178.755 ;
        RECT 69.085 178.545 69.255 178.755 ;
        RECT 71.945 178.735 72.015 178.755 ;
        RECT 69.545 178.545 69.715 178.735 ;
        RECT 71.385 178.545 71.555 178.735 ;
        RECT 71.845 178.565 72.015 178.735 ;
        RECT 75.525 178.545 75.695 178.735 ;
        RECT 76.040 178.595 76.160 178.705 ;
        RECT 76.445 178.565 76.615 178.755 ;
        RECT 79.660 178.545 79.830 178.735 ;
        RECT 80.130 178.545 80.300 178.735 ;
        RECT 83.340 178.565 83.510 178.755 ;
        RECT 84.725 178.545 84.895 178.735 ;
        RECT 85.185 178.545 85.355 178.755 ;
        RECT 89.050 178.565 89.220 178.755 ;
        RECT 90.705 178.565 90.875 178.755 ;
        RECT 91.165 178.565 91.335 178.755 ;
        RECT 92.545 178.545 92.715 178.735 ;
        RECT 98.065 178.545 98.235 178.735 ;
        RECT 101.285 178.565 101.455 178.755 ;
        RECT 101.740 178.545 101.910 178.735 ;
        RECT 103.125 178.545 103.295 178.735 ;
        RECT 104.505 178.545 104.675 178.735 ;
        RECT 104.970 178.545 105.140 178.735 ;
        RECT 105.425 178.565 105.595 178.755 ;
        RECT 109.105 178.565 109.275 178.755 ;
        RECT 109.620 178.595 109.740 178.705 ;
        RECT 110.025 178.545 110.195 178.755 ;
        RECT 113.890 178.545 114.060 178.735 ;
        RECT 116.465 178.545 116.635 178.735 ;
        RECT 116.925 178.545 117.095 178.735 ;
        RECT 120.145 178.565 120.315 178.755 ;
        RECT 120.605 178.545 120.775 178.755 ;
        RECT 121.985 178.565 122.155 178.755 ;
        RECT 123.420 178.595 123.540 178.705 ;
        RECT 126.125 178.545 126.295 178.755 ;
        RECT 127.505 178.545 127.675 178.755 ;
        RECT 14.665 177.735 16.035 178.545 ;
        RECT 16.045 177.735 19.715 178.545 ;
        RECT 19.725 177.735 25.235 178.545 ;
        RECT 25.255 177.635 26.605 178.545 ;
        RECT 26.635 177.635 27.985 178.545 ;
        RECT 28.005 177.865 37.195 178.545 ;
        RECT 28.005 177.635 28.925 177.865 ;
        RECT 31.755 177.645 32.685 177.865 ;
        RECT 37.215 177.675 37.645 178.460 ;
        RECT 37.895 177.865 41.795 178.545 ;
        RECT 42.835 177.865 46.300 178.545 ;
        RECT 40.865 177.635 41.795 177.865 ;
        RECT 45.380 177.635 46.300 177.865 ;
        RECT 46.600 177.635 50.075 178.545 ;
        RECT 50.195 177.865 53.660 178.545 ;
        RECT 52.740 177.635 53.660 177.865 ;
        RECT 53.765 177.865 62.955 178.545 ;
        RECT 53.765 177.635 54.685 177.865 ;
        RECT 57.515 177.645 58.445 177.865 ;
        RECT 62.975 177.675 63.405 178.460 ;
        RECT 63.425 177.765 64.795 178.545 ;
        RECT 64.805 177.735 67.555 178.545 ;
        RECT 67.565 177.865 69.395 178.545 ;
        RECT 69.405 177.865 71.235 178.545 ;
        RECT 71.245 177.865 73.075 178.545 ;
        RECT 67.565 177.635 68.910 177.865 ;
        RECT 69.890 177.635 71.235 177.865 ;
        RECT 71.730 177.635 73.075 177.865 ;
        RECT 73.115 177.635 75.835 178.545 ;
        RECT 76.500 177.635 79.975 178.545 ;
        RECT 79.985 177.635 83.460 178.545 ;
        RECT 83.665 177.735 85.035 178.545 ;
        RECT 85.155 177.865 88.620 178.545 ;
        RECT 87.700 177.635 88.620 177.865 ;
        RECT 88.735 177.675 89.165 178.460 ;
        RECT 89.185 177.735 92.855 178.545 ;
        RECT 92.865 177.735 98.375 178.545 ;
        RECT 98.580 177.635 102.055 178.545 ;
        RECT 102.065 177.765 103.435 178.545 ;
        RECT 103.445 177.735 104.815 178.545 ;
        RECT 104.825 177.635 108.300 178.545 ;
        RECT 108.505 177.735 110.335 178.545 ;
        RECT 110.575 177.865 114.475 178.545 ;
        RECT 113.545 177.635 114.475 177.865 ;
        RECT 114.495 177.675 114.925 178.460 ;
        RECT 114.945 177.735 116.775 178.545 ;
        RECT 116.785 177.765 118.155 178.545 ;
        RECT 118.165 177.735 120.915 178.545 ;
        RECT 120.925 177.735 126.435 178.545 ;
        RECT 126.445 177.735 127.815 178.545 ;
      LAYER nwell ;
        RECT 14.470 174.515 128.010 177.345 ;
      LAYER pwell ;
        RECT 14.665 173.315 16.035 174.125 ;
        RECT 16.045 173.315 18.795 174.125 ;
        RECT 18.805 173.315 24.315 174.125 ;
        RECT 24.335 173.400 24.765 174.185 ;
        RECT 25.705 173.315 27.075 174.095 ;
        RECT 29.740 173.995 30.660 174.225 ;
        RECT 27.195 173.315 30.660 173.995 ;
        RECT 30.765 173.995 31.695 174.225 ;
        RECT 30.765 173.315 34.665 173.995 ;
        RECT 35.560 173.315 39.035 174.225 ;
        RECT 39.045 173.315 42.520 174.225 ;
        RECT 42.920 173.315 46.395 174.225 ;
        RECT 49.060 173.995 49.980 174.225 ;
        RECT 46.515 173.315 49.980 173.995 ;
        RECT 50.095 173.400 50.525 174.185 ;
        RECT 50.545 173.315 53.295 174.125 ;
        RECT 56.505 173.995 57.435 174.225 ;
        RECT 53.535 173.315 57.435 173.995 ;
        RECT 57.445 173.995 58.365 174.225 ;
        RECT 61.195 173.995 62.125 174.215 ;
        RECT 57.445 173.315 66.635 173.995 ;
        RECT 66.645 173.315 68.475 174.125 ;
        RECT 68.485 173.315 71.095 174.225 ;
        RECT 71.245 173.995 72.590 174.225 ;
        RECT 71.245 173.315 73.075 173.995 ;
        RECT 73.085 173.315 75.835 174.125 ;
        RECT 75.855 173.400 76.285 174.185 ;
        RECT 77.225 173.315 80.895 174.125 ;
        RECT 80.905 173.315 84.380 174.225 ;
        RECT 85.045 173.315 90.555 174.125 ;
        RECT 90.565 173.315 96.075 174.125 ;
        RECT 96.085 173.315 101.595 174.125 ;
        RECT 101.615 173.400 102.045 174.185 ;
        RECT 102.065 173.315 103.895 174.125 ;
        RECT 104.100 173.315 107.575 174.225 ;
        RECT 107.585 173.315 111.060 174.225 ;
        RECT 111.265 173.315 112.635 174.125 ;
        RECT 112.645 173.315 118.155 174.125 ;
        RECT 118.175 173.315 119.525 174.225 ;
        RECT 119.545 173.315 120.915 174.125 ;
        RECT 120.925 173.315 126.435 174.125 ;
        RECT 126.445 173.315 127.815 174.125 ;
        RECT 14.805 173.105 14.975 173.315 ;
        RECT 16.645 173.150 16.805 173.260 ;
        RECT 18.485 173.125 18.655 173.315 ;
        RECT 20.325 173.105 20.495 173.295 ;
        RECT 24.005 173.125 24.175 173.315 ;
        RECT 25.385 173.160 25.545 173.270 ;
        RECT 25.845 173.105 26.015 173.295 ;
        RECT 26.765 173.125 26.935 173.315 ;
        RECT 27.225 173.125 27.395 173.315 ;
        RECT 31.180 173.125 31.350 173.315 ;
        RECT 31.365 173.105 31.535 173.295 ;
        RECT 35.100 173.155 35.220 173.265 ;
        RECT 36.885 173.105 37.055 173.295 ;
        RECT 37.810 173.105 37.980 173.295 ;
        RECT 38.720 173.125 38.890 173.315 ;
        RECT 39.190 173.125 39.360 173.315 ;
        RECT 41.540 173.155 41.660 173.265 ;
        RECT 42.865 173.105 43.035 173.295 ;
        RECT 43.785 173.150 43.945 173.260 ;
        RECT 44.250 173.105 44.420 173.295 ;
        RECT 46.080 173.125 46.250 173.315 ;
        RECT 46.545 173.125 46.715 173.315 ;
        RECT 47.930 173.105 48.100 173.295 ;
        RECT 51.610 173.105 51.780 173.295 ;
        RECT 52.985 173.125 53.155 173.315 ;
        RECT 56.205 173.105 56.375 173.295 ;
        RECT 56.850 173.125 57.020 173.315 ;
        RECT 59.885 173.105 60.055 173.295 ;
        RECT 61.265 173.105 61.435 173.295 ;
        RECT 61.725 173.105 61.895 173.295 ;
        RECT 63.620 173.155 63.740 173.265 ;
        RECT 65.405 173.105 65.575 173.295 ;
        RECT 66.325 173.125 66.495 173.315 ;
        RECT 68.165 173.125 68.335 173.315 ;
        RECT 68.630 173.125 68.800 173.315 ;
        RECT 70.925 173.105 71.095 173.295 ;
        RECT 72.765 173.125 72.935 173.315 ;
        RECT 75.525 173.125 75.695 173.315 ;
        RECT 76.445 173.105 76.615 173.295 ;
        RECT 76.905 173.160 77.065 173.270 ;
        RECT 80.585 173.125 80.755 173.315 ;
        RECT 81.050 173.125 81.220 173.315 ;
        RECT 81.965 173.105 82.135 173.295 ;
        RECT 82.430 173.105 82.600 173.295 ;
        RECT 84.780 173.155 84.900 173.265 ;
        RECT 85.185 173.105 85.355 173.295 ;
        RECT 89.380 173.155 89.500 173.265 ;
        RECT 89.785 173.105 89.955 173.295 ;
        RECT 90.245 173.125 90.415 173.315 ;
        RECT 95.765 173.125 95.935 173.315 ;
        RECT 99.905 173.105 100.075 173.295 ;
        RECT 100.825 173.150 100.985 173.260 ;
        RECT 101.285 173.125 101.455 173.315 ;
        RECT 103.585 173.125 103.755 173.315 ;
        RECT 106.345 173.105 106.515 173.295 ;
        RECT 107.260 173.125 107.430 173.315 ;
        RECT 107.730 173.295 107.900 173.315 ;
        RECT 107.725 173.125 107.900 173.295 ;
        RECT 107.725 173.105 107.895 173.125 ;
        RECT 111.400 173.105 111.570 173.295 ;
        RECT 112.325 173.125 112.495 173.315 ;
        RECT 112.785 173.105 112.955 173.295 ;
        RECT 113.245 173.105 113.415 173.295 ;
        RECT 115.545 173.150 115.705 173.260 ;
        RECT 117.845 173.125 118.015 173.315 ;
        RECT 118.305 173.125 118.475 173.315 ;
        RECT 120.605 173.125 120.775 173.315 ;
        RECT 124.745 173.105 124.915 173.295 ;
        RECT 126.125 173.105 126.295 173.315 ;
        RECT 127.505 173.105 127.675 173.315 ;
        RECT 14.665 172.295 16.035 173.105 ;
        RECT 16.965 172.295 20.635 173.105 ;
        RECT 20.645 172.295 26.155 173.105 ;
        RECT 26.165 172.295 31.675 173.105 ;
        RECT 31.685 172.295 37.195 173.105 ;
        RECT 37.215 172.235 37.645 173.020 ;
        RECT 37.665 172.195 41.140 173.105 ;
        RECT 41.805 172.325 43.175 173.105 ;
        RECT 44.105 172.195 47.580 173.105 ;
        RECT 47.785 172.195 51.260 173.105 ;
        RECT 51.465 172.195 54.940 173.105 ;
        RECT 55.145 172.295 56.515 173.105 ;
        RECT 56.525 172.295 60.195 173.105 ;
        RECT 60.215 172.195 61.565 173.105 ;
        RECT 61.585 172.325 62.955 173.105 ;
        RECT 62.975 172.235 63.405 173.020 ;
        RECT 63.885 172.295 65.715 173.105 ;
        RECT 65.725 172.295 71.235 173.105 ;
        RECT 71.245 172.295 76.755 173.105 ;
        RECT 76.765 172.295 82.275 173.105 ;
        RECT 82.285 172.195 84.895 173.105 ;
        RECT 85.155 172.425 88.620 173.105 ;
        RECT 87.700 172.195 88.620 172.425 ;
        RECT 88.735 172.235 89.165 173.020 ;
        RECT 89.655 172.195 91.005 173.105 ;
        RECT 91.025 172.425 100.215 173.105 ;
        RECT 91.025 172.195 91.945 172.425 ;
        RECT 94.775 172.205 95.705 172.425 ;
        RECT 101.145 172.295 106.655 173.105 ;
        RECT 106.675 172.195 108.025 173.105 ;
        RECT 108.240 172.195 111.715 173.105 ;
        RECT 111.725 172.295 113.095 173.105 ;
        RECT 113.115 172.195 114.465 173.105 ;
        RECT 114.495 172.235 114.925 173.020 ;
        RECT 115.865 172.425 125.055 173.105 ;
        RECT 115.865 172.195 116.785 172.425 ;
        RECT 119.615 172.205 120.545 172.425 ;
        RECT 125.065 172.295 126.435 173.105 ;
        RECT 126.445 172.295 127.815 173.105 ;
      LAYER nwell ;
        RECT 14.470 169.075 128.010 171.905 ;
      LAYER pwell ;
        RECT 14.665 167.875 16.035 168.685 ;
        RECT 16.045 167.875 18.795 168.685 ;
        RECT 18.805 167.875 24.315 168.685 ;
        RECT 24.335 167.960 24.765 168.745 ;
        RECT 25.245 167.875 27.075 168.685 ;
        RECT 27.095 167.875 28.445 168.785 ;
        RECT 28.925 167.875 32.595 168.685 ;
        RECT 32.615 167.875 33.965 168.785 ;
        RECT 33.985 167.875 35.355 168.685 ;
        RECT 35.450 167.875 44.555 168.555 ;
        RECT 44.565 167.875 50.075 168.685 ;
        RECT 50.095 167.960 50.525 168.745 ;
        RECT 50.545 167.875 51.915 168.685 ;
        RECT 51.925 167.875 57.435 168.685 ;
        RECT 57.445 167.875 62.955 168.685 ;
        RECT 62.965 167.875 68.475 168.685 ;
        RECT 68.485 168.555 69.830 168.785 ;
        RECT 70.325 168.555 71.670 168.785 ;
        RECT 68.485 167.875 70.315 168.555 ;
        RECT 70.325 167.875 72.155 168.555 ;
        RECT 72.165 167.875 75.835 168.685 ;
        RECT 75.855 167.960 76.285 168.745 ;
        RECT 79.505 168.555 80.435 168.785 ;
        RECT 76.535 167.875 80.435 168.555 ;
        RECT 80.815 168.675 81.735 168.785 ;
        RECT 80.815 168.555 83.150 168.675 ;
        RECT 87.815 168.555 88.735 168.775 ;
        RECT 80.815 167.875 90.095 168.555 ;
        RECT 90.105 167.875 91.475 168.685 ;
        RECT 94.685 168.555 95.615 168.785 ;
        RECT 91.715 167.875 95.615 168.555 ;
        RECT 96.085 167.875 97.455 168.655 ;
        RECT 97.925 167.875 101.595 168.685 ;
        RECT 101.615 167.960 102.045 168.745 ;
        RECT 102.985 168.555 103.905 168.785 ;
        RECT 106.735 168.555 107.665 168.775 ;
        RECT 112.645 168.555 113.575 168.785 ;
        RECT 116.880 168.555 117.800 168.785 ;
        RECT 102.985 167.875 112.175 168.555 ;
        RECT 112.645 167.875 116.545 168.555 ;
        RECT 116.880 167.875 120.345 168.555 ;
        RECT 120.465 167.875 121.835 168.655 ;
        RECT 121.845 167.875 123.675 168.555 ;
        RECT 123.685 167.875 126.435 168.685 ;
        RECT 126.445 167.875 127.815 168.685 ;
        RECT 14.805 167.665 14.975 167.875 ;
        RECT 17.565 167.665 17.735 167.855 ;
        RECT 18.485 167.685 18.655 167.875 ;
        RECT 23.085 167.665 23.255 167.855 ;
        RECT 23.545 167.665 23.715 167.855 ;
        RECT 24.005 167.685 24.175 167.875 ;
        RECT 24.980 167.715 25.100 167.825 ;
        RECT 26.765 167.685 26.935 167.875 ;
        RECT 27.225 167.685 27.395 167.875 ;
        RECT 28.660 167.715 28.780 167.825 ;
        RECT 32.285 167.685 32.455 167.875 ;
        RECT 33.665 167.665 33.835 167.875 ;
        RECT 35.045 167.685 35.215 167.875 ;
        RECT 36.885 167.665 37.055 167.855 ;
        RECT 37.805 167.665 37.975 167.855 ;
        RECT 39.185 167.665 39.355 167.855 ;
        RECT 44.245 167.685 44.415 167.875 ;
        RECT 46.085 167.665 46.255 167.855 ;
        RECT 47.005 167.710 47.165 167.820 ;
        RECT 49.765 167.685 49.935 167.875 ;
        RECT 51.605 167.685 51.775 167.875 ;
        RECT 56.205 167.665 56.375 167.855 ;
        RECT 57.125 167.685 57.295 167.875 ;
        RECT 62.645 167.855 62.815 167.875 ;
        RECT 58.045 167.665 58.215 167.855 ;
        RECT 59.425 167.665 59.595 167.855 ;
        RECT 59.940 167.715 60.060 167.825 ;
        RECT 62.640 167.685 62.815 167.855 ;
        RECT 62.640 167.665 62.810 167.685 ;
        RECT 64.945 167.665 65.115 167.855 ;
        RECT 67.705 167.665 67.875 167.855 ;
        RECT 68.165 167.665 68.335 167.875 ;
        RECT 70.005 167.685 70.175 167.875 ;
        RECT 70.925 167.665 71.095 167.855 ;
        RECT 71.845 167.685 72.015 167.875 ;
        RECT 75.065 167.665 75.235 167.855 ;
        RECT 75.525 167.685 75.695 167.875 ;
        RECT 79.850 167.685 80.020 167.875 ;
        RECT 84.725 167.665 84.895 167.855 ;
        RECT 86.105 167.665 86.275 167.855 ;
        RECT 87.485 167.665 87.655 167.855 ;
        RECT 88.405 167.710 88.565 167.820 ;
        RECT 89.380 167.715 89.500 167.825 ;
        RECT 89.785 167.685 89.955 167.875 ;
        RECT 91.165 167.685 91.335 167.875 ;
        RECT 93.005 167.665 93.175 167.855 ;
        RECT 95.030 167.685 95.200 167.875 ;
        RECT 95.820 167.715 95.940 167.825 ;
        RECT 96.225 167.685 96.395 167.875 ;
        RECT 96.870 167.665 97.040 167.855 ;
        RECT 97.660 167.715 97.780 167.825 ;
        RECT 101.285 167.685 101.455 167.875 ;
        RECT 102.665 167.720 102.825 167.830 ;
        RECT 106.805 167.665 106.975 167.855 ;
        RECT 107.265 167.665 107.435 167.855 ;
        RECT 110.945 167.665 111.115 167.855 ;
        RECT 111.865 167.685 112.035 167.875 ;
        RECT 112.380 167.715 112.500 167.825 ;
        RECT 113.060 167.685 113.230 167.875 ;
        RECT 115.545 167.710 115.705 167.820 ;
        RECT 120.145 167.685 120.315 167.875 ;
        RECT 120.605 167.685 120.775 167.875 ;
        RECT 123.365 167.685 123.535 167.875 ;
        RECT 124.745 167.665 124.915 167.855 ;
        RECT 126.125 167.665 126.295 167.875 ;
        RECT 127.505 167.665 127.675 167.875 ;
        RECT 14.665 166.855 16.035 167.665 ;
        RECT 16.045 166.855 17.875 167.665 ;
        RECT 17.885 166.855 23.395 167.665 ;
        RECT 23.405 166.985 32.595 167.665 ;
        RECT 27.915 166.765 28.845 166.985 ;
        RECT 31.675 166.755 32.595 166.985 ;
        RECT 32.605 166.885 33.975 167.665 ;
        RECT 33.985 166.755 37.145 167.665 ;
        RECT 37.215 166.795 37.645 167.580 ;
        RECT 37.675 166.755 39.025 167.665 ;
        RECT 39.155 166.985 42.620 167.665 ;
        RECT 41.700 166.755 42.620 166.985 ;
        RECT 42.820 166.985 46.285 167.665 ;
        RECT 47.325 166.985 56.515 167.665 ;
        RECT 42.820 166.755 43.740 166.985 ;
        RECT 47.325 166.755 48.245 166.985 ;
        RECT 51.075 166.765 52.005 166.985 ;
        RECT 56.525 166.855 58.355 167.665 ;
        RECT 58.375 166.755 59.725 167.665 ;
        RECT 60.345 166.755 62.955 167.665 ;
        RECT 62.975 166.795 63.405 167.580 ;
        RECT 63.425 166.855 65.255 167.665 ;
        RECT 65.275 166.985 68.015 167.665 ;
        RECT 68.025 166.985 70.765 167.665 ;
        RECT 70.785 166.755 73.505 167.665 ;
        RECT 73.545 166.855 75.375 167.665 ;
        RECT 75.755 166.985 85.035 167.665 ;
        RECT 75.755 166.865 78.090 166.985 ;
        RECT 75.755 166.755 76.675 166.865 ;
        RECT 82.755 166.765 83.675 166.985 ;
        RECT 85.055 166.755 86.405 167.665 ;
        RECT 86.435 166.755 87.785 167.665 ;
        RECT 88.735 166.795 89.165 167.580 ;
        RECT 89.645 166.855 93.315 167.665 ;
        RECT 93.555 166.985 97.455 167.665 ;
        RECT 96.525 166.755 97.455 166.985 ;
        RECT 97.835 166.985 107.115 167.665 ;
        RECT 107.235 166.985 110.700 167.665 ;
        RECT 110.915 166.985 114.380 167.665 ;
        RECT 97.835 166.865 100.170 166.985 ;
        RECT 97.835 166.755 98.755 166.865 ;
        RECT 104.835 166.765 105.755 166.985 ;
        RECT 109.780 166.755 110.700 166.985 ;
        RECT 113.460 166.755 114.380 166.985 ;
        RECT 114.495 166.795 114.925 167.580 ;
        RECT 115.865 166.985 125.055 167.665 ;
        RECT 115.865 166.755 116.785 166.985 ;
        RECT 119.615 166.765 120.545 166.985 ;
        RECT 125.065 166.855 126.435 167.665 ;
        RECT 126.445 166.855 127.815 167.665 ;
      LAYER nwell ;
        RECT 14.470 163.635 128.010 166.465 ;
      LAYER pwell ;
        RECT 14.665 162.435 16.035 163.245 ;
        RECT 16.045 162.435 18.795 163.245 ;
        RECT 18.805 162.435 24.315 163.245 ;
        RECT 24.335 162.520 24.765 163.305 ;
        RECT 25.705 162.435 27.075 163.215 ;
        RECT 31.595 163.115 32.525 163.335 ;
        RECT 35.355 163.115 36.275 163.345 ;
        RECT 27.085 162.435 36.275 163.115 ;
        RECT 36.285 163.115 37.205 163.345 ;
        RECT 40.035 163.115 40.965 163.335 ;
        RECT 49.060 163.115 49.980 163.345 ;
        RECT 36.285 162.435 45.475 163.115 ;
        RECT 46.515 162.435 49.980 163.115 ;
        RECT 50.095 162.520 50.525 163.305 ;
        RECT 50.555 162.435 51.905 163.345 ;
        RECT 51.925 162.435 53.755 163.245 ;
        RECT 53.765 162.435 55.135 163.215 ;
        RECT 55.145 163.115 56.065 163.345 ;
        RECT 58.895 163.115 59.825 163.335 ;
        RECT 55.145 162.435 64.335 163.115 ;
        RECT 64.485 162.435 67.095 163.345 ;
        RECT 67.115 162.435 69.855 163.115 ;
        RECT 70.325 162.435 75.835 163.245 ;
        RECT 75.855 162.520 76.285 163.305 ;
        RECT 76.305 162.435 78.135 163.245 ;
        RECT 81.345 163.115 82.275 163.345 ;
        RECT 78.375 162.435 82.275 163.115 ;
        RECT 82.285 162.435 83.655 163.215 ;
        RECT 83.665 162.435 85.495 163.245 ;
        RECT 85.505 162.435 86.875 163.215 ;
        RECT 86.885 162.435 92.395 163.245 ;
        RECT 92.490 162.435 101.595 163.115 ;
        RECT 101.615 162.520 102.045 163.305 ;
        RECT 105.265 163.115 106.195 163.345 ;
        RECT 102.295 162.435 106.195 163.115 ;
        RECT 106.665 163.115 107.595 163.345 ;
        RECT 106.665 162.435 110.565 163.115 ;
        RECT 110.945 162.435 113.555 163.345 ;
        RECT 113.565 163.115 114.485 163.345 ;
        RECT 117.315 163.115 118.245 163.335 ;
        RECT 113.565 162.435 122.755 163.115 ;
        RECT 122.765 162.435 124.135 163.215 ;
        RECT 124.605 162.435 126.435 163.245 ;
        RECT 126.445 162.435 127.815 163.245 ;
        RECT 14.805 162.225 14.975 162.435 ;
        RECT 17.565 162.225 17.735 162.415 ;
        RECT 18.485 162.245 18.655 162.435 ;
        RECT 24.005 162.245 24.175 162.435 ;
        RECT 25.385 162.280 25.545 162.390 ;
        RECT 26.765 162.245 26.935 162.435 ;
        RECT 27.225 162.225 27.395 162.435 ;
        RECT 27.960 162.225 28.130 162.415 ;
        RECT 32.745 162.225 32.915 162.415 ;
        RECT 33.480 162.225 33.650 162.415 ;
        RECT 37.860 162.275 37.980 162.385 ;
        RECT 39.645 162.225 39.815 162.415 ;
        RECT 40.105 162.225 40.275 162.415 ;
        RECT 44.060 162.225 44.230 162.415 ;
        RECT 45.165 162.245 45.335 162.435 ;
        RECT 46.085 162.280 46.245 162.390 ;
        RECT 46.545 162.245 46.715 162.435 ;
        RECT 48.845 162.225 49.015 162.415 ;
        RECT 49.580 162.225 49.750 162.415 ;
        RECT 51.605 162.245 51.775 162.435 ;
        RECT 53.445 162.245 53.615 162.435 ;
        RECT 53.905 162.245 54.075 162.435 ;
        RECT 56.850 162.225 57.020 162.415 ;
        RECT 57.640 162.275 57.760 162.385 ;
        RECT 59.425 162.225 59.595 162.415 ;
        RECT 59.885 162.225 60.055 162.415 ;
        RECT 62.645 162.225 62.815 162.415 ;
        RECT 64.025 162.245 64.195 162.435 ;
        RECT 64.485 162.225 64.655 162.415 ;
        RECT 66.325 162.225 66.495 162.415 ;
        RECT 66.780 162.245 66.950 162.435 ;
        RECT 68.165 162.225 68.335 162.415 ;
        RECT 68.625 162.225 68.795 162.415 ;
        RECT 69.545 162.245 69.715 162.435 ;
        RECT 70.060 162.275 70.180 162.385 ;
        RECT 70.465 162.225 70.635 162.415 ;
        RECT 72.360 162.275 72.480 162.385 ;
        RECT 75.065 162.225 75.235 162.415 ;
        RECT 75.525 162.245 75.695 162.435 ;
        RECT 77.825 162.245 77.995 162.435 ;
        RECT 80.585 162.225 80.755 162.415 ;
        RECT 81.690 162.245 81.860 162.435 ;
        RECT 81.965 162.225 82.135 162.415 ;
        RECT 82.425 162.245 82.595 162.435 ;
        RECT 85.185 162.245 85.355 162.435 ;
        RECT 85.645 162.245 85.815 162.435 ;
        RECT 85.830 162.225 86.000 162.415 ;
        RECT 86.565 162.225 86.735 162.415 ;
        RECT 88.405 162.270 88.565 162.380 ;
        RECT 89.380 162.275 89.500 162.385 ;
        RECT 92.085 162.245 92.255 162.435 ;
        RECT 98.985 162.225 99.155 162.415 ;
        RECT 101.285 162.245 101.455 162.435 ;
        RECT 102.205 162.225 102.375 162.415 ;
        RECT 102.665 162.225 102.835 162.415 ;
        RECT 105.610 162.245 105.780 162.435 ;
        RECT 106.400 162.275 106.520 162.385 ;
        RECT 106.805 162.225 106.975 162.415 ;
        RECT 107.080 162.245 107.250 162.435 ;
        RECT 113.240 162.245 113.410 162.435 ;
        RECT 113.890 162.225 114.060 162.415 ;
        RECT 118.490 162.225 118.660 162.415 ;
        RECT 119.225 162.225 119.395 162.415 ;
        RECT 120.660 162.275 120.780 162.385 ;
        RECT 121.065 162.225 121.235 162.415 ;
        RECT 122.445 162.385 122.615 162.435 ;
        RECT 122.445 162.275 122.620 162.385 ;
        RECT 122.445 162.245 122.615 162.275 ;
        RECT 123.825 162.245 123.995 162.435 ;
        RECT 124.340 162.275 124.460 162.385 ;
        RECT 126.125 162.225 126.295 162.435 ;
        RECT 127.505 162.225 127.675 162.435 ;
        RECT 14.665 161.415 16.035 162.225 ;
        RECT 16.045 161.415 17.875 162.225 ;
        RECT 18.255 161.545 27.535 162.225 ;
        RECT 27.545 161.545 31.445 162.225 ;
        RECT 18.255 161.425 20.590 161.545 ;
        RECT 18.255 161.315 19.175 161.425 ;
        RECT 25.255 161.325 26.175 161.545 ;
        RECT 27.545 161.315 28.475 161.545 ;
        RECT 31.685 161.415 33.055 162.225 ;
        RECT 33.065 161.545 36.965 162.225 ;
        RECT 33.065 161.315 33.995 161.545 ;
        RECT 37.215 161.355 37.645 162.140 ;
        RECT 38.125 161.415 39.955 162.225 ;
        RECT 40.075 161.545 43.540 162.225 ;
        RECT 42.620 161.315 43.540 161.545 ;
        RECT 43.645 161.545 47.545 162.225 ;
        RECT 43.645 161.315 44.575 161.545 ;
        RECT 47.785 161.445 49.155 162.225 ;
        RECT 49.165 161.545 53.065 162.225 ;
        RECT 53.535 161.545 57.435 162.225 ;
        RECT 49.165 161.315 50.095 161.545 ;
        RECT 56.505 161.315 57.435 161.545 ;
        RECT 57.905 161.415 59.735 162.225 ;
        RECT 59.745 161.445 61.115 162.225 ;
        RECT 61.125 161.415 62.955 162.225 ;
        RECT 62.975 161.355 63.405 162.140 ;
        RECT 63.425 161.415 64.795 162.225 ;
        RECT 64.805 161.545 66.635 162.225 ;
        RECT 66.645 161.545 68.475 162.225 ;
        RECT 68.485 161.545 70.315 162.225 ;
        RECT 70.325 161.545 72.155 162.225 ;
        RECT 64.805 161.315 66.150 161.545 ;
        RECT 66.645 161.315 67.990 161.545 ;
        RECT 68.970 161.315 70.315 161.545 ;
        RECT 70.810 161.315 72.155 161.545 ;
        RECT 72.625 161.415 75.375 162.225 ;
        RECT 75.385 161.415 80.895 162.225 ;
        RECT 80.915 161.315 82.265 162.225 ;
        RECT 82.515 161.545 86.415 162.225 ;
        RECT 85.485 161.315 86.415 161.545 ;
        RECT 86.425 161.445 87.795 162.225 ;
        RECT 88.735 161.355 89.165 162.140 ;
        RECT 90.015 161.545 99.295 162.225 ;
        RECT 90.015 161.425 92.350 161.545 ;
        RECT 90.015 161.315 90.935 161.425 ;
        RECT 97.015 161.325 97.935 161.545 ;
        RECT 99.305 161.315 102.465 162.225 ;
        RECT 102.635 161.545 106.100 162.225 ;
        RECT 106.775 161.545 110.240 162.225 ;
        RECT 110.575 161.545 114.475 162.225 ;
        RECT 105.180 161.315 106.100 161.545 ;
        RECT 109.320 161.315 110.240 161.545 ;
        RECT 113.545 161.315 114.475 161.545 ;
        RECT 114.495 161.355 114.925 162.140 ;
        RECT 115.175 161.545 119.075 162.225 ;
        RECT 118.145 161.315 119.075 161.545 ;
        RECT 119.095 161.315 120.445 162.225 ;
        RECT 120.925 161.445 122.295 162.225 ;
        RECT 122.765 161.415 126.435 162.225 ;
        RECT 126.445 161.415 127.815 162.225 ;
      LAYER nwell ;
        RECT 14.470 158.195 128.010 161.025 ;
      LAYER pwell ;
        RECT 14.665 156.995 16.035 157.805 ;
        RECT 16.045 156.995 17.415 157.805 ;
        RECT 17.435 156.995 18.785 157.905 ;
        RECT 18.815 156.995 20.165 157.905 ;
        RECT 23.385 157.675 24.315 157.905 ;
        RECT 20.415 156.995 24.315 157.675 ;
        RECT 24.335 157.080 24.765 157.865 ;
        RECT 24.785 156.995 26.155 157.775 ;
        RECT 26.165 156.995 27.995 157.805 ;
        RECT 30.660 157.675 31.580 157.905 ;
        RECT 34.340 157.675 35.260 157.905 ;
        RECT 28.115 156.995 31.580 157.675 ;
        RECT 31.795 156.995 35.260 157.675 ;
        RECT 35.365 156.995 39.035 157.805 ;
        RECT 39.240 156.995 42.715 157.905 ;
        RECT 42.920 156.995 46.395 157.905 ;
        RECT 49.060 157.675 49.980 157.905 ;
        RECT 46.515 156.995 49.980 157.675 ;
        RECT 50.095 157.080 50.525 157.865 ;
        RECT 50.545 156.995 54.020 157.905 ;
        RECT 54.685 156.995 60.195 157.805 ;
        RECT 60.215 156.995 61.565 157.905 ;
        RECT 61.725 156.995 64.335 157.905 ;
        RECT 64.805 156.995 68.475 157.805 ;
        RECT 68.970 157.675 70.315 157.905 ;
        RECT 70.810 157.675 72.155 157.905 ;
        RECT 68.485 156.995 70.315 157.675 ;
        RECT 70.325 156.995 72.155 157.675 ;
        RECT 72.360 156.995 75.835 157.905 ;
        RECT 75.855 157.080 76.285 157.865 ;
        RECT 76.960 156.995 80.435 157.905 ;
        RECT 81.275 157.795 82.195 157.905 ;
        RECT 81.275 157.675 83.610 157.795 ;
        RECT 88.275 157.675 89.195 157.895 ;
        RECT 81.275 156.995 90.555 157.675 ;
        RECT 91.025 156.995 92.855 157.805 ;
        RECT 92.875 156.995 94.225 157.905 ;
        RECT 94.705 156.995 96.535 157.805 ;
        RECT 96.545 156.995 97.915 157.775 ;
        RECT 97.925 156.995 99.755 157.805 ;
        RECT 99.775 156.995 101.125 157.905 ;
        RECT 101.615 157.080 102.045 157.865 ;
        RECT 102.525 156.995 104.355 157.805 ;
        RECT 104.365 156.995 105.735 157.775 ;
        RECT 105.745 156.995 107.115 157.775 ;
        RECT 108.045 156.995 111.520 157.905 ;
        RECT 112.645 156.995 116.315 157.805 ;
        RECT 118.980 157.675 119.900 157.905 ;
        RECT 116.435 156.995 119.900 157.675 ;
        RECT 120.925 156.995 126.435 157.805 ;
        RECT 126.445 156.995 127.815 157.805 ;
        RECT 14.805 156.785 14.975 156.995 ;
        RECT 16.645 156.830 16.805 156.940 ;
        RECT 17.105 156.805 17.275 156.995 ;
        RECT 18.485 156.805 18.655 156.995 ;
        RECT 18.945 156.805 19.115 156.995 ;
        RECT 23.730 156.805 23.900 156.995 ;
        RECT 24.925 156.805 25.095 156.995 ;
        RECT 26.305 156.785 26.475 156.975 ;
        RECT 27.685 156.785 27.855 156.995 ;
        RECT 28.145 156.805 28.315 156.995 ;
        RECT 29.065 156.785 29.235 156.975 ;
        RECT 31.825 156.805 31.995 156.995 ;
        RECT 32.745 156.785 32.915 156.975 ;
        RECT 36.610 156.785 36.780 156.975 ;
        RECT 37.860 156.835 37.980 156.945 ;
        RECT 38.725 156.805 38.895 156.995 ;
        RECT 39.645 156.785 39.815 156.975 ;
        RECT 40.110 156.785 40.280 156.975 ;
        RECT 42.400 156.805 42.570 156.995 ;
        RECT 43.790 156.785 43.960 156.975 ;
        RECT 46.080 156.805 46.250 156.995 ;
        RECT 46.545 156.805 46.715 156.995 ;
        RECT 47.470 156.785 47.640 156.975 ;
        RECT 50.690 156.805 50.860 156.995 ;
        RECT 51.200 156.835 51.320 156.945 ;
        RECT 52.985 156.785 53.155 156.975 ;
        RECT 54.420 156.835 54.540 156.945 ;
        RECT 59.885 156.805 60.055 156.995 ;
        RECT 61.265 156.805 61.435 156.995 ;
        RECT 62.645 156.785 62.815 156.975 ;
        RECT 63.620 156.835 63.740 156.945 ;
        RECT 64.020 156.805 64.190 156.995 ;
        RECT 64.540 156.835 64.660 156.945 ;
        RECT 65.405 156.785 65.575 156.975 ;
        RECT 68.165 156.805 68.335 156.995 ;
        RECT 68.625 156.805 68.795 156.995 ;
        RECT 70.465 156.805 70.635 156.995 ;
        RECT 74.605 156.785 74.775 156.975 ;
        RECT 75.520 156.805 75.690 156.995 ;
        RECT 76.445 156.945 76.615 156.975 ;
        RECT 76.445 156.835 76.620 156.945 ;
        RECT 76.445 156.785 76.615 156.835 ;
        RECT 76.910 156.785 77.080 156.975 ;
        RECT 80.120 156.805 80.290 156.995 ;
        RECT 80.590 156.785 80.760 156.975 ;
        RECT 84.725 156.830 84.885 156.940 ;
        RECT 88.405 156.785 88.575 156.975 ;
        RECT 90.245 156.805 90.415 156.995 ;
        RECT 90.760 156.835 90.880 156.945 ;
        RECT 91.625 156.785 91.795 156.975 ;
        RECT 92.545 156.805 92.715 156.995 ;
        RECT 93.005 156.805 93.175 156.995 ;
        RECT 94.440 156.835 94.560 156.945 ;
        RECT 96.225 156.805 96.395 156.995 ;
        RECT 96.685 156.805 96.855 156.995 ;
        RECT 97.145 156.785 97.315 156.975 ;
        RECT 99.445 156.805 99.615 156.995 ;
        RECT 99.905 156.805 100.075 156.995 ;
        RECT 100.820 156.785 100.990 156.975 ;
        RECT 101.340 156.835 101.460 156.945 ;
        RECT 102.260 156.835 102.380 156.945 ;
        RECT 103.125 156.785 103.295 156.975 ;
        RECT 103.590 156.785 103.760 156.975 ;
        RECT 104.045 156.805 104.215 156.995 ;
        RECT 105.425 156.805 105.595 156.995 ;
        RECT 105.885 156.805 106.055 156.995 ;
        RECT 107.725 156.840 107.885 156.950 ;
        RECT 108.190 156.805 108.360 156.995 ;
        RECT 110.480 156.785 110.650 156.975 ;
        RECT 112.325 156.840 112.485 156.950 ;
        RECT 114.165 156.785 114.335 156.975 ;
        RECT 116.005 156.785 116.175 156.995 ;
        RECT 116.465 156.975 116.635 156.995 ;
        RECT 116.465 156.805 116.640 156.975 ;
        RECT 116.470 156.785 116.640 156.805 ;
        RECT 120.605 156.785 120.775 156.975 ;
        RECT 126.125 156.785 126.295 156.995 ;
        RECT 127.505 156.785 127.675 156.995 ;
        RECT 14.665 155.975 16.035 156.785 ;
        RECT 17.335 156.105 26.615 156.785 ;
        RECT 17.335 155.985 19.670 156.105 ;
        RECT 17.335 155.875 18.255 155.985 ;
        RECT 24.335 155.885 25.255 156.105 ;
        RECT 26.625 156.005 27.995 156.785 ;
        RECT 28.005 155.975 29.375 156.785 ;
        RECT 29.385 155.975 33.055 156.785 ;
        RECT 33.295 156.105 37.195 156.785 ;
        RECT 36.265 155.875 37.195 156.105 ;
        RECT 37.215 155.915 37.645 156.700 ;
        RECT 38.125 155.975 39.955 156.785 ;
        RECT 39.965 155.875 43.440 156.785 ;
        RECT 43.645 155.875 47.120 156.785 ;
        RECT 47.325 155.875 50.800 156.785 ;
        RECT 51.465 155.975 53.295 156.785 ;
        RECT 53.675 156.105 62.955 156.785 ;
        RECT 53.675 155.985 56.010 156.105 ;
        RECT 53.675 155.875 54.595 155.985 ;
        RECT 60.675 155.885 61.595 156.105 ;
        RECT 62.975 155.915 63.405 156.700 ;
        RECT 63.885 155.975 65.715 156.785 ;
        RECT 65.810 156.105 74.915 156.785 ;
        RECT 74.925 155.975 76.755 156.785 ;
        RECT 76.765 155.875 80.240 156.785 ;
        RECT 80.445 155.875 83.920 156.785 ;
        RECT 85.045 155.975 88.715 156.785 ;
        RECT 88.735 155.915 89.165 156.700 ;
        RECT 89.185 155.975 91.935 156.785 ;
        RECT 91.945 155.975 97.455 156.785 ;
        RECT 97.660 155.875 101.135 156.785 ;
        RECT 101.605 155.975 103.435 156.785 ;
        RECT 103.445 155.875 106.920 156.785 ;
        RECT 107.320 155.875 110.795 156.785 ;
        RECT 110.805 155.975 114.475 156.785 ;
        RECT 114.495 155.915 114.925 156.700 ;
        RECT 114.945 155.975 116.315 156.785 ;
        RECT 116.325 155.875 118.935 156.785 ;
        RECT 119.085 155.975 120.915 156.785 ;
        RECT 120.925 155.975 126.435 156.785 ;
        RECT 126.445 155.975 127.815 156.785 ;
      LAYER nwell ;
        RECT 14.470 152.755 128.010 155.585 ;
      LAYER pwell ;
        RECT 14.665 151.555 16.035 152.365 ;
        RECT 16.505 151.555 20.175 152.365 ;
        RECT 23.385 152.235 24.315 152.465 ;
        RECT 20.415 151.555 24.315 152.235 ;
        RECT 24.335 151.640 24.765 152.425 ;
        RECT 24.785 151.555 26.155 152.365 ;
        RECT 26.165 151.555 29.835 152.365 ;
        RECT 30.215 152.355 31.135 152.465 ;
        RECT 30.215 152.235 32.550 152.355 ;
        RECT 37.215 152.235 38.135 152.455 ;
        RECT 30.215 151.555 39.495 152.235 ;
        RECT 39.505 151.555 42.980 152.465 ;
        RECT 43.185 151.555 44.555 152.365 ;
        RECT 44.565 151.555 50.075 152.365 ;
        RECT 50.095 151.640 50.525 152.425 ;
        RECT 51.465 151.555 56.975 152.365 ;
        RECT 56.995 151.555 58.345 152.465 ;
        RECT 58.735 152.355 59.655 152.465 ;
        RECT 58.735 152.235 61.070 152.355 ;
        RECT 65.735 152.235 66.655 152.455 ;
        RECT 58.735 151.555 68.015 152.235 ;
        RECT 68.485 151.555 71.235 152.365 ;
        RECT 71.730 152.235 73.075 152.465 ;
        RECT 71.245 151.555 73.075 152.235 ;
        RECT 73.085 151.555 75.805 152.465 ;
        RECT 75.855 151.640 76.285 152.425 ;
        RECT 77.225 151.555 80.895 152.365 ;
        RECT 80.905 151.555 86.415 152.365 ;
        RECT 86.795 152.355 87.715 152.465 ;
        RECT 86.795 152.235 89.130 152.355 ;
        RECT 93.795 152.235 94.715 152.455 ;
        RECT 86.795 151.555 96.075 152.235 ;
        RECT 96.085 151.555 101.595 152.365 ;
        RECT 101.615 151.640 102.045 152.425 ;
        RECT 102.525 152.265 103.470 152.465 ;
        RECT 102.525 151.585 105.275 152.265 ;
        RECT 102.525 151.555 103.470 151.585 ;
        RECT 14.805 151.345 14.975 151.555 ;
        RECT 16.240 151.395 16.360 151.505 ;
        RECT 19.865 151.365 20.035 151.555 ;
        RECT 23.730 151.365 23.900 151.555 ;
        RECT 25.845 151.345 26.015 151.555 ;
        RECT 27.225 151.345 27.395 151.535 ;
        RECT 29.525 151.365 29.695 151.555 ;
        RECT 32.745 151.345 32.915 151.535 ;
        RECT 33.205 151.345 33.375 151.535 ;
        RECT 35.505 151.345 35.675 151.535 ;
        RECT 35.965 151.345 36.135 151.535 ;
        RECT 39.185 151.365 39.355 151.555 ;
        RECT 39.650 151.365 39.820 151.555 ;
        RECT 41.025 151.345 41.195 151.535 ;
        RECT 41.490 151.345 41.660 151.535 ;
        RECT 44.245 151.365 44.415 151.555 ;
        RECT 48.385 151.345 48.555 151.535 ;
        RECT 14.665 150.535 16.035 151.345 ;
        RECT 16.875 150.665 26.155 151.345 ;
        RECT 16.875 150.545 19.210 150.665 ;
        RECT 16.875 150.435 17.795 150.545 ;
        RECT 23.875 150.445 24.795 150.665 ;
        RECT 26.165 150.535 27.535 151.345 ;
        RECT 27.545 150.535 33.055 151.345 ;
        RECT 33.075 150.435 34.425 151.345 ;
        RECT 34.445 150.535 35.815 151.345 ;
        RECT 35.825 150.565 37.195 151.345 ;
        RECT 37.215 150.475 37.645 151.260 ;
        RECT 37.665 150.535 41.335 151.345 ;
        RECT 41.345 150.435 44.820 151.345 ;
        RECT 45.025 150.535 48.695 151.345 ;
        RECT 48.850 151.315 49.020 151.535 ;
        RECT 49.765 151.365 49.935 151.555 ;
        RECT 51.145 151.400 51.305 151.510 ;
        RECT 51.610 151.345 51.780 151.535 ;
        RECT 56.665 151.345 56.835 151.555 ;
        RECT 57.125 151.365 57.295 151.555 ;
        RECT 60.530 151.345 60.700 151.535 ;
        RECT 61.320 151.395 61.440 151.505 ;
        RECT 62.645 151.345 62.815 151.535 ;
        RECT 63.620 151.395 63.740 151.505 ;
        RECT 64.025 151.345 64.195 151.535 ;
        RECT 65.460 151.395 65.580 151.505 ;
        RECT 67.245 151.345 67.415 151.535 ;
        RECT 67.705 151.345 67.875 151.555 ;
        RECT 68.220 151.395 68.340 151.505 ;
        RECT 70.925 151.345 71.095 151.555 ;
        RECT 71.385 151.365 71.555 151.555 ;
        RECT 73.225 151.365 73.395 151.555 ;
        RECT 73.685 151.345 73.855 151.535 ;
        RECT 74.605 151.390 74.765 151.500 ;
        RECT 75.065 151.345 75.235 151.535 ;
        RECT 76.905 151.400 77.065 151.510 ;
        RECT 50.510 151.315 51.455 151.345 ;
        RECT 48.705 150.635 51.455 151.315 ;
        RECT 50.510 150.435 51.455 150.635 ;
        RECT 51.465 150.435 54.940 151.345 ;
        RECT 55.145 150.535 56.975 151.345 ;
        RECT 57.215 150.665 61.115 151.345 ;
        RECT 60.185 150.435 61.115 150.665 ;
        RECT 61.585 150.565 62.955 151.345 ;
        RECT 62.975 150.475 63.405 151.260 ;
        RECT 63.885 150.565 65.255 151.345 ;
        RECT 65.725 150.535 67.555 151.345 ;
        RECT 67.565 150.665 69.395 151.345 ;
        RECT 68.050 150.435 69.395 150.665 ;
        RECT 69.405 150.665 71.235 151.345 ;
        RECT 71.255 150.665 73.995 151.345 ;
        RECT 74.925 150.665 77.665 151.345 ;
        RECT 77.685 151.315 78.630 151.345 ;
        RECT 80.120 151.315 80.290 151.535 ;
        RECT 80.585 151.505 80.755 151.555 ;
        RECT 80.585 151.395 80.760 151.505 ;
        RECT 80.585 151.365 80.755 151.395 ;
        RECT 84.265 151.345 84.435 151.535 ;
        RECT 86.105 151.365 86.275 151.555 ;
        RECT 88.130 151.345 88.300 151.535 ;
        RECT 89.380 151.395 89.500 151.505 ;
        RECT 90.705 151.345 90.875 151.535 ;
        RECT 91.625 151.390 91.785 151.500 ;
        RECT 92.085 151.345 92.255 151.535 ;
        RECT 94.385 151.345 94.555 151.535 ;
        RECT 95.765 151.365 95.935 151.555 ;
        RECT 96.225 151.345 96.395 151.535 ;
        RECT 101.285 151.365 101.455 151.555 ;
        RECT 102.260 151.395 102.380 151.505 ;
        RECT 104.960 151.365 105.130 151.585 ;
        RECT 105.285 151.555 108.760 152.465 ;
        RECT 108.965 151.555 112.440 152.465 ;
        RECT 113.105 151.555 118.615 152.365 ;
        RECT 118.635 151.555 119.985 152.465 ;
        RECT 120.465 151.555 121.835 152.335 ;
        RECT 122.765 151.555 126.435 152.365 ;
        RECT 126.445 151.555 127.815 152.365 ;
        RECT 105.430 151.535 105.600 151.555 ;
        RECT 105.425 151.365 105.600 151.535 ;
        RECT 105.425 151.345 105.595 151.365 ;
        RECT 106.805 151.345 106.975 151.535 ;
        RECT 107.270 151.345 107.440 151.535 ;
        RECT 109.110 151.365 109.280 151.555 ;
        RECT 110.945 151.345 111.115 151.535 ;
        RECT 112.840 151.395 112.960 151.505 ;
        RECT 115.545 151.390 115.705 151.500 ;
        RECT 118.305 151.365 118.475 151.555 ;
        RECT 119.685 151.365 119.855 151.555 ;
        RECT 120.200 151.395 120.320 151.505 ;
        RECT 120.605 151.365 120.775 151.555 ;
        RECT 122.445 151.400 122.605 151.510 ;
        RECT 124.745 151.345 124.915 151.535 ;
        RECT 126.125 151.345 126.295 151.555 ;
        RECT 127.505 151.345 127.675 151.555 ;
        RECT 69.405 150.435 70.750 150.665 ;
        RECT 77.685 150.635 80.435 151.315 ;
        RECT 77.685 150.435 78.630 150.635 ;
        RECT 80.905 150.535 84.575 151.345 ;
        RECT 84.815 150.665 88.715 151.345 ;
        RECT 87.785 150.435 88.715 150.665 ;
        RECT 88.735 150.475 89.165 151.260 ;
        RECT 89.655 150.435 91.005 151.345 ;
        RECT 91.945 150.565 93.315 151.345 ;
        RECT 93.335 150.435 94.685 151.345 ;
        RECT 94.705 150.535 96.535 151.345 ;
        RECT 96.545 150.665 105.735 151.345 ;
        RECT 96.545 150.435 97.465 150.665 ;
        RECT 100.295 150.445 101.225 150.665 ;
        RECT 105.745 150.535 107.115 151.345 ;
        RECT 107.125 150.435 110.600 151.345 ;
        RECT 110.915 150.665 114.380 151.345 ;
        RECT 113.460 150.435 114.380 150.665 ;
        RECT 114.495 150.475 114.925 151.260 ;
        RECT 115.865 150.665 125.055 151.345 ;
        RECT 115.865 150.435 116.785 150.665 ;
        RECT 119.615 150.445 120.545 150.665 ;
        RECT 125.065 150.535 126.435 151.345 ;
        RECT 126.445 150.535 127.815 151.345 ;
      LAYER nwell ;
        RECT 14.470 147.315 128.010 150.145 ;
      LAYER pwell ;
        RECT 14.665 146.115 16.035 146.925 ;
        RECT 16.505 146.115 20.175 146.925 ;
        RECT 23.385 146.795 24.315 147.025 ;
        RECT 20.415 146.115 24.315 146.795 ;
        RECT 24.335 146.200 24.765 146.985 ;
        RECT 24.785 146.115 26.155 146.895 ;
        RECT 26.165 146.115 27.995 146.925 ;
        RECT 28.005 146.115 29.375 146.895 ;
        RECT 29.385 146.795 30.315 147.025 ;
        RECT 29.385 146.115 33.285 146.795 ;
        RECT 33.985 146.115 35.815 146.925 ;
        RECT 36.020 146.115 39.495 147.025 ;
        RECT 39.505 146.115 42.980 147.025 ;
        RECT 43.645 146.115 47.315 146.925 ;
        RECT 49.130 146.825 50.075 147.025 ;
        RECT 47.325 146.145 50.075 146.825 ;
        RECT 50.095 146.200 50.525 146.985 ;
        RECT 14.805 145.905 14.975 146.115 ;
        RECT 16.240 145.955 16.360 146.065 ;
        RECT 19.405 145.905 19.575 146.095 ;
        RECT 19.865 145.905 20.035 146.115 ;
        RECT 21.245 145.905 21.415 146.095 ;
        RECT 23.730 145.925 23.900 146.115 ;
        RECT 25.845 145.925 26.015 146.115 ;
        RECT 27.685 145.925 27.855 146.115 ;
        RECT 28.145 145.925 28.315 146.115 ;
        RECT 29.800 145.925 29.970 146.115 ;
        RECT 31.825 145.905 31.995 146.095 ;
        RECT 33.205 145.905 33.375 146.095 ;
        RECT 33.720 145.955 33.840 146.065 ;
        RECT 35.505 145.925 35.675 146.115 ;
        RECT 36.885 145.905 37.055 146.095 ;
        RECT 37.860 145.955 37.980 146.065 ;
        RECT 39.180 145.925 39.350 146.115 ;
        RECT 39.650 145.925 39.820 146.115 ;
        RECT 40.565 145.905 40.735 146.095 ;
        RECT 41.025 145.905 41.195 146.095 ;
        RECT 43.380 145.955 43.500 146.065 ;
        RECT 47.005 145.925 47.175 146.115 ;
        RECT 47.470 145.925 47.640 146.145 ;
        RECT 49.130 146.115 50.075 146.145 ;
        RECT 51.005 146.115 52.375 146.895 ;
        RECT 53.305 146.115 56.780 147.025 ;
        RECT 56.985 146.115 59.735 146.925 ;
        RECT 62.945 146.795 63.875 147.025 ;
        RECT 59.975 146.115 63.875 146.795 ;
        RECT 63.885 146.115 65.255 146.925 ;
        RECT 65.265 146.115 70.775 146.925 ;
        RECT 70.785 146.795 72.130 147.025 ;
        RECT 73.110 146.795 74.455 147.025 ;
        RECT 70.785 146.115 72.615 146.795 ;
        RECT 72.625 146.115 74.455 146.795 ;
        RECT 74.465 146.115 75.835 146.925 ;
        RECT 75.855 146.200 76.285 146.985 ;
        RECT 76.500 146.115 79.975 147.025 ;
        RECT 79.985 146.115 83.460 147.025 ;
        RECT 83.665 146.115 85.035 146.925 ;
        RECT 85.415 146.915 86.335 147.025 ;
        RECT 85.415 146.795 87.750 146.915 ;
        RECT 92.415 146.795 93.335 147.015 ;
        RECT 85.415 146.115 94.695 146.795 ;
        RECT 95.175 146.115 96.525 147.025 ;
        RECT 99.745 146.795 100.675 147.025 ;
        RECT 96.775 146.115 100.675 146.795 ;
        RECT 101.615 146.200 102.045 146.985 ;
        RECT 102.065 146.115 103.435 146.895 ;
        RECT 103.905 146.825 104.850 147.025 ;
        RECT 103.905 146.145 106.655 146.825 ;
        RECT 103.905 146.115 104.850 146.145 ;
        RECT 50.740 145.955 50.860 146.065 ;
        RECT 51.605 145.905 51.775 146.095 ;
        RECT 52.065 145.925 52.235 146.115 ;
        RECT 52.340 145.905 52.510 146.095 ;
        RECT 52.985 145.960 53.145 146.070 ;
        RECT 53.450 145.925 53.620 146.115 ;
        RECT 56.260 145.955 56.380 146.065 ;
        RECT 58.045 145.905 58.215 146.095 ;
        RECT 58.505 145.905 58.675 146.095 ;
        RECT 59.425 145.925 59.595 146.115 ;
        RECT 59.940 145.955 60.060 146.065 ;
        RECT 62.645 145.905 62.815 146.095 ;
        RECT 63.290 145.925 63.460 146.115 ;
        RECT 63.620 145.955 63.740 146.065 ;
        RECT 64.945 145.925 65.115 146.115 ;
        RECT 67.430 145.905 67.600 146.095 ;
        RECT 68.220 145.955 68.340 146.065 ;
        RECT 70.465 145.925 70.635 146.115 ;
        RECT 72.305 145.925 72.475 146.115 ;
        RECT 72.765 145.925 72.935 146.115 ;
        RECT 73.685 145.905 73.855 146.095 ;
        RECT 75.525 145.925 75.695 146.115 ;
        RECT 79.660 146.095 79.830 146.115 ;
        RECT 79.205 145.905 79.375 146.095 ;
        RECT 79.660 145.925 79.840 146.095 ;
        RECT 80.130 145.925 80.300 146.115 ;
        RECT 82.480 145.955 82.600 146.065 ;
        RECT 14.665 145.095 16.035 145.905 ;
        RECT 16.045 145.095 19.715 145.905 ;
        RECT 19.735 144.995 21.085 145.905 ;
        RECT 21.115 144.995 22.465 145.905 ;
        RECT 22.855 145.225 32.135 145.905 ;
        RECT 22.855 145.105 25.190 145.225 ;
        RECT 22.855 144.995 23.775 145.105 ;
        RECT 29.855 145.005 30.775 145.225 ;
        RECT 32.145 145.095 33.515 145.905 ;
        RECT 33.525 145.095 37.195 145.905 ;
        RECT 37.215 145.035 37.645 145.820 ;
        RECT 38.125 145.095 40.875 145.905 ;
        RECT 40.895 144.995 42.245 145.905 ;
        RECT 42.635 145.225 51.915 145.905 ;
        RECT 51.925 145.225 55.825 145.905 ;
        RECT 42.635 145.105 44.970 145.225 ;
        RECT 42.635 144.995 43.555 145.105 ;
        RECT 49.635 145.005 50.555 145.225 ;
        RECT 51.925 144.995 52.855 145.225 ;
        RECT 56.525 145.095 58.355 145.905 ;
        RECT 58.375 144.995 59.725 145.905 ;
        RECT 60.205 145.095 62.955 145.905 ;
        RECT 62.975 145.035 63.405 145.820 ;
        RECT 64.115 145.225 68.015 145.905 ;
        RECT 67.085 144.995 68.015 145.225 ;
        RECT 68.485 145.095 73.995 145.905 ;
        RECT 74.005 145.095 79.515 145.905 ;
        RECT 79.670 145.875 79.840 145.925 ;
        RECT 84.265 145.905 84.435 146.095 ;
        RECT 84.725 145.925 84.895 146.115 ;
        RECT 88.130 145.905 88.300 146.095 ;
        RECT 89.785 145.950 89.945 146.060 ;
        RECT 90.245 145.905 90.415 146.095 ;
        RECT 91.680 145.955 91.800 146.065 ;
        RECT 93.465 145.905 93.635 146.095 ;
        RECT 93.925 145.905 94.095 146.095 ;
        RECT 94.385 145.925 94.555 146.115 ;
        RECT 94.900 145.955 95.020 146.065 ;
        RECT 95.305 145.925 95.475 146.115 ;
        RECT 97.660 145.955 97.780 146.065 ;
        RECT 100.090 145.925 100.260 146.115 ;
        RECT 101.285 145.905 101.455 146.095 ;
        RECT 102.205 145.925 102.375 146.115 ;
        RECT 103.640 145.955 103.760 146.065 ;
        RECT 106.340 145.925 106.510 146.145 ;
        RECT 106.665 146.115 110.140 147.025 ;
        RECT 110.345 146.115 112.175 146.925 ;
        RECT 115.385 146.795 116.315 147.025 ;
        RECT 112.415 146.115 116.315 146.795 ;
        RECT 116.695 146.915 117.615 147.025 ;
        RECT 116.695 146.795 119.030 146.915 ;
        RECT 123.695 146.795 124.615 147.015 ;
        RECT 116.695 146.115 125.975 146.795 ;
        RECT 126.445 146.115 127.815 146.925 ;
        RECT 106.810 146.095 106.980 146.115 ;
        RECT 106.805 145.925 106.980 146.095 ;
        RECT 106.805 145.905 106.975 145.925 ;
        RECT 81.330 145.875 82.275 145.905 ;
        RECT 79.525 145.195 82.275 145.875 ;
        RECT 81.330 144.995 82.275 145.195 ;
        RECT 82.745 145.095 84.575 145.905 ;
        RECT 84.815 145.225 88.715 145.905 ;
        RECT 87.785 144.995 88.715 145.225 ;
        RECT 88.735 145.035 89.165 145.820 ;
        RECT 90.105 145.125 91.475 145.905 ;
        RECT 91.945 145.095 93.775 145.905 ;
        RECT 93.895 145.225 97.360 145.905 ;
        RECT 96.440 144.995 97.360 145.225 ;
        RECT 97.925 145.095 101.595 145.905 ;
        RECT 101.605 145.095 107.115 145.905 ;
        RECT 107.270 145.875 107.440 146.095 ;
        RECT 110.030 145.905 110.200 146.095 ;
        RECT 111.865 145.925 112.035 146.115 ;
        RECT 114.165 145.950 114.325 146.060 ;
        RECT 115.140 145.955 115.260 146.065 ;
        RECT 115.730 145.925 115.900 146.115 ;
        RECT 118.950 145.905 119.120 146.095 ;
        RECT 119.685 145.905 119.855 146.095 ;
        RECT 121.120 145.955 121.240 146.065 ;
        RECT 121.525 145.905 121.695 146.095 ;
        RECT 125.665 145.925 125.835 146.115 ;
        RECT 126.125 146.065 126.295 146.095 ;
        RECT 126.125 145.955 126.300 146.065 ;
        RECT 126.125 145.905 126.295 145.955 ;
        RECT 127.505 145.905 127.675 146.115 ;
        RECT 108.930 145.875 109.875 145.905 ;
        RECT 107.125 145.195 109.875 145.875 ;
        RECT 108.930 144.995 109.875 145.195 ;
        RECT 109.885 144.995 113.360 145.905 ;
        RECT 114.495 145.035 114.925 145.820 ;
        RECT 115.635 145.225 119.535 145.905 ;
        RECT 118.605 144.995 119.535 145.225 ;
        RECT 119.555 144.995 120.905 145.905 ;
        RECT 121.385 145.125 122.755 145.905 ;
        RECT 122.765 145.095 126.435 145.905 ;
        RECT 126.445 145.095 127.815 145.905 ;
      LAYER nwell ;
        RECT 14.470 141.875 128.010 144.705 ;
      LAYER pwell ;
        RECT 14.665 140.675 16.035 141.485 ;
        RECT 16.045 140.675 18.795 141.485 ;
        RECT 18.805 140.675 24.315 141.485 ;
        RECT 24.335 140.760 24.765 141.545 ;
        RECT 25.245 140.675 28.915 141.485 ;
        RECT 28.925 140.675 34.435 141.485 ;
        RECT 34.445 141.385 35.390 141.585 ;
        RECT 34.445 140.705 37.195 141.385 ;
        RECT 34.445 140.675 35.390 140.705 ;
        RECT 14.805 140.465 14.975 140.675 ;
        RECT 18.485 140.485 18.655 140.675 ;
        RECT 24.005 140.485 24.175 140.675 ;
        RECT 24.980 140.515 25.100 140.625 ;
        RECT 25.385 140.465 25.555 140.655 ;
        RECT 28.145 140.465 28.315 140.655 ;
        RECT 28.605 140.485 28.775 140.675 ;
        RECT 33.665 140.465 33.835 140.655 ;
        RECT 34.125 140.485 34.295 140.675 ;
        RECT 36.880 140.485 37.050 140.705 ;
        RECT 38.125 140.675 41.795 141.485 ;
        RECT 41.805 140.675 47.315 141.485 ;
        RECT 47.325 141.385 48.270 141.585 ;
        RECT 47.325 140.705 50.075 141.385 ;
        RECT 50.095 140.760 50.525 141.545 ;
        RECT 47.325 140.675 48.270 140.705 ;
        RECT 37.805 140.520 37.965 140.630 ;
        RECT 38.265 140.510 38.425 140.620 ;
        RECT 34.145 140.465 34.295 140.485 ;
        RECT 14.665 139.655 16.035 140.465 ;
        RECT 16.415 139.785 25.695 140.465 ;
        RECT 16.415 139.665 18.750 139.785 ;
        RECT 16.415 139.555 17.335 139.665 ;
        RECT 23.415 139.565 24.335 139.785 ;
        RECT 25.705 139.655 28.455 140.465 ;
        RECT 28.465 139.655 33.975 140.465 ;
        RECT 34.145 139.645 36.075 140.465 ;
        RECT 38.585 140.435 39.530 140.465 ;
        RECT 41.020 140.435 41.190 140.655 ;
        RECT 41.485 140.625 41.655 140.675 ;
        RECT 41.485 140.515 41.660 140.625 ;
        RECT 41.485 140.485 41.655 140.515 ;
        RECT 44.245 140.465 44.415 140.655 ;
        RECT 47.005 140.485 47.175 140.675 ;
        RECT 49.760 140.655 49.930 140.705 ;
        RECT 50.545 140.675 52.375 141.485 ;
        RECT 52.385 140.675 55.860 141.585 ;
        RECT 58.720 141.355 59.640 141.585 ;
        RECT 56.175 140.675 59.640 141.355 ;
        RECT 59.745 141.355 60.665 141.585 ;
        RECT 63.495 141.355 64.425 141.575 ;
        RECT 59.745 140.675 68.935 141.355 ;
        RECT 68.945 140.675 70.315 141.455 ;
        RECT 70.325 140.675 71.695 141.485 ;
        RECT 71.715 140.675 73.065 141.585 ;
        RECT 73.085 140.675 75.835 141.485 ;
        RECT 75.855 140.760 76.285 141.545 ;
        RECT 76.765 140.675 79.515 141.485 ;
        RECT 79.525 140.675 85.035 141.485 ;
        RECT 85.045 140.675 90.555 141.485 ;
        RECT 90.565 140.675 96.075 141.485 ;
        RECT 96.085 140.675 101.595 141.485 ;
        RECT 101.615 140.760 102.045 141.545 ;
        RECT 102.065 140.675 104.815 141.485 ;
        RECT 104.825 140.675 110.335 141.485 ;
        RECT 110.345 140.675 115.855 141.485 ;
        RECT 119.065 141.355 119.995 141.585 ;
        RECT 116.095 140.675 119.995 141.355 ;
        RECT 120.015 140.675 121.365 141.585 ;
        RECT 121.385 140.675 122.755 141.485 ;
        RECT 122.765 140.675 126.435 141.485 ;
        RECT 126.445 140.675 127.815 141.485 ;
        RECT 49.760 140.485 49.935 140.655 ;
        RECT 52.065 140.485 52.235 140.675 ;
        RECT 52.530 140.485 52.700 140.675 ;
        RECT 49.765 140.465 49.935 140.485 ;
        RECT 55.285 140.465 55.455 140.655 ;
        RECT 55.745 140.465 55.915 140.655 ;
        RECT 56.205 140.485 56.375 140.675 ;
        RECT 57.180 140.515 57.300 140.625 ;
        RECT 58.965 140.465 59.135 140.655 ;
        RECT 59.430 140.465 59.600 140.655 ;
        RECT 63.620 140.515 63.740 140.625 ;
        RECT 64.030 140.465 64.200 140.655 ;
        RECT 68.625 140.485 68.795 140.675 ;
        RECT 70.005 140.485 70.175 140.675 ;
        RECT 71.385 140.485 71.555 140.675 ;
        RECT 72.765 140.485 72.935 140.675 ;
        RECT 75.525 140.485 75.695 140.675 ;
        RECT 76.500 140.515 76.620 140.625 ;
        RECT 76.905 140.465 77.075 140.655 ;
        RECT 77.420 140.515 77.540 140.625 ;
        RECT 79.205 140.465 79.375 140.675 ;
        RECT 79.670 140.465 79.840 140.655 ;
        RECT 84.265 140.465 84.435 140.655 ;
        RECT 84.725 140.485 84.895 140.675 ;
        RECT 88.130 140.465 88.300 140.655 ;
        RECT 89.325 140.465 89.495 140.655 ;
        RECT 90.245 140.485 90.415 140.675 ;
        RECT 92.085 140.465 92.255 140.655 ;
        RECT 95.765 140.485 95.935 140.675 ;
        RECT 97.605 140.465 97.775 140.655 ;
        RECT 101.285 140.485 101.455 140.675 ;
        RECT 104.505 140.485 104.675 140.675 ;
        RECT 107.265 140.465 107.435 140.655 ;
        RECT 107.780 140.515 107.900 140.625 ;
        RECT 109.565 140.465 109.735 140.655 ;
        RECT 110.025 140.485 110.195 140.675 ;
        RECT 113.240 140.465 113.410 140.655 ;
        RECT 114.165 140.510 114.325 140.620 ;
        RECT 115.140 140.515 115.260 140.625 ;
        RECT 115.545 140.465 115.715 140.675 ;
        RECT 119.410 140.485 119.580 140.675 ;
        RECT 120.145 140.485 120.315 140.675 ;
        RECT 122.445 140.485 122.615 140.675 ;
        RECT 126.125 140.465 126.295 140.675 ;
        RECT 127.505 140.465 127.675 140.675 ;
        RECT 35.125 139.555 36.075 139.645 ;
        RECT 37.215 139.595 37.645 140.380 ;
        RECT 38.585 139.755 41.335 140.435 ;
        RECT 38.585 139.555 39.530 139.755 ;
        RECT 41.805 139.655 44.555 140.465 ;
        RECT 44.565 139.655 50.075 140.465 ;
        RECT 50.085 139.655 55.595 140.465 ;
        RECT 55.615 139.555 56.965 140.465 ;
        RECT 57.445 139.655 59.275 140.465 ;
        RECT 59.285 139.555 62.760 140.465 ;
        RECT 62.975 139.595 63.405 140.380 ;
        RECT 63.885 139.555 67.360 140.465 ;
        RECT 67.935 139.785 77.215 140.465 ;
        RECT 67.935 139.665 70.270 139.785 ;
        RECT 67.935 139.555 68.855 139.665 ;
        RECT 74.935 139.565 75.855 139.785 ;
        RECT 77.685 139.655 79.515 140.465 ;
        RECT 79.525 139.555 83.000 140.465 ;
        RECT 83.205 139.655 84.575 140.465 ;
        RECT 84.815 139.785 88.715 140.465 ;
        RECT 87.785 139.555 88.715 139.785 ;
        RECT 88.735 139.595 89.165 140.380 ;
        RECT 89.185 139.685 90.555 140.465 ;
        RECT 90.565 139.655 92.395 140.465 ;
        RECT 92.405 139.655 97.915 140.465 ;
        RECT 98.295 139.785 107.575 140.465 ;
        RECT 98.295 139.665 100.630 139.785 ;
        RECT 98.295 139.555 99.215 139.665 ;
        RECT 105.295 139.565 106.215 139.785 ;
        RECT 108.045 139.655 109.875 140.465 ;
        RECT 110.080 139.555 113.555 140.465 ;
        RECT 114.495 139.595 114.925 140.380 ;
        RECT 115.415 139.555 116.765 140.465 ;
        RECT 117.155 139.785 126.435 140.465 ;
        RECT 117.155 139.665 119.490 139.785 ;
        RECT 117.155 139.555 118.075 139.665 ;
        RECT 124.155 139.565 125.075 139.785 ;
        RECT 126.445 139.655 127.815 140.465 ;
      LAYER nwell ;
        RECT 14.470 136.435 128.010 139.265 ;
      LAYER pwell ;
        RECT 14.665 135.235 16.035 136.045 ;
        RECT 16.505 135.235 20.175 136.045 ;
        RECT 20.185 135.915 21.115 136.145 ;
        RECT 20.185 135.235 24.085 135.915 ;
        RECT 24.335 135.320 24.765 136.105 ;
        RECT 24.785 135.235 28.455 136.045 ;
        RECT 28.465 135.915 29.395 136.145 ;
        RECT 33.745 136.055 34.695 136.145 ;
        RECT 28.465 135.235 32.365 135.915 ;
        RECT 32.765 135.235 34.695 136.055 ;
        RECT 34.905 135.945 35.850 136.145 ;
        RECT 37.665 135.945 38.610 136.145 ;
        RECT 34.905 135.265 37.655 135.945 ;
        RECT 37.665 135.265 40.415 135.945 ;
        RECT 34.905 135.235 35.850 135.265 ;
        RECT 14.805 135.025 14.975 135.235 ;
        RECT 16.240 135.075 16.360 135.185 ;
        RECT 17.565 135.025 17.735 135.215 ;
        RECT 18.025 135.025 18.195 135.215 ;
        RECT 19.405 135.025 19.575 135.215 ;
        RECT 19.865 135.045 20.035 135.235 ;
        RECT 20.600 135.045 20.770 135.235 ;
        RECT 28.145 135.045 28.315 135.235 ;
        RECT 28.880 135.045 29.050 135.235 ;
        RECT 32.765 135.215 32.915 135.235 ;
        RECT 29.985 135.025 30.155 135.215 ;
        RECT 30.500 135.075 30.620 135.185 ;
        RECT 30.905 135.045 31.075 135.215 ;
        RECT 32.745 135.045 32.915 135.215 ;
        RECT 30.925 135.025 31.075 135.045 ;
        RECT 36.610 135.025 36.780 135.215 ;
        RECT 37.340 135.045 37.510 135.265 ;
        RECT 37.665 135.235 38.610 135.265 ;
        RECT 39.185 135.025 39.355 135.215 ;
        RECT 14.665 134.215 16.035 135.025 ;
        RECT 16.515 134.115 17.865 135.025 ;
        RECT 17.885 134.245 19.255 135.025 ;
        RECT 19.275 134.115 20.625 135.025 ;
        RECT 21.015 134.345 30.295 135.025 ;
        RECT 21.015 134.225 23.350 134.345 ;
        RECT 21.015 134.115 21.935 134.225 ;
        RECT 28.015 134.125 28.935 134.345 ;
        RECT 30.925 134.205 32.855 135.025 ;
        RECT 33.295 134.345 37.195 135.025 ;
        RECT 31.905 134.115 32.855 134.205 ;
        RECT 36.265 134.115 37.195 134.345 ;
        RECT 37.215 134.155 37.645 134.940 ;
        RECT 37.665 134.215 39.495 135.025 ;
        RECT 39.650 134.995 39.820 135.215 ;
        RECT 40.100 135.045 40.270 135.265 ;
        RECT 40.885 135.235 43.635 136.045 ;
        RECT 43.645 135.945 44.590 136.145 ;
        RECT 43.645 135.265 46.395 135.945 ;
        RECT 43.645 135.235 44.590 135.265 ;
        RECT 40.620 135.075 40.740 135.185 ;
        RECT 41.310 134.995 42.255 135.025 ;
        RECT 42.410 134.995 42.580 135.215 ;
        RECT 43.325 135.045 43.495 135.235 ;
        RECT 45.170 135.025 45.340 135.215 ;
        RECT 46.080 135.045 46.250 135.265 ;
        RECT 46.405 135.235 49.880 136.145 ;
        RECT 50.095 135.320 50.525 136.105 ;
        RECT 50.545 135.235 53.295 136.045 ;
        RECT 56.505 135.915 57.435 136.145 ;
        RECT 53.535 135.235 57.435 135.915 ;
        RECT 57.905 135.235 59.275 136.015 ;
        RECT 59.285 135.235 61.115 136.045 ;
        RECT 61.125 135.235 64.600 136.145 ;
        RECT 67.460 135.915 68.380 136.145 ;
        RECT 64.915 135.235 68.380 135.915 ;
        RECT 68.485 135.235 71.695 136.145 ;
        RECT 72.165 135.235 75.835 136.045 ;
        RECT 75.855 135.320 76.285 136.105 ;
        RECT 77.225 135.945 78.170 136.145 ;
        RECT 77.225 135.265 79.975 135.945 ;
        RECT 77.225 135.235 78.170 135.265 ;
        RECT 46.550 135.045 46.720 135.235 ;
        RECT 48.850 135.025 49.020 135.215 ;
        RECT 52.985 135.045 53.155 135.235 ;
        RECT 56.850 135.045 57.020 135.235 ;
        RECT 57.640 135.075 57.760 135.185 ;
        RECT 58.045 135.045 58.215 135.235 ;
        RECT 60.805 135.045 60.975 135.235 ;
        RECT 61.270 135.045 61.440 135.235 ;
        RECT 61.725 135.025 61.895 135.215 ;
        RECT 62.645 135.070 62.805 135.180 ;
        RECT 63.570 135.025 63.740 135.215 ;
        RECT 64.945 135.045 65.115 135.235 ;
        RECT 67.705 135.070 67.865 135.180 ;
        RECT 68.625 135.045 68.795 135.235 ;
        RECT 71.900 135.075 72.020 135.185 ;
        RECT 73.225 135.025 73.395 135.215 ;
        RECT 75.525 135.045 75.695 135.235 ;
        RECT 76.905 135.080 77.065 135.190 ;
        RECT 78.745 135.025 78.915 135.215 ;
        RECT 44.070 134.995 45.015 135.025 ;
        RECT 39.505 134.315 42.255 134.995 ;
        RECT 42.265 134.315 45.015 134.995 ;
        RECT 41.310 134.115 42.255 134.315 ;
        RECT 44.070 134.115 45.015 134.315 ;
        RECT 45.025 134.115 48.500 135.025 ;
        RECT 48.705 134.115 52.180 135.025 ;
        RECT 52.755 134.345 62.035 135.025 ;
        RECT 52.755 134.225 55.090 134.345 ;
        RECT 52.755 134.115 53.675 134.225 ;
        RECT 59.755 134.125 60.675 134.345 ;
        RECT 62.975 134.155 63.405 134.940 ;
        RECT 63.425 134.115 66.900 135.025 ;
        RECT 68.025 134.215 73.535 135.025 ;
        RECT 73.545 134.215 79.055 135.025 ;
        RECT 79.210 134.995 79.380 135.215 ;
        RECT 79.660 135.045 79.830 135.265 ;
        RECT 79.985 135.235 83.460 136.145 ;
        RECT 84.035 136.035 84.955 136.145 ;
        RECT 84.035 135.915 86.370 136.035 ;
        RECT 91.035 135.915 91.955 136.135 ;
        RECT 93.325 135.915 94.255 136.145 ;
        RECT 84.035 135.235 93.315 135.915 ;
        RECT 93.325 135.235 97.225 135.915 ;
        RECT 98.120 135.235 101.595 136.145 ;
        RECT 101.615 135.320 102.045 136.105 ;
        RECT 106.185 135.915 107.115 136.145 ;
        RECT 103.215 135.235 107.115 135.915 ;
        RECT 107.125 135.235 108.495 136.015 ;
        RECT 112.625 135.915 113.555 136.145 ;
        RECT 109.655 135.235 113.555 135.915 ;
        RECT 113.935 136.035 114.855 136.145 ;
        RECT 113.935 135.915 116.270 136.035 ;
        RECT 120.935 135.915 121.855 136.135 ;
        RECT 113.935 135.235 123.215 135.915 ;
        RECT 123.225 135.235 124.595 136.015 ;
        RECT 124.605 135.235 126.435 136.045 ;
        RECT 126.445 135.235 127.815 136.045 ;
        RECT 80.130 135.045 80.300 135.235 ;
        RECT 87.025 135.025 87.195 135.215 ;
        RECT 88.405 135.025 88.575 135.215 ;
        RECT 93.005 135.045 93.175 135.235 ;
        RECT 93.740 135.045 93.910 135.235 ;
        RECT 97.660 135.075 97.780 135.185 ;
        RECT 98.525 135.025 98.695 135.215 ;
        RECT 80.870 134.995 81.815 135.025 ;
        RECT 79.065 134.315 81.815 134.995 ;
        RECT 80.870 134.115 81.815 134.315 ;
        RECT 81.825 134.215 87.335 135.025 ;
        RECT 87.355 134.115 88.705 135.025 ;
        RECT 88.735 134.155 89.165 134.940 ;
        RECT 89.555 134.345 98.835 135.025 ;
        RECT 98.845 134.995 99.790 135.025 ;
        RECT 101.280 134.995 101.450 135.235 ;
        RECT 102.665 135.025 102.835 135.215 ;
        RECT 103.180 135.075 103.300 135.185 ;
        RECT 89.555 134.225 91.890 134.345 ;
        RECT 89.555 134.115 90.475 134.225 ;
        RECT 96.555 134.125 97.475 134.345 ;
        RECT 98.845 134.315 101.595 134.995 ;
        RECT 98.845 134.115 99.790 134.315 ;
        RECT 101.615 134.115 102.965 135.025 ;
        RECT 103.445 134.995 104.390 135.025 ;
        RECT 105.880 134.995 106.050 135.215 ;
        RECT 106.350 135.025 106.520 135.215 ;
        RECT 106.530 135.045 106.700 135.235 ;
        RECT 108.185 135.045 108.355 135.235 ;
        RECT 109.105 135.080 109.265 135.190 ;
        RECT 103.445 134.315 106.195 134.995 ;
        RECT 103.445 134.115 104.390 134.315 ;
        RECT 106.205 134.115 109.680 135.025 ;
        RECT 109.885 134.995 110.830 135.025 ;
        RECT 112.320 134.995 112.490 135.215 ;
        RECT 112.970 135.045 113.140 135.235 ;
        RECT 114.165 135.025 114.335 135.215 ;
        RECT 115.140 135.075 115.260 135.185 ;
        RECT 118.765 135.025 118.935 135.215 ;
        RECT 119.225 135.025 119.395 135.215 ;
        RECT 120.660 135.075 120.780 135.185 ;
        RECT 122.905 135.045 123.075 135.235 ;
        RECT 123.365 135.045 123.535 135.235 ;
        RECT 126.125 135.025 126.295 135.235 ;
        RECT 127.505 135.025 127.675 135.235 ;
        RECT 109.885 134.315 112.635 134.995 ;
        RECT 109.885 134.115 110.830 134.315 ;
        RECT 112.645 134.215 114.475 135.025 ;
        RECT 114.495 134.155 114.925 134.940 ;
        RECT 115.405 134.215 119.075 135.025 ;
        RECT 119.085 134.245 120.455 135.025 ;
        RECT 120.925 134.215 126.435 135.025 ;
        RECT 126.445 134.215 127.815 135.025 ;
      LAYER nwell ;
        RECT 14.470 130.995 128.010 133.825 ;
      LAYER pwell ;
        RECT 14.665 129.795 16.035 130.605 ;
        RECT 16.505 129.795 20.175 130.605 ;
        RECT 23.385 130.475 24.315 130.705 ;
        RECT 20.415 129.795 24.315 130.475 ;
        RECT 24.335 129.880 24.765 130.665 ;
        RECT 25.245 129.795 28.915 130.605 ;
        RECT 30.675 130.595 31.595 130.705 ;
        RECT 28.925 129.795 30.295 130.575 ;
        RECT 30.675 130.475 33.010 130.595 ;
        RECT 37.675 130.475 38.595 130.695 ;
        RECT 30.675 129.795 39.955 130.475 ;
        RECT 40.050 129.795 49.155 130.475 ;
        RECT 50.095 129.880 50.525 130.665 ;
        RECT 51.005 129.795 54.675 130.605 ;
        RECT 54.685 129.795 60.195 130.605 ;
        RECT 60.205 129.795 65.715 130.605 ;
        RECT 68.925 130.475 69.855 130.705 ;
        RECT 71.905 130.615 72.855 130.705 ;
        RECT 65.955 129.795 69.855 130.475 ;
        RECT 69.865 129.795 71.695 130.475 ;
        RECT 71.905 129.795 73.835 130.615 ;
        RECT 74.005 129.795 75.835 130.475 ;
        RECT 75.855 129.880 76.285 130.665 ;
        RECT 78.805 130.615 79.755 130.705 ;
        RECT 76.765 129.795 78.595 130.605 ;
        RECT 78.805 129.795 80.735 130.615 ;
        RECT 80.905 129.795 83.655 130.605 ;
        RECT 83.665 129.795 89.175 130.605 ;
        RECT 89.195 129.795 90.545 130.705 ;
        RECT 90.585 129.795 101.595 130.705 ;
        RECT 101.615 129.880 102.045 130.665 ;
        RECT 110.085 130.615 111.035 130.705 ;
        RECT 102.525 129.795 104.355 130.605 ;
        RECT 104.365 129.795 109.875 130.605 ;
        RECT 110.085 129.795 112.015 130.615 ;
        RECT 112.645 129.795 115.395 130.605 ;
        RECT 115.405 129.795 120.915 130.605 ;
        RECT 120.925 129.795 126.435 130.605 ;
        RECT 126.445 129.795 127.815 130.605 ;
        RECT 14.805 129.585 14.975 129.795 ;
        RECT 16.240 129.635 16.360 129.745 ;
        RECT 17.105 129.585 17.275 129.775 ;
        RECT 19.865 129.605 20.035 129.795 ;
        RECT 23.730 129.605 23.900 129.795 ;
        RECT 24.980 129.635 25.100 129.745 ;
        RECT 26.765 129.585 26.935 129.775 ;
        RECT 27.685 129.630 27.845 129.740 ;
        RECT 28.605 129.605 28.775 129.795 ;
        RECT 29.985 129.605 30.155 129.795 ;
        RECT 33.205 129.585 33.375 129.775 ;
        RECT 33.665 129.585 33.835 129.775 ;
        RECT 35.100 129.635 35.220 129.745 ;
        RECT 36.885 129.585 37.055 129.775 ;
        RECT 38.265 129.630 38.425 129.740 ;
        RECT 39.645 129.585 39.815 129.795 ;
        RECT 40.105 129.605 40.275 129.775 ;
        RECT 42.405 129.605 42.575 129.775 ;
        RECT 40.125 129.585 40.275 129.605 ;
        RECT 42.425 129.585 42.575 129.605 ;
        RECT 47.005 129.585 47.175 129.775 ;
        RECT 47.465 129.605 47.635 129.775 ;
        RECT 48.845 129.605 49.015 129.795 ;
        RECT 49.765 129.640 49.925 129.750 ;
        RECT 50.685 129.745 50.855 129.775 ;
        RECT 50.685 129.635 50.860 129.745 ;
        RECT 47.485 129.585 47.635 129.605 ;
        RECT 50.685 129.585 50.855 129.635 ;
        RECT 54.365 129.585 54.535 129.795 ;
        RECT 58.230 129.585 58.400 129.775 ;
        RECT 59.020 129.635 59.140 129.745 ;
        RECT 59.885 129.605 60.055 129.795 ;
        RECT 62.645 129.585 62.815 129.775 ;
        RECT 64.485 129.585 64.655 129.775 ;
        RECT 65.405 129.605 65.575 129.795 ;
        RECT 69.270 129.605 69.440 129.795 ;
        RECT 71.385 129.605 71.555 129.795 ;
        RECT 73.685 129.775 73.835 129.795 ;
        RECT 73.685 129.605 73.855 129.775 ;
        RECT 74.145 129.585 74.315 129.795 ;
        RECT 74.605 129.605 74.775 129.775 ;
        RECT 76.500 129.635 76.620 129.745 ;
        RECT 76.905 129.605 77.075 129.775 ;
        RECT 78.285 129.605 78.455 129.795 ;
        RECT 80.585 129.775 80.735 129.795 ;
        RECT 80.585 129.605 80.755 129.775 ;
        RECT 74.625 129.585 74.775 129.605 ;
        RECT 76.925 129.585 77.075 129.605 ;
        RECT 82.610 129.585 82.780 129.775 ;
        RECT 83.345 129.605 83.515 129.795 ;
        RECT 85.185 129.605 85.355 129.775 ;
        RECT 85.185 129.585 85.335 129.605 ;
        RECT 87.025 129.585 87.195 129.775 ;
        RECT 87.485 129.585 87.655 129.775 ;
        RECT 88.865 129.605 89.035 129.795 ;
        RECT 89.325 129.745 89.495 129.795 ;
        RECT 89.325 129.635 89.500 129.745 ;
        RECT 89.325 129.605 89.495 129.635 ;
        RECT 90.060 129.585 90.230 129.775 ;
        RECT 93.980 129.635 94.100 129.745 ;
        RECT 94.385 129.585 94.555 129.775 ;
        RECT 95.765 129.585 95.935 129.775 ;
        RECT 101.280 129.605 101.450 129.795 ;
        RECT 102.260 129.635 102.380 129.745 ;
        RECT 104.045 129.605 104.215 129.795 ;
        RECT 106.805 129.605 106.975 129.775 ;
        RECT 109.105 129.605 109.275 129.775 ;
        RECT 109.565 129.605 109.735 129.795 ;
        RECT 111.865 129.775 112.015 129.795 ;
        RECT 111.865 129.605 112.035 129.775 ;
        RECT 112.380 129.635 112.500 129.745 ;
        RECT 113.705 129.605 113.875 129.775 ;
        RECT 115.085 129.745 115.255 129.795 ;
        RECT 114.220 129.635 114.340 129.745 ;
        RECT 115.085 129.635 115.260 129.745 ;
        RECT 115.085 129.605 115.255 129.635 ;
        RECT 106.805 129.585 106.955 129.605 ;
        RECT 109.105 129.585 109.255 129.605 ;
        RECT 14.665 128.775 16.035 129.585 ;
        RECT 16.045 128.775 17.415 129.585 ;
        RECT 17.795 128.905 27.075 129.585 ;
        RECT 17.795 128.785 20.130 128.905 ;
        RECT 17.795 128.675 18.715 128.785 ;
        RECT 24.795 128.685 25.715 128.905 ;
        RECT 28.005 128.775 33.515 129.585 ;
        RECT 33.535 128.675 34.885 129.585 ;
        RECT 35.365 128.775 37.195 129.585 ;
        RECT 37.215 128.715 37.645 129.500 ;
        RECT 38.585 128.805 39.955 129.585 ;
        RECT 40.125 128.765 42.055 129.585 ;
        RECT 42.425 128.765 44.355 129.585 ;
        RECT 45.225 128.775 47.315 129.585 ;
        RECT 47.485 128.765 49.415 129.585 ;
        RECT 49.625 128.775 50.995 129.585 ;
        RECT 51.005 128.775 54.675 129.585 ;
        RECT 54.915 128.905 58.815 129.585 ;
        RECT 41.105 128.675 42.055 128.765 ;
        RECT 43.405 128.675 44.355 128.765 ;
        RECT 48.465 128.675 49.415 128.765 ;
        RECT 57.885 128.675 58.815 128.905 ;
        RECT 59.285 128.775 62.955 129.585 ;
        RECT 62.975 128.715 63.405 129.500 ;
        RECT 63.425 128.775 64.795 129.585 ;
        RECT 65.175 128.905 74.455 129.585 ;
        RECT 65.175 128.785 67.510 128.905 ;
        RECT 65.175 128.675 66.095 128.785 ;
        RECT 72.175 128.685 73.095 128.905 ;
        RECT 74.625 128.765 76.555 129.585 ;
        RECT 76.925 128.765 78.855 129.585 ;
        RECT 79.295 128.905 83.195 129.585 ;
        RECT 75.605 128.675 76.555 128.765 ;
        RECT 77.905 128.675 78.855 128.765 ;
        RECT 82.265 128.675 83.195 128.905 ;
        RECT 83.405 128.765 85.335 129.585 ;
        RECT 85.505 128.775 87.335 129.585 ;
        RECT 87.345 128.805 88.715 129.585 ;
        RECT 83.405 128.675 84.355 128.765 ;
        RECT 88.735 128.715 89.165 129.500 ;
        RECT 89.645 128.905 93.545 129.585 ;
        RECT 89.645 128.675 90.575 128.905 ;
        RECT 94.245 128.805 95.615 129.585 ;
        RECT 95.625 128.905 104.730 129.585 ;
        RECT 105.025 128.765 106.955 129.585 ;
        RECT 107.325 128.765 109.255 129.585 ;
        RECT 109.585 129.585 109.735 129.605 ;
        RECT 113.705 129.585 113.855 129.605 ;
        RECT 117.845 129.585 118.015 129.775 ;
        RECT 118.305 129.585 118.475 129.775 ;
        RECT 119.685 129.585 119.855 129.775 ;
        RECT 120.605 129.605 120.775 129.795 ;
        RECT 126.125 129.585 126.295 129.795 ;
        RECT 127.505 129.585 127.675 129.795 ;
        RECT 109.585 128.765 111.515 129.585 ;
        RECT 105.025 128.675 105.975 128.765 ;
        RECT 107.325 128.675 108.275 128.765 ;
        RECT 110.565 128.675 111.515 128.765 ;
        RECT 111.925 128.765 113.855 129.585 ;
        RECT 111.925 128.675 112.875 128.765 ;
        RECT 114.495 128.715 114.925 129.500 ;
        RECT 115.405 128.775 118.155 129.585 ;
        RECT 118.175 128.675 119.525 129.585 ;
        RECT 119.545 128.805 120.915 129.585 ;
        RECT 120.925 128.775 126.435 129.585 ;
        RECT 126.445 128.775 127.815 129.585 ;
      LAYER nwell ;
        RECT 14.470 125.555 128.010 128.385 ;
      LAYER pwell ;
        RECT 14.665 124.355 16.035 125.165 ;
        RECT 16.045 124.355 17.415 125.165 ;
        RECT 17.425 124.355 21.095 125.165 ;
        RECT 21.115 124.355 22.465 125.265 ;
        RECT 22.945 124.355 24.315 125.135 ;
        RECT 24.335 124.440 24.765 125.225 ;
        RECT 37.885 125.175 38.835 125.265 ;
        RECT 25.705 124.355 31.215 125.165 ;
        RECT 31.225 124.355 36.735 125.165 ;
        RECT 36.905 124.355 38.835 125.175 ;
        RECT 40.625 125.175 41.575 125.265 ;
        RECT 43.865 125.175 44.815 125.265 ;
        RECT 39.045 124.355 40.415 125.165 ;
        RECT 40.625 124.355 42.555 125.175 ;
        RECT 14.805 124.145 14.975 124.355 ;
        RECT 17.105 124.145 17.275 124.355 ;
        RECT 20.785 124.165 20.955 124.355 ;
        RECT 22.165 124.165 22.335 124.355 ;
        RECT 22.625 124.305 22.795 124.335 ;
        RECT 22.625 124.195 22.800 124.305 ;
        RECT 22.625 124.145 22.795 124.195 ;
        RECT 23.085 124.165 23.255 124.355 ;
        RECT 25.385 124.200 25.545 124.310 ;
        RECT 26.490 124.145 26.660 124.335 ;
        RECT 27.280 124.195 27.400 124.305 ;
        RECT 30.905 124.165 31.075 124.355 ;
        RECT 32.745 124.145 32.915 124.335 ;
        RECT 36.425 124.165 36.595 124.355 ;
        RECT 36.905 124.335 37.055 124.355 ;
        RECT 36.610 124.145 36.780 124.335 ;
        RECT 36.885 124.165 37.055 124.335 ;
        RECT 37.860 124.195 37.980 124.305 ;
        RECT 40.105 124.165 40.275 124.355 ;
        RECT 42.405 124.335 42.555 124.355 ;
        RECT 42.885 124.355 44.815 125.175 ;
        RECT 45.225 125.175 46.175 125.265 ;
        RECT 45.225 124.355 47.155 125.175 ;
        RECT 47.335 124.355 50.075 125.035 ;
        RECT 50.095 124.440 50.525 125.225 ;
        RECT 50.545 124.355 52.375 125.165 ;
        RECT 52.385 124.355 57.895 125.165 ;
        RECT 57.905 124.355 59.275 125.135 ;
        RECT 62.485 125.035 63.415 125.265 ;
        RECT 59.515 124.355 63.415 125.035 ;
        RECT 63.425 124.355 64.795 125.165 ;
        RECT 64.805 124.355 68.475 125.165 ;
        RECT 68.495 124.355 69.845 125.265 ;
        RECT 70.325 124.355 71.695 125.135 ;
        RECT 72.625 124.355 75.365 125.035 ;
        RECT 75.855 124.440 76.285 125.225 ;
        RECT 76.305 124.355 78.135 125.165 ;
        RECT 78.515 125.155 79.435 125.265 ;
        RECT 78.515 125.035 80.850 125.155 ;
        RECT 85.515 125.035 86.435 125.255 ;
        RECT 78.515 124.355 87.795 125.035 ;
        RECT 87.805 124.355 89.635 125.165 ;
        RECT 91.005 125.035 91.925 125.255 ;
        RECT 98.005 125.155 98.925 125.265 ;
        RECT 100.445 125.175 101.395 125.265 ;
        RECT 96.590 125.035 98.925 125.155 ;
        RECT 89.645 124.355 98.925 125.035 ;
        RECT 99.465 124.355 101.395 125.175 ;
        RECT 101.615 124.440 102.045 125.225 ;
        RECT 102.065 124.355 105.735 125.165 ;
        RECT 105.745 124.355 111.255 125.165 ;
        RECT 114.465 125.035 115.395 125.265 ;
        RECT 111.495 124.355 115.395 125.035 ;
        RECT 115.775 125.155 116.695 125.265 ;
        RECT 115.775 125.035 118.110 125.155 ;
        RECT 122.775 125.035 123.695 125.255 ;
        RECT 115.775 124.355 125.055 125.035 ;
        RECT 125.065 124.355 126.435 125.165 ;
        RECT 126.445 124.355 127.815 125.165 ;
        RECT 42.885 124.335 43.035 124.355 ;
        RECT 41.485 124.145 41.655 124.335 ;
        RECT 42.405 124.165 42.575 124.335 ;
        RECT 42.865 124.165 43.035 124.335 ;
        RECT 47.005 124.335 47.155 124.355 ;
        RECT 47.005 124.145 47.175 124.335 ;
        RECT 49.765 124.165 49.935 124.355 ;
        RECT 52.065 124.165 52.235 124.355 ;
        RECT 52.525 124.145 52.695 124.335 ;
        RECT 57.585 124.165 57.755 124.355 ;
        RECT 58.045 124.165 58.215 124.355 ;
        RECT 62.185 124.145 62.355 124.335 ;
        RECT 62.700 124.195 62.820 124.305 ;
        RECT 62.830 124.165 63.000 124.355 ;
        RECT 63.620 124.195 63.740 124.305 ;
        RECT 64.485 124.165 64.655 124.355 ;
        RECT 67.430 124.145 67.600 124.335 ;
        RECT 68.165 124.165 68.335 124.355 ;
        RECT 69.545 124.165 69.715 124.355 ;
        RECT 70.060 124.195 70.180 124.305 ;
        RECT 70.465 124.145 70.635 124.355 ;
        RECT 72.305 124.200 72.465 124.310 ;
        RECT 72.765 124.165 72.935 124.355 ;
        RECT 75.580 124.195 75.700 124.305 ;
        RECT 75.985 124.145 76.155 124.335 ;
        RECT 77.825 124.165 77.995 124.355 ;
        RECT 81.505 124.145 81.675 124.335 ;
        RECT 82.885 124.145 83.055 124.335 ;
        RECT 83.400 124.195 83.520 124.305 ;
        RECT 83.805 124.145 83.975 124.335 ;
        RECT 87.485 124.165 87.655 124.355 ;
        RECT 88.405 124.145 88.575 124.335 ;
        RECT 89.325 124.165 89.495 124.355 ;
        RECT 89.785 124.165 89.955 124.355 ;
        RECT 99.465 124.335 99.615 124.355 ;
        RECT 92.545 124.145 92.715 124.335 ;
        RECT 93.005 124.145 93.175 124.335 ;
        RECT 95.305 124.145 95.475 124.335 ;
        RECT 98.985 124.145 99.155 124.335 ;
        RECT 99.445 124.165 99.615 124.335 ;
        RECT 104.505 124.145 104.675 124.335 ;
        RECT 105.425 124.165 105.595 124.355 ;
        RECT 110.025 124.145 110.195 124.335 ;
        RECT 110.945 124.165 111.115 124.355 ;
        RECT 113.890 124.145 114.060 124.335 ;
        RECT 114.810 124.165 114.980 124.355 ;
        RECT 115.140 124.195 115.260 124.305 ;
        RECT 124.745 124.145 124.915 124.355 ;
        RECT 126.125 124.145 126.295 124.355 ;
        RECT 127.505 124.145 127.675 124.355 ;
        RECT 14.665 123.335 16.035 124.145 ;
        RECT 16.045 123.335 17.415 124.145 ;
        RECT 17.425 123.335 22.935 124.145 ;
        RECT 23.175 123.465 27.075 124.145 ;
        RECT 26.145 123.235 27.075 123.465 ;
        RECT 27.545 123.335 33.055 124.145 ;
        RECT 33.295 123.465 37.195 124.145 ;
        RECT 36.265 123.235 37.195 123.465 ;
        RECT 37.215 123.275 37.645 124.060 ;
        RECT 38.125 123.335 41.795 124.145 ;
        RECT 41.805 123.335 47.315 124.145 ;
        RECT 47.325 123.335 52.835 124.145 ;
        RECT 53.215 123.465 62.495 124.145 ;
        RECT 53.215 123.345 55.550 123.465 ;
        RECT 53.215 123.235 54.135 123.345 ;
        RECT 60.215 123.245 61.135 123.465 ;
        RECT 62.975 123.275 63.405 124.060 ;
        RECT 64.115 123.465 68.015 124.145 ;
        RECT 67.085 123.235 68.015 123.465 ;
        RECT 68.025 123.335 70.775 124.145 ;
        RECT 70.785 123.335 76.295 124.145 ;
        RECT 76.305 123.335 81.815 124.145 ;
        RECT 81.835 123.235 83.185 124.145 ;
        RECT 83.665 123.365 85.035 124.145 ;
        RECT 85.045 123.335 88.715 124.145 ;
        RECT 88.735 123.275 89.165 124.060 ;
        RECT 89.185 123.335 92.855 124.145 ;
        RECT 92.875 123.235 94.225 124.145 ;
        RECT 94.245 123.335 95.615 124.145 ;
        RECT 95.625 123.335 99.295 124.145 ;
        RECT 99.305 123.335 104.815 124.145 ;
        RECT 104.825 123.335 110.335 124.145 ;
        RECT 110.575 123.465 114.475 124.145 ;
        RECT 113.545 123.235 114.475 123.465 ;
        RECT 114.495 123.275 114.925 124.060 ;
        RECT 115.775 123.465 125.055 124.145 ;
        RECT 115.775 123.345 118.110 123.465 ;
        RECT 115.775 123.235 116.695 123.345 ;
        RECT 122.775 123.245 123.695 123.465 ;
        RECT 125.065 123.335 126.435 124.145 ;
        RECT 126.445 123.335 127.815 124.145 ;
      LAYER nwell ;
        RECT 14.470 120.115 128.010 122.945 ;
      LAYER pwell ;
        RECT 14.665 118.915 16.035 119.725 ;
        RECT 16.505 118.915 20.175 119.725 ;
        RECT 20.185 119.595 21.115 119.825 ;
        RECT 20.185 118.915 24.085 119.595 ;
        RECT 24.335 119.000 24.765 119.785 ;
        RECT 24.785 118.915 26.155 119.725 ;
        RECT 26.165 118.915 27.535 119.695 ;
        RECT 27.545 118.915 30.295 119.725 ;
        RECT 30.675 119.715 31.595 119.825 ;
        RECT 30.675 119.595 33.010 119.715 ;
        RECT 37.675 119.595 38.595 119.815 ;
        RECT 39.965 119.595 40.895 119.825 ;
        RECT 30.675 118.915 39.955 119.595 ;
        RECT 39.965 118.915 43.865 119.595 ;
        RECT 44.565 118.915 45.935 119.695 ;
        RECT 49.145 119.595 50.075 119.825 ;
        RECT 46.175 118.915 50.075 119.595 ;
        RECT 50.095 119.000 50.525 119.785 ;
        RECT 50.555 118.915 51.905 119.825 ;
        RECT 51.925 118.915 53.295 119.725 ;
        RECT 53.445 118.915 56.055 119.825 ;
        RECT 56.995 118.915 58.345 119.825 ;
        RECT 59.655 119.715 60.575 119.825 ;
        RECT 59.655 119.595 61.990 119.715 ;
        RECT 66.655 119.595 67.575 119.815 ;
        RECT 59.655 118.915 68.935 119.595 ;
        RECT 68.945 118.915 70.315 119.695 ;
        RECT 70.785 118.915 74.455 119.725 ;
        RECT 74.475 118.915 75.825 119.825 ;
        RECT 75.855 119.000 76.285 119.785 ;
        RECT 79.965 119.595 80.895 119.825 ;
        RECT 76.995 118.915 80.895 119.595 ;
        RECT 80.905 118.915 82.275 119.695 ;
        RECT 82.295 118.915 83.645 119.825 ;
        RECT 84.125 118.915 85.495 119.695 ;
        RECT 85.505 118.915 91.015 119.725 ;
        RECT 91.025 119.595 91.955 119.825 ;
        RECT 91.025 118.915 94.925 119.595 ;
        RECT 95.625 118.915 97.455 119.725 ;
        RECT 100.665 119.595 101.595 119.825 ;
        RECT 97.695 118.915 101.595 119.595 ;
        RECT 101.615 119.000 102.045 119.785 ;
        RECT 102.065 118.915 103.435 119.725 ;
        RECT 103.455 118.915 104.805 119.825 ;
        RECT 108.025 119.595 108.955 119.825 ;
        RECT 105.055 118.915 108.955 119.595 ;
        RECT 109.335 119.715 110.255 119.825 ;
        RECT 109.335 119.595 111.670 119.715 ;
        RECT 116.335 119.595 117.255 119.815 ;
        RECT 109.335 118.915 118.615 119.595 ;
        RECT 118.635 118.915 119.985 119.825 ;
        RECT 120.465 118.915 121.835 119.695 ;
        RECT 122.765 118.915 126.435 119.725 ;
        RECT 126.445 118.915 127.815 119.725 ;
        RECT 14.805 118.705 14.975 118.915 ;
        RECT 16.240 118.755 16.360 118.865 ;
        RECT 17.565 118.705 17.735 118.895 ;
        RECT 19.865 118.725 20.035 118.915 ;
        RECT 20.600 118.725 20.770 118.915 ;
        RECT 25.845 118.725 26.015 118.915 ;
        RECT 27.225 118.705 27.395 118.915 ;
        RECT 27.685 118.705 27.855 118.895 ;
        RECT 29.985 118.725 30.155 118.915 ;
        RECT 39.645 118.725 39.815 118.915 ;
        RECT 40.380 118.725 40.550 118.915 ;
        RECT 44.300 118.755 44.420 118.865 ;
        RECT 45.625 118.725 45.795 118.915 ;
        RECT 47.005 118.705 47.175 118.895 ;
        RECT 49.490 118.725 49.660 118.915 ;
        RECT 50.685 118.725 50.855 118.915 ;
        RECT 52.985 118.725 53.155 118.915 ;
        RECT 55.740 118.725 55.910 118.915 ;
        RECT 56.665 118.705 56.835 118.895 ;
        RECT 57.585 118.750 57.745 118.860 ;
        RECT 58.045 118.725 58.215 118.915 ;
        RECT 58.965 118.760 59.125 118.870 ;
        RECT 61.265 118.705 61.435 118.895 ;
        RECT 61.725 118.705 61.895 118.895 ;
        RECT 68.625 118.725 68.795 118.915 ;
        RECT 70.005 118.725 70.175 118.915 ;
        RECT 70.520 118.755 70.640 118.865 ;
        RECT 72.765 118.705 72.935 118.895 ;
        RECT 74.145 118.725 74.315 118.915 ;
        RECT 74.605 118.725 74.775 118.915 ;
        RECT 76.500 118.755 76.620 118.865 ;
        RECT 80.310 118.725 80.480 118.915 ;
        RECT 81.965 118.725 82.135 118.915 ;
        RECT 82.425 118.705 82.595 118.895 ;
        RECT 83.160 118.705 83.330 118.895 ;
        RECT 83.345 118.725 83.515 118.915 ;
        RECT 83.860 118.755 83.980 118.865 ;
        RECT 84.265 118.725 84.435 118.915 ;
        RECT 87.080 118.755 87.200 118.865 ;
        RECT 87.485 118.705 87.655 118.895 ;
        RECT 89.325 118.705 89.495 118.895 ;
        RECT 90.705 118.705 90.875 118.915 ;
        RECT 91.440 118.725 91.610 118.915 ;
        RECT 92.545 118.750 92.705 118.860 ;
        RECT 95.360 118.755 95.480 118.865 ;
        RECT 97.145 118.725 97.315 118.915 ;
        RECT 101.010 118.725 101.180 118.915 ;
        RECT 102.205 118.705 102.375 118.895 ;
        RECT 103.125 118.725 103.295 118.915 ;
        RECT 103.585 118.725 103.755 118.915 ;
        RECT 108.370 118.725 108.540 118.915 ;
        RECT 111.865 118.705 112.035 118.895 ;
        RECT 112.785 118.750 112.945 118.860 ;
        RECT 114.165 118.705 114.335 118.895 ;
        RECT 115.140 118.755 115.260 118.865 ;
        RECT 115.545 118.705 115.715 118.895 ;
        RECT 116.980 118.755 117.100 118.865 ;
        RECT 118.305 118.725 118.475 118.915 ;
        RECT 118.765 118.725 118.935 118.915 ;
        RECT 120.200 118.755 120.320 118.865 ;
        RECT 120.605 118.705 120.775 118.915 ;
        RECT 122.445 118.760 122.605 118.870 ;
        RECT 126.125 118.705 126.295 118.915 ;
        RECT 127.505 118.705 127.675 118.915 ;
        RECT 14.665 117.895 16.035 118.705 ;
        RECT 16.515 117.795 17.865 118.705 ;
        RECT 18.255 118.025 27.535 118.705 ;
        RECT 27.545 118.025 36.825 118.705 ;
        RECT 18.255 117.905 20.590 118.025 ;
        RECT 18.255 117.795 19.175 117.905 ;
        RECT 25.255 117.805 26.175 118.025 ;
        RECT 28.905 117.805 29.825 118.025 ;
        RECT 34.490 117.905 36.825 118.025 ;
        RECT 35.905 117.795 36.825 117.905 ;
        RECT 37.215 117.835 37.645 118.620 ;
        RECT 38.035 118.025 47.315 118.705 ;
        RECT 47.695 118.025 56.975 118.705 ;
        RECT 38.035 117.905 40.370 118.025 ;
        RECT 38.035 117.795 38.955 117.905 ;
        RECT 45.035 117.805 45.955 118.025 ;
        RECT 47.695 117.905 50.030 118.025 ;
        RECT 47.695 117.795 48.615 117.905 ;
        RECT 54.695 117.805 55.615 118.025 ;
        RECT 57.905 117.895 61.575 118.705 ;
        RECT 61.595 117.795 62.945 118.705 ;
        RECT 62.975 117.835 63.405 118.620 ;
        RECT 63.795 118.025 73.075 118.705 ;
        RECT 73.455 118.025 82.735 118.705 ;
        RECT 82.745 118.025 86.645 118.705 ;
        RECT 63.795 117.905 66.130 118.025 ;
        RECT 63.795 117.795 64.715 117.905 ;
        RECT 70.795 117.805 71.715 118.025 ;
        RECT 73.455 117.905 75.790 118.025 ;
        RECT 73.455 117.795 74.375 117.905 ;
        RECT 80.455 117.805 81.375 118.025 ;
        RECT 82.745 117.795 83.675 118.025 ;
        RECT 87.345 117.925 88.715 118.705 ;
        RECT 88.735 117.835 89.165 118.620 ;
        RECT 89.195 117.795 90.545 118.705 ;
        RECT 90.575 117.795 91.925 118.705 ;
        RECT 93.235 118.025 102.515 118.705 ;
        RECT 102.895 118.025 112.175 118.705 ;
        RECT 93.235 117.905 95.570 118.025 ;
        RECT 93.235 117.795 94.155 117.905 ;
        RECT 100.235 117.805 101.155 118.025 ;
        RECT 102.895 117.905 105.230 118.025 ;
        RECT 102.895 117.795 103.815 117.905 ;
        RECT 109.895 117.805 110.815 118.025 ;
        RECT 113.115 117.795 114.465 118.705 ;
        RECT 114.495 117.835 114.925 118.620 ;
        RECT 115.405 117.925 116.775 118.705 ;
        RECT 117.245 117.895 120.915 118.705 ;
        RECT 120.925 117.895 126.435 118.705 ;
        RECT 126.445 117.895 127.815 118.705 ;
      LAYER nwell ;
        RECT 14.470 114.675 128.010 117.505 ;
      LAYER pwell ;
        RECT 14.665 113.475 16.035 114.285 ;
        RECT 16.045 113.475 17.415 114.285 ;
        RECT 17.425 113.475 21.095 114.285 ;
        RECT 21.105 113.475 22.475 114.255 ;
        RECT 22.495 113.475 23.845 114.385 ;
        RECT 24.335 113.560 24.765 114.345 ;
        RECT 26.145 114.155 27.065 114.375 ;
        RECT 33.145 114.275 34.065 114.385 ;
        RECT 31.730 114.155 34.065 114.275 ;
        RECT 24.785 113.475 34.065 114.155 ;
        RECT 34.915 113.475 36.265 114.385 ;
        RECT 36.745 113.475 38.115 114.255 ;
        RECT 39.045 113.475 40.415 114.255 ;
        RECT 40.425 113.475 44.095 114.285 ;
        RECT 44.115 113.475 45.465 114.385 ;
        RECT 45.485 114.155 46.415 114.385 ;
        RECT 45.485 113.475 49.385 114.155 ;
        RECT 50.095 113.560 50.525 114.345 ;
        RECT 50.545 113.475 52.375 114.285 ;
        RECT 52.385 113.475 53.755 114.255 ;
        RECT 53.765 113.475 55.135 114.285 ;
        RECT 55.145 113.475 60.655 114.285 ;
        RECT 60.665 113.475 66.175 114.285 ;
        RECT 66.195 113.475 67.545 114.385 ;
        RECT 68.025 113.475 69.395 114.255 ;
        RECT 70.325 113.475 75.835 114.285 ;
        RECT 75.855 113.560 76.285 114.345 ;
        RECT 77.595 114.275 78.515 114.385 ;
        RECT 77.595 114.155 79.930 114.275 ;
        RECT 84.595 114.155 85.515 114.375 ;
        RECT 88.705 114.155 89.625 114.375 ;
        RECT 95.705 114.275 96.625 114.385 ;
        RECT 94.290 114.155 96.625 114.275 ;
        RECT 77.595 113.475 86.875 114.155 ;
        RECT 87.345 113.475 96.625 114.155 ;
        RECT 97.465 113.475 100.215 114.285 ;
        RECT 100.225 113.475 101.595 114.255 ;
        RECT 101.615 113.560 102.045 114.345 ;
        RECT 102.525 113.475 108.035 114.285 ;
        RECT 108.045 113.475 109.415 114.255 ;
        RECT 109.425 113.475 111.255 114.285 ;
        RECT 114.465 114.155 115.395 114.385 ;
        RECT 111.495 113.475 115.395 114.155 ;
        RECT 115.405 113.475 120.915 114.285 ;
        RECT 120.925 113.475 126.435 114.285 ;
        RECT 126.445 113.475 127.815 114.285 ;
        RECT 14.805 113.265 14.975 113.475 ;
        RECT 17.105 113.285 17.275 113.475 ;
        RECT 20.785 113.285 20.955 113.475 ;
        RECT 21.245 113.285 21.415 113.475 ;
        RECT 23.545 113.285 23.715 113.475 ;
        RECT 24.060 113.315 24.180 113.425 ;
        RECT 24.925 113.285 25.095 113.475 ;
        RECT 26.305 113.265 26.475 113.455 ;
        RECT 28.145 113.265 28.315 113.455 ;
        RECT 33.665 113.265 33.835 113.455 ;
        RECT 34.640 113.315 34.760 113.425 ;
        RECT 35.045 113.265 35.215 113.455 ;
        RECT 35.965 113.285 36.135 113.475 ;
        RECT 36.480 113.315 36.600 113.425 ;
        RECT 36.885 113.265 37.055 113.475 ;
        RECT 37.860 113.315 37.980 113.425 ;
        RECT 38.725 113.320 38.885 113.430 ;
        RECT 40.105 113.285 40.275 113.475 ;
        RECT 43.785 113.285 43.955 113.475 ;
        RECT 45.165 113.285 45.335 113.475 ;
        RECT 45.900 113.285 46.070 113.475 ;
        RECT 47.005 113.265 47.175 113.455 ;
        RECT 47.925 113.310 48.085 113.420 ;
        RECT 49.820 113.315 49.940 113.425 ;
        RECT 51.605 113.265 51.775 113.455 ;
        RECT 52.065 113.285 52.235 113.475 ;
        RECT 52.525 113.285 52.695 113.475 ;
        RECT 54.825 113.285 54.995 113.475 ;
        RECT 57.125 113.265 57.295 113.455 ;
        RECT 60.345 113.285 60.515 113.475 ;
        RECT 62.645 113.265 62.815 113.455 ;
        RECT 63.620 113.315 63.740 113.425 ;
        RECT 65.865 113.285 66.035 113.475 ;
        RECT 66.325 113.285 66.495 113.475 ;
        RECT 67.760 113.315 67.880 113.425 ;
        RECT 68.165 113.285 68.335 113.475 ;
        RECT 69.085 113.265 69.255 113.455 ;
        RECT 70.005 113.320 70.165 113.430 ;
        RECT 74.605 113.265 74.775 113.455 ;
        RECT 75.525 113.285 75.695 113.475 ;
        RECT 76.905 113.320 77.065 113.430 ;
        RECT 80.125 113.265 80.295 113.455 ;
        RECT 81.505 113.265 81.675 113.455 ;
        RECT 82.885 113.265 83.055 113.455 ;
        RECT 86.565 113.285 86.735 113.475 ;
        RECT 87.080 113.315 87.200 113.425 ;
        RECT 87.485 113.285 87.655 113.475 ;
        RECT 88.405 113.265 88.575 113.455 ;
        RECT 92.545 113.265 92.715 113.455 ;
        RECT 93.005 113.265 93.175 113.455 ;
        RECT 97.200 113.315 97.320 113.425 ;
        RECT 99.905 113.285 100.075 113.475 ;
        RECT 101.285 113.285 101.455 113.475 ;
        RECT 102.260 113.315 102.380 113.425 ;
        RECT 103.125 113.285 103.295 113.455 ;
        RECT 107.725 113.285 107.895 113.475 ;
        RECT 108.185 113.285 108.355 113.475 ;
        RECT 108.645 113.265 108.815 113.455 ;
        RECT 110.945 113.285 111.115 113.475 ;
        RECT 114.165 113.265 114.335 113.455 ;
        RECT 114.810 113.285 114.980 113.475 ;
        RECT 115.545 113.310 115.705 113.420 ;
        RECT 119.225 113.265 119.395 113.455 ;
        RECT 119.685 113.265 119.855 113.455 ;
        RECT 120.605 113.285 120.775 113.475 ;
        RECT 121.985 113.265 122.155 113.455 ;
        RECT 123.365 113.265 123.535 113.455 ;
        RECT 126.125 113.265 126.295 113.475 ;
        RECT 127.505 113.265 127.675 113.475 ;
        RECT 14.665 112.455 16.035 113.265 ;
        RECT 16.245 112.585 26.615 113.265 ;
        RECT 16.245 112.355 18.455 112.585 ;
        RECT 21.175 112.365 22.105 112.585 ;
        RECT 26.625 112.455 28.455 113.265 ;
        RECT 28.465 112.455 33.975 113.265 ;
        RECT 33.995 112.355 35.345 113.265 ;
        RECT 35.365 112.455 37.195 113.265 ;
        RECT 37.215 112.395 37.645 113.180 ;
        RECT 38.210 112.585 47.315 113.265 ;
        RECT 48.245 112.455 51.915 113.265 ;
        RECT 51.925 112.455 57.435 113.265 ;
        RECT 57.445 112.455 62.955 113.265 ;
        RECT 62.975 112.395 63.405 113.180 ;
        RECT 63.885 112.455 69.395 113.265 ;
        RECT 69.405 112.455 74.915 113.265 ;
        RECT 74.925 112.455 80.435 113.265 ;
        RECT 80.455 112.355 81.805 113.265 ;
        RECT 81.825 112.455 83.195 113.265 ;
        RECT 83.205 112.455 88.715 113.265 ;
        RECT 88.735 112.395 89.165 113.180 ;
        RECT 89.185 112.455 92.855 113.265 ;
        RECT 92.865 112.585 101.970 113.265 ;
        RECT 102.065 112.585 103.020 113.265 ;
        RECT 103.445 112.455 108.955 113.265 ;
        RECT 108.965 112.455 114.475 113.265 ;
        RECT 114.495 112.395 114.925 113.180 ;
        RECT 115.865 112.455 119.535 113.265 ;
        RECT 119.555 112.355 120.905 113.265 ;
        RECT 120.925 112.485 122.295 113.265 ;
        RECT 122.305 112.485 123.675 113.265 ;
        RECT 123.685 112.455 126.435 113.265 ;
        RECT 126.445 112.455 127.815 113.265 ;
      LAYER nwell ;
        RECT 14.470 109.235 128.010 112.065 ;
      LAYER pwell ;
        RECT 14.665 108.035 16.035 108.845 ;
        RECT 16.965 108.035 20.635 108.845 ;
        RECT 20.655 108.035 22.005 108.945 ;
        RECT 22.955 108.035 24.305 108.945 ;
        RECT 24.335 108.120 24.765 108.905 ;
        RECT 24.785 108.035 27.535 108.845 ;
        RECT 27.545 108.035 28.915 108.815 ;
        RECT 28.925 108.035 30.755 108.845 ;
        RECT 30.775 108.035 32.125 108.945 ;
        RECT 32.145 108.035 33.515 108.815 ;
        RECT 34.445 108.035 35.815 108.815 ;
        RECT 36.285 108.035 39.035 108.845 ;
        RECT 39.045 108.035 44.555 108.845 ;
        RECT 44.565 108.035 50.075 108.845 ;
        RECT 50.095 108.120 50.525 108.905 ;
        RECT 51.005 108.035 52.375 108.815 ;
        RECT 53.305 108.035 56.975 108.845 ;
        RECT 56.985 108.035 58.355 108.815 ;
        RECT 58.365 108.035 59.735 108.845 ;
        RECT 59.745 108.035 62.355 108.945 ;
        RECT 62.965 108.035 64.795 108.845 ;
        RECT 64.815 108.035 66.165 108.945 ;
        RECT 66.645 108.035 68.475 108.845 ;
        RECT 68.485 108.035 69.855 108.815 ;
        RECT 70.325 108.035 75.835 108.845 ;
        RECT 75.855 108.120 76.285 108.905 ;
        RECT 76.315 108.035 77.665 108.945 ;
        RECT 77.695 108.035 79.045 108.945 ;
        RECT 79.985 108.035 82.595 108.945 ;
        RECT 82.745 108.035 84.115 108.815 ;
        RECT 84.585 108.035 87.335 108.845 ;
        RECT 87.355 108.035 88.705 108.945 ;
        RECT 88.725 108.035 92.395 108.845 ;
        RECT 92.415 108.035 93.765 108.945 ;
        RECT 93.785 108.035 95.155 108.815 ;
        RECT 95.165 108.035 96.535 108.845 ;
        RECT 96.545 108.035 100.215 108.845 ;
        RECT 100.225 108.035 101.595 108.815 ;
        RECT 101.615 108.120 102.045 108.905 ;
        RECT 102.525 108.035 106.195 108.845 ;
        RECT 106.205 108.035 107.575 108.815 ;
        RECT 107.585 108.035 108.955 108.845 ;
        RECT 108.975 108.035 110.325 108.945 ;
        RECT 110.345 108.035 111.715 108.815 ;
        RECT 111.725 108.035 113.095 108.815 ;
        RECT 113.105 108.035 114.475 108.845 ;
        RECT 114.495 108.035 115.845 108.945 ;
        RECT 120.375 108.715 121.305 108.935 ;
        RECT 124.025 108.715 126.235 108.945 ;
        RECT 115.865 108.035 126.235 108.715 ;
        RECT 126.445 108.035 127.815 108.845 ;
        RECT 14.805 107.825 14.975 108.035 ;
        RECT 16.645 107.880 16.805 107.990 ;
        RECT 20.325 107.845 20.495 108.035 ;
        RECT 21.705 107.845 21.875 108.035 ;
        RECT 22.625 107.880 22.785 107.990 ;
        RECT 24.005 107.845 24.175 108.035 ;
        RECT 26.305 107.825 26.475 108.015 ;
        RECT 27.225 107.845 27.395 108.035 ;
        RECT 28.605 107.845 28.775 108.035 ;
        RECT 30.445 107.845 30.615 108.035 ;
        RECT 31.825 107.845 31.995 108.035 ;
        RECT 33.205 107.845 33.375 108.035 ;
        RECT 34.125 107.880 34.285 107.990 ;
        RECT 35.505 107.845 35.675 108.035 ;
        RECT 36.020 107.875 36.140 107.985 ;
        RECT 36.885 107.825 37.055 108.015 ;
        RECT 38.725 107.825 38.895 108.035 ;
        RECT 39.240 107.875 39.360 107.985 ;
        RECT 40.565 107.825 40.735 108.015 ;
        RECT 41.945 107.825 42.115 108.015 ;
        RECT 43.325 107.825 43.495 108.015 ;
        RECT 43.840 107.875 43.960 107.985 ;
        RECT 44.245 107.845 44.415 108.035 ;
        RECT 45.165 107.825 45.335 108.015 ;
        RECT 45.625 107.825 45.795 108.015 ;
        RECT 49.765 107.845 49.935 108.035 ;
        RECT 50.740 107.875 50.860 107.985 ;
        RECT 51.145 107.845 51.315 108.035 ;
        RECT 52.985 107.880 53.145 107.990 ;
        RECT 56.665 107.845 56.835 108.035 ;
        RECT 57.125 107.825 57.295 108.035 ;
        RECT 58.505 107.825 58.675 108.015 ;
        RECT 59.425 107.845 59.595 108.035 ;
        RECT 59.890 108.015 60.060 108.035 ;
        RECT 59.885 107.845 60.060 108.015 ;
        RECT 59.885 107.825 60.055 107.845 ;
        RECT 60.345 107.825 60.515 108.015 ;
        RECT 61.725 107.825 61.895 108.015 ;
        RECT 62.700 107.875 62.820 107.985 ;
        RECT 64.485 107.845 64.655 108.035 ;
        RECT 64.945 107.845 65.115 108.035 ;
        RECT 66.380 107.875 66.500 107.985 ;
        RECT 68.165 107.845 68.335 108.035 ;
        RECT 68.625 107.845 68.795 108.035 ;
        RECT 70.060 107.875 70.180 107.985 ;
        RECT 73.685 107.825 73.855 108.015 ;
        RECT 74.605 107.870 74.765 107.980 ;
        RECT 75.065 107.825 75.235 108.015 ;
        RECT 75.525 107.845 75.695 108.035 ;
        RECT 77.365 107.845 77.535 108.035 ;
        RECT 78.745 107.845 78.915 108.035 ;
        RECT 79.665 107.880 79.825 107.990 ;
        RECT 80.130 107.845 80.300 108.035 ;
        RECT 82.885 107.845 83.055 108.035 ;
        RECT 84.320 107.875 84.440 107.985 ;
        RECT 86.565 107.825 86.735 108.015 ;
        RECT 87.025 107.985 87.195 108.035 ;
        RECT 87.025 107.875 87.200 107.985 ;
        RECT 87.025 107.845 87.195 107.875 ;
        RECT 87.485 107.825 87.655 108.035 ;
        RECT 92.085 107.845 92.255 108.035 ;
        RECT 92.545 107.845 92.715 108.035 ;
        RECT 93.925 107.845 94.095 108.035 ;
        RECT 96.225 107.845 96.395 108.035 ;
        RECT 99.445 107.825 99.615 108.015 ;
        RECT 99.905 107.845 100.075 108.035 ;
        RECT 100.825 107.825 100.995 108.015 ;
        RECT 101.285 107.845 101.455 108.035 ;
        RECT 102.205 107.985 102.375 108.015 ;
        RECT 102.205 107.875 102.380 107.985 ;
        RECT 102.205 107.825 102.375 107.875 ;
        RECT 102.665 107.825 102.835 108.015 ;
        RECT 105.885 107.845 106.055 108.035 ;
        RECT 106.345 107.845 106.515 108.035 ;
        RECT 108.645 107.845 108.815 108.035 ;
        RECT 110.025 107.845 110.195 108.035 ;
        RECT 110.485 107.845 110.655 108.035 ;
        RECT 111.865 107.845 112.035 108.035 ;
        RECT 114.165 107.825 114.335 108.035 ;
        RECT 114.625 107.845 114.795 108.035 ;
        RECT 115.545 107.870 115.705 107.980 ;
        RECT 116.005 107.825 116.175 108.035 ;
        RECT 127.505 107.825 127.675 108.035 ;
        RECT 14.665 107.015 16.035 107.825 ;
        RECT 16.245 107.145 26.615 107.825 ;
        RECT 26.825 107.145 37.195 107.825 ;
        RECT 16.245 106.915 18.455 107.145 ;
        RECT 21.175 106.925 22.105 107.145 ;
        RECT 26.825 106.915 29.035 107.145 ;
        RECT 31.755 106.925 32.685 107.145 ;
        RECT 37.215 106.955 37.645 107.740 ;
        RECT 37.665 107.045 39.035 107.825 ;
        RECT 39.515 106.915 40.865 107.825 ;
        RECT 40.885 107.015 42.255 107.825 ;
        RECT 42.265 107.045 43.635 107.825 ;
        RECT 44.115 106.915 45.465 107.825 ;
        RECT 45.485 107.045 46.855 107.825 ;
        RECT 47.065 107.145 57.435 107.825 ;
        RECT 47.065 106.915 49.275 107.145 ;
        RECT 51.995 106.925 52.925 107.145 ;
        RECT 57.455 106.915 58.805 107.825 ;
        RECT 58.825 107.015 60.195 107.825 ;
        RECT 60.215 106.915 61.565 107.825 ;
        RECT 61.585 107.045 62.955 107.825 ;
        RECT 62.975 106.955 63.405 107.740 ;
        RECT 63.625 107.145 73.995 107.825 ;
        RECT 63.625 106.915 65.835 107.145 ;
        RECT 68.555 106.925 69.485 107.145 ;
        RECT 74.925 107.045 76.295 107.825 ;
        RECT 76.505 107.145 86.875 107.825 ;
        RECT 76.505 106.915 78.715 107.145 ;
        RECT 81.435 106.925 82.365 107.145 ;
        RECT 87.345 107.045 88.715 107.825 ;
        RECT 88.735 106.955 89.165 107.740 ;
        RECT 89.385 107.145 99.755 107.825 ;
        RECT 89.385 106.915 91.595 107.145 ;
        RECT 94.315 106.925 95.245 107.145 ;
        RECT 99.775 106.915 101.125 107.825 ;
        RECT 101.145 107.015 102.515 107.825 ;
        RECT 102.535 106.915 103.885 107.825 ;
        RECT 104.105 107.145 114.475 107.825 ;
        RECT 104.105 106.915 106.315 107.145 ;
        RECT 109.035 106.925 109.965 107.145 ;
        RECT 114.495 106.955 114.925 107.740 ;
        RECT 115.865 107.145 126.235 107.825 ;
        RECT 120.375 106.925 121.305 107.145 ;
        RECT 124.025 106.915 126.235 107.145 ;
        RECT 126.445 107.015 127.815 107.825 ;
      LAYER nwell ;
        RECT 14.470 103.795 128.010 106.625 ;
      LAYER pwell ;
        RECT 14.665 102.595 16.035 103.405 ;
        RECT 16.045 102.595 18.795 103.405 ;
        RECT 18.805 102.595 24.315 103.405 ;
        RECT 24.335 102.680 24.765 103.465 ;
        RECT 24.785 102.595 27.535 103.405 ;
        RECT 27.555 102.595 28.905 103.505 ;
        RECT 33.435 103.275 34.365 103.495 ;
        RECT 37.085 103.275 39.295 103.505 ;
        RECT 28.925 102.595 39.295 103.275 ;
        RECT 39.705 103.275 41.915 103.505 ;
        RECT 44.635 103.275 45.565 103.495 ;
        RECT 39.705 102.595 50.075 103.275 ;
        RECT 50.095 102.680 50.525 103.465 ;
        RECT 51.475 102.595 52.825 103.505 ;
        RECT 53.045 103.275 55.255 103.505 ;
        RECT 57.975 103.275 58.905 103.495 ;
        RECT 63.625 103.275 65.835 103.505 ;
        RECT 68.555 103.275 69.485 103.495 ;
        RECT 53.045 102.595 63.415 103.275 ;
        RECT 63.625 102.595 73.995 103.275 ;
        RECT 74.005 102.595 75.835 103.405 ;
        RECT 75.855 102.680 76.285 103.465 ;
        RECT 76.505 103.275 78.715 103.505 ;
        RECT 81.435 103.275 82.365 103.495 ;
        RECT 87.085 103.275 89.295 103.505 ;
        RECT 92.015 103.275 92.945 103.495 ;
        RECT 76.505 102.595 86.875 103.275 ;
        RECT 87.085 102.595 97.455 103.275 ;
        RECT 97.925 102.595 101.595 103.405 ;
        RECT 101.615 102.680 102.045 103.465 ;
        RECT 102.265 103.275 104.475 103.505 ;
        RECT 107.195 103.275 108.125 103.495 ;
        RECT 117.155 103.275 118.085 103.495 ;
        RECT 120.805 103.275 123.015 103.505 ;
        RECT 102.265 102.595 112.635 103.275 ;
        RECT 112.645 102.595 123.015 103.275 ;
        RECT 123.225 102.595 125.055 103.405 ;
        RECT 125.065 102.595 126.435 103.375 ;
        RECT 126.445 102.595 127.815 103.405 ;
        RECT 14.805 102.385 14.975 102.595 ;
        RECT 18.485 102.385 18.655 102.595 ;
        RECT 24.005 102.385 24.175 102.595 ;
        RECT 27.225 102.405 27.395 102.595 ;
        RECT 27.685 102.405 27.855 102.595 ;
        RECT 29.065 102.405 29.235 102.595 ;
        RECT 35.045 102.385 35.215 102.575 ;
        RECT 36.885 102.385 37.055 102.575 ;
        RECT 38.725 102.385 38.895 102.575 ;
        RECT 44.245 102.385 44.415 102.575 ;
        RECT 49.765 102.385 49.935 102.595 ;
        RECT 51.145 102.440 51.305 102.550 ;
        RECT 51.605 102.385 51.775 102.575 ;
        RECT 52.525 102.405 52.695 102.595 ;
        RECT 57.125 102.385 57.295 102.575 ;
        RECT 62.645 102.385 62.815 102.575 ;
        RECT 63.105 102.405 63.275 102.595 ;
        RECT 64.485 102.385 64.655 102.575 ;
        RECT 70.005 102.385 70.175 102.575 ;
        RECT 73.685 102.405 73.855 102.595 ;
        RECT 75.525 102.385 75.695 102.595 ;
        RECT 77.365 102.385 77.535 102.575 ;
        RECT 82.885 102.385 83.055 102.575 ;
        RECT 86.565 102.405 86.735 102.595 ;
        RECT 88.405 102.385 88.575 102.575 ;
        RECT 90.705 102.385 90.875 102.575 ;
        RECT 97.145 102.405 97.315 102.595 ;
        RECT 97.660 102.435 97.780 102.545 ;
        RECT 101.285 102.385 101.455 102.595 ;
        RECT 103.125 102.385 103.295 102.575 ;
        RECT 108.645 102.385 108.815 102.575 ;
        RECT 112.325 102.405 112.495 102.595 ;
        RECT 112.785 102.405 112.955 102.595 ;
        RECT 114.165 102.385 114.335 102.575 ;
        RECT 115.545 102.430 115.705 102.540 ;
        RECT 119.225 102.385 119.395 102.575 ;
        RECT 119.685 102.385 119.855 102.575 ;
        RECT 124.745 102.405 124.915 102.595 ;
        RECT 126.115 102.575 126.285 102.595 ;
        RECT 126.115 102.405 126.295 102.575 ;
        RECT 126.125 102.385 126.295 102.405 ;
        RECT 127.505 102.385 127.675 102.595 ;
        RECT 14.665 101.575 16.035 102.385 ;
        RECT 16.045 101.575 18.795 102.385 ;
        RECT 18.805 101.575 24.315 102.385 ;
        RECT 24.335 101.515 24.765 102.300 ;
        RECT 24.985 101.705 35.355 102.385 ;
        RECT 24.985 101.475 27.195 101.705 ;
        RECT 29.915 101.485 30.845 101.705 ;
        RECT 35.365 101.575 37.195 102.385 ;
        RECT 37.215 101.515 37.645 102.300 ;
        RECT 37.665 101.575 39.035 102.385 ;
        RECT 39.045 101.575 44.555 102.385 ;
        RECT 44.565 101.575 50.075 102.385 ;
        RECT 50.095 101.515 50.525 102.300 ;
        RECT 50.545 101.575 51.915 102.385 ;
        RECT 51.925 101.575 57.435 102.385 ;
        RECT 57.445 101.575 62.955 102.385 ;
        RECT 62.975 101.515 63.405 102.300 ;
        RECT 63.425 101.575 64.795 102.385 ;
        RECT 64.805 101.575 70.315 102.385 ;
        RECT 70.325 101.575 75.835 102.385 ;
        RECT 75.855 101.515 76.285 102.300 ;
        RECT 76.305 101.575 77.675 102.385 ;
        RECT 77.685 101.575 83.195 102.385 ;
        RECT 83.205 101.575 88.715 102.385 ;
        RECT 88.735 101.515 89.165 102.300 ;
        RECT 89.185 101.575 91.015 102.385 ;
        RECT 91.225 101.705 101.595 102.385 ;
        RECT 91.225 101.475 93.435 101.705 ;
        RECT 96.155 101.485 97.085 101.705 ;
        RECT 101.615 101.515 102.045 102.300 ;
        RECT 102.065 101.575 103.435 102.385 ;
        RECT 103.445 101.575 108.955 102.385 ;
        RECT 108.965 101.575 114.475 102.385 ;
        RECT 114.495 101.515 114.925 102.300 ;
        RECT 115.865 101.575 119.535 102.385 ;
        RECT 119.555 101.475 120.905 102.385 ;
        RECT 120.925 101.575 126.435 102.385 ;
        RECT 126.445 101.575 127.815 102.385 ;
      LAYER nwell ;
        RECT 14.470 99.580 128.010 101.185 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 14.660 211.205 127.820 211.375 ;
        RECT 14.745 210.455 15.955 211.205 ;
        RECT 14.745 209.915 15.265 210.455 ;
        RECT 16.125 210.435 18.715 211.205 ;
        RECT 18.890 210.660 24.235 211.205 ;
        RECT 15.435 209.745 15.955 210.285 ;
        RECT 14.745 208.655 15.955 209.745 ;
        RECT 16.125 209.745 17.335 210.265 ;
        RECT 17.505 209.915 18.715 210.435 ;
        RECT 16.125 208.655 18.715 209.745 ;
        RECT 20.480 209.090 20.830 210.340 ;
        RECT 22.310 209.830 22.650 210.660 ;
        RECT 24.405 210.480 24.695 211.205 ;
        RECT 24.865 210.455 26.075 211.205 ;
        RECT 26.250 210.660 31.595 211.205 ;
        RECT 31.770 210.660 37.115 211.205 ;
        RECT 18.890 208.655 24.235 209.090 ;
        RECT 24.405 208.655 24.695 209.820 ;
        RECT 24.865 209.745 25.385 210.285 ;
        RECT 25.555 209.915 26.075 210.455 ;
        RECT 24.865 208.655 26.075 209.745 ;
        RECT 27.840 209.090 28.190 210.340 ;
        RECT 29.670 209.830 30.010 210.660 ;
        RECT 33.360 209.090 33.710 210.340 ;
        RECT 35.190 209.830 35.530 210.660 ;
        RECT 37.285 210.480 37.575 211.205 ;
        RECT 37.745 210.455 38.955 211.205 ;
        RECT 39.130 210.660 44.475 211.205 ;
        RECT 44.650 210.660 49.995 211.205 ;
        RECT 26.250 208.655 31.595 209.090 ;
        RECT 31.770 208.655 37.115 209.090 ;
        RECT 37.285 208.655 37.575 209.820 ;
        RECT 37.745 209.745 38.265 210.285 ;
        RECT 38.435 209.915 38.955 210.455 ;
        RECT 37.745 208.655 38.955 209.745 ;
        RECT 40.720 209.090 41.070 210.340 ;
        RECT 42.550 209.830 42.890 210.660 ;
        RECT 46.240 209.090 46.590 210.340 ;
        RECT 48.070 209.830 48.410 210.660 ;
        RECT 50.165 210.480 50.455 211.205 ;
        RECT 50.625 210.455 51.835 211.205 ;
        RECT 52.010 210.660 57.355 211.205 ;
        RECT 57.530 210.660 62.875 211.205 ;
        RECT 39.130 208.655 44.475 209.090 ;
        RECT 44.650 208.655 49.995 209.090 ;
        RECT 50.165 208.655 50.455 209.820 ;
        RECT 50.625 209.745 51.145 210.285 ;
        RECT 51.315 209.915 51.835 210.455 ;
        RECT 50.625 208.655 51.835 209.745 ;
        RECT 53.600 209.090 53.950 210.340 ;
        RECT 55.430 209.830 55.770 210.660 ;
        RECT 59.120 209.090 59.470 210.340 ;
        RECT 60.950 209.830 61.290 210.660 ;
        RECT 63.045 210.480 63.335 211.205 ;
        RECT 63.505 210.455 64.715 211.205 ;
        RECT 64.890 210.660 70.235 211.205 ;
        RECT 70.410 210.660 75.755 211.205 ;
        RECT 52.010 208.655 57.355 209.090 ;
        RECT 57.530 208.655 62.875 209.090 ;
        RECT 63.045 208.655 63.335 209.820 ;
        RECT 63.505 209.745 64.025 210.285 ;
        RECT 64.195 209.915 64.715 210.455 ;
        RECT 63.505 208.655 64.715 209.745 ;
        RECT 66.480 209.090 66.830 210.340 ;
        RECT 68.310 209.830 68.650 210.660 ;
        RECT 72.000 209.090 72.350 210.340 ;
        RECT 73.830 209.830 74.170 210.660 ;
        RECT 75.925 210.480 76.215 211.205 ;
        RECT 76.385 210.455 77.595 211.205 ;
        RECT 77.770 210.660 83.115 211.205 ;
        RECT 83.290 210.660 88.635 211.205 ;
        RECT 64.890 208.655 70.235 209.090 ;
        RECT 70.410 208.655 75.755 209.090 ;
        RECT 75.925 208.655 76.215 209.820 ;
        RECT 76.385 209.745 76.905 210.285 ;
        RECT 77.075 209.915 77.595 210.455 ;
        RECT 76.385 208.655 77.595 209.745 ;
        RECT 79.360 209.090 79.710 210.340 ;
        RECT 81.190 209.830 81.530 210.660 ;
        RECT 84.880 209.090 85.230 210.340 ;
        RECT 86.710 209.830 87.050 210.660 ;
        RECT 88.805 210.480 89.095 211.205 ;
        RECT 89.265 210.455 90.475 211.205 ;
        RECT 90.650 210.660 95.995 211.205 ;
        RECT 96.170 210.660 101.515 211.205 ;
        RECT 77.770 208.655 83.115 209.090 ;
        RECT 83.290 208.655 88.635 209.090 ;
        RECT 88.805 208.655 89.095 209.820 ;
        RECT 89.265 209.745 89.785 210.285 ;
        RECT 89.955 209.915 90.475 210.455 ;
        RECT 89.265 208.655 90.475 209.745 ;
        RECT 92.240 209.090 92.590 210.340 ;
        RECT 94.070 209.830 94.410 210.660 ;
        RECT 97.760 209.090 98.110 210.340 ;
        RECT 99.590 209.830 99.930 210.660 ;
        RECT 101.685 210.480 101.975 211.205 ;
        RECT 102.145 210.455 103.355 211.205 ;
        RECT 103.530 210.660 108.875 211.205 ;
        RECT 109.050 210.660 114.395 211.205 ;
        RECT 90.650 208.655 95.995 209.090 ;
        RECT 96.170 208.655 101.515 209.090 ;
        RECT 101.685 208.655 101.975 209.820 ;
        RECT 102.145 209.745 102.665 210.285 ;
        RECT 102.835 209.915 103.355 210.455 ;
        RECT 102.145 208.655 103.355 209.745 ;
        RECT 105.120 209.090 105.470 210.340 ;
        RECT 106.950 209.830 107.290 210.660 ;
        RECT 110.640 209.090 110.990 210.340 ;
        RECT 112.470 209.830 112.810 210.660 ;
        RECT 114.565 210.480 114.855 211.205 ;
        RECT 115.490 210.660 120.835 211.205 ;
        RECT 121.010 210.660 126.355 211.205 ;
        RECT 103.530 208.655 108.875 209.090 ;
        RECT 109.050 208.655 114.395 209.090 ;
        RECT 114.565 208.655 114.855 209.820 ;
        RECT 117.080 209.090 117.430 210.340 ;
        RECT 118.910 209.830 119.250 210.660 ;
        RECT 122.600 209.090 122.950 210.340 ;
        RECT 124.430 209.830 124.770 210.660 ;
        RECT 126.525 210.455 127.735 211.205 ;
        RECT 126.525 209.745 127.045 210.285 ;
        RECT 127.215 209.915 127.735 210.455 ;
        RECT 115.490 208.655 120.835 209.090 ;
        RECT 121.010 208.655 126.355 209.090 ;
        RECT 126.525 208.655 127.735 209.745 ;
        RECT 14.660 208.485 127.820 208.655 ;
        RECT 14.745 207.395 15.955 208.485 ;
        RECT 14.745 206.685 15.265 207.225 ;
        RECT 15.435 206.855 15.955 207.395 ;
        RECT 16.125 207.395 18.715 208.485 ;
        RECT 18.890 208.050 24.235 208.485 ;
        RECT 16.125 206.875 17.335 207.395 ;
        RECT 17.505 206.705 18.715 207.225 ;
        RECT 20.480 206.800 20.830 208.050 ;
        RECT 24.405 207.320 24.695 208.485 ;
        RECT 25.325 207.395 27.915 208.485 ;
        RECT 28.090 208.050 33.435 208.485 ;
        RECT 33.610 208.050 38.955 208.485 ;
        RECT 39.130 208.050 44.475 208.485 ;
        RECT 44.650 208.050 49.995 208.485 ;
        RECT 14.745 205.935 15.955 206.685 ;
        RECT 16.125 205.935 18.715 206.705 ;
        RECT 22.310 206.480 22.650 207.310 ;
        RECT 25.325 206.875 26.535 207.395 ;
        RECT 26.705 206.705 27.915 207.225 ;
        RECT 29.680 206.800 30.030 208.050 ;
        RECT 18.890 205.935 24.235 206.480 ;
        RECT 24.405 205.935 24.695 206.660 ;
        RECT 25.325 205.935 27.915 206.705 ;
        RECT 31.510 206.480 31.850 207.310 ;
        RECT 35.200 206.800 35.550 208.050 ;
        RECT 37.030 206.480 37.370 207.310 ;
        RECT 40.720 206.800 41.070 208.050 ;
        RECT 42.550 206.480 42.890 207.310 ;
        RECT 46.240 206.800 46.590 208.050 ;
        RECT 50.165 207.320 50.455 208.485 ;
        RECT 50.630 208.050 55.975 208.485 ;
        RECT 56.150 208.050 61.495 208.485 ;
        RECT 61.670 208.050 67.015 208.485 ;
        RECT 67.190 208.050 72.535 208.485 ;
        RECT 48.070 206.480 48.410 207.310 ;
        RECT 52.220 206.800 52.570 208.050 ;
        RECT 28.090 205.935 33.435 206.480 ;
        RECT 33.610 205.935 38.955 206.480 ;
        RECT 39.130 205.935 44.475 206.480 ;
        RECT 44.650 205.935 49.995 206.480 ;
        RECT 50.165 205.935 50.455 206.660 ;
        RECT 54.050 206.480 54.390 207.310 ;
        RECT 57.740 206.800 58.090 208.050 ;
        RECT 59.570 206.480 59.910 207.310 ;
        RECT 63.260 206.800 63.610 208.050 ;
        RECT 65.090 206.480 65.430 207.310 ;
        RECT 68.780 206.800 69.130 208.050 ;
        RECT 72.745 207.345 72.975 208.485 ;
        RECT 73.145 207.335 73.475 208.315 ;
        RECT 73.645 207.345 73.855 208.485 ;
        RECT 74.175 207.555 74.345 208.315 ;
        RECT 74.560 207.725 74.890 208.485 ;
        RECT 74.175 207.385 74.890 207.555 ;
        RECT 75.060 207.410 75.315 208.315 ;
        RECT 70.610 206.480 70.950 207.310 ;
        RECT 72.725 206.925 73.055 207.175 ;
        RECT 50.630 205.935 55.975 206.480 ;
        RECT 56.150 205.935 61.495 206.480 ;
        RECT 61.670 205.935 67.015 206.480 ;
        RECT 67.190 205.935 72.535 206.480 ;
        RECT 72.745 205.935 72.975 206.755 ;
        RECT 73.225 206.735 73.475 207.335 ;
        RECT 74.085 206.835 74.440 207.205 ;
        RECT 74.720 207.175 74.890 207.385 ;
        RECT 74.720 206.845 74.975 207.175 ;
        RECT 73.145 206.105 73.475 206.735 ;
        RECT 73.645 205.935 73.855 206.755 ;
        RECT 74.720 206.655 74.890 206.845 ;
        RECT 75.145 206.680 75.315 207.410 ;
        RECT 75.490 207.335 75.750 208.485 ;
        RECT 75.925 207.320 76.215 208.485 ;
        RECT 77.325 207.975 77.625 208.485 ;
        RECT 77.795 207.975 78.175 208.145 ;
        RECT 78.755 207.975 79.385 208.485 ;
        RECT 77.795 207.805 77.965 207.975 ;
        RECT 79.555 207.805 79.885 208.315 ;
        RECT 80.055 207.975 80.355 208.485 ;
        RECT 77.305 207.605 77.965 207.805 ;
        RECT 78.135 207.635 80.355 207.805 ;
        RECT 74.175 206.485 74.890 206.655 ;
        RECT 74.175 206.105 74.345 206.485 ;
        RECT 74.560 205.935 74.890 206.315 ;
        RECT 75.060 206.105 75.315 206.680 ;
        RECT 75.490 205.935 75.750 206.775 ;
        RECT 77.305 206.675 77.475 207.605 ;
        RECT 78.135 207.435 78.305 207.635 ;
        RECT 77.645 207.265 78.305 207.435 ;
        RECT 78.475 207.295 80.015 207.465 ;
        RECT 77.645 206.845 77.815 207.265 ;
        RECT 78.475 207.095 78.645 207.295 ;
        RECT 78.045 206.925 78.645 207.095 ;
        RECT 78.815 206.925 79.510 207.125 ;
        RECT 79.770 206.845 80.015 207.295 ;
        RECT 78.135 206.675 79.045 206.755 ;
        RECT 75.925 205.935 76.215 206.660 ;
        RECT 77.305 206.195 77.625 206.675 ;
        RECT 77.795 206.585 79.045 206.675 ;
        RECT 77.795 206.505 78.305 206.585 ;
        RECT 77.795 206.105 78.025 206.505 ;
        RECT 78.195 205.935 78.545 206.325 ;
        RECT 78.715 206.105 79.045 206.585 ;
        RECT 79.215 205.935 79.385 206.755 ;
        RECT 80.185 206.675 80.355 207.635 ;
        RECT 81.445 207.395 84.955 208.485 ;
        RECT 85.130 208.050 90.475 208.485 ;
        RECT 90.650 208.050 95.995 208.485 ;
        RECT 96.170 208.050 101.515 208.485 ;
        RECT 81.445 206.875 83.135 207.395 ;
        RECT 83.305 206.705 84.955 207.225 ;
        RECT 86.720 206.800 87.070 208.050 ;
        RECT 79.890 206.130 80.355 206.675 ;
        RECT 81.445 205.935 84.955 206.705 ;
        RECT 88.550 206.480 88.890 207.310 ;
        RECT 92.240 206.800 92.590 208.050 ;
        RECT 94.070 206.480 94.410 207.310 ;
        RECT 97.760 206.800 98.110 208.050 ;
        RECT 101.685 207.320 101.975 208.485 ;
        RECT 102.605 207.395 104.275 208.485 ;
        RECT 104.450 208.050 109.795 208.485 ;
        RECT 109.970 208.050 115.315 208.485 ;
        RECT 115.490 208.050 120.835 208.485 ;
        RECT 121.010 208.050 126.355 208.485 ;
        RECT 99.590 206.480 99.930 207.310 ;
        RECT 102.605 206.875 103.355 207.395 ;
        RECT 103.525 206.705 104.275 207.225 ;
        RECT 106.040 206.800 106.390 208.050 ;
        RECT 85.130 205.935 90.475 206.480 ;
        RECT 90.650 205.935 95.995 206.480 ;
        RECT 96.170 205.935 101.515 206.480 ;
        RECT 101.685 205.935 101.975 206.660 ;
        RECT 102.605 205.935 104.275 206.705 ;
        RECT 107.870 206.480 108.210 207.310 ;
        RECT 111.560 206.800 111.910 208.050 ;
        RECT 113.390 206.480 113.730 207.310 ;
        RECT 117.080 206.800 117.430 208.050 ;
        RECT 118.910 206.480 119.250 207.310 ;
        RECT 122.600 206.800 122.950 208.050 ;
        RECT 126.525 207.395 127.735 208.485 ;
        RECT 124.430 206.480 124.770 207.310 ;
        RECT 126.525 206.855 127.045 207.395 ;
        RECT 127.215 206.685 127.735 207.225 ;
        RECT 104.450 205.935 109.795 206.480 ;
        RECT 109.970 205.935 115.315 206.480 ;
        RECT 115.490 205.935 120.835 206.480 ;
        RECT 121.010 205.935 126.355 206.480 ;
        RECT 126.525 205.935 127.735 206.685 ;
        RECT 14.660 205.765 127.820 205.935 ;
        RECT 14.745 205.015 15.955 205.765 ;
        RECT 14.745 204.475 15.265 205.015 ;
        RECT 17.045 204.995 20.555 205.765 ;
        RECT 20.730 205.220 26.075 205.765 ;
        RECT 26.250 205.220 31.595 205.765 ;
        RECT 31.770 205.220 37.115 205.765 ;
        RECT 15.435 204.305 15.955 204.845 ;
        RECT 14.745 203.215 15.955 204.305 ;
        RECT 17.045 204.305 18.735 204.825 ;
        RECT 18.905 204.475 20.555 204.995 ;
        RECT 17.045 203.215 20.555 204.305 ;
        RECT 22.320 203.650 22.670 204.900 ;
        RECT 24.150 204.390 24.490 205.220 ;
        RECT 27.840 203.650 28.190 204.900 ;
        RECT 29.670 204.390 30.010 205.220 ;
        RECT 33.360 203.650 33.710 204.900 ;
        RECT 35.190 204.390 35.530 205.220 ;
        RECT 37.285 205.040 37.575 205.765 ;
        RECT 38.205 204.995 40.795 205.765 ;
        RECT 40.970 205.220 46.315 205.765 ;
        RECT 46.490 205.220 51.835 205.765 ;
        RECT 52.010 205.220 57.355 205.765 ;
        RECT 57.530 205.220 62.875 205.765 ;
        RECT 20.730 203.215 26.075 203.650 ;
        RECT 26.250 203.215 31.595 203.650 ;
        RECT 31.770 203.215 37.115 203.650 ;
        RECT 37.285 203.215 37.575 204.380 ;
        RECT 38.205 204.305 39.415 204.825 ;
        RECT 39.585 204.475 40.795 204.995 ;
        RECT 38.205 203.215 40.795 204.305 ;
        RECT 42.560 203.650 42.910 204.900 ;
        RECT 44.390 204.390 44.730 205.220 ;
        RECT 48.080 203.650 48.430 204.900 ;
        RECT 49.910 204.390 50.250 205.220 ;
        RECT 53.600 203.650 53.950 204.900 ;
        RECT 55.430 204.390 55.770 205.220 ;
        RECT 59.120 203.650 59.470 204.900 ;
        RECT 60.950 204.390 61.290 205.220 ;
        RECT 63.045 205.040 63.335 205.765 ;
        RECT 63.505 205.015 64.715 205.765 ;
        RECT 40.970 203.215 46.315 203.650 ;
        RECT 46.490 203.215 51.835 203.650 ;
        RECT 52.010 203.215 57.355 203.650 ;
        RECT 57.530 203.215 62.875 203.650 ;
        RECT 63.045 203.215 63.335 204.380 ;
        RECT 63.505 204.305 64.025 204.845 ;
        RECT 64.195 204.475 64.715 205.015 ;
        RECT 64.945 204.945 65.155 205.765 ;
        RECT 65.325 204.965 65.655 205.595 ;
        RECT 65.325 204.365 65.575 204.965 ;
        RECT 65.825 204.945 66.055 205.765 ;
        RECT 67.225 204.945 67.455 205.765 ;
        RECT 67.625 204.965 67.955 205.595 ;
        RECT 65.745 204.525 66.075 204.775 ;
        RECT 67.205 204.525 67.535 204.775 ;
        RECT 67.705 204.365 67.955 204.965 ;
        RECT 68.125 204.945 68.335 205.765 ;
        RECT 68.570 205.055 68.825 205.585 ;
        RECT 68.995 205.305 69.300 205.765 ;
        RECT 69.545 205.385 70.615 205.555 ;
        RECT 63.505 203.215 64.715 204.305 ;
        RECT 64.945 203.215 65.155 204.355 ;
        RECT 65.325 203.385 65.655 204.365 ;
        RECT 65.825 203.215 66.055 204.355 ;
        RECT 67.225 203.215 67.455 204.355 ;
        RECT 67.625 203.385 67.955 204.365 ;
        RECT 68.570 204.405 68.780 205.055 ;
        RECT 69.545 205.030 69.865 205.385 ;
        RECT 69.540 204.855 69.865 205.030 ;
        RECT 68.950 204.555 69.865 204.855 ;
        RECT 70.035 204.815 70.275 205.215 ;
        RECT 70.445 205.155 70.615 205.385 ;
        RECT 70.785 205.325 70.975 205.765 ;
        RECT 71.145 205.315 72.095 205.595 ;
        RECT 72.315 205.405 72.665 205.575 ;
        RECT 70.445 204.985 70.975 205.155 ;
        RECT 68.950 204.525 69.690 204.555 ;
        RECT 68.125 203.215 68.335 204.355 ;
        RECT 68.570 203.525 68.825 204.405 ;
        RECT 68.995 203.215 69.300 204.355 ;
        RECT 69.520 203.935 69.690 204.525 ;
        RECT 70.035 204.445 70.575 204.815 ;
        RECT 70.755 204.705 70.975 204.985 ;
        RECT 71.145 204.535 71.315 205.315 ;
        RECT 70.910 204.365 71.315 204.535 ;
        RECT 71.485 204.525 71.835 205.145 ;
        RECT 70.910 204.275 71.080 204.365 ;
        RECT 72.005 204.355 72.215 205.145 ;
        RECT 69.860 204.105 71.080 204.275 ;
        RECT 71.540 204.195 72.215 204.355 ;
        RECT 69.520 203.765 70.320 203.935 ;
        RECT 69.640 203.215 69.970 203.595 ;
        RECT 70.150 203.475 70.320 203.765 ;
        RECT 70.910 203.725 71.080 204.105 ;
        RECT 71.250 204.185 72.215 204.195 ;
        RECT 72.405 205.015 72.665 205.405 ;
        RECT 72.875 205.305 73.205 205.765 ;
        RECT 74.080 205.375 74.935 205.545 ;
        RECT 75.140 205.375 75.635 205.545 ;
        RECT 75.805 205.405 76.135 205.765 ;
        RECT 72.405 204.325 72.575 205.015 ;
        RECT 72.745 204.665 72.915 204.845 ;
        RECT 73.085 204.835 73.875 205.085 ;
        RECT 74.080 204.665 74.250 205.375 ;
        RECT 74.420 204.865 74.775 205.085 ;
        RECT 72.745 204.495 74.435 204.665 ;
        RECT 71.250 203.895 71.710 204.185 ;
        RECT 72.405 204.155 73.905 204.325 ;
        RECT 72.405 204.015 72.575 204.155 ;
        RECT 72.015 203.845 72.575 204.015 ;
        RECT 70.490 203.215 70.740 203.675 ;
        RECT 70.910 203.385 71.780 203.725 ;
        RECT 72.015 203.385 72.185 203.845 ;
        RECT 73.020 203.815 74.095 203.985 ;
        RECT 72.355 203.215 72.725 203.675 ;
        RECT 73.020 203.475 73.190 203.815 ;
        RECT 73.360 203.215 73.690 203.645 ;
        RECT 73.925 203.475 74.095 203.815 ;
        RECT 74.265 203.715 74.435 204.495 ;
        RECT 74.605 204.275 74.775 204.865 ;
        RECT 74.945 204.465 75.295 205.085 ;
        RECT 74.605 203.885 75.070 204.275 ;
        RECT 75.465 204.015 75.635 205.375 ;
        RECT 75.805 204.185 76.265 205.235 ;
        RECT 75.240 203.845 75.635 204.015 ;
        RECT 75.240 203.715 75.410 203.845 ;
        RECT 74.265 203.385 74.945 203.715 ;
        RECT 75.160 203.385 75.410 203.715 ;
        RECT 75.580 203.215 75.830 203.675 ;
        RECT 76.000 203.400 76.325 204.185 ;
        RECT 76.495 203.385 76.665 205.505 ;
        RECT 76.835 205.385 77.165 205.765 ;
        RECT 77.335 205.215 77.590 205.505 ;
        RECT 76.840 205.045 77.590 205.215 ;
        RECT 77.770 205.055 78.025 205.585 ;
        RECT 78.195 205.305 78.500 205.765 ;
        RECT 78.745 205.385 79.815 205.555 ;
        RECT 76.840 204.055 77.070 205.045 ;
        RECT 77.240 204.225 77.590 204.875 ;
        RECT 77.770 204.405 77.980 205.055 ;
        RECT 78.745 205.030 79.065 205.385 ;
        RECT 78.740 204.855 79.065 205.030 ;
        RECT 78.150 204.555 79.065 204.855 ;
        RECT 79.235 204.815 79.475 205.215 ;
        RECT 79.645 205.155 79.815 205.385 ;
        RECT 79.985 205.325 80.175 205.765 ;
        RECT 80.345 205.315 81.295 205.595 ;
        RECT 81.515 205.405 81.865 205.575 ;
        RECT 79.645 204.985 80.175 205.155 ;
        RECT 78.150 204.525 78.890 204.555 ;
        RECT 76.840 203.885 77.590 204.055 ;
        RECT 76.835 203.215 77.165 203.715 ;
        RECT 77.335 203.385 77.590 203.885 ;
        RECT 77.770 203.525 78.025 204.405 ;
        RECT 78.195 203.215 78.500 204.355 ;
        RECT 78.720 203.935 78.890 204.525 ;
        RECT 79.235 204.445 79.775 204.815 ;
        RECT 79.955 204.705 80.175 204.985 ;
        RECT 80.345 204.535 80.515 205.315 ;
        RECT 80.110 204.365 80.515 204.535 ;
        RECT 80.685 204.525 81.035 205.145 ;
        RECT 80.110 204.275 80.280 204.365 ;
        RECT 81.205 204.355 81.415 205.145 ;
        RECT 79.060 204.105 80.280 204.275 ;
        RECT 80.740 204.195 81.415 204.355 ;
        RECT 78.720 203.765 79.520 203.935 ;
        RECT 78.840 203.215 79.170 203.595 ;
        RECT 79.350 203.475 79.520 203.765 ;
        RECT 80.110 203.725 80.280 204.105 ;
        RECT 80.450 204.185 81.415 204.195 ;
        RECT 81.605 205.015 81.865 205.405 ;
        RECT 82.075 205.305 82.405 205.765 ;
        RECT 83.280 205.375 84.135 205.545 ;
        RECT 84.340 205.375 84.835 205.545 ;
        RECT 85.005 205.405 85.335 205.765 ;
        RECT 81.605 204.325 81.775 205.015 ;
        RECT 81.945 204.665 82.115 204.845 ;
        RECT 82.285 204.835 83.075 205.085 ;
        RECT 83.280 204.665 83.450 205.375 ;
        RECT 83.620 204.865 83.975 205.085 ;
        RECT 81.945 204.495 83.635 204.665 ;
        RECT 80.450 203.895 80.910 204.185 ;
        RECT 81.605 204.155 83.105 204.325 ;
        RECT 81.605 204.015 81.775 204.155 ;
        RECT 81.215 203.845 81.775 204.015 ;
        RECT 79.690 203.215 79.940 203.675 ;
        RECT 80.110 203.385 80.980 203.725 ;
        RECT 81.215 203.385 81.385 203.845 ;
        RECT 82.220 203.815 83.295 203.985 ;
        RECT 81.555 203.215 81.925 203.675 ;
        RECT 82.220 203.475 82.390 203.815 ;
        RECT 82.560 203.215 82.890 203.645 ;
        RECT 83.125 203.475 83.295 203.815 ;
        RECT 83.465 203.715 83.635 204.495 ;
        RECT 83.805 204.275 83.975 204.865 ;
        RECT 84.145 204.465 84.495 205.085 ;
        RECT 83.805 203.885 84.270 204.275 ;
        RECT 84.665 204.015 84.835 205.375 ;
        RECT 85.005 204.185 85.465 205.235 ;
        RECT 84.440 203.845 84.835 204.015 ;
        RECT 84.440 203.715 84.610 203.845 ;
        RECT 83.465 203.385 84.145 203.715 ;
        RECT 84.360 203.385 84.610 203.715 ;
        RECT 84.780 203.215 85.030 203.675 ;
        RECT 85.200 203.400 85.525 204.185 ;
        RECT 85.695 203.385 85.865 205.505 ;
        RECT 86.035 205.385 86.365 205.765 ;
        RECT 86.535 205.215 86.790 205.505 ;
        RECT 86.040 205.045 86.790 205.215 ;
        RECT 86.040 204.055 86.270 205.045 ;
        RECT 86.965 204.995 88.635 205.765 ;
        RECT 88.805 205.040 89.095 205.765 ;
        RECT 89.725 204.995 92.315 205.765 ;
        RECT 92.490 205.220 97.835 205.765 ;
        RECT 98.010 205.220 103.355 205.765 ;
        RECT 103.530 205.220 108.875 205.765 ;
        RECT 109.050 205.220 114.395 205.765 ;
        RECT 86.440 204.225 86.790 204.875 ;
        RECT 86.965 204.305 87.715 204.825 ;
        RECT 87.885 204.475 88.635 204.995 ;
        RECT 86.040 203.885 86.790 204.055 ;
        RECT 86.035 203.215 86.365 203.715 ;
        RECT 86.535 203.385 86.790 203.885 ;
        RECT 86.965 203.215 88.635 204.305 ;
        RECT 88.805 203.215 89.095 204.380 ;
        RECT 89.725 204.305 90.935 204.825 ;
        RECT 91.105 204.475 92.315 204.995 ;
        RECT 89.725 203.215 92.315 204.305 ;
        RECT 94.080 203.650 94.430 204.900 ;
        RECT 95.910 204.390 96.250 205.220 ;
        RECT 99.600 203.650 99.950 204.900 ;
        RECT 101.430 204.390 101.770 205.220 ;
        RECT 105.120 203.650 105.470 204.900 ;
        RECT 106.950 204.390 107.290 205.220 ;
        RECT 110.640 203.650 110.990 204.900 ;
        RECT 112.470 204.390 112.810 205.220 ;
        RECT 114.565 205.040 114.855 205.765 ;
        RECT 115.490 205.220 120.835 205.765 ;
        RECT 121.010 205.220 126.355 205.765 ;
        RECT 92.490 203.215 97.835 203.650 ;
        RECT 98.010 203.215 103.355 203.650 ;
        RECT 103.530 203.215 108.875 203.650 ;
        RECT 109.050 203.215 114.395 203.650 ;
        RECT 114.565 203.215 114.855 204.380 ;
        RECT 117.080 203.650 117.430 204.900 ;
        RECT 118.910 204.390 119.250 205.220 ;
        RECT 122.600 203.650 122.950 204.900 ;
        RECT 124.430 204.390 124.770 205.220 ;
        RECT 126.525 205.015 127.735 205.765 ;
        RECT 126.525 204.305 127.045 204.845 ;
        RECT 127.215 204.475 127.735 205.015 ;
        RECT 115.490 203.215 120.835 203.650 ;
        RECT 121.010 203.215 126.355 203.650 ;
        RECT 126.525 203.215 127.735 204.305 ;
        RECT 14.660 203.045 127.820 203.215 ;
        RECT 14.745 201.955 15.955 203.045 ;
        RECT 14.745 201.245 15.265 201.785 ;
        RECT 15.435 201.415 15.955 201.955 ;
        RECT 16.125 201.955 18.715 203.045 ;
        RECT 18.890 202.610 24.235 203.045 ;
        RECT 16.125 201.435 17.335 201.955 ;
        RECT 17.505 201.265 18.715 201.785 ;
        RECT 20.480 201.360 20.830 202.610 ;
        RECT 24.405 201.880 24.695 203.045 ;
        RECT 25.325 201.955 27.915 203.045 ;
        RECT 28.090 202.610 33.435 203.045 ;
        RECT 33.610 202.610 38.955 203.045 ;
        RECT 39.130 202.610 44.475 203.045 ;
        RECT 44.650 202.610 49.995 203.045 ;
        RECT 14.745 200.495 15.955 201.245 ;
        RECT 16.125 200.495 18.715 201.265 ;
        RECT 22.310 201.040 22.650 201.870 ;
        RECT 25.325 201.435 26.535 201.955 ;
        RECT 26.705 201.265 27.915 201.785 ;
        RECT 29.680 201.360 30.030 202.610 ;
        RECT 18.890 200.495 24.235 201.040 ;
        RECT 24.405 200.495 24.695 201.220 ;
        RECT 25.325 200.495 27.915 201.265 ;
        RECT 31.510 201.040 31.850 201.870 ;
        RECT 35.200 201.360 35.550 202.610 ;
        RECT 37.030 201.040 37.370 201.870 ;
        RECT 40.720 201.360 41.070 202.610 ;
        RECT 42.550 201.040 42.890 201.870 ;
        RECT 46.240 201.360 46.590 202.610 ;
        RECT 50.165 201.880 50.455 203.045 ;
        RECT 50.625 201.955 54.135 203.045 ;
        RECT 54.310 202.610 59.655 203.045 ;
        RECT 48.070 201.040 48.410 201.870 ;
        RECT 50.625 201.435 52.315 201.955 ;
        RECT 52.485 201.265 54.135 201.785 ;
        RECT 55.900 201.360 56.250 202.610 ;
        RECT 59.830 202.375 60.085 202.875 ;
        RECT 60.255 202.545 60.585 203.045 ;
        RECT 59.830 202.205 60.580 202.375 ;
        RECT 28.090 200.495 33.435 201.040 ;
        RECT 33.610 200.495 38.955 201.040 ;
        RECT 39.130 200.495 44.475 201.040 ;
        RECT 44.650 200.495 49.995 201.040 ;
        RECT 50.165 200.495 50.455 201.220 ;
        RECT 50.625 200.495 54.135 201.265 ;
        RECT 57.730 201.040 58.070 201.870 ;
        RECT 59.830 201.385 60.180 202.035 ;
        RECT 60.350 201.215 60.580 202.205 ;
        RECT 59.830 201.045 60.580 201.215 ;
        RECT 54.310 200.495 59.655 201.040 ;
        RECT 59.830 200.755 60.085 201.045 ;
        RECT 60.255 200.495 60.585 200.875 ;
        RECT 60.755 200.755 60.925 202.875 ;
        RECT 61.095 202.075 61.420 202.860 ;
        RECT 61.590 202.585 61.840 203.045 ;
        RECT 62.010 202.545 62.260 202.875 ;
        RECT 62.475 202.545 63.155 202.875 ;
        RECT 62.010 202.415 62.180 202.545 ;
        RECT 61.785 202.245 62.180 202.415 ;
        RECT 61.155 201.025 61.615 202.075 ;
        RECT 61.785 200.885 61.955 202.245 ;
        RECT 62.350 201.985 62.815 202.375 ;
        RECT 62.125 201.175 62.475 201.795 ;
        RECT 62.645 201.395 62.815 201.985 ;
        RECT 62.985 201.765 63.155 202.545 ;
        RECT 63.325 202.445 63.495 202.785 ;
        RECT 63.730 202.615 64.060 203.045 ;
        RECT 64.230 202.445 64.400 202.785 ;
        RECT 64.695 202.585 65.065 203.045 ;
        RECT 63.325 202.275 64.400 202.445 ;
        RECT 65.235 202.415 65.405 202.875 ;
        RECT 65.640 202.535 66.510 202.875 ;
        RECT 66.680 202.585 66.930 203.045 ;
        RECT 64.845 202.245 65.405 202.415 ;
        RECT 64.845 202.105 65.015 202.245 ;
        RECT 63.515 201.935 65.015 202.105 ;
        RECT 65.710 202.075 66.170 202.365 ;
        RECT 62.985 201.595 64.675 201.765 ;
        RECT 62.645 201.175 63.000 201.395 ;
        RECT 63.170 200.885 63.340 201.595 ;
        RECT 63.545 201.175 64.335 201.425 ;
        RECT 64.505 201.415 64.675 201.595 ;
        RECT 64.845 201.245 65.015 201.935 ;
        RECT 61.285 200.495 61.615 200.855 ;
        RECT 61.785 200.715 62.280 200.885 ;
        RECT 62.485 200.715 63.340 200.885 ;
        RECT 64.215 200.495 64.545 200.955 ;
        RECT 64.755 200.855 65.015 201.245 ;
        RECT 65.205 202.065 66.170 202.075 ;
        RECT 66.340 202.155 66.510 202.535 ;
        RECT 67.100 202.495 67.270 202.785 ;
        RECT 67.450 202.665 67.780 203.045 ;
        RECT 67.100 202.325 67.900 202.495 ;
        RECT 65.205 201.905 65.880 202.065 ;
        RECT 66.340 201.985 67.560 202.155 ;
        RECT 65.205 201.115 65.415 201.905 ;
        RECT 66.340 201.895 66.510 201.985 ;
        RECT 65.585 201.115 65.935 201.735 ;
        RECT 66.105 201.725 66.510 201.895 ;
        RECT 66.105 200.945 66.275 201.725 ;
        RECT 66.445 201.275 66.665 201.555 ;
        RECT 66.845 201.445 67.385 201.815 ;
        RECT 67.730 201.705 67.900 202.325 ;
        RECT 68.075 201.985 68.245 203.045 ;
        RECT 68.455 202.035 68.745 202.875 ;
        RECT 68.915 202.205 69.085 203.045 ;
        RECT 69.295 202.035 69.545 202.875 ;
        RECT 69.755 202.205 69.925 203.045 ;
        RECT 68.455 201.865 70.180 202.035 ;
        RECT 66.445 201.105 66.975 201.275 ;
        RECT 64.755 200.685 65.105 200.855 ;
        RECT 65.325 200.665 66.275 200.945 ;
        RECT 66.445 200.495 66.635 200.935 ;
        RECT 66.805 200.875 66.975 201.105 ;
        RECT 67.145 201.045 67.385 201.445 ;
        RECT 67.555 201.695 67.900 201.705 ;
        RECT 67.555 201.485 69.585 201.695 ;
        RECT 67.555 201.230 67.880 201.485 ;
        RECT 69.770 201.315 70.180 201.865 ;
        RECT 67.555 200.875 67.875 201.230 ;
        RECT 66.805 200.705 67.875 200.875 ;
        RECT 68.075 200.495 68.245 201.305 ;
        RECT 68.415 201.145 70.180 201.315 ;
        RECT 70.405 201.905 70.665 202.875 ;
        RECT 70.860 202.635 71.190 203.045 ;
        RECT 71.390 202.455 71.560 202.875 ;
        RECT 71.775 202.635 72.445 203.045 ;
        RECT 72.680 202.455 72.850 202.875 ;
        RECT 73.155 202.605 73.485 203.045 ;
        RECT 70.835 202.285 72.850 202.455 ;
        RECT 73.655 202.425 73.830 202.875 ;
        RECT 74.090 202.620 74.425 203.045 ;
        RECT 74.595 202.440 74.780 202.845 ;
        RECT 70.405 201.215 70.575 201.905 ;
        RECT 70.835 201.735 71.005 202.285 ;
        RECT 70.745 201.405 71.005 201.735 ;
        RECT 68.415 200.665 68.745 201.145 ;
        RECT 68.915 200.495 69.085 200.965 ;
        RECT 69.255 200.665 69.585 201.145 ;
        RECT 69.755 200.495 69.925 200.965 ;
        RECT 70.405 200.750 70.745 201.215 ;
        RECT 71.175 201.075 71.515 202.105 ;
        RECT 71.705 201.005 71.975 202.105 ;
        RECT 70.410 200.705 70.745 200.750 ;
        RECT 70.915 200.495 71.245 200.875 ;
        RECT 71.705 200.835 72.015 201.005 ;
        RECT 71.705 200.830 71.975 200.835 ;
        RECT 72.200 200.830 72.480 202.105 ;
        RECT 72.680 200.995 72.850 202.285 ;
        RECT 73.200 202.255 73.830 202.425 ;
        RECT 74.115 202.265 74.780 202.440 ;
        RECT 74.985 202.265 75.315 203.045 ;
        RECT 73.200 201.735 73.370 202.255 ;
        RECT 73.020 201.405 73.370 201.735 ;
        RECT 73.550 201.405 73.915 202.085 ;
        RECT 73.200 201.235 73.370 201.405 ;
        RECT 74.115 201.235 74.455 202.265 ;
        RECT 75.485 202.075 75.755 202.845 ;
        RECT 74.625 201.905 75.755 202.075 ;
        RECT 74.625 201.405 74.875 201.905 ;
        RECT 73.200 201.065 73.830 201.235 ;
        RECT 74.115 201.065 74.800 201.235 ;
        RECT 75.055 201.155 75.415 201.735 ;
        RECT 72.680 200.665 72.910 200.995 ;
        RECT 73.155 200.495 73.485 200.875 ;
        RECT 73.655 200.665 73.830 201.065 ;
        RECT 74.090 200.495 74.425 200.895 ;
        RECT 74.595 200.665 74.800 201.065 ;
        RECT 75.585 200.995 75.755 201.905 ;
        RECT 75.925 201.880 76.215 203.045 ;
        RECT 76.845 202.175 77.120 202.875 ;
        RECT 77.290 202.500 77.545 203.045 ;
        RECT 77.715 202.535 78.195 202.875 ;
        RECT 78.370 202.490 78.975 203.045 ;
        RECT 78.360 202.390 78.975 202.490 ;
        RECT 78.360 202.365 78.545 202.390 ;
        RECT 75.010 200.495 75.285 200.975 ;
        RECT 75.495 200.665 75.755 200.995 ;
        RECT 75.925 200.495 76.215 201.220 ;
        RECT 76.845 201.145 77.015 202.175 ;
        RECT 77.290 202.045 78.045 202.295 ;
        RECT 78.215 202.120 78.545 202.365 ;
        RECT 77.290 202.010 78.060 202.045 ;
        RECT 77.290 202.000 78.075 202.010 ;
        RECT 77.185 201.985 78.080 202.000 ;
        RECT 77.185 201.970 78.100 201.985 ;
        RECT 77.185 201.960 78.120 201.970 ;
        RECT 77.185 201.950 78.145 201.960 ;
        RECT 77.185 201.920 78.215 201.950 ;
        RECT 77.185 201.890 78.235 201.920 ;
        RECT 77.185 201.860 78.255 201.890 ;
        RECT 77.185 201.835 78.285 201.860 ;
        RECT 77.185 201.800 78.320 201.835 ;
        RECT 77.185 201.795 78.350 201.800 ;
        RECT 77.185 201.400 77.415 201.795 ;
        RECT 77.960 201.790 78.350 201.795 ;
        RECT 77.985 201.780 78.350 201.790 ;
        RECT 78.000 201.775 78.350 201.780 ;
        RECT 78.015 201.770 78.350 201.775 ;
        RECT 78.715 201.770 78.975 202.220 ;
        RECT 78.015 201.765 78.975 201.770 ;
        RECT 78.025 201.755 78.975 201.765 ;
        RECT 78.035 201.750 78.975 201.755 ;
        RECT 78.045 201.740 78.975 201.750 ;
        RECT 78.050 201.730 78.975 201.740 ;
        RECT 78.055 201.725 78.975 201.730 ;
        RECT 78.065 201.710 78.975 201.725 ;
        RECT 78.070 201.695 78.975 201.710 ;
        RECT 78.080 201.670 78.975 201.695 ;
        RECT 77.585 201.200 77.915 201.625 ;
        RECT 77.665 201.175 77.915 201.200 ;
        RECT 76.845 200.665 77.105 201.145 ;
        RECT 77.275 200.495 77.525 201.035 ;
        RECT 77.695 200.715 77.915 201.175 ;
        RECT 78.085 201.600 78.975 201.670 ;
        RECT 79.610 201.855 79.865 202.735 ;
        RECT 80.035 201.905 80.340 203.045 ;
        RECT 80.680 202.665 81.010 203.045 ;
        RECT 81.190 202.495 81.360 202.785 ;
        RECT 81.530 202.585 81.780 203.045 ;
        RECT 80.560 202.325 81.360 202.495 ;
        RECT 81.950 202.535 82.820 202.875 ;
        RECT 78.085 200.875 78.255 201.600 ;
        RECT 78.425 201.045 78.975 201.430 ;
        RECT 79.610 201.205 79.820 201.855 ;
        RECT 80.560 201.735 80.730 202.325 ;
        RECT 81.950 202.155 82.120 202.535 ;
        RECT 83.055 202.415 83.225 202.875 ;
        RECT 83.395 202.585 83.765 203.045 ;
        RECT 84.060 202.445 84.230 202.785 ;
        RECT 84.400 202.615 84.730 203.045 ;
        RECT 84.965 202.445 85.135 202.785 ;
        RECT 80.900 201.985 82.120 202.155 ;
        RECT 82.290 202.075 82.750 202.365 ;
        RECT 83.055 202.245 83.615 202.415 ;
        RECT 84.060 202.275 85.135 202.445 ;
        RECT 85.305 202.545 85.985 202.875 ;
        RECT 86.200 202.545 86.450 202.875 ;
        RECT 86.620 202.585 86.870 203.045 ;
        RECT 83.445 202.105 83.615 202.245 ;
        RECT 82.290 202.065 83.255 202.075 ;
        RECT 81.950 201.895 82.120 201.985 ;
        RECT 82.580 201.905 83.255 202.065 ;
        RECT 79.990 201.705 80.730 201.735 ;
        RECT 79.990 201.405 80.905 201.705 ;
        RECT 80.580 201.230 80.905 201.405 ;
        RECT 78.085 200.705 78.975 200.875 ;
        RECT 79.610 200.675 79.865 201.205 ;
        RECT 80.035 200.495 80.340 200.955 ;
        RECT 80.585 200.875 80.905 201.230 ;
        RECT 81.075 201.445 81.615 201.815 ;
        RECT 81.950 201.725 82.355 201.895 ;
        RECT 81.075 201.045 81.315 201.445 ;
        RECT 81.795 201.275 82.015 201.555 ;
        RECT 81.485 201.105 82.015 201.275 ;
        RECT 81.485 200.875 81.655 201.105 ;
        RECT 82.185 200.945 82.355 201.725 ;
        RECT 82.525 201.115 82.875 201.735 ;
        RECT 83.045 201.115 83.255 201.905 ;
        RECT 83.445 201.935 84.945 202.105 ;
        RECT 83.445 201.245 83.615 201.935 ;
        RECT 85.305 201.765 85.475 202.545 ;
        RECT 86.280 202.415 86.450 202.545 ;
        RECT 83.785 201.595 85.475 201.765 ;
        RECT 85.645 201.985 86.110 202.375 ;
        RECT 86.280 202.245 86.675 202.415 ;
        RECT 83.785 201.415 83.955 201.595 ;
        RECT 80.585 200.705 81.655 200.875 ;
        RECT 81.825 200.495 82.015 200.935 ;
        RECT 82.185 200.665 83.135 200.945 ;
        RECT 83.445 200.855 83.705 201.245 ;
        RECT 84.125 201.175 84.915 201.425 ;
        RECT 83.355 200.685 83.705 200.855 ;
        RECT 83.915 200.495 84.245 200.955 ;
        RECT 85.120 200.885 85.290 201.595 ;
        RECT 85.645 201.395 85.815 201.985 ;
        RECT 85.460 201.175 85.815 201.395 ;
        RECT 85.985 201.175 86.335 201.795 ;
        RECT 86.505 200.885 86.675 202.245 ;
        RECT 87.040 202.075 87.365 202.860 ;
        RECT 86.845 201.025 87.305 202.075 ;
        RECT 85.120 200.715 85.975 200.885 ;
        RECT 86.180 200.715 86.675 200.885 ;
        RECT 86.845 200.495 87.175 200.855 ;
        RECT 87.535 200.755 87.705 202.875 ;
        RECT 87.875 202.545 88.205 203.045 ;
        RECT 88.375 202.375 88.630 202.875 ;
        RECT 87.880 202.205 88.630 202.375 ;
        RECT 87.880 201.215 88.110 202.205 ;
        RECT 88.280 201.385 88.630 202.035 ;
        RECT 88.805 201.955 90.475 203.045 ;
        RECT 90.650 202.610 95.995 203.045 ;
        RECT 96.170 202.610 101.515 203.045 ;
        RECT 88.805 201.435 89.555 201.955 ;
        RECT 89.725 201.265 90.475 201.785 ;
        RECT 92.240 201.360 92.590 202.610 ;
        RECT 87.880 201.045 88.630 201.215 ;
        RECT 87.875 200.495 88.205 200.875 ;
        RECT 88.375 200.755 88.630 201.045 ;
        RECT 88.805 200.495 90.475 201.265 ;
        RECT 94.070 201.040 94.410 201.870 ;
        RECT 97.760 201.360 98.110 202.610 ;
        RECT 101.685 201.880 101.975 203.045 ;
        RECT 102.605 201.955 104.275 203.045 ;
        RECT 104.450 202.610 109.795 203.045 ;
        RECT 109.970 202.610 115.315 203.045 ;
        RECT 115.490 202.610 120.835 203.045 ;
        RECT 121.010 202.610 126.355 203.045 ;
        RECT 99.590 201.040 99.930 201.870 ;
        RECT 102.605 201.435 103.355 201.955 ;
        RECT 103.525 201.265 104.275 201.785 ;
        RECT 106.040 201.360 106.390 202.610 ;
        RECT 90.650 200.495 95.995 201.040 ;
        RECT 96.170 200.495 101.515 201.040 ;
        RECT 101.685 200.495 101.975 201.220 ;
        RECT 102.605 200.495 104.275 201.265 ;
        RECT 107.870 201.040 108.210 201.870 ;
        RECT 111.560 201.360 111.910 202.610 ;
        RECT 113.390 201.040 113.730 201.870 ;
        RECT 117.080 201.360 117.430 202.610 ;
        RECT 118.910 201.040 119.250 201.870 ;
        RECT 122.600 201.360 122.950 202.610 ;
        RECT 126.525 201.955 127.735 203.045 ;
        RECT 124.430 201.040 124.770 201.870 ;
        RECT 126.525 201.415 127.045 201.955 ;
        RECT 127.215 201.245 127.735 201.785 ;
        RECT 104.450 200.495 109.795 201.040 ;
        RECT 109.970 200.495 115.315 201.040 ;
        RECT 115.490 200.495 120.835 201.040 ;
        RECT 121.010 200.495 126.355 201.040 ;
        RECT 126.525 200.495 127.735 201.245 ;
        RECT 14.660 200.325 127.820 200.495 ;
        RECT 14.745 199.575 15.955 200.325 ;
        RECT 14.745 199.035 15.265 199.575 ;
        RECT 17.045 199.555 20.555 200.325 ;
        RECT 20.730 199.780 26.075 200.325 ;
        RECT 26.250 199.780 31.595 200.325 ;
        RECT 31.770 199.780 37.115 200.325 ;
        RECT 15.435 198.865 15.955 199.405 ;
        RECT 14.745 197.775 15.955 198.865 ;
        RECT 17.045 198.865 18.735 199.385 ;
        RECT 18.905 199.035 20.555 199.555 ;
        RECT 17.045 197.775 20.555 198.865 ;
        RECT 22.320 198.210 22.670 199.460 ;
        RECT 24.150 198.950 24.490 199.780 ;
        RECT 27.840 198.210 28.190 199.460 ;
        RECT 29.670 198.950 30.010 199.780 ;
        RECT 33.360 198.210 33.710 199.460 ;
        RECT 35.190 198.950 35.530 199.780 ;
        RECT 37.285 199.600 37.575 200.325 ;
        RECT 38.205 199.555 40.795 200.325 ;
        RECT 40.970 199.780 46.315 200.325 ;
        RECT 46.490 199.780 51.835 200.325 ;
        RECT 52.010 199.780 57.355 200.325 ;
        RECT 57.530 199.780 62.875 200.325 ;
        RECT 20.730 197.775 26.075 198.210 ;
        RECT 26.250 197.775 31.595 198.210 ;
        RECT 31.770 197.775 37.115 198.210 ;
        RECT 37.285 197.775 37.575 198.940 ;
        RECT 38.205 198.865 39.415 199.385 ;
        RECT 39.585 199.035 40.795 199.555 ;
        RECT 38.205 197.775 40.795 198.865 ;
        RECT 42.560 198.210 42.910 199.460 ;
        RECT 44.390 198.950 44.730 199.780 ;
        RECT 48.080 198.210 48.430 199.460 ;
        RECT 49.910 198.950 50.250 199.780 ;
        RECT 53.600 198.210 53.950 199.460 ;
        RECT 55.430 198.950 55.770 199.780 ;
        RECT 59.120 198.210 59.470 199.460 ;
        RECT 60.950 198.950 61.290 199.780 ;
        RECT 63.045 199.600 63.335 200.325 ;
        RECT 63.965 199.555 67.475 200.325 ;
        RECT 40.970 197.775 46.315 198.210 ;
        RECT 46.490 197.775 51.835 198.210 ;
        RECT 52.010 197.775 57.355 198.210 ;
        RECT 57.530 197.775 62.875 198.210 ;
        RECT 63.045 197.775 63.335 198.940 ;
        RECT 63.965 198.865 65.655 199.385 ;
        RECT 65.825 199.035 67.475 199.555 ;
        RECT 67.645 199.650 67.905 200.155 ;
        RECT 68.085 199.945 68.415 200.325 ;
        RECT 68.595 199.775 68.765 200.155 ;
        RECT 69.030 199.925 69.365 200.325 ;
        RECT 63.965 197.775 67.475 198.865 ;
        RECT 67.645 198.850 67.815 199.650 ;
        RECT 68.100 199.605 68.765 199.775 ;
        RECT 69.535 199.755 69.740 200.155 ;
        RECT 69.950 199.845 70.225 200.325 ;
        RECT 70.435 199.825 70.695 200.155 ;
        RECT 68.100 199.350 68.270 199.605 ;
        RECT 69.055 199.585 69.740 199.755 ;
        RECT 67.985 199.020 68.270 199.350 ;
        RECT 68.505 199.055 68.835 199.425 ;
        RECT 68.100 198.875 68.270 199.020 ;
        RECT 67.645 197.945 67.915 198.850 ;
        RECT 68.100 198.705 68.765 198.875 ;
        RECT 68.085 197.775 68.415 198.535 ;
        RECT 68.595 197.945 68.765 198.705 ;
        RECT 69.055 198.555 69.395 199.585 ;
        RECT 69.565 198.915 69.815 199.415 ;
        RECT 69.995 199.085 70.355 199.665 ;
        RECT 70.525 198.915 70.695 199.825 ;
        RECT 69.565 198.745 70.695 198.915 ;
        RECT 69.055 198.380 69.720 198.555 ;
        RECT 69.030 197.775 69.365 198.200 ;
        RECT 69.535 197.975 69.720 198.380 ;
        RECT 69.925 197.775 70.255 198.555 ;
        RECT 70.425 197.975 70.695 198.745 ;
        RECT 70.865 197.945 71.125 200.155 ;
        RECT 71.295 199.945 71.625 200.325 ;
        RECT 71.835 199.415 72.030 199.990 ;
        RECT 72.300 199.415 72.485 199.995 ;
        RECT 71.295 198.495 71.465 199.415 ;
        RECT 71.775 199.085 72.030 199.415 ;
        RECT 72.255 199.085 72.485 199.415 ;
        RECT 72.735 199.985 74.215 200.155 ;
        RECT 72.735 199.085 72.905 199.985 ;
        RECT 73.075 199.485 73.625 199.815 ;
        RECT 73.815 199.655 74.215 199.985 ;
        RECT 74.395 199.945 74.725 200.325 ;
        RECT 75.035 199.825 75.295 200.155 ;
        RECT 71.835 198.775 72.030 199.085 ;
        RECT 72.300 198.775 72.485 199.085 ;
        RECT 73.075 198.495 73.245 199.485 ;
        RECT 73.815 199.175 73.985 199.655 ;
        RECT 74.565 199.465 74.775 199.645 ;
        RECT 74.155 199.295 74.775 199.465 ;
        RECT 71.295 198.325 73.245 198.495 ;
        RECT 73.415 199.005 73.985 199.175 ;
        RECT 75.125 199.125 75.295 199.825 ;
        RECT 73.415 198.495 73.585 199.005 ;
        RECT 74.165 198.955 75.295 199.125 ;
        RECT 74.165 198.835 74.335 198.955 ;
        RECT 73.755 198.665 74.335 198.835 ;
        RECT 73.415 198.325 74.155 198.495 ;
        RECT 74.605 198.455 74.955 198.785 ;
        RECT 71.295 197.775 71.625 198.155 ;
        RECT 72.050 197.945 72.220 198.325 ;
        RECT 72.480 197.775 72.810 198.155 ;
        RECT 73.005 197.945 73.175 198.325 ;
        RECT 73.385 197.775 73.715 198.155 ;
        RECT 73.965 197.945 74.155 198.325 ;
        RECT 75.125 198.275 75.295 198.955 ;
        RECT 74.395 197.775 74.725 198.155 ;
        RECT 75.035 197.945 75.295 198.275 ;
        RECT 75.465 199.585 75.850 200.155 ;
        RECT 76.020 199.865 76.345 200.325 ;
        RECT 76.865 199.695 77.145 200.155 ;
        RECT 75.465 198.915 75.745 199.585 ;
        RECT 76.020 199.525 77.145 199.695 ;
        RECT 76.020 199.415 76.470 199.525 ;
        RECT 75.915 199.085 76.470 199.415 ;
        RECT 77.335 199.355 77.735 200.155 ;
        RECT 78.135 199.865 78.405 200.325 ;
        RECT 78.575 199.695 78.860 200.155 ;
        RECT 75.465 197.945 75.850 198.915 ;
        RECT 76.020 198.625 76.470 199.085 ;
        RECT 76.640 198.795 77.735 199.355 ;
        RECT 76.020 198.405 77.145 198.625 ;
        RECT 76.020 197.775 76.345 198.235 ;
        RECT 76.865 197.945 77.145 198.405 ;
        RECT 77.335 197.945 77.735 198.795 ;
        RECT 77.905 199.525 78.860 199.695 ;
        RECT 79.180 199.585 79.795 200.155 ;
        RECT 79.965 199.815 80.180 200.325 ;
        RECT 80.410 199.815 80.690 200.145 ;
        RECT 80.870 199.815 81.110 200.325 ;
        RECT 77.905 198.625 78.115 199.525 ;
        RECT 78.285 198.795 78.975 199.355 ;
        RECT 77.905 198.405 78.860 198.625 ;
        RECT 78.135 197.775 78.405 198.235 ;
        RECT 78.575 197.945 78.860 198.405 ;
        RECT 79.180 198.565 79.495 199.585 ;
        RECT 79.665 198.915 79.835 199.415 ;
        RECT 80.085 199.085 80.350 199.645 ;
        RECT 80.520 198.915 80.690 199.815 ;
        RECT 80.860 199.085 81.215 199.645 ;
        RECT 81.445 199.525 82.140 200.155 ;
        RECT 82.345 199.525 82.655 200.325 ;
        RECT 82.915 199.775 83.085 200.155 ;
        RECT 83.265 199.945 83.595 200.325 ;
        RECT 82.915 199.605 83.580 199.775 ;
        RECT 83.775 199.650 84.035 200.155 ;
        RECT 81.465 199.085 81.800 199.335 ;
        RECT 81.970 198.925 82.140 199.525 ;
        RECT 82.310 199.085 82.645 199.355 ;
        RECT 82.845 199.055 83.175 199.425 ;
        RECT 83.410 199.350 83.580 199.605 ;
        RECT 83.410 199.020 83.695 199.350 ;
        RECT 79.665 198.745 81.090 198.915 ;
        RECT 79.180 197.945 79.715 198.565 ;
        RECT 79.885 197.775 80.215 198.575 ;
        RECT 80.700 198.570 81.090 198.745 ;
        RECT 81.445 197.775 81.705 198.915 ;
        RECT 81.875 197.945 82.205 198.925 ;
        RECT 82.375 197.775 82.655 198.915 ;
        RECT 83.410 198.875 83.580 199.020 ;
        RECT 82.915 198.705 83.580 198.875 ;
        RECT 83.865 198.850 84.035 199.650 ;
        RECT 84.245 199.505 84.475 200.325 ;
        RECT 84.645 199.525 84.975 200.155 ;
        RECT 84.225 199.085 84.555 199.335 ;
        RECT 84.725 198.925 84.975 199.525 ;
        RECT 85.145 199.505 85.355 200.325 ;
        RECT 85.645 199.505 85.855 200.325 ;
        RECT 86.025 199.525 86.355 200.155 ;
        RECT 82.915 197.945 83.085 198.705 ;
        RECT 83.265 197.775 83.595 198.535 ;
        RECT 83.765 197.945 84.035 198.850 ;
        RECT 84.245 197.775 84.475 198.915 ;
        RECT 84.645 197.945 84.975 198.925 ;
        RECT 86.025 198.925 86.275 199.525 ;
        RECT 86.525 199.505 86.755 200.325 ;
        RECT 86.965 199.555 88.635 200.325 ;
        RECT 88.805 199.600 89.095 200.325 ;
        RECT 89.725 199.555 91.395 200.325 ;
        RECT 91.570 199.780 96.915 200.325 ;
        RECT 86.445 199.085 86.775 199.335 ;
        RECT 85.145 197.775 85.355 198.915 ;
        RECT 85.645 197.775 85.855 198.915 ;
        RECT 86.025 197.945 86.355 198.925 ;
        RECT 86.525 197.775 86.755 198.915 ;
        RECT 86.965 198.865 87.715 199.385 ;
        RECT 87.885 199.035 88.635 199.555 ;
        RECT 86.965 197.775 88.635 198.865 ;
        RECT 88.805 197.775 89.095 198.940 ;
        RECT 89.725 198.865 90.475 199.385 ;
        RECT 90.645 199.035 91.395 199.555 ;
        RECT 89.725 197.775 91.395 198.865 ;
        RECT 93.160 198.210 93.510 199.460 ;
        RECT 94.990 198.950 95.330 199.780 ;
        RECT 97.090 199.615 97.345 200.145 ;
        RECT 97.515 199.865 97.820 200.325 ;
        RECT 98.065 199.945 99.135 200.115 ;
        RECT 97.090 198.965 97.300 199.615 ;
        RECT 98.065 199.590 98.385 199.945 ;
        RECT 98.060 199.415 98.385 199.590 ;
        RECT 97.470 199.115 98.385 199.415 ;
        RECT 98.555 199.375 98.795 199.775 ;
        RECT 98.965 199.715 99.135 199.945 ;
        RECT 99.305 199.885 99.495 200.325 ;
        RECT 99.665 199.875 100.615 200.155 ;
        RECT 100.835 199.965 101.185 200.135 ;
        RECT 98.965 199.545 99.495 199.715 ;
        RECT 97.470 199.085 98.210 199.115 ;
        RECT 91.570 197.775 96.915 198.210 ;
        RECT 97.090 198.085 97.345 198.965 ;
        RECT 97.515 197.775 97.820 198.915 ;
        RECT 98.040 198.495 98.210 199.085 ;
        RECT 98.555 199.005 99.095 199.375 ;
        RECT 99.275 199.265 99.495 199.545 ;
        RECT 99.665 199.095 99.835 199.875 ;
        RECT 99.430 198.925 99.835 199.095 ;
        RECT 100.005 199.085 100.355 199.705 ;
        RECT 99.430 198.835 99.600 198.925 ;
        RECT 100.525 198.915 100.735 199.705 ;
        RECT 98.380 198.665 99.600 198.835 ;
        RECT 100.060 198.755 100.735 198.915 ;
        RECT 98.040 198.325 98.840 198.495 ;
        RECT 98.160 197.775 98.490 198.155 ;
        RECT 98.670 198.035 98.840 198.325 ;
        RECT 99.430 198.285 99.600 198.665 ;
        RECT 99.770 198.745 100.735 198.755 ;
        RECT 100.925 199.575 101.185 199.965 ;
        RECT 101.395 199.865 101.725 200.325 ;
        RECT 102.600 199.935 103.455 200.105 ;
        RECT 103.660 199.935 104.155 200.105 ;
        RECT 104.325 199.965 104.655 200.325 ;
        RECT 100.925 198.885 101.095 199.575 ;
        RECT 101.265 199.225 101.435 199.405 ;
        RECT 101.605 199.395 102.395 199.645 ;
        RECT 102.600 199.225 102.770 199.935 ;
        RECT 102.940 199.425 103.295 199.645 ;
        RECT 101.265 199.055 102.955 199.225 ;
        RECT 99.770 198.455 100.230 198.745 ;
        RECT 100.925 198.715 102.425 198.885 ;
        RECT 100.925 198.575 101.095 198.715 ;
        RECT 100.535 198.405 101.095 198.575 ;
        RECT 99.010 197.775 99.260 198.235 ;
        RECT 99.430 197.945 100.300 198.285 ;
        RECT 100.535 197.945 100.705 198.405 ;
        RECT 101.540 198.375 102.615 198.545 ;
        RECT 100.875 197.775 101.245 198.235 ;
        RECT 101.540 198.035 101.710 198.375 ;
        RECT 101.880 197.775 102.210 198.205 ;
        RECT 102.445 198.035 102.615 198.375 ;
        RECT 102.785 198.275 102.955 199.055 ;
        RECT 103.125 198.835 103.295 199.425 ;
        RECT 103.465 199.025 103.815 199.645 ;
        RECT 103.125 198.445 103.590 198.835 ;
        RECT 103.985 198.575 104.155 199.935 ;
        RECT 104.325 198.745 104.785 199.795 ;
        RECT 103.760 198.405 104.155 198.575 ;
        RECT 103.760 198.275 103.930 198.405 ;
        RECT 102.785 197.945 103.465 198.275 ;
        RECT 103.680 197.945 103.930 198.275 ;
        RECT 104.100 197.775 104.350 198.235 ;
        RECT 104.520 197.960 104.845 198.745 ;
        RECT 105.015 197.945 105.185 200.065 ;
        RECT 105.355 199.945 105.685 200.325 ;
        RECT 105.855 199.775 106.110 200.065 ;
        RECT 105.360 199.605 106.110 199.775 ;
        RECT 105.360 198.615 105.590 199.605 ;
        RECT 106.285 199.555 108.875 200.325 ;
        RECT 109.050 199.780 114.395 200.325 ;
        RECT 105.760 198.785 106.110 199.435 ;
        RECT 106.285 198.865 107.495 199.385 ;
        RECT 107.665 199.035 108.875 199.555 ;
        RECT 105.360 198.445 106.110 198.615 ;
        RECT 105.355 197.775 105.685 198.275 ;
        RECT 105.855 197.945 106.110 198.445 ;
        RECT 106.285 197.775 108.875 198.865 ;
        RECT 110.640 198.210 110.990 199.460 ;
        RECT 112.470 198.950 112.810 199.780 ;
        RECT 114.565 199.600 114.855 200.325 ;
        RECT 115.490 199.780 120.835 200.325 ;
        RECT 121.010 199.780 126.355 200.325 ;
        RECT 109.050 197.775 114.395 198.210 ;
        RECT 114.565 197.775 114.855 198.940 ;
        RECT 117.080 198.210 117.430 199.460 ;
        RECT 118.910 198.950 119.250 199.780 ;
        RECT 122.600 198.210 122.950 199.460 ;
        RECT 124.430 198.950 124.770 199.780 ;
        RECT 126.525 199.575 127.735 200.325 ;
        RECT 126.525 198.865 127.045 199.405 ;
        RECT 127.215 199.035 127.735 199.575 ;
        RECT 115.490 197.775 120.835 198.210 ;
        RECT 121.010 197.775 126.355 198.210 ;
        RECT 126.525 197.775 127.735 198.865 ;
        RECT 14.660 197.605 127.820 197.775 ;
        RECT 14.745 196.515 15.955 197.605 ;
        RECT 14.745 195.805 15.265 196.345 ;
        RECT 15.435 195.975 15.955 196.515 ;
        RECT 16.125 196.515 18.715 197.605 ;
        RECT 18.890 197.170 24.235 197.605 ;
        RECT 16.125 195.995 17.335 196.515 ;
        RECT 17.505 195.825 18.715 196.345 ;
        RECT 20.480 195.920 20.830 197.170 ;
        RECT 24.405 196.440 24.695 197.605 ;
        RECT 25.325 196.515 27.915 197.605 ;
        RECT 28.090 197.170 33.435 197.605 ;
        RECT 33.610 197.170 38.955 197.605 ;
        RECT 39.130 197.170 44.475 197.605 ;
        RECT 44.650 197.170 49.995 197.605 ;
        RECT 14.745 195.055 15.955 195.805 ;
        RECT 16.125 195.055 18.715 195.825 ;
        RECT 22.310 195.600 22.650 196.430 ;
        RECT 25.325 195.995 26.535 196.515 ;
        RECT 26.705 195.825 27.915 196.345 ;
        RECT 29.680 195.920 30.030 197.170 ;
        RECT 18.890 195.055 24.235 195.600 ;
        RECT 24.405 195.055 24.695 195.780 ;
        RECT 25.325 195.055 27.915 195.825 ;
        RECT 31.510 195.600 31.850 196.430 ;
        RECT 35.200 195.920 35.550 197.170 ;
        RECT 37.030 195.600 37.370 196.430 ;
        RECT 40.720 195.920 41.070 197.170 ;
        RECT 42.550 195.600 42.890 196.430 ;
        RECT 46.240 195.920 46.590 197.170 ;
        RECT 50.165 196.440 50.455 197.605 ;
        RECT 51.085 196.515 52.755 197.605 ;
        RECT 48.070 195.600 48.410 196.430 ;
        RECT 51.085 195.995 51.835 196.515 ;
        RECT 52.985 196.465 53.195 197.605 ;
        RECT 53.365 196.455 53.695 197.435 ;
        RECT 53.865 196.465 54.095 197.605 ;
        RECT 54.420 196.975 54.705 197.435 ;
        RECT 54.875 197.145 55.145 197.605 ;
        RECT 54.420 196.755 55.375 196.975 ;
        RECT 52.005 195.825 52.755 196.345 ;
        RECT 28.090 195.055 33.435 195.600 ;
        RECT 33.610 195.055 38.955 195.600 ;
        RECT 39.130 195.055 44.475 195.600 ;
        RECT 44.650 195.055 49.995 195.600 ;
        RECT 50.165 195.055 50.455 195.780 ;
        RECT 51.085 195.055 52.755 195.825 ;
        RECT 52.985 195.055 53.195 195.875 ;
        RECT 53.365 195.855 53.615 196.455 ;
        RECT 53.785 196.045 54.115 196.295 ;
        RECT 54.305 196.025 54.995 196.585 ;
        RECT 53.365 195.225 53.695 195.855 ;
        RECT 53.865 195.055 54.095 195.875 ;
        RECT 55.165 195.855 55.375 196.755 ;
        RECT 54.420 195.685 55.375 195.855 ;
        RECT 55.545 196.585 55.945 197.435 ;
        RECT 56.135 196.975 56.415 197.435 ;
        RECT 56.935 197.145 57.260 197.605 ;
        RECT 56.135 196.755 57.260 196.975 ;
        RECT 55.545 196.025 56.640 196.585 ;
        RECT 56.810 196.295 57.260 196.755 ;
        RECT 57.430 196.465 57.815 197.435 ;
        RECT 57.990 197.170 63.335 197.605 ;
        RECT 63.510 197.170 68.855 197.605 ;
        RECT 54.420 195.225 54.705 195.685 ;
        RECT 54.875 195.055 55.145 195.515 ;
        RECT 55.545 195.225 55.945 196.025 ;
        RECT 56.810 195.965 57.365 196.295 ;
        RECT 56.810 195.855 57.260 195.965 ;
        RECT 56.135 195.685 57.260 195.855 ;
        RECT 57.535 195.795 57.815 196.465 ;
        RECT 59.580 195.920 59.930 197.170 ;
        RECT 56.135 195.225 56.415 195.685 ;
        RECT 56.935 195.055 57.260 195.515 ;
        RECT 57.430 195.225 57.815 195.795 ;
        RECT 61.410 195.600 61.750 196.430 ;
        RECT 65.100 195.920 65.450 197.170 ;
        RECT 69.025 196.735 69.300 197.435 ;
        RECT 69.470 197.060 69.725 197.605 ;
        RECT 69.895 197.095 70.375 197.435 ;
        RECT 70.550 197.050 71.155 197.605 ;
        RECT 70.540 196.950 71.155 197.050 ;
        RECT 70.540 196.925 70.725 196.950 ;
        RECT 66.930 195.600 67.270 196.430 ;
        RECT 69.025 195.705 69.195 196.735 ;
        RECT 69.470 196.605 70.225 196.855 ;
        RECT 70.395 196.680 70.725 196.925 ;
        RECT 69.470 196.570 70.240 196.605 ;
        RECT 69.470 196.560 70.255 196.570 ;
        RECT 69.365 196.545 70.260 196.560 ;
        RECT 69.365 196.530 70.280 196.545 ;
        RECT 69.365 196.520 70.300 196.530 ;
        RECT 69.365 196.510 70.325 196.520 ;
        RECT 69.365 196.480 70.395 196.510 ;
        RECT 69.365 196.450 70.415 196.480 ;
        RECT 69.365 196.420 70.435 196.450 ;
        RECT 69.365 196.395 70.465 196.420 ;
        RECT 69.365 196.360 70.500 196.395 ;
        RECT 69.365 196.355 70.530 196.360 ;
        RECT 69.365 195.960 69.595 196.355 ;
        RECT 70.140 196.350 70.530 196.355 ;
        RECT 70.165 196.340 70.530 196.350 ;
        RECT 70.180 196.335 70.530 196.340 ;
        RECT 70.195 196.330 70.530 196.335 ;
        RECT 70.895 196.330 71.155 196.780 ;
        RECT 70.195 196.325 71.155 196.330 ;
        RECT 70.205 196.315 71.155 196.325 ;
        RECT 70.215 196.310 71.155 196.315 ;
        RECT 70.225 196.300 71.155 196.310 ;
        RECT 70.230 196.290 71.155 196.300 ;
        RECT 70.235 196.285 71.155 196.290 ;
        RECT 70.245 196.270 71.155 196.285 ;
        RECT 70.250 196.255 71.155 196.270 ;
        RECT 70.260 196.230 71.155 196.255 ;
        RECT 69.765 195.760 70.095 196.185 ;
        RECT 57.990 195.055 63.335 195.600 ;
        RECT 63.510 195.055 68.855 195.600 ;
        RECT 69.025 195.225 69.285 195.705 ;
        RECT 69.455 195.055 69.705 195.595 ;
        RECT 69.875 195.275 70.095 195.760 ;
        RECT 70.265 196.160 71.155 196.230 ;
        RECT 71.335 196.545 71.665 197.395 ;
        RECT 70.265 195.435 70.435 196.160 ;
        RECT 70.605 195.605 71.155 195.990 ;
        RECT 71.335 195.780 71.525 196.545 ;
        RECT 71.835 196.465 72.085 197.605 ;
        RECT 72.275 196.965 72.525 197.385 ;
        RECT 72.755 197.135 73.085 197.605 ;
        RECT 73.315 196.965 73.565 197.385 ;
        RECT 72.275 196.795 73.565 196.965 ;
        RECT 73.745 196.965 74.075 197.395 ;
        RECT 73.745 196.795 74.200 196.965 ;
        RECT 72.265 196.295 72.480 196.625 ;
        RECT 71.695 195.965 72.005 196.295 ;
        RECT 72.175 195.965 72.480 196.295 ;
        RECT 72.655 195.965 72.940 196.625 ;
        RECT 73.135 195.965 73.400 196.625 ;
        RECT 73.615 195.965 73.860 196.625 ;
        RECT 71.835 195.795 72.005 195.965 ;
        RECT 74.030 195.795 74.200 196.795 ;
        RECT 74.545 196.515 75.755 197.605 ;
        RECT 74.545 195.975 75.065 196.515 ;
        RECT 75.925 196.440 76.215 197.605 ;
        RECT 76.385 196.515 79.895 197.605 ;
        RECT 80.070 197.170 85.415 197.605 ;
        RECT 75.235 195.805 75.755 196.345 ;
        RECT 76.385 195.995 78.075 196.515 ;
        RECT 78.245 195.825 79.895 196.345 ;
        RECT 81.660 195.920 82.010 197.170 ;
        RECT 85.960 196.625 86.215 197.295 ;
        RECT 86.395 196.805 86.680 197.605 ;
        RECT 86.860 196.885 87.190 197.395 ;
        RECT 70.265 195.265 71.155 195.435 ;
        RECT 71.335 195.270 71.665 195.780 ;
        RECT 71.835 195.625 74.200 195.795 ;
        RECT 71.835 195.055 72.165 195.455 ;
        RECT 73.215 195.285 73.545 195.625 ;
        RECT 73.715 195.055 74.045 195.455 ;
        RECT 74.545 195.055 75.755 195.805 ;
        RECT 75.925 195.055 76.215 195.780 ;
        RECT 76.385 195.055 79.895 195.825 ;
        RECT 83.490 195.600 83.830 196.430 ;
        RECT 85.960 195.765 86.140 196.625 ;
        RECT 86.860 196.295 87.110 196.885 ;
        RECT 87.460 196.735 87.630 197.345 ;
        RECT 87.800 196.915 88.130 197.605 ;
        RECT 88.360 197.055 88.600 197.345 ;
        RECT 88.800 197.225 89.220 197.605 ;
        RECT 89.400 197.135 90.030 197.385 ;
        RECT 90.500 197.225 90.830 197.605 ;
        RECT 89.400 197.055 89.570 197.135 ;
        RECT 91.000 197.055 91.170 197.345 ;
        RECT 91.350 197.225 91.730 197.605 ;
        RECT 91.970 197.220 92.800 197.390 ;
        RECT 88.360 196.885 89.570 197.055 ;
        RECT 86.310 195.965 87.110 196.295 ;
        RECT 80.070 195.055 85.415 195.600 ;
        RECT 85.960 195.565 86.215 195.765 ;
        RECT 85.875 195.395 86.215 195.565 ;
        RECT 85.960 195.235 86.215 195.395 ;
        RECT 86.395 195.055 86.680 195.515 ;
        RECT 86.860 195.315 87.110 195.965 ;
        RECT 87.310 196.715 87.630 196.735 ;
        RECT 87.310 196.545 89.230 196.715 ;
        RECT 87.310 195.650 87.500 196.545 ;
        RECT 89.400 196.375 89.570 196.885 ;
        RECT 89.740 196.625 90.260 196.935 ;
        RECT 87.670 196.205 89.570 196.375 ;
        RECT 87.670 196.145 88.000 196.205 ;
        RECT 88.150 195.975 88.480 196.035 ;
        RECT 87.820 195.705 88.480 195.975 ;
        RECT 87.310 195.320 87.630 195.650 ;
        RECT 87.810 195.055 88.470 195.535 ;
        RECT 88.670 195.445 88.840 196.205 ;
        RECT 89.740 196.035 89.920 196.445 ;
        RECT 89.010 195.865 89.340 195.985 ;
        RECT 90.090 195.865 90.260 196.625 ;
        RECT 89.010 195.695 90.260 195.865 ;
        RECT 90.430 196.805 91.800 197.055 ;
        RECT 90.430 196.035 90.620 196.805 ;
        RECT 91.550 196.545 91.800 196.805 ;
        RECT 90.790 196.375 91.040 196.535 ;
        RECT 91.970 196.375 92.140 197.220 ;
        RECT 93.035 196.935 93.205 197.435 ;
        RECT 93.375 197.105 93.705 197.605 ;
        RECT 92.310 196.545 92.810 196.925 ;
        RECT 93.035 196.765 93.730 196.935 ;
        RECT 90.790 196.205 92.140 196.375 ;
        RECT 91.720 196.165 92.140 196.205 ;
        RECT 90.430 195.695 90.850 196.035 ;
        RECT 91.140 195.705 91.550 196.035 ;
        RECT 88.670 195.275 89.520 195.445 ;
        RECT 90.080 195.055 90.400 195.515 ;
        RECT 90.600 195.265 90.850 195.695 ;
        RECT 91.140 195.055 91.550 195.495 ;
        RECT 91.720 195.435 91.890 196.165 ;
        RECT 92.060 195.615 92.410 195.985 ;
        RECT 92.590 195.675 92.810 196.545 ;
        RECT 92.980 195.975 93.390 196.595 ;
        RECT 93.560 195.795 93.730 196.765 ;
        RECT 93.035 195.605 93.730 195.795 ;
        RECT 91.720 195.235 92.735 195.435 ;
        RECT 93.035 195.275 93.205 195.605 ;
        RECT 93.375 195.055 93.705 195.435 ;
        RECT 93.920 195.315 94.145 197.435 ;
        RECT 94.315 197.105 94.645 197.605 ;
        RECT 94.815 196.935 94.985 197.435 ;
        RECT 94.320 196.765 94.985 196.935 ;
        RECT 94.320 195.775 94.550 196.765 ;
        RECT 94.720 195.945 95.070 196.595 ;
        RECT 95.245 196.515 97.835 197.605 ;
        RECT 98.120 196.975 98.405 197.435 ;
        RECT 98.575 197.145 98.845 197.605 ;
        RECT 98.120 196.755 99.075 196.975 ;
        RECT 95.245 195.995 96.455 196.515 ;
        RECT 96.625 195.825 97.835 196.345 ;
        RECT 98.005 196.025 98.695 196.585 ;
        RECT 98.865 195.855 99.075 196.755 ;
        RECT 94.320 195.605 94.985 195.775 ;
        RECT 94.315 195.055 94.645 195.435 ;
        RECT 94.815 195.315 94.985 195.605 ;
        RECT 95.245 195.055 97.835 195.825 ;
        RECT 98.120 195.685 99.075 195.855 ;
        RECT 99.245 196.585 99.645 197.435 ;
        RECT 99.835 196.975 100.115 197.435 ;
        RECT 100.635 197.145 100.960 197.605 ;
        RECT 99.835 196.755 100.960 196.975 ;
        RECT 99.245 196.025 100.340 196.585 ;
        RECT 100.510 196.295 100.960 196.755 ;
        RECT 101.130 196.465 101.515 197.435 ;
        RECT 98.120 195.225 98.405 195.685 ;
        RECT 98.575 195.055 98.845 195.515 ;
        RECT 99.245 195.225 99.645 196.025 ;
        RECT 100.510 195.965 101.065 196.295 ;
        RECT 100.510 195.855 100.960 195.965 ;
        RECT 99.835 195.685 100.960 195.855 ;
        RECT 101.235 195.795 101.515 196.465 ;
        RECT 101.685 196.440 101.975 197.605 ;
        RECT 102.145 196.515 104.735 197.605 ;
        RECT 104.910 197.170 110.255 197.605 ;
        RECT 102.145 195.995 103.355 196.515 ;
        RECT 103.525 195.825 104.735 196.345 ;
        RECT 106.500 195.920 106.850 197.170 ;
        RECT 99.835 195.225 100.115 195.685 ;
        RECT 100.635 195.055 100.960 195.515 ;
        RECT 101.130 195.225 101.515 195.795 ;
        RECT 101.685 195.055 101.975 195.780 ;
        RECT 102.145 195.055 104.735 195.825 ;
        RECT 108.330 195.600 108.670 196.430 ;
        RECT 110.430 196.415 110.685 197.295 ;
        RECT 110.855 196.465 111.160 197.605 ;
        RECT 111.500 197.225 111.830 197.605 ;
        RECT 112.010 197.055 112.180 197.345 ;
        RECT 112.350 197.145 112.600 197.605 ;
        RECT 111.380 196.885 112.180 197.055 ;
        RECT 112.770 197.095 113.640 197.435 ;
        RECT 110.430 195.765 110.640 196.415 ;
        RECT 111.380 196.295 111.550 196.885 ;
        RECT 112.770 196.715 112.940 197.095 ;
        RECT 113.875 196.975 114.045 197.435 ;
        RECT 114.215 197.145 114.585 197.605 ;
        RECT 114.880 197.005 115.050 197.345 ;
        RECT 115.220 197.175 115.550 197.605 ;
        RECT 115.785 197.005 115.955 197.345 ;
        RECT 111.720 196.545 112.940 196.715 ;
        RECT 113.110 196.635 113.570 196.925 ;
        RECT 113.875 196.805 114.435 196.975 ;
        RECT 114.880 196.835 115.955 197.005 ;
        RECT 116.125 197.105 116.805 197.435 ;
        RECT 117.020 197.105 117.270 197.435 ;
        RECT 117.440 197.145 117.690 197.605 ;
        RECT 114.265 196.665 114.435 196.805 ;
        RECT 113.110 196.625 114.075 196.635 ;
        RECT 112.770 196.455 112.940 196.545 ;
        RECT 113.400 196.465 114.075 196.625 ;
        RECT 110.810 196.265 111.550 196.295 ;
        RECT 110.810 195.965 111.725 196.265 ;
        RECT 111.400 195.790 111.725 195.965 ;
        RECT 104.910 195.055 110.255 195.600 ;
        RECT 110.430 195.235 110.685 195.765 ;
        RECT 110.855 195.055 111.160 195.515 ;
        RECT 111.405 195.435 111.725 195.790 ;
        RECT 111.895 196.005 112.435 196.375 ;
        RECT 112.770 196.285 113.175 196.455 ;
        RECT 111.895 195.605 112.135 196.005 ;
        RECT 112.615 195.835 112.835 196.115 ;
        RECT 112.305 195.665 112.835 195.835 ;
        RECT 112.305 195.435 112.475 195.665 ;
        RECT 113.005 195.505 113.175 196.285 ;
        RECT 113.345 195.675 113.695 196.295 ;
        RECT 113.865 195.675 114.075 196.465 ;
        RECT 114.265 196.495 115.765 196.665 ;
        RECT 114.265 195.805 114.435 196.495 ;
        RECT 116.125 196.325 116.295 197.105 ;
        RECT 117.100 196.975 117.270 197.105 ;
        RECT 114.605 196.155 116.295 196.325 ;
        RECT 116.465 196.545 116.930 196.935 ;
        RECT 117.100 196.805 117.495 196.975 ;
        RECT 114.605 195.975 114.775 196.155 ;
        RECT 111.405 195.265 112.475 195.435 ;
        RECT 112.645 195.055 112.835 195.495 ;
        RECT 113.005 195.225 113.955 195.505 ;
        RECT 114.265 195.415 114.525 195.805 ;
        RECT 114.945 195.735 115.735 195.985 ;
        RECT 114.175 195.245 114.525 195.415 ;
        RECT 114.735 195.055 115.065 195.515 ;
        RECT 115.940 195.445 116.110 196.155 ;
        RECT 116.465 195.955 116.635 196.545 ;
        RECT 116.280 195.735 116.635 195.955 ;
        RECT 116.805 195.735 117.155 196.355 ;
        RECT 117.325 195.445 117.495 196.805 ;
        RECT 117.860 196.635 118.185 197.420 ;
        RECT 117.665 195.585 118.125 196.635 ;
        RECT 115.940 195.275 116.795 195.445 ;
        RECT 117.000 195.275 117.495 195.445 ;
        RECT 117.665 195.055 117.995 195.415 ;
        RECT 118.355 195.315 118.525 197.435 ;
        RECT 118.695 197.105 119.025 197.605 ;
        RECT 119.195 196.935 119.450 197.435 ;
        RECT 118.700 196.765 119.450 196.935 ;
        RECT 118.700 195.775 118.930 196.765 ;
        RECT 119.100 195.945 119.450 196.595 ;
        RECT 119.625 196.515 120.835 197.605 ;
        RECT 121.010 197.170 126.355 197.605 ;
        RECT 119.625 195.975 120.145 196.515 ;
        RECT 120.315 195.805 120.835 196.345 ;
        RECT 122.600 195.920 122.950 197.170 ;
        RECT 126.525 196.515 127.735 197.605 ;
        RECT 118.700 195.605 119.450 195.775 ;
        RECT 118.695 195.055 119.025 195.435 ;
        RECT 119.195 195.315 119.450 195.605 ;
        RECT 119.625 195.055 120.835 195.805 ;
        RECT 124.430 195.600 124.770 196.430 ;
        RECT 126.525 195.975 127.045 196.515 ;
        RECT 127.215 195.805 127.735 196.345 ;
        RECT 121.010 195.055 126.355 195.600 ;
        RECT 126.525 195.055 127.735 195.805 ;
        RECT 14.660 194.885 127.820 195.055 ;
        RECT 14.745 194.135 15.955 194.885 ;
        RECT 14.745 193.595 15.265 194.135 ;
        RECT 17.045 194.115 20.555 194.885 ;
        RECT 20.730 194.340 26.075 194.885 ;
        RECT 26.250 194.340 31.595 194.885 ;
        RECT 31.770 194.340 37.115 194.885 ;
        RECT 15.435 193.425 15.955 193.965 ;
        RECT 14.745 192.335 15.955 193.425 ;
        RECT 17.045 193.425 18.735 193.945 ;
        RECT 18.905 193.595 20.555 194.115 ;
        RECT 17.045 192.335 20.555 193.425 ;
        RECT 22.320 192.770 22.670 194.020 ;
        RECT 24.150 193.510 24.490 194.340 ;
        RECT 27.840 192.770 28.190 194.020 ;
        RECT 29.670 193.510 30.010 194.340 ;
        RECT 33.360 192.770 33.710 194.020 ;
        RECT 35.190 193.510 35.530 194.340 ;
        RECT 37.285 194.160 37.575 194.885 ;
        RECT 38.665 194.115 42.175 194.885 ;
        RECT 42.350 194.340 47.695 194.885 ;
        RECT 20.730 192.335 26.075 192.770 ;
        RECT 26.250 192.335 31.595 192.770 ;
        RECT 31.770 192.335 37.115 192.770 ;
        RECT 37.285 192.335 37.575 193.500 ;
        RECT 38.665 193.425 40.355 193.945 ;
        RECT 40.525 193.595 42.175 194.115 ;
        RECT 38.665 192.335 42.175 193.425 ;
        RECT 43.940 192.770 44.290 194.020 ;
        RECT 45.770 193.510 46.110 194.340 ;
        RECT 47.925 194.065 48.135 194.885 ;
        RECT 48.305 194.085 48.635 194.715 ;
        RECT 48.305 193.485 48.555 194.085 ;
        RECT 48.805 194.065 49.035 194.885 ;
        RECT 49.250 194.335 49.505 194.625 ;
        RECT 49.675 194.505 50.005 194.885 ;
        RECT 49.250 194.165 50.000 194.335 ;
        RECT 48.725 193.645 49.055 193.895 ;
        RECT 42.350 192.335 47.695 192.770 ;
        RECT 47.925 192.335 48.135 193.475 ;
        RECT 48.305 192.505 48.635 193.485 ;
        RECT 48.805 192.335 49.035 193.475 ;
        RECT 49.250 193.345 49.600 193.995 ;
        RECT 49.770 193.175 50.000 194.165 ;
        RECT 49.250 193.005 50.000 193.175 ;
        RECT 49.250 192.505 49.505 193.005 ;
        RECT 49.675 192.335 50.005 192.835 ;
        RECT 50.175 192.505 50.345 194.625 ;
        RECT 50.705 194.525 51.035 194.885 ;
        RECT 51.205 194.495 51.700 194.665 ;
        RECT 51.905 194.495 52.760 194.665 ;
        RECT 50.575 193.305 51.035 194.355 ;
        RECT 50.515 192.520 50.840 193.305 ;
        RECT 51.205 193.135 51.375 194.495 ;
        RECT 51.545 193.585 51.895 194.205 ;
        RECT 52.065 193.985 52.420 194.205 ;
        RECT 52.065 193.395 52.235 193.985 ;
        RECT 52.590 193.785 52.760 194.495 ;
        RECT 53.635 194.425 53.965 194.885 ;
        RECT 54.175 194.525 54.525 194.695 ;
        RECT 52.965 193.955 53.755 194.205 ;
        RECT 54.175 194.135 54.435 194.525 ;
        RECT 54.745 194.435 55.695 194.715 ;
        RECT 55.865 194.445 56.055 194.885 ;
        RECT 56.225 194.505 57.295 194.675 ;
        RECT 53.925 193.785 54.095 193.965 ;
        RECT 51.205 192.965 51.600 193.135 ;
        RECT 51.770 193.005 52.235 193.395 ;
        RECT 52.405 193.615 54.095 193.785 ;
        RECT 51.430 192.835 51.600 192.965 ;
        RECT 52.405 192.835 52.575 193.615 ;
        RECT 54.265 193.445 54.435 194.135 ;
        RECT 52.935 193.275 54.435 193.445 ;
        RECT 54.625 193.475 54.835 194.265 ;
        RECT 55.005 193.645 55.355 194.265 ;
        RECT 55.525 193.655 55.695 194.435 ;
        RECT 56.225 194.275 56.395 194.505 ;
        RECT 55.865 194.105 56.395 194.275 ;
        RECT 55.865 193.825 56.085 194.105 ;
        RECT 56.565 193.935 56.805 194.335 ;
        RECT 55.525 193.485 55.930 193.655 ;
        RECT 56.265 193.565 56.805 193.935 ;
        RECT 56.975 194.150 57.295 194.505 ;
        RECT 57.540 194.425 57.845 194.885 ;
        RECT 58.015 194.175 58.270 194.705 ;
        RECT 56.975 193.975 57.300 194.150 ;
        RECT 56.975 193.675 57.890 193.975 ;
        RECT 57.150 193.645 57.890 193.675 ;
        RECT 54.625 193.315 55.300 193.475 ;
        RECT 55.760 193.395 55.930 193.485 ;
        RECT 54.625 193.305 55.590 193.315 ;
        RECT 54.265 193.135 54.435 193.275 ;
        RECT 51.010 192.335 51.260 192.795 ;
        RECT 51.430 192.505 51.680 192.835 ;
        RECT 51.895 192.505 52.575 192.835 ;
        RECT 52.745 192.935 53.820 193.105 ;
        RECT 54.265 192.965 54.825 193.135 ;
        RECT 55.130 193.015 55.590 193.305 ;
        RECT 55.760 193.225 56.980 193.395 ;
        RECT 52.745 192.595 52.915 192.935 ;
        RECT 53.150 192.335 53.480 192.765 ;
        RECT 53.650 192.595 53.820 192.935 ;
        RECT 54.115 192.335 54.485 192.795 ;
        RECT 54.655 192.505 54.825 192.965 ;
        RECT 55.760 192.845 55.930 193.225 ;
        RECT 57.150 193.055 57.320 193.645 ;
        RECT 58.060 193.525 58.270 194.175 ;
        RECT 59.365 194.115 62.875 194.885 ;
        RECT 63.045 194.160 63.335 194.885 ;
        RECT 63.505 194.115 65.175 194.885 ;
        RECT 55.060 192.505 55.930 192.845 ;
        RECT 56.520 192.885 57.320 193.055 ;
        RECT 56.100 192.335 56.350 192.795 ;
        RECT 56.520 192.595 56.690 192.885 ;
        RECT 56.870 192.335 57.200 192.715 ;
        RECT 57.540 192.335 57.845 193.475 ;
        RECT 58.015 192.645 58.270 193.525 ;
        RECT 59.365 193.425 61.055 193.945 ;
        RECT 61.225 193.595 62.875 194.115 ;
        RECT 59.365 192.335 62.875 193.425 ;
        RECT 63.045 192.335 63.335 193.500 ;
        RECT 63.505 193.425 64.255 193.945 ;
        RECT 64.425 193.595 65.175 194.115 ;
        RECT 65.405 194.065 65.615 194.885 ;
        RECT 65.785 194.085 66.115 194.715 ;
        RECT 65.785 193.485 66.035 194.085 ;
        RECT 66.285 194.065 66.515 194.885 ;
        RECT 67.185 194.115 68.855 194.885 ;
        RECT 66.205 193.645 66.535 193.895 ;
        RECT 63.505 192.335 65.175 193.425 ;
        RECT 65.405 192.335 65.615 193.475 ;
        RECT 65.785 192.505 66.115 193.485 ;
        RECT 66.285 192.335 66.515 193.475 ;
        RECT 67.185 193.425 67.935 193.945 ;
        RECT 68.105 193.595 68.855 194.115 ;
        RECT 69.025 194.065 69.285 194.885 ;
        RECT 69.455 194.065 69.785 194.485 ;
        RECT 69.965 194.315 70.225 194.715 ;
        RECT 70.395 194.485 70.725 194.885 ;
        RECT 70.895 194.315 71.065 194.665 ;
        RECT 71.235 194.485 71.610 194.885 ;
        RECT 69.965 194.145 71.630 194.315 ;
        RECT 71.800 194.210 72.075 194.555 ;
        RECT 69.535 193.975 69.785 194.065 ;
        RECT 71.460 193.975 71.630 194.145 ;
        RECT 69.030 193.645 69.365 193.895 ;
        RECT 69.535 193.645 70.250 193.975 ;
        RECT 70.465 193.645 71.290 193.975 ;
        RECT 71.460 193.645 71.735 193.975 ;
        RECT 67.185 192.335 68.855 193.425 ;
        RECT 69.025 192.335 69.285 193.475 ;
        RECT 69.535 193.085 69.705 193.645 ;
        RECT 69.965 193.185 70.295 193.475 ;
        RECT 70.465 193.355 70.710 193.645 ;
        RECT 71.460 193.475 71.630 193.645 ;
        RECT 71.905 193.475 72.075 194.210 ;
        RECT 70.970 193.305 71.630 193.475 ;
        RECT 70.970 193.185 71.140 193.305 ;
        RECT 69.965 193.015 71.140 193.185 ;
        RECT 69.525 192.515 71.140 192.845 ;
        RECT 71.310 192.335 71.590 193.135 ;
        RECT 71.800 192.505 72.075 193.475 ;
        RECT 72.245 194.210 72.520 194.555 ;
        RECT 72.710 194.485 73.085 194.885 ;
        RECT 73.255 194.315 73.425 194.665 ;
        RECT 73.595 194.485 73.925 194.885 ;
        RECT 74.095 194.315 74.355 194.715 ;
        RECT 72.245 193.475 72.415 194.210 ;
        RECT 72.690 194.145 74.355 194.315 ;
        RECT 72.690 193.975 72.860 194.145 ;
        RECT 74.535 194.065 74.865 194.485 ;
        RECT 75.035 194.065 75.295 194.885 ;
        RECT 75.465 194.115 78.975 194.885 ;
        RECT 79.150 194.340 84.495 194.885 ;
        RECT 74.535 193.975 74.785 194.065 ;
        RECT 72.585 193.645 72.860 193.975 ;
        RECT 73.030 193.645 73.855 193.975 ;
        RECT 74.070 193.645 74.785 193.975 ;
        RECT 74.955 193.645 75.290 193.895 ;
        RECT 72.690 193.475 72.860 193.645 ;
        RECT 72.245 192.505 72.520 193.475 ;
        RECT 72.690 193.305 73.350 193.475 ;
        RECT 73.610 193.355 73.855 193.645 ;
        RECT 73.180 193.185 73.350 193.305 ;
        RECT 74.025 193.185 74.355 193.475 ;
        RECT 72.730 192.335 73.010 193.135 ;
        RECT 73.180 193.015 74.355 193.185 ;
        RECT 74.615 193.085 74.785 193.645 ;
        RECT 73.180 192.515 74.795 192.845 ;
        RECT 75.035 192.335 75.295 193.475 ;
        RECT 75.465 193.425 77.155 193.945 ;
        RECT 77.325 193.595 78.975 194.115 ;
        RECT 75.465 192.335 78.975 193.425 ;
        RECT 80.740 192.770 81.090 194.020 ;
        RECT 82.570 193.510 82.910 194.340 ;
        RECT 84.940 194.075 85.185 194.680 ;
        RECT 85.405 194.350 85.915 194.885 ;
        RECT 84.665 193.905 85.895 194.075 ;
        RECT 84.665 193.095 85.005 193.905 ;
        RECT 85.175 193.340 85.925 193.530 ;
        RECT 79.150 192.335 84.495 192.770 ;
        RECT 84.665 192.685 85.180 193.095 ;
        RECT 85.415 192.335 85.585 193.095 ;
        RECT 85.755 192.675 85.925 193.340 ;
        RECT 86.095 193.355 86.285 194.715 ;
        RECT 86.455 193.865 86.730 194.715 ;
        RECT 86.920 194.350 87.450 194.715 ;
        RECT 87.875 194.485 88.205 194.885 ;
        RECT 87.275 194.315 87.450 194.350 ;
        RECT 86.455 193.695 86.735 193.865 ;
        RECT 86.455 193.555 86.730 193.695 ;
        RECT 86.935 193.355 87.105 194.155 ;
        RECT 86.095 193.185 87.105 193.355 ;
        RECT 87.275 194.145 88.205 194.315 ;
        RECT 88.375 194.145 88.630 194.715 ;
        RECT 88.805 194.160 89.095 194.885 ;
        RECT 87.275 193.015 87.445 194.145 ;
        RECT 88.035 193.975 88.205 194.145 ;
        RECT 86.320 192.845 87.445 193.015 ;
        RECT 87.615 193.645 87.810 193.975 ;
        RECT 88.035 193.645 88.290 193.975 ;
        RECT 87.615 192.675 87.785 193.645 ;
        RECT 88.460 193.475 88.630 194.145 ;
        RECT 89.325 194.065 89.535 194.885 ;
        RECT 89.705 194.085 90.035 194.715 ;
        RECT 85.755 192.505 87.785 192.675 ;
        RECT 87.955 192.335 88.125 193.475 ;
        RECT 88.295 192.505 88.630 193.475 ;
        RECT 88.805 192.335 89.095 193.500 ;
        RECT 89.705 193.485 89.955 194.085 ;
        RECT 90.205 194.065 90.435 194.885 ;
        RECT 90.645 194.115 93.235 194.885 ;
        RECT 90.125 193.645 90.455 193.895 ;
        RECT 89.325 192.335 89.535 193.475 ;
        RECT 89.705 192.505 90.035 193.485 ;
        RECT 90.205 192.335 90.435 193.475 ;
        RECT 90.645 193.425 91.855 193.945 ;
        RECT 92.025 193.595 93.235 194.115 ;
        RECT 93.445 194.065 93.675 194.885 ;
        RECT 93.845 194.085 94.175 194.715 ;
        RECT 93.425 193.645 93.755 193.895 ;
        RECT 93.925 193.485 94.175 194.085 ;
        RECT 94.345 194.065 94.555 194.885 ;
        RECT 94.785 194.375 95.090 194.885 ;
        RECT 94.785 193.645 95.100 194.205 ;
        RECT 95.270 193.895 95.520 194.705 ;
        RECT 95.690 194.360 95.950 194.885 ;
        RECT 96.130 193.895 96.380 194.705 ;
        RECT 96.550 194.325 96.810 194.885 ;
        RECT 96.980 194.235 97.240 194.690 ;
        RECT 97.410 194.405 97.670 194.885 ;
        RECT 97.840 194.235 98.100 194.690 ;
        RECT 98.270 194.405 98.530 194.885 ;
        RECT 98.700 194.235 98.960 194.690 ;
        RECT 99.130 194.405 99.375 194.885 ;
        RECT 99.545 194.235 99.820 194.690 ;
        RECT 99.990 194.405 100.235 194.885 ;
        RECT 100.405 194.235 100.665 194.690 ;
        RECT 100.845 194.405 101.095 194.885 ;
        RECT 101.265 194.235 101.525 194.690 ;
        RECT 101.705 194.405 101.955 194.885 ;
        RECT 102.125 194.235 102.385 194.690 ;
        RECT 102.565 194.405 102.825 194.885 ;
        RECT 102.995 194.235 103.255 194.690 ;
        RECT 103.425 194.405 103.725 194.885 ;
        RECT 96.980 194.205 103.725 194.235 ;
        RECT 96.980 194.065 103.755 194.205 ;
        RECT 103.985 194.135 105.195 194.885 ;
        RECT 102.560 194.035 103.755 194.065 ;
        RECT 95.270 193.645 102.390 193.895 ;
        RECT 90.645 192.335 93.235 193.425 ;
        RECT 93.445 192.335 93.675 193.475 ;
        RECT 93.845 192.505 94.175 193.485 ;
        RECT 94.345 192.335 94.555 193.475 ;
        RECT 94.795 192.335 95.090 193.145 ;
        RECT 95.270 192.505 95.515 193.645 ;
        RECT 95.690 192.335 95.950 193.145 ;
        RECT 96.130 192.510 96.380 193.645 ;
        RECT 102.560 193.475 103.725 194.035 ;
        RECT 96.980 193.250 103.725 193.475 ;
        RECT 103.985 193.425 104.505 193.965 ;
        RECT 104.675 193.595 105.195 194.135 ;
        RECT 105.365 194.115 108.875 194.885 ;
        RECT 105.365 193.425 107.055 193.945 ;
        RECT 107.225 193.595 108.875 194.115 ;
        RECT 109.085 194.065 109.315 194.885 ;
        RECT 109.485 194.085 109.815 194.715 ;
        RECT 109.065 193.645 109.395 193.895 ;
        RECT 109.565 193.485 109.815 194.085 ;
        RECT 109.985 194.065 110.195 194.885 ;
        RECT 110.700 194.075 110.945 194.680 ;
        RECT 111.165 194.350 111.675 194.885 ;
        RECT 96.980 193.235 102.385 193.250 ;
        RECT 96.550 192.340 96.810 193.135 ;
        RECT 96.980 192.510 97.240 193.235 ;
        RECT 97.410 192.340 97.670 193.065 ;
        RECT 97.840 192.510 98.100 193.235 ;
        RECT 98.270 192.340 98.530 193.065 ;
        RECT 98.700 192.510 98.960 193.235 ;
        RECT 99.130 192.340 99.390 193.065 ;
        RECT 99.560 192.510 99.820 193.235 ;
        RECT 99.990 192.340 100.235 193.065 ;
        RECT 100.405 192.510 100.665 193.235 ;
        RECT 100.850 192.340 101.095 193.065 ;
        RECT 101.265 192.510 101.525 193.235 ;
        RECT 101.710 192.340 101.955 193.065 ;
        RECT 102.125 192.510 102.385 193.235 ;
        RECT 102.570 192.340 102.825 193.065 ;
        RECT 102.995 192.510 103.285 193.250 ;
        RECT 96.550 192.335 102.825 192.340 ;
        RECT 103.455 192.335 103.725 193.080 ;
        RECT 103.985 192.335 105.195 193.425 ;
        RECT 105.365 192.335 108.875 193.425 ;
        RECT 109.085 192.335 109.315 193.475 ;
        RECT 109.485 192.505 109.815 193.485 ;
        RECT 110.425 193.905 111.655 194.075 ;
        RECT 109.985 192.335 110.195 193.475 ;
        RECT 110.425 193.095 110.765 193.905 ;
        RECT 110.935 193.340 111.685 193.530 ;
        RECT 110.425 192.685 110.940 193.095 ;
        RECT 111.175 192.335 111.345 193.095 ;
        RECT 111.515 192.675 111.685 193.340 ;
        RECT 111.855 193.355 112.045 194.715 ;
        RECT 112.215 194.545 112.490 194.715 ;
        RECT 112.215 194.375 112.495 194.545 ;
        RECT 112.215 193.555 112.490 194.375 ;
        RECT 112.680 194.350 113.210 194.715 ;
        RECT 113.635 194.485 113.965 194.885 ;
        RECT 113.035 194.315 113.210 194.350 ;
        RECT 112.695 193.355 112.865 194.155 ;
        RECT 111.855 193.185 112.865 193.355 ;
        RECT 113.035 194.145 113.965 194.315 ;
        RECT 114.135 194.145 114.390 194.715 ;
        RECT 114.565 194.160 114.855 194.885 ;
        RECT 113.035 193.015 113.205 194.145 ;
        RECT 113.795 193.975 113.965 194.145 ;
        RECT 112.080 192.845 113.205 193.015 ;
        RECT 113.375 193.645 113.570 193.975 ;
        RECT 113.795 193.645 114.050 193.975 ;
        RECT 113.375 192.675 113.545 193.645 ;
        RECT 114.220 193.475 114.390 194.145 ;
        RECT 115.085 194.065 115.295 194.885 ;
        RECT 115.465 194.085 115.795 194.715 ;
        RECT 111.515 192.505 113.545 192.675 ;
        RECT 113.715 192.335 113.885 193.475 ;
        RECT 114.055 192.505 114.390 193.475 ;
        RECT 114.565 192.335 114.855 193.500 ;
        RECT 115.465 193.485 115.715 194.085 ;
        RECT 115.965 194.065 116.195 194.885 ;
        RECT 117.325 194.115 120.835 194.885 ;
        RECT 121.010 194.340 126.355 194.885 ;
        RECT 115.885 193.645 116.215 193.895 ;
        RECT 115.085 192.335 115.295 193.475 ;
        RECT 115.465 192.505 115.795 193.485 ;
        RECT 115.965 192.335 116.195 193.475 ;
        RECT 117.325 193.425 119.015 193.945 ;
        RECT 119.185 193.595 120.835 194.115 ;
        RECT 117.325 192.335 120.835 193.425 ;
        RECT 122.600 192.770 122.950 194.020 ;
        RECT 124.430 193.510 124.770 194.340 ;
        RECT 126.525 194.135 127.735 194.885 ;
        RECT 126.525 193.425 127.045 193.965 ;
        RECT 127.215 193.595 127.735 194.135 ;
        RECT 121.010 192.335 126.355 192.770 ;
        RECT 126.525 192.335 127.735 193.425 ;
        RECT 14.660 192.165 127.820 192.335 ;
        RECT 14.745 191.075 15.955 192.165 ;
        RECT 14.745 190.365 15.265 190.905 ;
        RECT 15.435 190.535 15.955 191.075 ;
        RECT 16.125 191.075 18.715 192.165 ;
        RECT 18.890 191.730 24.235 192.165 ;
        RECT 16.125 190.555 17.335 191.075 ;
        RECT 17.505 190.385 18.715 190.905 ;
        RECT 20.480 190.480 20.830 191.730 ;
        RECT 24.405 191.000 24.695 192.165 ;
        RECT 25.330 191.730 30.675 192.165 ;
        RECT 30.850 191.730 36.195 192.165 ;
        RECT 14.745 189.615 15.955 190.365 ;
        RECT 16.125 189.615 18.715 190.385 ;
        RECT 22.310 190.160 22.650 190.990 ;
        RECT 26.920 190.480 27.270 191.730 ;
        RECT 18.890 189.615 24.235 190.160 ;
        RECT 24.405 189.615 24.695 190.340 ;
        RECT 28.750 190.160 29.090 190.990 ;
        RECT 32.440 190.480 32.790 191.730 ;
        RECT 36.740 191.185 36.995 191.855 ;
        RECT 37.175 191.365 37.460 192.165 ;
        RECT 37.640 191.445 37.970 191.955 ;
        RECT 36.740 191.145 36.920 191.185 ;
        RECT 34.270 190.160 34.610 190.990 ;
        RECT 36.655 190.975 36.920 191.145 ;
        RECT 36.740 190.325 36.920 190.975 ;
        RECT 37.640 190.855 37.890 191.445 ;
        RECT 38.240 191.295 38.410 191.905 ;
        RECT 38.580 191.475 38.910 192.165 ;
        RECT 39.140 191.615 39.380 191.905 ;
        RECT 39.580 191.785 40.000 192.165 ;
        RECT 40.180 191.695 40.810 191.945 ;
        RECT 41.280 191.785 41.610 192.165 ;
        RECT 40.180 191.615 40.350 191.695 ;
        RECT 41.780 191.615 41.950 191.905 ;
        RECT 42.130 191.785 42.510 192.165 ;
        RECT 42.750 191.780 43.580 191.950 ;
        RECT 39.140 191.445 40.350 191.615 ;
        RECT 37.090 190.525 37.890 190.855 ;
        RECT 25.330 189.615 30.675 190.160 ;
        RECT 30.850 189.615 36.195 190.160 ;
        RECT 36.740 189.795 36.995 190.325 ;
        RECT 37.175 189.615 37.460 190.075 ;
        RECT 37.640 189.875 37.890 190.525 ;
        RECT 38.090 191.275 38.410 191.295 ;
        RECT 38.090 191.105 40.010 191.275 ;
        RECT 38.090 190.210 38.280 191.105 ;
        RECT 40.180 190.935 40.350 191.445 ;
        RECT 40.520 191.185 41.040 191.495 ;
        RECT 38.450 190.765 40.350 190.935 ;
        RECT 38.450 190.705 38.780 190.765 ;
        RECT 38.930 190.535 39.260 190.595 ;
        RECT 38.600 190.265 39.260 190.535 ;
        RECT 38.090 189.880 38.410 190.210 ;
        RECT 38.590 189.615 39.250 190.095 ;
        RECT 39.450 190.005 39.620 190.765 ;
        RECT 40.520 190.595 40.700 191.005 ;
        RECT 39.790 190.425 40.120 190.545 ;
        RECT 40.870 190.425 41.040 191.185 ;
        RECT 39.790 190.255 41.040 190.425 ;
        RECT 41.210 191.365 42.580 191.615 ;
        RECT 41.210 190.595 41.400 191.365 ;
        RECT 42.330 191.105 42.580 191.365 ;
        RECT 41.570 190.935 41.820 191.095 ;
        RECT 42.750 190.935 42.920 191.780 ;
        RECT 43.815 191.495 43.985 191.995 ;
        RECT 44.155 191.665 44.485 192.165 ;
        RECT 43.090 191.105 43.590 191.485 ;
        RECT 43.815 191.325 44.510 191.495 ;
        RECT 41.570 190.765 42.920 190.935 ;
        RECT 42.500 190.725 42.920 190.765 ;
        RECT 41.210 190.255 41.630 190.595 ;
        RECT 41.920 190.265 42.330 190.595 ;
        RECT 39.450 189.835 40.300 190.005 ;
        RECT 40.860 189.615 41.180 190.075 ;
        RECT 41.380 189.825 41.630 190.255 ;
        RECT 41.920 189.615 42.330 190.055 ;
        RECT 42.500 189.995 42.670 190.725 ;
        RECT 42.840 190.175 43.190 190.545 ;
        RECT 43.370 190.235 43.590 191.105 ;
        RECT 43.760 190.535 44.170 191.155 ;
        RECT 44.340 190.355 44.510 191.325 ;
        RECT 43.815 190.165 44.510 190.355 ;
        RECT 42.500 189.795 43.515 189.995 ;
        RECT 43.815 189.835 43.985 190.165 ;
        RECT 44.155 189.615 44.485 189.995 ;
        RECT 44.700 189.875 44.925 191.995 ;
        RECT 45.095 191.665 45.425 192.165 ;
        RECT 45.595 191.495 45.765 191.995 ;
        RECT 45.100 191.325 45.765 191.495 ;
        RECT 46.025 191.405 46.540 191.815 ;
        RECT 46.775 191.405 46.945 192.165 ;
        RECT 47.115 191.825 49.145 191.995 ;
        RECT 45.100 190.335 45.330 191.325 ;
        RECT 45.500 190.505 45.850 191.155 ;
        RECT 46.025 190.595 46.365 191.405 ;
        RECT 47.115 191.160 47.285 191.825 ;
        RECT 47.680 191.485 48.805 191.655 ;
        RECT 46.535 190.970 47.285 191.160 ;
        RECT 47.455 191.145 48.465 191.315 ;
        RECT 46.025 190.425 47.255 190.595 ;
        RECT 45.100 190.165 45.765 190.335 ;
        RECT 45.095 189.615 45.425 189.995 ;
        RECT 45.595 189.875 45.765 190.165 ;
        RECT 46.300 189.820 46.545 190.425 ;
        RECT 46.765 189.615 47.275 190.150 ;
        RECT 47.455 189.785 47.645 191.145 ;
        RECT 47.815 190.805 48.090 190.945 ;
        RECT 47.815 190.635 48.095 190.805 ;
        RECT 47.815 189.785 48.090 190.635 ;
        RECT 48.295 190.345 48.465 191.145 ;
        RECT 48.635 190.355 48.805 191.485 ;
        RECT 48.975 190.855 49.145 191.825 ;
        RECT 49.315 191.025 49.485 192.165 ;
        RECT 49.655 191.025 49.990 191.995 ;
        RECT 48.975 190.525 49.170 190.855 ;
        RECT 49.395 190.525 49.650 190.855 ;
        RECT 49.395 190.355 49.565 190.525 ;
        RECT 49.820 190.355 49.990 191.025 ;
        RECT 50.165 191.000 50.455 192.165 ;
        RECT 51.085 191.090 51.355 191.995 ;
        RECT 51.525 191.405 51.855 192.165 ;
        RECT 52.035 191.235 52.205 191.995 ;
        RECT 48.635 190.185 49.565 190.355 ;
        RECT 48.635 190.150 48.810 190.185 ;
        RECT 48.280 189.785 48.810 190.150 ;
        RECT 49.235 189.615 49.565 190.015 ;
        RECT 49.735 189.785 49.990 190.355 ;
        RECT 50.165 189.615 50.455 190.340 ;
        RECT 51.085 190.290 51.255 191.090 ;
        RECT 51.540 191.065 52.205 191.235 ;
        RECT 51.540 190.920 51.710 191.065 ;
        RECT 51.425 190.590 51.710 190.920 ;
        RECT 52.470 190.975 52.725 191.855 ;
        RECT 52.895 191.025 53.200 192.165 ;
        RECT 53.540 191.785 53.870 192.165 ;
        RECT 54.050 191.615 54.220 191.905 ;
        RECT 54.390 191.705 54.640 192.165 ;
        RECT 53.420 191.445 54.220 191.615 ;
        RECT 54.810 191.655 55.680 191.995 ;
        RECT 51.540 190.335 51.710 190.590 ;
        RECT 51.945 190.515 52.275 190.885 ;
        RECT 51.085 189.785 51.345 190.290 ;
        RECT 51.540 190.165 52.205 190.335 ;
        RECT 51.525 189.615 51.855 189.995 ;
        RECT 52.035 189.785 52.205 190.165 ;
        RECT 52.470 190.325 52.680 190.975 ;
        RECT 53.420 190.855 53.590 191.445 ;
        RECT 54.810 191.275 54.980 191.655 ;
        RECT 55.915 191.535 56.085 191.995 ;
        RECT 56.255 191.705 56.625 192.165 ;
        RECT 56.920 191.565 57.090 191.905 ;
        RECT 57.260 191.735 57.590 192.165 ;
        RECT 57.825 191.565 57.995 191.905 ;
        RECT 53.760 191.105 54.980 191.275 ;
        RECT 55.150 191.195 55.610 191.485 ;
        RECT 55.915 191.365 56.475 191.535 ;
        RECT 56.920 191.395 57.995 191.565 ;
        RECT 58.165 191.665 58.845 191.995 ;
        RECT 59.060 191.665 59.310 191.995 ;
        RECT 59.480 191.705 59.730 192.165 ;
        RECT 56.305 191.225 56.475 191.365 ;
        RECT 55.150 191.185 56.115 191.195 ;
        RECT 54.810 191.015 54.980 191.105 ;
        RECT 55.440 191.025 56.115 191.185 ;
        RECT 52.850 190.825 53.590 190.855 ;
        RECT 52.850 190.525 53.765 190.825 ;
        RECT 53.440 190.350 53.765 190.525 ;
        RECT 52.470 189.795 52.725 190.325 ;
        RECT 52.895 189.615 53.200 190.075 ;
        RECT 53.445 189.995 53.765 190.350 ;
        RECT 53.935 190.565 54.475 190.935 ;
        RECT 54.810 190.845 55.215 191.015 ;
        RECT 53.935 190.165 54.175 190.565 ;
        RECT 54.655 190.395 54.875 190.675 ;
        RECT 54.345 190.225 54.875 190.395 ;
        RECT 54.345 189.995 54.515 190.225 ;
        RECT 55.045 190.065 55.215 190.845 ;
        RECT 55.385 190.235 55.735 190.855 ;
        RECT 55.905 190.235 56.115 191.025 ;
        RECT 56.305 191.055 57.805 191.225 ;
        RECT 56.305 190.365 56.475 191.055 ;
        RECT 58.165 190.885 58.335 191.665 ;
        RECT 59.140 191.535 59.310 191.665 ;
        RECT 56.645 190.715 58.335 190.885 ;
        RECT 58.505 191.105 58.970 191.495 ;
        RECT 59.140 191.365 59.535 191.535 ;
        RECT 56.645 190.535 56.815 190.715 ;
        RECT 53.445 189.825 54.515 189.995 ;
        RECT 54.685 189.615 54.875 190.055 ;
        RECT 55.045 189.785 55.995 190.065 ;
        RECT 56.305 189.975 56.565 190.365 ;
        RECT 56.985 190.295 57.775 190.545 ;
        RECT 56.215 189.805 56.565 189.975 ;
        RECT 56.775 189.615 57.105 190.075 ;
        RECT 57.980 190.005 58.150 190.715 ;
        RECT 58.505 190.515 58.675 191.105 ;
        RECT 58.320 190.295 58.675 190.515 ;
        RECT 58.845 190.295 59.195 190.915 ;
        RECT 59.365 190.005 59.535 191.365 ;
        RECT 59.900 191.195 60.225 191.980 ;
        RECT 59.705 190.145 60.165 191.195 ;
        RECT 57.980 189.835 58.835 190.005 ;
        RECT 59.040 189.835 59.535 190.005 ;
        RECT 59.705 189.615 60.035 189.975 ;
        RECT 60.395 189.875 60.565 191.995 ;
        RECT 60.735 191.665 61.065 192.165 ;
        RECT 61.235 191.495 61.490 191.995 ;
        RECT 60.740 191.325 61.490 191.495 ;
        RECT 60.740 190.335 60.970 191.325 ;
        RECT 61.140 190.505 61.490 191.155 ;
        RECT 61.715 191.025 61.965 192.165 ;
        RECT 62.135 190.975 62.385 191.855 ;
        RECT 62.555 191.025 62.860 192.165 ;
        RECT 63.200 191.785 63.530 192.165 ;
        RECT 63.710 191.615 63.880 191.905 ;
        RECT 64.050 191.705 64.300 192.165 ;
        RECT 63.080 191.445 63.880 191.615 ;
        RECT 64.470 191.655 65.340 191.995 ;
        RECT 60.740 190.165 61.490 190.335 ;
        RECT 60.735 189.615 61.065 189.995 ;
        RECT 61.235 189.875 61.490 190.165 ;
        RECT 61.715 189.615 61.965 190.370 ;
        RECT 62.135 190.325 62.340 190.975 ;
        RECT 63.080 190.855 63.250 191.445 ;
        RECT 64.470 191.275 64.640 191.655 ;
        RECT 65.575 191.535 65.745 191.995 ;
        RECT 65.915 191.705 66.285 192.165 ;
        RECT 66.580 191.565 66.750 191.905 ;
        RECT 66.920 191.735 67.250 192.165 ;
        RECT 67.485 191.565 67.655 191.905 ;
        RECT 63.420 191.105 64.640 191.275 ;
        RECT 64.810 191.195 65.270 191.485 ;
        RECT 65.575 191.365 66.135 191.535 ;
        RECT 66.580 191.395 67.655 191.565 ;
        RECT 67.825 191.665 68.505 191.995 ;
        RECT 68.720 191.665 68.970 191.995 ;
        RECT 69.140 191.705 69.390 192.165 ;
        RECT 65.965 191.225 66.135 191.365 ;
        RECT 64.810 191.185 65.775 191.195 ;
        RECT 64.470 191.015 64.640 191.105 ;
        RECT 65.100 191.025 65.775 191.185 ;
        RECT 62.510 190.825 63.250 190.855 ;
        RECT 62.510 190.525 63.425 190.825 ;
        RECT 63.100 190.350 63.425 190.525 ;
        RECT 62.135 189.795 62.385 190.325 ;
        RECT 62.555 189.615 62.860 190.075 ;
        RECT 63.105 189.995 63.425 190.350 ;
        RECT 63.595 190.565 64.135 190.935 ;
        RECT 64.470 190.845 64.875 191.015 ;
        RECT 63.595 190.165 63.835 190.565 ;
        RECT 64.315 190.395 64.535 190.675 ;
        RECT 64.005 190.225 64.535 190.395 ;
        RECT 64.005 189.995 64.175 190.225 ;
        RECT 64.705 190.065 64.875 190.845 ;
        RECT 65.045 190.235 65.395 190.855 ;
        RECT 65.565 190.235 65.775 191.025 ;
        RECT 65.965 191.055 67.465 191.225 ;
        RECT 65.965 190.365 66.135 191.055 ;
        RECT 67.825 190.885 67.995 191.665 ;
        RECT 68.800 191.535 68.970 191.665 ;
        RECT 66.305 190.715 67.995 190.885 ;
        RECT 68.165 191.105 68.630 191.495 ;
        RECT 68.800 191.365 69.195 191.535 ;
        RECT 66.305 190.535 66.475 190.715 ;
        RECT 63.105 189.825 64.175 189.995 ;
        RECT 64.345 189.615 64.535 190.055 ;
        RECT 64.705 189.785 65.655 190.065 ;
        RECT 65.965 189.975 66.225 190.365 ;
        RECT 66.645 190.295 67.435 190.545 ;
        RECT 65.875 189.805 66.225 189.975 ;
        RECT 66.435 189.615 66.765 190.075 ;
        RECT 67.640 190.005 67.810 190.715 ;
        RECT 68.165 190.515 68.335 191.105 ;
        RECT 67.980 190.295 68.335 190.515 ;
        RECT 68.505 190.295 68.855 190.915 ;
        RECT 69.025 190.005 69.195 191.365 ;
        RECT 69.560 191.195 69.885 191.980 ;
        RECT 69.365 190.145 69.825 191.195 ;
        RECT 67.640 189.835 68.495 190.005 ;
        RECT 68.700 189.835 69.195 190.005 ;
        RECT 69.365 189.615 69.695 189.975 ;
        RECT 70.055 189.875 70.225 191.995 ;
        RECT 70.395 191.665 70.725 192.165 ;
        RECT 70.895 191.495 71.150 191.995 ;
        RECT 71.345 191.655 71.645 192.165 ;
        RECT 71.815 191.655 72.195 191.825 ;
        RECT 72.775 191.655 73.405 192.165 ;
        RECT 70.400 191.325 71.150 191.495 ;
        RECT 71.815 191.485 71.985 191.655 ;
        RECT 73.575 191.485 73.905 191.995 ;
        RECT 74.075 191.655 74.375 192.165 ;
        RECT 70.400 190.335 70.630 191.325 ;
        RECT 71.325 191.285 71.985 191.485 ;
        RECT 72.155 191.315 74.375 191.485 ;
        RECT 70.800 190.505 71.150 191.155 ;
        RECT 71.325 190.355 71.495 191.285 ;
        RECT 72.155 191.115 72.325 191.315 ;
        RECT 71.665 190.945 72.325 191.115 ;
        RECT 72.495 190.975 74.035 191.145 ;
        RECT 71.665 190.525 71.835 190.945 ;
        RECT 72.495 190.775 72.665 190.975 ;
        RECT 72.065 190.605 72.665 190.775 ;
        RECT 72.835 190.605 73.530 190.805 ;
        RECT 73.790 190.525 74.035 190.975 ;
        RECT 72.155 190.355 73.065 190.435 ;
        RECT 70.400 190.165 71.150 190.335 ;
        RECT 70.395 189.615 70.725 189.995 ;
        RECT 70.895 189.875 71.150 190.165 ;
        RECT 71.325 189.875 71.645 190.355 ;
        RECT 71.815 190.265 73.065 190.355 ;
        RECT 71.815 190.185 72.325 190.265 ;
        RECT 71.815 189.785 72.045 190.185 ;
        RECT 72.215 189.615 72.565 190.005 ;
        RECT 72.735 189.785 73.065 190.265 ;
        RECT 73.235 189.615 73.405 190.435 ;
        RECT 74.205 190.355 74.375 191.315 ;
        RECT 74.545 191.075 75.755 192.165 ;
        RECT 74.545 190.535 75.065 191.075 ;
        RECT 75.925 191.000 76.215 192.165 ;
        RECT 76.385 191.025 76.645 192.165 ;
        RECT 76.815 191.195 77.145 191.995 ;
        RECT 77.315 191.365 77.485 192.165 ;
        RECT 77.685 191.195 78.015 191.995 ;
        RECT 78.215 191.365 78.495 192.165 ;
        RECT 76.815 191.025 78.095 191.195 ;
        RECT 75.235 190.365 75.755 190.905 ;
        RECT 76.410 190.525 76.695 190.855 ;
        RECT 76.895 190.525 77.275 190.855 ;
        RECT 77.445 190.525 77.755 190.855 ;
        RECT 73.910 189.810 74.375 190.355 ;
        RECT 74.545 189.615 75.755 190.365 ;
        RECT 75.925 189.615 76.215 190.340 ;
        RECT 76.390 189.615 76.725 190.355 ;
        RECT 76.895 189.830 77.110 190.525 ;
        RECT 77.445 190.355 77.650 190.525 ;
        RECT 77.925 190.355 78.095 191.025 ;
        RECT 78.275 190.525 78.515 191.195 ;
        RECT 79.605 191.075 83.115 192.165 ;
        RECT 83.660 191.185 83.915 191.855 ;
        RECT 84.095 191.365 84.380 192.165 ;
        RECT 84.560 191.445 84.890 191.955 ;
        RECT 79.605 190.555 81.295 191.075 ;
        RECT 81.465 190.385 83.115 190.905 ;
        RECT 77.300 189.830 77.650 190.355 ;
        RECT 77.820 189.785 78.515 190.355 ;
        RECT 79.605 189.615 83.115 190.385 ;
        RECT 83.660 190.325 83.840 191.185 ;
        RECT 84.560 190.855 84.810 191.445 ;
        RECT 85.160 191.295 85.330 191.905 ;
        RECT 85.500 191.475 85.830 192.165 ;
        RECT 86.060 191.615 86.300 191.905 ;
        RECT 86.500 191.785 86.920 192.165 ;
        RECT 87.100 191.695 87.730 191.945 ;
        RECT 88.200 191.785 88.530 192.165 ;
        RECT 87.100 191.615 87.270 191.695 ;
        RECT 88.700 191.615 88.870 191.905 ;
        RECT 89.050 191.785 89.430 192.165 ;
        RECT 89.670 191.780 90.500 191.950 ;
        RECT 86.060 191.445 87.270 191.615 ;
        RECT 84.010 190.525 84.810 190.855 ;
        RECT 83.660 190.125 83.915 190.325 ;
        RECT 83.575 189.955 83.915 190.125 ;
        RECT 83.660 189.795 83.915 189.955 ;
        RECT 84.095 189.615 84.380 190.075 ;
        RECT 84.560 189.875 84.810 190.525 ;
        RECT 85.010 191.275 85.330 191.295 ;
        RECT 85.010 191.105 86.930 191.275 ;
        RECT 85.010 190.210 85.200 191.105 ;
        RECT 87.100 190.935 87.270 191.445 ;
        RECT 87.440 191.185 87.960 191.495 ;
        RECT 85.370 190.765 87.270 190.935 ;
        RECT 85.370 190.705 85.700 190.765 ;
        RECT 85.850 190.535 86.180 190.595 ;
        RECT 85.520 190.265 86.180 190.535 ;
        RECT 85.010 189.880 85.330 190.210 ;
        RECT 85.510 189.615 86.170 190.095 ;
        RECT 86.370 190.005 86.540 190.765 ;
        RECT 87.440 190.595 87.620 191.005 ;
        RECT 86.710 190.425 87.040 190.545 ;
        RECT 87.790 190.425 87.960 191.185 ;
        RECT 86.710 190.255 87.960 190.425 ;
        RECT 88.130 191.365 89.500 191.615 ;
        RECT 88.130 190.595 88.320 191.365 ;
        RECT 89.250 191.105 89.500 191.365 ;
        RECT 88.490 190.935 88.740 191.095 ;
        RECT 89.670 190.935 89.840 191.780 ;
        RECT 90.735 191.495 90.905 191.995 ;
        RECT 91.075 191.665 91.405 192.165 ;
        RECT 90.010 191.105 90.510 191.485 ;
        RECT 90.735 191.325 91.430 191.495 ;
        RECT 88.490 190.765 89.840 190.935 ;
        RECT 89.420 190.725 89.840 190.765 ;
        RECT 88.130 190.255 88.550 190.595 ;
        RECT 88.840 190.265 89.250 190.595 ;
        RECT 86.370 189.835 87.220 190.005 ;
        RECT 87.780 189.615 88.100 190.075 ;
        RECT 88.300 189.825 88.550 190.255 ;
        RECT 88.840 189.615 89.250 190.055 ;
        RECT 89.420 189.995 89.590 190.725 ;
        RECT 89.760 190.175 90.110 190.545 ;
        RECT 90.290 190.235 90.510 191.105 ;
        RECT 90.680 190.535 91.090 191.155 ;
        RECT 91.260 190.355 91.430 191.325 ;
        RECT 90.735 190.165 91.430 190.355 ;
        RECT 89.420 189.795 90.435 189.995 ;
        RECT 90.735 189.835 90.905 190.165 ;
        RECT 91.075 189.615 91.405 189.995 ;
        RECT 91.620 189.875 91.845 191.995 ;
        RECT 92.015 191.665 92.345 192.165 ;
        RECT 92.515 191.495 92.685 191.995 ;
        RECT 92.020 191.325 92.685 191.495 ;
        RECT 92.020 190.335 92.250 191.325 ;
        RECT 93.035 191.235 93.205 191.995 ;
        RECT 93.385 191.405 93.715 192.165 ;
        RECT 92.420 190.505 92.770 191.155 ;
        RECT 93.035 191.065 93.700 191.235 ;
        RECT 93.885 191.090 94.155 191.995 ;
        RECT 94.325 191.330 94.710 192.165 ;
        RECT 94.880 191.160 95.140 191.965 ;
        RECT 95.310 191.330 95.570 192.165 ;
        RECT 95.740 191.160 95.995 191.965 ;
        RECT 96.170 191.330 96.430 192.165 ;
        RECT 96.600 191.160 96.855 191.965 ;
        RECT 97.030 191.330 97.375 192.165 ;
        RECT 97.545 191.405 98.060 191.815 ;
        RECT 98.295 191.405 98.465 192.165 ;
        RECT 98.635 191.825 100.665 191.995 ;
        RECT 93.530 190.920 93.700 191.065 ;
        RECT 92.965 190.515 93.295 190.885 ;
        RECT 93.530 190.590 93.815 190.920 ;
        RECT 93.530 190.335 93.700 190.590 ;
        RECT 92.020 190.165 92.685 190.335 ;
        RECT 92.015 189.615 92.345 189.995 ;
        RECT 92.515 189.875 92.685 190.165 ;
        RECT 93.035 190.165 93.700 190.335 ;
        RECT 93.985 190.290 94.155 191.090 ;
        RECT 93.035 189.785 93.205 190.165 ;
        RECT 93.385 189.615 93.715 189.995 ;
        RECT 93.895 189.785 94.155 190.290 ;
        RECT 94.325 190.990 97.355 191.160 ;
        RECT 94.325 190.425 94.625 190.990 ;
        RECT 94.800 190.595 97.015 190.820 ;
        RECT 97.185 190.425 97.355 190.990 ;
        RECT 97.545 190.595 97.885 191.405 ;
        RECT 98.635 191.160 98.805 191.825 ;
        RECT 99.200 191.485 100.325 191.655 ;
        RECT 98.055 190.970 98.805 191.160 ;
        RECT 98.975 191.145 99.985 191.315 ;
        RECT 97.545 190.425 98.775 190.595 ;
        RECT 94.325 190.255 97.355 190.425 ;
        RECT 94.845 189.615 95.145 190.085 ;
        RECT 95.315 189.810 95.570 190.255 ;
        RECT 95.740 189.615 96.000 190.085 ;
        RECT 96.170 189.810 96.430 190.255 ;
        RECT 96.600 189.615 96.895 190.085 ;
        RECT 97.820 189.820 98.065 190.425 ;
        RECT 98.285 189.615 98.795 190.150 ;
        RECT 98.975 189.785 99.165 191.145 ;
        RECT 99.335 190.805 99.610 190.945 ;
        RECT 99.335 190.635 99.615 190.805 ;
        RECT 99.335 189.785 99.610 190.635 ;
        RECT 99.815 190.345 99.985 191.145 ;
        RECT 100.155 190.355 100.325 191.485 ;
        RECT 100.495 190.855 100.665 191.825 ;
        RECT 100.835 191.025 101.005 192.165 ;
        RECT 101.175 191.025 101.510 191.995 ;
        RECT 100.495 190.525 100.690 190.855 ;
        RECT 100.915 190.525 101.170 190.855 ;
        RECT 100.915 190.355 101.085 190.525 ;
        RECT 101.340 190.355 101.510 191.025 ;
        RECT 101.685 191.000 101.975 192.165 ;
        RECT 102.235 191.235 102.405 191.995 ;
        RECT 102.585 191.405 102.915 192.165 ;
        RECT 102.235 191.065 102.900 191.235 ;
        RECT 103.085 191.090 103.355 191.995 ;
        RECT 102.730 190.920 102.900 191.065 ;
        RECT 102.165 190.515 102.495 190.885 ;
        RECT 102.730 190.590 103.015 190.920 ;
        RECT 100.155 190.185 101.085 190.355 ;
        RECT 100.155 190.150 100.330 190.185 ;
        RECT 99.800 189.785 100.330 190.150 ;
        RECT 100.755 189.615 101.085 190.015 ;
        RECT 101.255 189.785 101.510 190.355 ;
        RECT 101.685 189.615 101.975 190.340 ;
        RECT 102.730 190.335 102.900 190.590 ;
        RECT 102.235 190.165 102.900 190.335 ;
        RECT 103.185 190.290 103.355 191.090 ;
        RECT 103.525 191.075 104.735 192.165 ;
        RECT 104.905 191.405 105.420 191.815 ;
        RECT 105.655 191.405 105.825 192.165 ;
        RECT 105.995 191.825 108.025 191.995 ;
        RECT 103.525 190.535 104.045 191.075 ;
        RECT 104.215 190.365 104.735 190.905 ;
        RECT 104.905 190.595 105.245 191.405 ;
        RECT 105.995 191.160 106.165 191.825 ;
        RECT 106.560 191.485 107.685 191.655 ;
        RECT 105.415 190.970 106.165 191.160 ;
        RECT 106.335 191.145 107.345 191.315 ;
        RECT 104.905 190.425 106.135 190.595 ;
        RECT 102.235 189.785 102.405 190.165 ;
        RECT 102.585 189.615 102.915 189.995 ;
        RECT 103.095 189.785 103.355 190.290 ;
        RECT 103.525 189.615 104.735 190.365 ;
        RECT 105.180 189.820 105.425 190.425 ;
        RECT 105.645 189.615 106.155 190.150 ;
        RECT 106.335 189.785 106.525 191.145 ;
        RECT 106.695 190.805 106.970 190.945 ;
        RECT 106.695 190.635 106.975 190.805 ;
        RECT 106.695 189.785 106.970 190.635 ;
        RECT 107.175 190.345 107.345 191.145 ;
        RECT 107.515 190.355 107.685 191.485 ;
        RECT 107.855 190.855 108.025 191.825 ;
        RECT 108.195 191.025 108.365 192.165 ;
        RECT 108.535 191.025 108.870 191.995 ;
        RECT 107.855 190.525 108.050 190.855 ;
        RECT 108.275 190.525 108.530 190.855 ;
        RECT 108.275 190.355 108.445 190.525 ;
        RECT 108.700 190.355 108.870 191.025 ;
        RECT 107.515 190.185 108.445 190.355 ;
        RECT 107.515 190.150 107.690 190.185 ;
        RECT 107.160 189.785 107.690 190.150 ;
        RECT 108.115 189.615 108.445 190.015 ;
        RECT 108.615 189.785 108.870 190.355 ;
        RECT 109.050 190.975 109.305 191.855 ;
        RECT 109.475 191.025 109.780 192.165 ;
        RECT 110.120 191.785 110.450 192.165 ;
        RECT 110.630 191.615 110.800 191.905 ;
        RECT 110.970 191.705 111.220 192.165 ;
        RECT 110.000 191.445 110.800 191.615 ;
        RECT 111.390 191.655 112.260 191.995 ;
        RECT 109.050 190.325 109.260 190.975 ;
        RECT 110.000 190.855 110.170 191.445 ;
        RECT 111.390 191.275 111.560 191.655 ;
        RECT 112.495 191.535 112.665 191.995 ;
        RECT 112.835 191.705 113.205 192.165 ;
        RECT 113.500 191.565 113.670 191.905 ;
        RECT 113.840 191.735 114.170 192.165 ;
        RECT 114.405 191.565 114.575 191.905 ;
        RECT 110.340 191.105 111.560 191.275 ;
        RECT 111.730 191.195 112.190 191.485 ;
        RECT 112.495 191.365 113.055 191.535 ;
        RECT 113.500 191.395 114.575 191.565 ;
        RECT 114.745 191.665 115.425 191.995 ;
        RECT 115.640 191.665 115.890 191.995 ;
        RECT 116.060 191.705 116.310 192.165 ;
        RECT 112.885 191.225 113.055 191.365 ;
        RECT 111.730 191.185 112.695 191.195 ;
        RECT 111.390 191.015 111.560 191.105 ;
        RECT 112.020 191.025 112.695 191.185 ;
        RECT 109.430 190.825 110.170 190.855 ;
        RECT 109.430 190.525 110.345 190.825 ;
        RECT 110.020 190.350 110.345 190.525 ;
        RECT 109.050 189.795 109.305 190.325 ;
        RECT 109.475 189.615 109.780 190.075 ;
        RECT 110.025 189.995 110.345 190.350 ;
        RECT 110.515 190.565 111.055 190.935 ;
        RECT 111.390 190.845 111.795 191.015 ;
        RECT 110.515 190.165 110.755 190.565 ;
        RECT 111.235 190.395 111.455 190.675 ;
        RECT 110.925 190.225 111.455 190.395 ;
        RECT 110.925 189.995 111.095 190.225 ;
        RECT 111.625 190.065 111.795 190.845 ;
        RECT 111.965 190.235 112.315 190.855 ;
        RECT 112.485 190.235 112.695 191.025 ;
        RECT 112.885 191.055 114.385 191.225 ;
        RECT 112.885 190.365 113.055 191.055 ;
        RECT 114.745 190.885 114.915 191.665 ;
        RECT 115.720 191.535 115.890 191.665 ;
        RECT 113.225 190.715 114.915 190.885 ;
        RECT 115.085 191.105 115.550 191.495 ;
        RECT 115.720 191.365 116.115 191.535 ;
        RECT 113.225 190.535 113.395 190.715 ;
        RECT 110.025 189.825 111.095 189.995 ;
        RECT 111.265 189.615 111.455 190.055 ;
        RECT 111.625 189.785 112.575 190.065 ;
        RECT 112.885 189.975 113.145 190.365 ;
        RECT 113.565 190.295 114.355 190.545 ;
        RECT 112.795 189.805 113.145 189.975 ;
        RECT 113.355 189.615 113.685 190.075 ;
        RECT 114.560 190.005 114.730 190.715 ;
        RECT 115.085 190.515 115.255 191.105 ;
        RECT 114.900 190.295 115.255 190.515 ;
        RECT 115.425 190.295 115.775 190.915 ;
        RECT 115.945 190.005 116.115 191.365 ;
        RECT 116.480 191.195 116.805 191.980 ;
        RECT 116.285 190.145 116.745 191.195 ;
        RECT 114.560 189.835 115.415 190.005 ;
        RECT 115.620 189.835 116.115 190.005 ;
        RECT 116.285 189.615 116.615 189.975 ;
        RECT 116.975 189.875 117.145 191.995 ;
        RECT 117.315 191.665 117.645 192.165 ;
        RECT 117.815 191.495 118.070 191.995 ;
        RECT 117.320 191.325 118.070 191.495 ;
        RECT 117.320 190.335 117.550 191.325 ;
        RECT 117.720 190.505 118.070 191.155 ;
        RECT 118.245 191.090 118.515 191.995 ;
        RECT 118.685 191.405 119.015 192.165 ;
        RECT 119.195 191.235 119.365 191.995 ;
        RECT 117.320 190.165 118.070 190.335 ;
        RECT 117.315 189.615 117.645 189.995 ;
        RECT 117.815 189.875 118.070 190.165 ;
        RECT 118.245 190.290 118.415 191.090 ;
        RECT 118.700 191.065 119.365 191.235 ;
        RECT 119.625 191.075 120.835 192.165 ;
        RECT 121.010 191.730 126.355 192.165 ;
        RECT 118.700 190.920 118.870 191.065 ;
        RECT 118.585 190.590 118.870 190.920 ;
        RECT 118.700 190.335 118.870 190.590 ;
        RECT 119.105 190.515 119.435 190.885 ;
        RECT 119.625 190.535 120.145 191.075 ;
        RECT 120.315 190.365 120.835 190.905 ;
        RECT 122.600 190.480 122.950 191.730 ;
        RECT 126.525 191.075 127.735 192.165 ;
        RECT 118.245 189.785 118.505 190.290 ;
        RECT 118.700 190.165 119.365 190.335 ;
        RECT 118.685 189.615 119.015 189.995 ;
        RECT 119.195 189.785 119.365 190.165 ;
        RECT 119.625 189.615 120.835 190.365 ;
        RECT 124.430 190.160 124.770 190.990 ;
        RECT 126.525 190.535 127.045 191.075 ;
        RECT 127.215 190.365 127.735 190.905 ;
        RECT 121.010 189.615 126.355 190.160 ;
        RECT 126.525 189.615 127.735 190.365 ;
        RECT 14.660 189.445 127.820 189.615 ;
        RECT 14.745 188.695 15.955 189.445 ;
        RECT 14.745 188.155 15.265 188.695 ;
        RECT 16.585 188.675 18.255 189.445 ;
        RECT 18.430 188.900 23.775 189.445 ;
        RECT 23.950 188.900 29.295 189.445 ;
        RECT 15.435 187.985 15.955 188.525 ;
        RECT 14.745 186.895 15.955 187.985 ;
        RECT 16.585 187.985 17.335 188.505 ;
        RECT 17.505 188.155 18.255 188.675 ;
        RECT 16.585 186.895 18.255 187.985 ;
        RECT 20.020 187.330 20.370 188.580 ;
        RECT 21.850 188.070 22.190 188.900 ;
        RECT 25.540 187.330 25.890 188.580 ;
        RECT 27.370 188.070 27.710 188.900 ;
        RECT 29.525 188.625 29.735 189.445 ;
        RECT 29.905 188.645 30.235 189.275 ;
        RECT 29.905 188.045 30.155 188.645 ;
        RECT 30.405 188.625 30.635 189.445 ;
        RECT 30.845 188.695 32.055 189.445 ;
        RECT 30.325 188.205 30.655 188.455 ;
        RECT 18.430 186.895 23.775 187.330 ;
        RECT 23.950 186.895 29.295 187.330 ;
        RECT 29.525 186.895 29.735 188.035 ;
        RECT 29.905 187.065 30.235 188.045 ;
        RECT 30.405 186.895 30.635 188.035 ;
        RECT 30.845 187.985 31.365 188.525 ;
        RECT 31.535 188.155 32.055 188.695 ;
        RECT 32.225 188.675 35.735 189.445 ;
        RECT 32.225 187.985 33.915 188.505 ;
        RECT 34.085 188.155 35.735 188.675 ;
        RECT 35.945 188.625 36.175 189.445 ;
        RECT 36.345 188.645 36.675 189.275 ;
        RECT 35.925 188.205 36.255 188.455 ;
        RECT 36.425 188.045 36.675 188.645 ;
        RECT 36.845 188.625 37.055 189.445 ;
        RECT 37.285 188.720 37.575 189.445 ;
        RECT 37.750 188.735 38.005 189.265 ;
        RECT 38.175 188.985 38.480 189.445 ;
        RECT 38.725 189.065 39.795 189.235 ;
        RECT 37.750 188.085 37.960 188.735 ;
        RECT 38.725 188.710 39.045 189.065 ;
        RECT 38.720 188.535 39.045 188.710 ;
        RECT 38.130 188.235 39.045 188.535 ;
        RECT 39.215 188.495 39.455 188.895 ;
        RECT 39.625 188.835 39.795 189.065 ;
        RECT 39.965 189.005 40.155 189.445 ;
        RECT 40.325 188.995 41.275 189.275 ;
        RECT 41.495 189.085 41.845 189.255 ;
        RECT 39.625 188.665 40.155 188.835 ;
        RECT 38.130 188.205 38.870 188.235 ;
        RECT 30.845 186.895 32.055 187.985 ;
        RECT 32.225 186.895 35.735 187.985 ;
        RECT 35.945 186.895 36.175 188.035 ;
        RECT 36.345 187.065 36.675 188.045 ;
        RECT 36.845 186.895 37.055 188.035 ;
        RECT 37.285 186.895 37.575 188.060 ;
        RECT 37.750 187.205 38.005 188.085 ;
        RECT 38.175 186.895 38.480 188.035 ;
        RECT 38.700 187.615 38.870 188.205 ;
        RECT 39.215 188.125 39.755 188.495 ;
        RECT 39.935 188.385 40.155 188.665 ;
        RECT 40.325 188.215 40.495 188.995 ;
        RECT 40.090 188.045 40.495 188.215 ;
        RECT 40.665 188.205 41.015 188.825 ;
        RECT 40.090 187.955 40.260 188.045 ;
        RECT 41.185 188.035 41.395 188.825 ;
        RECT 39.040 187.785 40.260 187.955 ;
        RECT 40.720 187.875 41.395 188.035 ;
        RECT 38.700 187.445 39.500 187.615 ;
        RECT 38.820 186.895 39.150 187.275 ;
        RECT 39.330 187.155 39.500 187.445 ;
        RECT 40.090 187.405 40.260 187.785 ;
        RECT 40.430 187.865 41.395 187.875 ;
        RECT 41.585 188.695 41.845 189.085 ;
        RECT 42.055 188.985 42.385 189.445 ;
        RECT 43.260 189.055 44.115 189.225 ;
        RECT 44.320 189.055 44.815 189.225 ;
        RECT 44.985 189.085 45.315 189.445 ;
        RECT 41.585 188.005 41.755 188.695 ;
        RECT 41.925 188.345 42.095 188.525 ;
        RECT 42.265 188.515 43.055 188.765 ;
        RECT 43.260 188.345 43.430 189.055 ;
        RECT 43.600 188.545 43.955 188.765 ;
        RECT 41.925 188.175 43.615 188.345 ;
        RECT 40.430 187.575 40.890 187.865 ;
        RECT 41.585 187.835 43.085 188.005 ;
        RECT 41.585 187.695 41.755 187.835 ;
        RECT 41.195 187.525 41.755 187.695 ;
        RECT 39.670 186.895 39.920 187.355 ;
        RECT 40.090 187.065 40.960 187.405 ;
        RECT 41.195 187.065 41.365 187.525 ;
        RECT 42.200 187.495 43.275 187.665 ;
        RECT 41.535 186.895 41.905 187.355 ;
        RECT 42.200 187.155 42.370 187.495 ;
        RECT 42.540 186.895 42.870 187.325 ;
        RECT 43.105 187.155 43.275 187.495 ;
        RECT 43.445 187.395 43.615 188.175 ;
        RECT 43.785 187.955 43.955 188.545 ;
        RECT 44.125 188.145 44.475 188.765 ;
        RECT 43.785 187.565 44.250 187.955 ;
        RECT 44.645 187.695 44.815 189.055 ;
        RECT 44.985 187.865 45.445 188.915 ;
        RECT 44.420 187.525 44.815 187.695 ;
        RECT 44.420 187.395 44.590 187.525 ;
        RECT 43.445 187.065 44.125 187.395 ;
        RECT 44.340 187.065 44.590 187.395 ;
        RECT 44.760 186.895 45.010 187.355 ;
        RECT 45.180 187.080 45.505 187.865 ;
        RECT 45.675 187.065 45.845 189.185 ;
        RECT 46.015 189.065 46.345 189.445 ;
        RECT 46.515 188.895 46.770 189.185 ;
        RECT 47.035 188.965 47.335 189.445 ;
        RECT 46.020 188.725 46.770 188.895 ;
        RECT 47.505 188.795 47.765 189.250 ;
        RECT 47.935 188.965 48.195 189.445 ;
        RECT 48.375 188.795 48.635 189.250 ;
        RECT 48.805 188.965 49.055 189.445 ;
        RECT 49.235 188.795 49.495 189.250 ;
        RECT 49.665 188.965 49.915 189.445 ;
        RECT 50.095 188.795 50.355 189.250 ;
        RECT 50.525 188.965 50.770 189.445 ;
        RECT 50.940 188.795 51.215 189.250 ;
        RECT 51.385 188.965 51.630 189.445 ;
        RECT 51.800 188.795 52.060 189.250 ;
        RECT 52.230 188.965 52.490 189.445 ;
        RECT 52.660 188.795 52.920 189.250 ;
        RECT 53.090 188.965 53.350 189.445 ;
        RECT 53.520 188.795 53.780 189.250 ;
        RECT 53.950 188.885 54.210 189.445 ;
        RECT 46.020 187.735 46.250 188.725 ;
        RECT 47.035 188.625 53.780 188.795 ;
        RECT 46.420 187.905 46.770 188.555 ;
        RECT 47.035 188.035 48.200 188.625 ;
        RECT 54.380 188.455 54.630 189.265 ;
        RECT 54.810 188.920 55.070 189.445 ;
        RECT 55.240 188.455 55.490 189.265 ;
        RECT 55.670 188.935 55.975 189.445 ;
        RECT 48.370 188.205 55.490 188.455 ;
        RECT 55.660 188.205 55.975 188.765 ;
        RECT 56.420 188.635 56.665 189.240 ;
        RECT 56.885 188.910 57.395 189.445 ;
        RECT 56.145 188.465 57.375 188.635 ;
        RECT 47.035 187.810 53.780 188.035 ;
        RECT 46.020 187.565 46.770 187.735 ;
        RECT 46.015 186.895 46.345 187.395 ;
        RECT 46.515 187.065 46.770 187.565 ;
        RECT 47.035 186.895 47.305 187.640 ;
        RECT 47.475 187.070 47.765 187.810 ;
        RECT 48.375 187.795 53.780 187.810 ;
        RECT 47.935 186.900 48.190 187.625 ;
        RECT 48.375 187.070 48.635 187.795 ;
        RECT 48.805 186.900 49.050 187.625 ;
        RECT 49.235 187.070 49.495 187.795 ;
        RECT 49.665 186.900 49.910 187.625 ;
        RECT 50.095 187.070 50.355 187.795 ;
        RECT 50.525 186.900 50.770 187.625 ;
        RECT 50.940 187.070 51.200 187.795 ;
        RECT 51.370 186.900 51.630 187.625 ;
        RECT 51.800 187.070 52.060 187.795 ;
        RECT 52.230 186.900 52.490 187.625 ;
        RECT 52.660 187.070 52.920 187.795 ;
        RECT 53.090 186.900 53.350 187.625 ;
        RECT 53.520 187.070 53.780 187.795 ;
        RECT 53.950 186.900 54.210 187.695 ;
        RECT 54.380 187.070 54.630 188.205 ;
        RECT 47.935 186.895 54.210 186.900 ;
        RECT 54.810 186.895 55.070 187.705 ;
        RECT 55.245 187.065 55.490 188.205 ;
        RECT 55.670 186.895 55.965 187.705 ;
        RECT 56.145 187.655 56.485 188.465 ;
        RECT 56.655 187.900 57.405 188.090 ;
        RECT 56.145 187.245 56.660 187.655 ;
        RECT 56.895 186.895 57.065 187.655 ;
        RECT 57.235 187.235 57.405 187.900 ;
        RECT 57.575 187.915 57.765 189.275 ;
        RECT 57.935 189.105 58.210 189.275 ;
        RECT 57.935 188.935 58.215 189.105 ;
        RECT 57.935 188.115 58.210 188.935 ;
        RECT 58.400 188.910 58.930 189.275 ;
        RECT 59.355 189.045 59.685 189.445 ;
        RECT 58.755 188.875 58.930 188.910 ;
        RECT 58.415 187.915 58.585 188.715 ;
        RECT 57.575 187.745 58.585 187.915 ;
        RECT 58.755 188.705 59.685 188.875 ;
        RECT 59.855 188.705 60.110 189.275 ;
        RECT 58.755 187.575 58.925 188.705 ;
        RECT 59.515 188.535 59.685 188.705 ;
        RECT 57.800 187.405 58.925 187.575 ;
        RECT 59.095 188.205 59.290 188.535 ;
        RECT 59.515 188.205 59.770 188.535 ;
        RECT 59.095 187.235 59.265 188.205 ;
        RECT 59.940 188.035 60.110 188.705 ;
        RECT 57.235 187.065 59.265 187.235 ;
        RECT 59.435 186.895 59.605 188.035 ;
        RECT 59.775 187.065 60.110 188.035 ;
        RECT 60.285 188.770 60.545 189.275 ;
        RECT 60.725 189.065 61.055 189.445 ;
        RECT 61.235 188.895 61.405 189.275 ;
        RECT 60.285 187.970 60.455 188.770 ;
        RECT 60.740 188.725 61.405 188.895 ;
        RECT 60.740 188.470 60.910 188.725 ;
        RECT 61.665 188.695 62.875 189.445 ;
        RECT 63.045 188.720 63.335 189.445 ;
        RECT 64.080 188.815 64.365 189.275 ;
        RECT 64.535 188.985 64.805 189.445 ;
        RECT 60.625 188.140 60.910 188.470 ;
        RECT 61.145 188.175 61.475 188.545 ;
        RECT 60.740 187.995 60.910 188.140 ;
        RECT 60.285 187.065 60.555 187.970 ;
        RECT 60.740 187.825 61.405 187.995 ;
        RECT 60.725 186.895 61.055 187.655 ;
        RECT 61.235 187.065 61.405 187.825 ;
        RECT 61.665 187.985 62.185 188.525 ;
        RECT 62.355 188.155 62.875 188.695 ;
        RECT 64.080 188.645 65.035 188.815 ;
        RECT 61.665 186.895 62.875 187.985 ;
        RECT 63.045 186.895 63.335 188.060 ;
        RECT 63.965 187.915 64.655 188.475 ;
        RECT 64.825 187.745 65.035 188.645 ;
        RECT 64.080 187.525 65.035 187.745 ;
        RECT 65.205 188.475 65.605 189.275 ;
        RECT 65.795 188.815 66.075 189.275 ;
        RECT 66.595 188.985 66.920 189.445 ;
        RECT 65.795 188.645 66.920 188.815 ;
        RECT 67.090 188.705 67.475 189.275 ;
        RECT 66.470 188.535 66.920 188.645 ;
        RECT 65.205 187.915 66.300 188.475 ;
        RECT 66.470 188.205 67.025 188.535 ;
        RECT 64.080 187.065 64.365 187.525 ;
        RECT 64.535 186.895 64.805 187.355 ;
        RECT 65.205 187.065 65.605 187.915 ;
        RECT 66.470 187.745 66.920 188.205 ;
        RECT 67.195 188.035 67.475 188.705 ;
        RECT 67.645 188.675 70.235 189.445 ;
        RECT 70.410 188.900 75.755 189.445 ;
        RECT 75.930 188.900 81.275 189.445 ;
        RECT 81.450 188.900 86.795 189.445 ;
        RECT 65.795 187.525 66.920 187.745 ;
        RECT 65.795 187.065 66.075 187.525 ;
        RECT 66.595 186.895 66.920 187.355 ;
        RECT 67.090 187.065 67.475 188.035 ;
        RECT 67.645 187.985 68.855 188.505 ;
        RECT 69.025 188.155 70.235 188.675 ;
        RECT 67.645 186.895 70.235 187.985 ;
        RECT 72.000 187.330 72.350 188.580 ;
        RECT 73.830 188.070 74.170 188.900 ;
        RECT 77.520 187.330 77.870 188.580 ;
        RECT 79.350 188.070 79.690 188.900 ;
        RECT 83.040 187.330 83.390 188.580 ;
        RECT 84.870 188.070 85.210 188.900 ;
        RECT 87.025 188.625 87.235 189.445 ;
        RECT 87.405 188.645 87.735 189.275 ;
        RECT 87.405 188.045 87.655 188.645 ;
        RECT 87.905 188.625 88.135 189.445 ;
        RECT 88.805 188.720 89.095 189.445 ;
        RECT 89.355 188.895 89.525 189.275 ;
        RECT 89.705 189.065 90.035 189.445 ;
        RECT 89.355 188.725 90.020 188.895 ;
        RECT 90.215 188.770 90.475 189.275 ;
        RECT 87.825 188.205 88.155 188.455 ;
        RECT 89.285 188.175 89.615 188.545 ;
        RECT 89.850 188.470 90.020 188.725 ;
        RECT 89.850 188.140 90.135 188.470 ;
        RECT 70.410 186.895 75.755 187.330 ;
        RECT 75.930 186.895 81.275 187.330 ;
        RECT 81.450 186.895 86.795 187.330 ;
        RECT 87.025 186.895 87.235 188.035 ;
        RECT 87.405 187.065 87.735 188.045 ;
        RECT 87.905 186.895 88.135 188.035 ;
        RECT 88.805 186.895 89.095 188.060 ;
        RECT 89.850 187.995 90.020 188.140 ;
        RECT 89.355 187.825 90.020 187.995 ;
        RECT 90.305 187.970 90.475 188.770 ;
        RECT 90.645 188.675 92.315 189.445 ;
        RECT 92.490 188.900 97.835 189.445 ;
        RECT 89.355 187.065 89.525 187.825 ;
        RECT 89.705 186.895 90.035 187.655 ;
        RECT 90.205 187.065 90.475 187.970 ;
        RECT 90.645 187.985 91.395 188.505 ;
        RECT 91.565 188.155 92.315 188.675 ;
        RECT 90.645 186.895 92.315 187.985 ;
        RECT 94.080 187.330 94.430 188.580 ;
        RECT 95.910 188.070 96.250 188.900 ;
        RECT 98.010 188.735 98.265 189.265 ;
        RECT 98.435 188.985 98.740 189.445 ;
        RECT 98.985 189.065 100.055 189.235 ;
        RECT 98.010 188.085 98.220 188.735 ;
        RECT 98.985 188.710 99.305 189.065 ;
        RECT 98.980 188.535 99.305 188.710 ;
        RECT 98.390 188.235 99.305 188.535 ;
        RECT 99.475 188.495 99.715 188.895 ;
        RECT 99.885 188.835 100.055 189.065 ;
        RECT 100.225 189.005 100.415 189.445 ;
        RECT 100.585 188.995 101.535 189.275 ;
        RECT 101.755 189.085 102.105 189.255 ;
        RECT 99.885 188.665 100.415 188.835 ;
        RECT 98.390 188.205 99.130 188.235 ;
        RECT 92.490 186.895 97.835 187.330 ;
        RECT 98.010 187.205 98.265 188.085 ;
        RECT 98.435 186.895 98.740 188.035 ;
        RECT 98.960 187.615 99.130 188.205 ;
        RECT 99.475 188.125 100.015 188.495 ;
        RECT 100.195 188.385 100.415 188.665 ;
        RECT 100.585 188.215 100.755 188.995 ;
        RECT 100.350 188.045 100.755 188.215 ;
        RECT 100.925 188.205 101.275 188.825 ;
        RECT 100.350 187.955 100.520 188.045 ;
        RECT 101.445 188.035 101.655 188.825 ;
        RECT 99.300 187.785 100.520 187.955 ;
        RECT 100.980 187.875 101.655 188.035 ;
        RECT 98.960 187.445 99.760 187.615 ;
        RECT 99.080 186.895 99.410 187.275 ;
        RECT 99.590 187.155 99.760 187.445 ;
        RECT 100.350 187.405 100.520 187.785 ;
        RECT 100.690 187.865 101.655 187.875 ;
        RECT 101.845 188.695 102.105 189.085 ;
        RECT 102.315 188.985 102.645 189.445 ;
        RECT 103.520 189.055 104.375 189.225 ;
        RECT 104.580 189.055 105.075 189.225 ;
        RECT 105.245 189.085 105.575 189.445 ;
        RECT 101.845 188.005 102.015 188.695 ;
        RECT 102.185 188.345 102.355 188.525 ;
        RECT 102.525 188.515 103.315 188.765 ;
        RECT 103.520 188.345 103.690 189.055 ;
        RECT 103.860 188.545 104.215 188.765 ;
        RECT 102.185 188.175 103.875 188.345 ;
        RECT 100.690 187.575 101.150 187.865 ;
        RECT 101.845 187.835 103.345 188.005 ;
        RECT 101.845 187.695 102.015 187.835 ;
        RECT 101.455 187.525 102.015 187.695 ;
        RECT 99.930 186.895 100.180 187.355 ;
        RECT 100.350 187.065 101.220 187.405 ;
        RECT 101.455 187.065 101.625 187.525 ;
        RECT 102.460 187.495 103.535 187.665 ;
        RECT 101.795 186.895 102.165 187.355 ;
        RECT 102.460 187.155 102.630 187.495 ;
        RECT 102.800 186.895 103.130 187.325 ;
        RECT 103.365 187.155 103.535 187.495 ;
        RECT 103.705 187.395 103.875 188.175 ;
        RECT 104.045 187.955 104.215 188.545 ;
        RECT 104.385 188.145 104.735 188.765 ;
        RECT 104.045 187.565 104.510 187.955 ;
        RECT 104.905 187.695 105.075 189.055 ;
        RECT 105.245 187.865 105.705 188.915 ;
        RECT 104.680 187.525 105.075 187.695 ;
        RECT 104.680 187.395 104.850 187.525 ;
        RECT 103.705 187.065 104.385 187.395 ;
        RECT 104.600 187.065 104.850 187.395 ;
        RECT 105.020 186.895 105.270 187.355 ;
        RECT 105.440 187.080 105.765 187.865 ;
        RECT 105.935 187.065 106.105 189.185 ;
        RECT 106.275 189.065 106.605 189.445 ;
        RECT 106.775 188.895 107.030 189.185 ;
        RECT 106.280 188.725 107.030 188.895 ;
        RECT 106.280 187.735 106.510 188.725 ;
        RECT 107.205 188.705 107.590 189.275 ;
        RECT 107.760 188.985 108.085 189.445 ;
        RECT 108.605 188.815 108.885 189.275 ;
        RECT 106.680 187.905 107.030 188.555 ;
        RECT 107.205 188.035 107.485 188.705 ;
        RECT 107.760 188.645 108.885 188.815 ;
        RECT 107.760 188.535 108.210 188.645 ;
        RECT 107.655 188.205 108.210 188.535 ;
        RECT 109.075 188.475 109.475 189.275 ;
        RECT 109.875 188.985 110.145 189.445 ;
        RECT 110.315 188.815 110.600 189.275 ;
        RECT 106.280 187.565 107.030 187.735 ;
        RECT 106.275 186.895 106.605 187.395 ;
        RECT 106.775 187.065 107.030 187.565 ;
        RECT 107.205 187.065 107.590 188.035 ;
        RECT 107.760 187.745 108.210 188.205 ;
        RECT 108.380 187.915 109.475 188.475 ;
        RECT 107.760 187.525 108.885 187.745 ;
        RECT 107.760 186.895 108.085 187.355 ;
        RECT 108.605 187.065 108.885 187.525 ;
        RECT 109.075 187.065 109.475 187.915 ;
        RECT 109.645 188.645 110.600 188.815 ;
        RECT 111.345 188.675 113.015 189.445 ;
        RECT 113.275 188.895 113.445 189.275 ;
        RECT 113.625 189.065 113.955 189.445 ;
        RECT 113.275 188.725 113.940 188.895 ;
        RECT 114.135 188.770 114.395 189.275 ;
        RECT 109.645 187.745 109.855 188.645 ;
        RECT 110.025 187.915 110.715 188.475 ;
        RECT 111.345 187.985 112.095 188.505 ;
        RECT 112.265 188.155 113.015 188.675 ;
        RECT 113.205 188.175 113.535 188.545 ;
        RECT 113.770 188.470 113.940 188.725 ;
        RECT 113.770 188.140 114.055 188.470 ;
        RECT 113.770 187.995 113.940 188.140 ;
        RECT 109.645 187.525 110.600 187.745 ;
        RECT 109.875 186.895 110.145 187.355 ;
        RECT 110.315 187.065 110.600 187.525 ;
        RECT 111.345 186.895 113.015 187.985 ;
        RECT 113.275 187.825 113.940 187.995 ;
        RECT 114.225 187.970 114.395 188.770 ;
        RECT 114.565 188.720 114.855 189.445 ;
        RECT 115.490 188.900 120.835 189.445 ;
        RECT 121.010 188.900 126.355 189.445 ;
        RECT 113.275 187.065 113.445 187.825 ;
        RECT 113.625 186.895 113.955 187.655 ;
        RECT 114.125 187.065 114.395 187.970 ;
        RECT 114.565 186.895 114.855 188.060 ;
        RECT 117.080 187.330 117.430 188.580 ;
        RECT 118.910 188.070 119.250 188.900 ;
        RECT 122.600 187.330 122.950 188.580 ;
        RECT 124.430 188.070 124.770 188.900 ;
        RECT 126.525 188.695 127.735 189.445 ;
        RECT 126.525 187.985 127.045 188.525 ;
        RECT 127.215 188.155 127.735 188.695 ;
        RECT 115.490 186.895 120.835 187.330 ;
        RECT 121.010 186.895 126.355 187.330 ;
        RECT 126.525 186.895 127.735 187.985 ;
        RECT 14.660 186.725 127.820 186.895 ;
        RECT 14.745 185.635 15.955 186.725 ;
        RECT 14.745 184.925 15.265 185.465 ;
        RECT 15.435 185.095 15.955 185.635 ;
        RECT 16.125 185.635 18.715 186.725 ;
        RECT 18.890 186.290 24.235 186.725 ;
        RECT 16.125 185.115 17.335 185.635 ;
        RECT 17.505 184.945 18.715 185.465 ;
        RECT 20.480 185.040 20.830 186.290 ;
        RECT 24.405 185.560 24.695 186.725 ;
        RECT 24.865 185.635 26.075 186.725 ;
        RECT 14.745 184.175 15.955 184.925 ;
        RECT 16.125 184.175 18.715 184.945 ;
        RECT 22.310 184.720 22.650 185.550 ;
        RECT 24.865 185.095 25.385 185.635 ;
        RECT 26.250 185.535 26.505 186.415 ;
        RECT 26.675 185.585 26.980 186.725 ;
        RECT 27.320 186.345 27.650 186.725 ;
        RECT 27.830 186.175 28.000 186.465 ;
        RECT 28.170 186.265 28.420 186.725 ;
        RECT 27.200 186.005 28.000 186.175 ;
        RECT 28.590 186.215 29.460 186.555 ;
        RECT 25.555 184.925 26.075 185.465 ;
        RECT 18.890 184.175 24.235 184.720 ;
        RECT 24.405 184.175 24.695 184.900 ;
        RECT 24.865 184.175 26.075 184.925 ;
        RECT 26.250 184.885 26.460 185.535 ;
        RECT 27.200 185.415 27.370 186.005 ;
        RECT 28.590 185.835 28.760 186.215 ;
        RECT 29.695 186.095 29.865 186.555 ;
        RECT 30.035 186.265 30.405 186.725 ;
        RECT 30.700 186.125 30.870 186.465 ;
        RECT 31.040 186.295 31.370 186.725 ;
        RECT 31.605 186.125 31.775 186.465 ;
        RECT 27.540 185.665 28.760 185.835 ;
        RECT 28.930 185.755 29.390 186.045 ;
        RECT 29.695 185.925 30.255 186.095 ;
        RECT 30.700 185.955 31.775 186.125 ;
        RECT 31.945 186.225 32.625 186.555 ;
        RECT 32.840 186.225 33.090 186.555 ;
        RECT 33.260 186.265 33.510 186.725 ;
        RECT 30.085 185.785 30.255 185.925 ;
        RECT 28.930 185.745 29.895 185.755 ;
        RECT 28.590 185.575 28.760 185.665 ;
        RECT 29.220 185.585 29.895 185.745 ;
        RECT 26.630 185.385 27.370 185.415 ;
        RECT 26.630 185.085 27.545 185.385 ;
        RECT 27.220 184.910 27.545 185.085 ;
        RECT 26.250 184.355 26.505 184.885 ;
        RECT 26.675 184.175 26.980 184.635 ;
        RECT 27.225 184.555 27.545 184.910 ;
        RECT 27.715 185.125 28.255 185.495 ;
        RECT 28.590 185.405 28.995 185.575 ;
        RECT 27.715 184.725 27.955 185.125 ;
        RECT 28.435 184.955 28.655 185.235 ;
        RECT 28.125 184.785 28.655 184.955 ;
        RECT 28.125 184.555 28.295 184.785 ;
        RECT 28.825 184.625 28.995 185.405 ;
        RECT 29.165 184.795 29.515 185.415 ;
        RECT 29.685 184.795 29.895 185.585 ;
        RECT 30.085 185.615 31.585 185.785 ;
        RECT 30.085 184.925 30.255 185.615 ;
        RECT 31.945 185.445 32.115 186.225 ;
        RECT 32.920 186.095 33.090 186.225 ;
        RECT 30.425 185.275 32.115 185.445 ;
        RECT 32.285 185.665 32.750 186.055 ;
        RECT 32.920 185.925 33.315 186.095 ;
        RECT 30.425 185.095 30.595 185.275 ;
        RECT 27.225 184.385 28.295 184.555 ;
        RECT 28.465 184.175 28.655 184.615 ;
        RECT 28.825 184.345 29.775 184.625 ;
        RECT 30.085 184.535 30.345 184.925 ;
        RECT 30.765 184.855 31.555 185.105 ;
        RECT 29.995 184.365 30.345 184.535 ;
        RECT 30.555 184.175 30.885 184.635 ;
        RECT 31.760 184.565 31.930 185.275 ;
        RECT 32.285 185.075 32.455 185.665 ;
        RECT 32.100 184.855 32.455 185.075 ;
        RECT 32.625 184.855 32.975 185.475 ;
        RECT 33.145 184.565 33.315 185.925 ;
        RECT 33.680 185.755 34.005 186.540 ;
        RECT 33.485 184.705 33.945 185.755 ;
        RECT 31.760 184.395 32.615 184.565 ;
        RECT 32.820 184.395 33.315 184.565 ;
        RECT 33.485 184.175 33.815 184.535 ;
        RECT 34.175 184.435 34.345 186.555 ;
        RECT 34.515 186.225 34.845 186.725 ;
        RECT 35.015 186.055 35.270 186.555 ;
        RECT 34.520 185.885 35.270 186.055 ;
        RECT 34.520 184.895 34.750 185.885 ;
        RECT 34.920 185.065 35.270 185.715 ;
        RECT 35.905 185.635 38.495 186.725 ;
        RECT 35.905 185.115 37.115 185.635 ;
        RECT 38.705 185.585 38.935 186.725 ;
        RECT 39.105 185.575 39.435 186.555 ;
        RECT 39.605 185.585 39.815 186.725 ;
        RECT 40.045 185.965 40.560 186.375 ;
        RECT 40.795 185.965 40.965 186.725 ;
        RECT 41.135 186.385 43.165 186.555 ;
        RECT 37.285 184.945 38.495 185.465 ;
        RECT 38.685 185.165 39.015 185.415 ;
        RECT 34.520 184.725 35.270 184.895 ;
        RECT 34.515 184.175 34.845 184.555 ;
        RECT 35.015 184.435 35.270 184.725 ;
        RECT 35.905 184.175 38.495 184.945 ;
        RECT 38.705 184.175 38.935 184.995 ;
        RECT 39.185 184.975 39.435 185.575 ;
        RECT 40.045 185.155 40.385 185.965 ;
        RECT 41.135 185.720 41.305 186.385 ;
        RECT 41.700 186.045 42.825 186.215 ;
        RECT 40.555 185.530 41.305 185.720 ;
        RECT 41.475 185.705 42.485 185.875 ;
        RECT 39.105 184.345 39.435 184.975 ;
        RECT 39.605 184.175 39.815 184.995 ;
        RECT 40.045 184.985 41.275 185.155 ;
        RECT 40.320 184.380 40.565 184.985 ;
        RECT 40.785 184.175 41.295 184.710 ;
        RECT 41.475 184.345 41.665 185.705 ;
        RECT 41.835 184.685 42.110 185.505 ;
        RECT 42.315 184.905 42.485 185.705 ;
        RECT 42.655 184.915 42.825 186.045 ;
        RECT 42.995 185.415 43.165 186.385 ;
        RECT 43.335 185.585 43.505 186.725 ;
        RECT 43.675 185.585 44.010 186.555 ;
        RECT 42.995 185.085 43.190 185.415 ;
        RECT 43.415 185.085 43.670 185.415 ;
        RECT 43.415 184.915 43.585 185.085 ;
        RECT 43.840 184.915 44.010 185.585 ;
        RECT 42.655 184.745 43.585 184.915 ;
        RECT 42.655 184.710 42.830 184.745 ;
        RECT 41.835 184.515 42.115 184.685 ;
        RECT 41.835 184.345 42.110 184.515 ;
        RECT 42.300 184.345 42.830 184.710 ;
        RECT 43.255 184.175 43.585 184.575 ;
        RECT 43.755 184.345 44.010 184.915 ;
        RECT 44.190 185.585 44.525 186.555 ;
        RECT 44.695 185.585 44.865 186.725 ;
        RECT 45.035 186.385 47.065 186.555 ;
        RECT 44.190 184.915 44.360 185.585 ;
        RECT 45.035 185.415 45.205 186.385 ;
        RECT 44.530 185.085 44.785 185.415 ;
        RECT 45.010 185.085 45.205 185.415 ;
        RECT 45.375 186.045 46.500 186.215 ;
        RECT 44.615 184.915 44.785 185.085 ;
        RECT 45.375 184.915 45.545 186.045 ;
        RECT 44.190 184.345 44.445 184.915 ;
        RECT 44.615 184.745 45.545 184.915 ;
        RECT 45.715 185.705 46.725 185.875 ;
        RECT 45.715 184.905 45.885 185.705 ;
        RECT 45.370 184.710 45.545 184.745 ;
        RECT 44.615 184.175 44.945 184.575 ;
        RECT 45.370 184.345 45.900 184.710 ;
        RECT 46.090 184.685 46.365 185.505 ;
        RECT 46.085 184.515 46.365 184.685 ;
        RECT 46.090 184.345 46.365 184.515 ;
        RECT 46.535 184.345 46.725 185.705 ;
        RECT 46.895 185.720 47.065 186.385 ;
        RECT 47.235 185.965 47.405 186.725 ;
        RECT 47.640 185.965 48.155 186.375 ;
        RECT 46.895 185.530 47.645 185.720 ;
        RECT 47.815 185.155 48.155 185.965 ;
        RECT 48.825 185.585 49.055 186.725 ;
        RECT 49.225 185.575 49.555 186.555 ;
        RECT 49.725 185.585 49.935 186.725 ;
        RECT 48.805 185.165 49.135 185.415 ;
        RECT 46.925 184.985 48.155 185.155 ;
        RECT 46.905 184.175 47.415 184.710 ;
        RECT 47.635 184.380 47.880 184.985 ;
        RECT 48.825 184.175 49.055 184.995 ;
        RECT 49.305 184.975 49.555 185.575 ;
        RECT 50.165 185.560 50.455 186.725 ;
        RECT 50.630 185.535 50.885 186.415 ;
        RECT 51.055 185.585 51.360 186.725 ;
        RECT 51.700 186.345 52.030 186.725 ;
        RECT 52.210 186.175 52.380 186.465 ;
        RECT 52.550 186.265 52.800 186.725 ;
        RECT 51.580 186.005 52.380 186.175 ;
        RECT 52.970 186.215 53.840 186.555 ;
        RECT 49.225 184.345 49.555 184.975 ;
        RECT 49.725 184.175 49.935 184.995 ;
        RECT 50.165 184.175 50.455 184.900 ;
        RECT 50.630 184.885 50.840 185.535 ;
        RECT 51.580 185.415 51.750 186.005 ;
        RECT 52.970 185.835 53.140 186.215 ;
        RECT 54.075 186.095 54.245 186.555 ;
        RECT 54.415 186.265 54.785 186.725 ;
        RECT 55.080 186.125 55.250 186.465 ;
        RECT 55.420 186.295 55.750 186.725 ;
        RECT 55.985 186.125 56.155 186.465 ;
        RECT 51.920 185.665 53.140 185.835 ;
        RECT 53.310 185.755 53.770 186.045 ;
        RECT 54.075 185.925 54.635 186.095 ;
        RECT 55.080 185.955 56.155 186.125 ;
        RECT 56.325 186.225 57.005 186.555 ;
        RECT 57.220 186.225 57.470 186.555 ;
        RECT 57.640 186.265 57.890 186.725 ;
        RECT 54.465 185.785 54.635 185.925 ;
        RECT 53.310 185.745 54.275 185.755 ;
        RECT 52.970 185.575 53.140 185.665 ;
        RECT 53.600 185.585 54.275 185.745 ;
        RECT 51.010 185.385 51.750 185.415 ;
        RECT 51.010 185.085 51.925 185.385 ;
        RECT 51.600 184.910 51.925 185.085 ;
        RECT 50.630 184.355 50.885 184.885 ;
        RECT 51.055 184.175 51.360 184.635 ;
        RECT 51.605 184.555 51.925 184.910 ;
        RECT 52.095 185.125 52.635 185.495 ;
        RECT 52.970 185.405 53.375 185.575 ;
        RECT 52.095 184.725 52.335 185.125 ;
        RECT 52.815 184.955 53.035 185.235 ;
        RECT 52.505 184.785 53.035 184.955 ;
        RECT 52.505 184.555 52.675 184.785 ;
        RECT 53.205 184.625 53.375 185.405 ;
        RECT 53.545 184.795 53.895 185.415 ;
        RECT 54.065 184.795 54.275 185.585 ;
        RECT 54.465 185.615 55.965 185.785 ;
        RECT 54.465 184.925 54.635 185.615 ;
        RECT 56.325 185.445 56.495 186.225 ;
        RECT 57.300 186.095 57.470 186.225 ;
        RECT 54.805 185.275 56.495 185.445 ;
        RECT 56.665 185.665 57.130 186.055 ;
        RECT 57.300 185.925 57.695 186.095 ;
        RECT 54.805 185.095 54.975 185.275 ;
        RECT 51.605 184.385 52.675 184.555 ;
        RECT 52.845 184.175 53.035 184.615 ;
        RECT 53.205 184.345 54.155 184.625 ;
        RECT 54.465 184.535 54.725 184.925 ;
        RECT 55.145 184.855 55.935 185.105 ;
        RECT 54.375 184.365 54.725 184.535 ;
        RECT 54.935 184.175 55.265 184.635 ;
        RECT 56.140 184.565 56.310 185.275 ;
        RECT 56.665 185.075 56.835 185.665 ;
        RECT 56.480 184.855 56.835 185.075 ;
        RECT 57.005 184.855 57.355 185.475 ;
        RECT 57.525 184.565 57.695 185.925 ;
        RECT 58.060 185.755 58.385 186.540 ;
        RECT 57.865 184.705 58.325 185.755 ;
        RECT 56.140 184.395 56.995 184.565 ;
        RECT 57.200 184.395 57.695 184.565 ;
        RECT 57.865 184.175 58.195 184.535 ;
        RECT 58.555 184.435 58.725 186.555 ;
        RECT 58.895 186.225 59.225 186.725 ;
        RECT 59.395 186.055 59.650 186.555 ;
        RECT 60.290 186.290 65.635 186.725 ;
        RECT 65.810 186.290 71.155 186.725 ;
        RECT 58.900 185.885 59.650 186.055 ;
        RECT 58.900 184.895 59.130 185.885 ;
        RECT 59.300 185.065 59.650 185.715 ;
        RECT 61.880 185.040 62.230 186.290 ;
        RECT 58.900 184.725 59.650 184.895 ;
        RECT 58.895 184.175 59.225 184.555 ;
        RECT 59.395 184.435 59.650 184.725 ;
        RECT 63.710 184.720 64.050 185.550 ;
        RECT 67.400 185.040 67.750 186.290 ;
        RECT 69.230 184.720 69.570 185.550 ;
        RECT 60.290 184.175 65.635 184.720 ;
        RECT 65.810 184.175 71.155 184.720 ;
        RECT 71.325 184.345 71.585 186.555 ;
        RECT 71.755 186.345 72.085 186.725 ;
        RECT 72.510 186.175 72.680 186.555 ;
        RECT 72.940 186.345 73.270 186.725 ;
        RECT 73.465 186.175 73.635 186.555 ;
        RECT 73.845 186.345 74.175 186.725 ;
        RECT 74.425 186.175 74.615 186.555 ;
        RECT 74.855 186.345 75.185 186.725 ;
        RECT 75.495 186.225 75.755 186.555 ;
        RECT 71.755 186.005 73.705 186.175 ;
        RECT 71.755 185.085 71.925 186.005 ;
        RECT 72.295 185.415 72.490 185.725 ;
        RECT 72.760 185.415 72.945 185.725 ;
        RECT 72.235 185.085 72.490 185.415 ;
        RECT 72.715 185.085 72.945 185.415 ;
        RECT 71.755 184.175 72.085 184.555 ;
        RECT 72.295 184.510 72.490 185.085 ;
        RECT 72.760 184.505 72.945 185.085 ;
        RECT 73.195 184.515 73.365 185.415 ;
        RECT 73.535 185.015 73.705 186.005 ;
        RECT 73.875 186.005 74.615 186.175 ;
        RECT 73.875 185.495 74.045 186.005 ;
        RECT 74.215 185.665 74.795 185.835 ;
        RECT 75.065 185.715 75.415 186.045 ;
        RECT 74.625 185.545 74.795 185.665 ;
        RECT 75.585 185.545 75.755 186.225 ;
        RECT 75.925 185.560 76.215 186.725 ;
        RECT 76.385 185.635 78.975 186.725 ;
        RECT 79.150 186.290 84.495 186.725 ;
        RECT 73.875 185.325 74.445 185.495 ;
        RECT 74.625 185.375 75.755 185.545 ;
        RECT 73.535 184.685 74.085 185.015 ;
        RECT 74.275 184.845 74.445 185.325 ;
        RECT 74.615 185.035 75.235 185.205 ;
        RECT 75.025 184.855 75.235 185.035 ;
        RECT 74.275 184.515 74.675 184.845 ;
        RECT 75.585 184.675 75.755 185.375 ;
        RECT 76.385 185.115 77.595 185.635 ;
        RECT 77.765 184.945 78.975 185.465 ;
        RECT 80.740 185.040 81.090 186.290 ;
        RECT 84.665 185.965 85.180 186.375 ;
        RECT 85.415 185.965 85.585 186.725 ;
        RECT 85.755 186.385 87.785 186.555 ;
        RECT 73.195 184.345 74.675 184.515 ;
        RECT 74.855 184.175 75.185 184.555 ;
        RECT 75.495 184.345 75.755 184.675 ;
        RECT 75.925 184.175 76.215 184.900 ;
        RECT 76.385 184.175 78.975 184.945 ;
        RECT 82.570 184.720 82.910 185.550 ;
        RECT 84.665 185.155 85.005 185.965 ;
        RECT 85.755 185.720 85.925 186.385 ;
        RECT 86.320 186.045 87.445 186.215 ;
        RECT 85.175 185.530 85.925 185.720 ;
        RECT 86.095 185.705 87.105 185.875 ;
        RECT 84.665 184.985 85.895 185.155 ;
        RECT 79.150 184.175 84.495 184.720 ;
        RECT 84.940 184.380 85.185 184.985 ;
        RECT 85.405 184.175 85.915 184.710 ;
        RECT 86.095 184.345 86.285 185.705 ;
        RECT 86.455 184.685 86.730 185.505 ;
        RECT 86.935 184.905 87.105 185.705 ;
        RECT 87.275 184.915 87.445 186.045 ;
        RECT 87.615 185.415 87.785 186.385 ;
        RECT 87.955 185.585 88.125 186.725 ;
        RECT 88.295 185.585 88.630 186.555 ;
        RECT 88.810 186.290 94.155 186.725 ;
        RECT 87.615 185.085 87.810 185.415 ;
        RECT 88.035 185.085 88.290 185.415 ;
        RECT 88.035 184.915 88.205 185.085 ;
        RECT 88.460 184.915 88.630 185.585 ;
        RECT 90.400 185.040 90.750 186.290 ;
        RECT 94.440 186.095 94.725 186.555 ;
        RECT 94.895 186.265 95.165 186.725 ;
        RECT 94.440 185.875 95.395 186.095 ;
        RECT 87.275 184.745 88.205 184.915 ;
        RECT 87.275 184.710 87.450 184.745 ;
        RECT 86.455 184.515 86.735 184.685 ;
        RECT 86.455 184.345 86.730 184.515 ;
        RECT 86.920 184.345 87.450 184.710 ;
        RECT 87.875 184.175 88.205 184.575 ;
        RECT 88.375 184.345 88.630 184.915 ;
        RECT 92.230 184.720 92.570 185.550 ;
        RECT 94.325 185.145 95.015 185.705 ;
        RECT 95.185 184.975 95.395 185.875 ;
        RECT 94.440 184.805 95.395 184.975 ;
        RECT 95.565 185.705 95.965 186.555 ;
        RECT 96.155 186.095 96.435 186.555 ;
        RECT 96.955 186.265 97.280 186.725 ;
        RECT 96.155 185.875 97.280 186.095 ;
        RECT 95.565 185.145 96.660 185.705 ;
        RECT 96.830 185.415 97.280 185.875 ;
        RECT 97.450 185.585 97.835 186.555 ;
        RECT 99.015 185.795 99.185 186.555 ;
        RECT 99.365 185.965 99.695 186.725 ;
        RECT 99.015 185.625 99.680 185.795 ;
        RECT 99.865 185.650 100.135 186.555 ;
        RECT 88.810 184.175 94.155 184.720 ;
        RECT 94.440 184.345 94.725 184.805 ;
        RECT 94.895 184.175 95.165 184.635 ;
        RECT 95.565 184.345 95.965 185.145 ;
        RECT 96.830 185.085 97.385 185.415 ;
        RECT 96.830 184.975 97.280 185.085 ;
        RECT 96.155 184.805 97.280 184.975 ;
        RECT 97.555 184.915 97.835 185.585 ;
        RECT 99.510 185.480 99.680 185.625 ;
        RECT 98.945 185.075 99.275 185.445 ;
        RECT 99.510 185.150 99.795 185.480 ;
        RECT 96.155 184.345 96.435 184.805 ;
        RECT 96.955 184.175 97.280 184.635 ;
        RECT 97.450 184.345 97.835 184.915 ;
        RECT 99.510 184.895 99.680 185.150 ;
        RECT 99.015 184.725 99.680 184.895 ;
        RECT 99.965 184.850 100.135 185.650 ;
        RECT 100.345 185.585 100.575 186.725 ;
        RECT 100.745 185.575 101.075 186.555 ;
        RECT 101.245 185.585 101.455 186.725 ;
        RECT 100.325 185.165 100.655 185.415 ;
        RECT 99.015 184.345 99.185 184.725 ;
        RECT 99.365 184.175 99.695 184.555 ;
        RECT 99.875 184.345 100.135 184.850 ;
        RECT 100.345 184.175 100.575 184.995 ;
        RECT 100.825 184.975 101.075 185.575 ;
        RECT 101.685 185.560 101.975 186.725 ;
        RECT 102.605 185.585 102.990 186.555 ;
        RECT 103.160 186.265 103.485 186.725 ;
        RECT 104.005 186.095 104.285 186.555 ;
        RECT 103.160 185.875 104.285 186.095 ;
        RECT 100.745 184.345 101.075 184.975 ;
        RECT 101.245 184.175 101.455 184.995 ;
        RECT 102.605 184.915 102.885 185.585 ;
        RECT 103.160 185.415 103.610 185.875 ;
        RECT 104.475 185.705 104.875 186.555 ;
        RECT 105.275 186.265 105.545 186.725 ;
        RECT 105.715 186.095 106.000 186.555 ;
        RECT 103.055 185.085 103.610 185.415 ;
        RECT 103.780 185.145 104.875 185.705 ;
        RECT 103.160 184.975 103.610 185.085 ;
        RECT 101.685 184.175 101.975 184.900 ;
        RECT 102.605 184.345 102.990 184.915 ;
        RECT 103.160 184.805 104.285 184.975 ;
        RECT 103.160 184.175 103.485 184.635 ;
        RECT 104.005 184.345 104.285 184.805 ;
        RECT 104.475 184.345 104.875 185.145 ;
        RECT 105.045 185.875 106.000 186.095 ;
        RECT 106.860 186.095 107.145 186.555 ;
        RECT 107.315 186.265 107.585 186.725 ;
        RECT 106.860 185.875 107.815 186.095 ;
        RECT 105.045 184.975 105.255 185.875 ;
        RECT 105.425 185.145 106.115 185.705 ;
        RECT 106.745 185.145 107.435 185.705 ;
        RECT 107.605 184.975 107.815 185.875 ;
        RECT 105.045 184.805 106.000 184.975 ;
        RECT 105.275 184.175 105.545 184.635 ;
        RECT 105.715 184.345 106.000 184.805 ;
        RECT 106.860 184.805 107.815 184.975 ;
        RECT 107.985 185.705 108.385 186.555 ;
        RECT 108.575 186.095 108.855 186.555 ;
        RECT 109.375 186.265 109.700 186.725 ;
        RECT 108.575 185.875 109.700 186.095 ;
        RECT 107.985 185.145 109.080 185.705 ;
        RECT 109.250 185.415 109.700 185.875 ;
        RECT 109.870 185.585 110.255 186.555 ;
        RECT 110.540 186.095 110.825 186.555 ;
        RECT 110.995 186.265 111.265 186.725 ;
        RECT 110.540 185.875 111.495 186.095 ;
        RECT 106.860 184.345 107.145 184.805 ;
        RECT 107.315 184.175 107.585 184.635 ;
        RECT 107.985 184.345 108.385 185.145 ;
        RECT 109.250 185.085 109.805 185.415 ;
        RECT 109.250 184.975 109.700 185.085 ;
        RECT 108.575 184.805 109.700 184.975 ;
        RECT 109.975 184.915 110.255 185.585 ;
        RECT 110.425 185.145 111.115 185.705 ;
        RECT 111.285 184.975 111.495 185.875 ;
        RECT 108.575 184.345 108.855 184.805 ;
        RECT 109.375 184.175 109.700 184.635 ;
        RECT 109.870 184.345 110.255 184.915 ;
        RECT 110.540 184.805 111.495 184.975 ;
        RECT 111.665 185.705 112.065 186.555 ;
        RECT 112.255 186.095 112.535 186.555 ;
        RECT 113.055 186.265 113.380 186.725 ;
        RECT 112.255 185.875 113.380 186.095 ;
        RECT 111.665 185.145 112.760 185.705 ;
        RECT 112.930 185.415 113.380 185.875 ;
        RECT 113.550 185.585 113.935 186.555 ;
        RECT 110.540 184.345 110.825 184.805 ;
        RECT 110.995 184.175 111.265 184.635 ;
        RECT 111.665 184.345 112.065 185.145 ;
        RECT 112.930 185.085 113.485 185.415 ;
        RECT 112.930 184.975 113.380 185.085 ;
        RECT 112.255 184.805 113.380 184.975 ;
        RECT 113.655 184.915 113.935 185.585 ;
        RECT 114.105 185.635 115.315 186.725 ;
        RECT 115.490 186.290 120.835 186.725 ;
        RECT 121.010 186.290 126.355 186.725 ;
        RECT 114.105 185.095 114.625 185.635 ;
        RECT 114.795 184.925 115.315 185.465 ;
        RECT 117.080 185.040 117.430 186.290 ;
        RECT 112.255 184.345 112.535 184.805 ;
        RECT 113.055 184.175 113.380 184.635 ;
        RECT 113.550 184.345 113.935 184.915 ;
        RECT 114.105 184.175 115.315 184.925 ;
        RECT 118.910 184.720 119.250 185.550 ;
        RECT 122.600 185.040 122.950 186.290 ;
        RECT 126.525 185.635 127.735 186.725 ;
        RECT 124.430 184.720 124.770 185.550 ;
        RECT 126.525 185.095 127.045 185.635 ;
        RECT 127.215 184.925 127.735 185.465 ;
        RECT 115.490 184.175 120.835 184.720 ;
        RECT 121.010 184.175 126.355 184.720 ;
        RECT 126.525 184.175 127.735 184.925 ;
        RECT 14.660 184.005 127.820 184.175 ;
        RECT 14.745 183.255 15.955 184.005 ;
        RECT 16.590 183.460 21.935 184.005 ;
        RECT 14.745 182.715 15.265 183.255 ;
        RECT 15.435 182.545 15.955 183.085 ;
        RECT 14.745 181.455 15.955 182.545 ;
        RECT 18.180 181.890 18.530 183.140 ;
        RECT 20.010 182.630 20.350 183.460 ;
        RECT 22.195 183.455 22.365 183.835 ;
        RECT 22.545 183.625 22.875 184.005 ;
        RECT 22.195 183.285 22.860 183.455 ;
        RECT 23.055 183.330 23.315 183.835 ;
        RECT 22.125 182.735 22.455 183.105 ;
        RECT 22.690 183.030 22.860 183.285 ;
        RECT 22.690 182.700 22.975 183.030 ;
        RECT 22.690 182.555 22.860 182.700 ;
        RECT 22.195 182.385 22.860 182.555 ;
        RECT 23.145 182.530 23.315 183.330 ;
        RECT 16.590 181.455 21.935 181.890 ;
        RECT 22.195 181.625 22.365 182.385 ;
        RECT 22.545 181.455 22.875 182.215 ;
        RECT 23.045 181.625 23.315 182.530 ;
        RECT 23.485 183.265 23.870 183.835 ;
        RECT 24.040 183.545 24.365 184.005 ;
        RECT 24.885 183.375 25.165 183.835 ;
        RECT 23.485 182.595 23.765 183.265 ;
        RECT 24.040 183.205 25.165 183.375 ;
        RECT 24.040 183.095 24.490 183.205 ;
        RECT 23.935 182.765 24.490 183.095 ;
        RECT 25.355 183.035 25.755 183.835 ;
        RECT 26.155 183.545 26.425 184.005 ;
        RECT 26.595 183.375 26.880 183.835 ;
        RECT 23.485 181.625 23.870 182.595 ;
        RECT 24.040 182.305 24.490 182.765 ;
        RECT 24.660 182.475 25.755 183.035 ;
        RECT 24.040 182.085 25.165 182.305 ;
        RECT 24.040 181.455 24.365 181.915 ;
        RECT 24.885 181.625 25.165 182.085 ;
        RECT 25.355 181.625 25.755 182.475 ;
        RECT 25.925 183.205 26.880 183.375 ;
        RECT 27.280 183.375 27.565 183.835 ;
        RECT 27.735 183.545 28.005 184.005 ;
        RECT 27.280 183.205 28.235 183.375 ;
        RECT 25.925 182.305 26.135 183.205 ;
        RECT 26.305 182.475 26.995 183.035 ;
        RECT 27.165 182.475 27.855 183.035 ;
        RECT 28.025 182.305 28.235 183.205 ;
        RECT 25.925 182.085 26.880 182.305 ;
        RECT 26.155 181.455 26.425 181.915 ;
        RECT 26.595 181.625 26.880 182.085 ;
        RECT 27.280 182.085 28.235 182.305 ;
        RECT 28.405 183.035 28.805 183.835 ;
        RECT 28.995 183.375 29.275 183.835 ;
        RECT 29.795 183.545 30.120 184.005 ;
        RECT 28.995 183.205 30.120 183.375 ;
        RECT 30.290 183.265 30.675 183.835 ;
        RECT 29.670 183.095 30.120 183.205 ;
        RECT 28.405 182.475 29.500 183.035 ;
        RECT 29.670 182.765 30.225 183.095 ;
        RECT 27.280 181.625 27.565 182.085 ;
        RECT 27.735 181.455 28.005 181.915 ;
        RECT 28.405 181.625 28.805 182.475 ;
        RECT 29.670 182.305 30.120 182.765 ;
        RECT 30.395 182.595 30.675 183.265 ;
        RECT 28.995 182.085 30.120 182.305 ;
        RECT 28.995 181.625 29.275 182.085 ;
        RECT 29.795 181.455 30.120 181.915 ;
        RECT 30.290 181.625 30.675 182.595 ;
        RECT 30.850 183.265 31.105 183.835 ;
        RECT 31.275 183.605 31.605 184.005 ;
        RECT 32.030 183.470 32.560 183.835 ;
        RECT 32.030 183.435 32.205 183.470 ;
        RECT 31.275 183.265 32.205 183.435 ;
        RECT 32.750 183.325 33.025 183.835 ;
        RECT 30.850 182.595 31.020 183.265 ;
        RECT 31.275 183.095 31.445 183.265 ;
        RECT 31.190 182.765 31.445 183.095 ;
        RECT 31.670 182.765 31.865 183.095 ;
        RECT 30.850 181.625 31.185 182.595 ;
        RECT 31.355 181.455 31.525 182.595 ;
        RECT 31.695 181.795 31.865 182.765 ;
        RECT 32.035 182.135 32.205 183.265 ;
        RECT 32.375 182.475 32.545 183.275 ;
        RECT 32.745 183.155 33.025 183.325 ;
        RECT 32.750 182.675 33.025 183.155 ;
        RECT 33.195 182.475 33.385 183.835 ;
        RECT 33.565 183.470 34.075 184.005 ;
        RECT 34.295 183.195 34.540 183.800 ;
        RECT 35.445 183.235 37.115 184.005 ;
        RECT 37.285 183.280 37.575 184.005 ;
        RECT 37.860 183.375 38.145 183.835 ;
        RECT 38.315 183.545 38.585 184.005 ;
        RECT 33.585 183.025 34.815 183.195 ;
        RECT 32.375 182.305 33.385 182.475 ;
        RECT 33.555 182.460 34.305 182.650 ;
        RECT 32.035 181.965 33.160 182.135 ;
        RECT 33.555 181.795 33.725 182.460 ;
        RECT 34.475 182.215 34.815 183.025 ;
        RECT 31.695 181.625 33.725 181.795 ;
        RECT 33.895 181.455 34.065 182.215 ;
        RECT 34.300 181.805 34.815 182.215 ;
        RECT 35.445 182.545 36.195 183.065 ;
        RECT 36.365 182.715 37.115 183.235 ;
        RECT 37.860 183.205 38.815 183.375 ;
        RECT 35.445 181.455 37.115 182.545 ;
        RECT 37.285 181.455 37.575 182.620 ;
        RECT 37.745 182.475 38.435 183.035 ;
        RECT 38.605 182.305 38.815 183.205 ;
        RECT 37.860 182.085 38.815 182.305 ;
        RECT 38.985 183.035 39.385 183.835 ;
        RECT 39.575 183.375 39.855 183.835 ;
        RECT 40.375 183.545 40.700 184.005 ;
        RECT 39.575 183.205 40.700 183.375 ;
        RECT 40.870 183.265 41.255 183.835 ;
        RECT 40.250 183.095 40.700 183.205 ;
        RECT 38.985 182.475 40.080 183.035 ;
        RECT 40.250 182.765 40.805 183.095 ;
        RECT 37.860 181.625 38.145 182.085 ;
        RECT 38.315 181.455 38.585 181.915 ;
        RECT 38.985 181.625 39.385 182.475 ;
        RECT 40.250 182.305 40.700 182.765 ;
        RECT 40.975 182.595 41.255 183.265 ;
        RECT 41.540 183.375 41.825 183.835 ;
        RECT 41.995 183.545 42.265 184.005 ;
        RECT 41.540 183.205 42.495 183.375 ;
        RECT 39.575 182.085 40.700 182.305 ;
        RECT 39.575 181.625 39.855 182.085 ;
        RECT 40.375 181.455 40.700 181.915 ;
        RECT 40.870 181.625 41.255 182.595 ;
        RECT 41.425 182.475 42.115 183.035 ;
        RECT 42.285 182.305 42.495 183.205 ;
        RECT 41.540 182.085 42.495 182.305 ;
        RECT 42.665 183.035 43.065 183.835 ;
        RECT 43.255 183.375 43.535 183.835 ;
        RECT 44.055 183.545 44.380 184.005 ;
        RECT 43.255 183.205 44.380 183.375 ;
        RECT 44.550 183.265 44.935 183.835 ;
        RECT 43.930 183.095 44.380 183.205 ;
        RECT 42.665 182.475 43.760 183.035 ;
        RECT 43.930 182.765 44.485 183.095 ;
        RECT 41.540 181.625 41.825 182.085 ;
        RECT 41.995 181.455 42.265 181.915 ;
        RECT 42.665 181.625 43.065 182.475 ;
        RECT 43.930 182.305 44.380 182.765 ;
        RECT 44.655 182.595 44.935 183.265 ;
        RECT 45.220 183.375 45.505 183.835 ;
        RECT 45.675 183.545 45.945 184.005 ;
        RECT 45.220 183.205 46.175 183.375 ;
        RECT 43.255 182.085 44.380 182.305 ;
        RECT 43.255 181.625 43.535 182.085 ;
        RECT 44.055 181.455 44.380 181.915 ;
        RECT 44.550 181.625 44.935 182.595 ;
        RECT 45.105 182.475 45.795 183.035 ;
        RECT 45.965 182.305 46.175 183.205 ;
        RECT 45.220 182.085 46.175 182.305 ;
        RECT 46.345 183.035 46.745 183.835 ;
        RECT 46.935 183.375 47.215 183.835 ;
        RECT 47.735 183.545 48.060 184.005 ;
        RECT 46.935 183.205 48.060 183.375 ;
        RECT 48.230 183.265 48.615 183.835 ;
        RECT 47.610 183.095 48.060 183.205 ;
        RECT 46.345 182.475 47.440 183.035 ;
        RECT 47.610 182.765 48.165 183.095 ;
        RECT 45.220 181.625 45.505 182.085 ;
        RECT 45.675 181.455 45.945 181.915 ;
        RECT 46.345 181.625 46.745 182.475 ;
        RECT 47.610 182.305 48.060 182.765 ;
        RECT 48.335 182.595 48.615 183.265 ;
        RECT 46.935 182.085 48.060 182.305 ;
        RECT 46.935 181.625 47.215 182.085 ;
        RECT 47.735 181.455 48.060 181.915 ;
        RECT 48.230 181.625 48.615 182.595 ;
        RECT 48.785 183.330 49.045 183.835 ;
        RECT 49.225 183.625 49.555 184.005 ;
        RECT 49.735 183.455 49.905 183.835 ;
        RECT 48.785 182.530 48.955 183.330 ;
        RECT 49.240 183.285 49.905 183.455 ;
        RECT 50.165 183.330 50.425 183.835 ;
        RECT 50.605 183.625 50.935 184.005 ;
        RECT 51.115 183.455 51.285 183.835 ;
        RECT 49.240 183.030 49.410 183.285 ;
        RECT 49.125 182.700 49.410 183.030 ;
        RECT 49.645 182.735 49.975 183.105 ;
        RECT 49.240 182.555 49.410 182.700 ;
        RECT 48.785 181.625 49.055 182.530 ;
        RECT 49.240 182.385 49.905 182.555 ;
        RECT 49.225 181.455 49.555 182.215 ;
        RECT 49.735 181.625 49.905 182.385 ;
        RECT 50.165 182.530 50.335 183.330 ;
        RECT 50.620 183.285 51.285 183.455 ;
        RECT 51.635 183.455 51.805 183.835 ;
        RECT 51.985 183.625 52.315 184.005 ;
        RECT 51.635 183.285 52.300 183.455 ;
        RECT 52.495 183.330 52.755 183.835 ;
        RECT 53.025 183.540 53.275 184.005 ;
        RECT 53.445 183.365 53.615 183.835 ;
        RECT 53.865 183.545 54.035 184.005 ;
        RECT 54.285 183.365 54.455 183.835 ;
        RECT 54.705 183.545 54.875 184.005 ;
        RECT 55.125 183.365 55.295 183.835 ;
        RECT 55.665 183.545 55.930 184.005 ;
        RECT 50.620 183.030 50.790 183.285 ;
        RECT 50.505 182.700 50.790 183.030 ;
        RECT 51.025 182.735 51.355 183.105 ;
        RECT 51.565 182.735 51.895 183.105 ;
        RECT 52.130 183.030 52.300 183.285 ;
        RECT 50.620 182.555 50.790 182.700 ;
        RECT 52.130 182.700 52.415 183.030 ;
        RECT 52.130 182.555 52.300 182.700 ;
        RECT 50.165 181.625 50.435 182.530 ;
        RECT 50.620 182.385 51.285 182.555 ;
        RECT 50.605 181.455 50.935 182.215 ;
        RECT 51.115 181.625 51.285 182.385 ;
        RECT 51.635 182.385 52.300 182.555 ;
        RECT 52.585 182.530 52.755 183.330 ;
        RECT 51.635 181.625 51.805 182.385 ;
        RECT 51.985 181.455 52.315 182.215 ;
        RECT 52.485 181.625 52.755 182.530 ;
        RECT 52.925 183.185 55.295 183.365 ;
        RECT 56.605 183.235 59.195 184.005 ;
        RECT 52.925 182.595 53.275 183.185 ;
        RECT 53.445 182.765 55.955 183.015 ;
        RECT 52.925 182.425 55.375 182.595 ;
        RECT 52.925 182.405 53.695 182.425 ;
        RECT 53.025 181.455 53.195 181.915 ;
        RECT 53.365 181.625 53.695 182.405 ;
        RECT 53.865 181.455 54.035 182.255 ;
        RECT 54.205 181.625 54.535 182.425 ;
        RECT 54.705 181.455 54.875 182.255 ;
        RECT 55.045 181.625 55.375 182.425 ;
        RECT 55.635 181.455 55.930 182.595 ;
        RECT 56.605 182.545 57.815 183.065 ;
        RECT 57.985 182.715 59.195 183.235 ;
        RECT 59.425 183.185 59.635 184.005 ;
        RECT 59.805 183.205 60.135 183.835 ;
        RECT 59.805 182.605 60.055 183.205 ;
        RECT 60.305 183.185 60.535 184.005 ;
        RECT 61.205 183.235 62.875 184.005 ;
        RECT 63.045 183.280 63.335 184.005 ;
        RECT 63.965 183.235 66.555 184.005 ;
        RECT 66.995 183.610 67.325 184.005 ;
        RECT 67.495 183.435 67.695 183.790 ;
        RECT 67.865 183.605 68.195 184.005 ;
        RECT 68.365 183.435 68.565 183.780 ;
        RECT 60.225 182.765 60.555 183.015 ;
        RECT 56.605 181.455 59.195 182.545 ;
        RECT 59.425 181.455 59.635 182.595 ;
        RECT 59.805 181.625 60.135 182.605 ;
        RECT 60.305 181.455 60.535 182.595 ;
        RECT 61.205 182.545 61.955 183.065 ;
        RECT 62.125 182.715 62.875 183.235 ;
        RECT 61.205 181.455 62.875 182.545 ;
        RECT 63.045 181.455 63.335 182.620 ;
        RECT 63.965 182.545 65.175 183.065 ;
        RECT 65.345 182.715 66.555 183.235 ;
        RECT 66.725 183.265 68.565 183.435 ;
        RECT 68.735 183.265 69.065 184.005 ;
        RECT 69.300 183.435 69.470 183.685 ;
        RECT 69.300 183.265 69.775 183.435 ;
        RECT 63.965 181.455 66.555 182.545 ;
        RECT 66.725 181.640 66.985 183.265 ;
        RECT 67.165 182.295 67.385 183.095 ;
        RECT 67.625 182.475 67.925 183.095 ;
        RECT 68.095 182.475 68.425 183.095 ;
        RECT 68.595 182.475 68.915 183.095 ;
        RECT 69.085 182.475 69.435 183.095 ;
        RECT 69.605 182.295 69.775 183.265 ;
        RECT 69.945 183.185 70.205 184.005 ;
        RECT 70.375 183.365 70.705 183.835 ;
        RECT 70.875 183.535 71.045 184.005 ;
        RECT 71.215 183.365 71.545 183.835 ;
        RECT 71.715 183.535 72.440 184.005 ;
        RECT 72.610 183.365 72.940 183.835 ;
        RECT 73.110 183.535 73.280 184.005 ;
        RECT 73.450 183.365 73.780 183.835 ;
        RECT 70.375 183.185 73.780 183.365 ;
        RECT 73.950 183.195 74.155 184.005 ;
        RECT 73.575 183.015 73.780 183.185 ;
        RECT 74.325 183.185 74.680 183.710 ;
        RECT 74.850 183.265 75.100 184.005 ;
        RECT 75.770 183.435 75.940 183.685 ;
        RECT 75.465 183.265 75.940 183.435 ;
        RECT 76.175 183.265 76.505 184.005 ;
        RECT 76.675 183.435 76.875 183.780 ;
        RECT 77.045 183.605 77.375 184.005 ;
        RECT 77.545 183.435 77.745 183.790 ;
        RECT 77.915 183.610 78.245 184.005 ;
        RECT 76.675 183.265 78.515 183.435 ;
        RECT 74.325 183.015 74.495 183.185 ;
        RECT 69.960 182.805 71.100 183.015 ;
        RECT 71.280 182.805 72.495 183.015 ;
        RECT 72.675 182.805 73.395 183.015 ;
        RECT 73.575 182.635 73.895 183.015 ;
        RECT 74.180 182.845 74.495 183.015 ;
        RECT 67.165 182.085 69.775 182.295 ;
        RECT 69.945 182.465 71.965 182.635 ;
        RECT 68.735 181.455 69.065 181.905 ;
        RECT 69.945 181.625 70.285 182.465 ;
        RECT 70.455 181.455 70.665 182.295 ;
        RECT 70.835 181.625 71.085 182.465 ;
        RECT 71.255 181.795 71.465 182.295 ;
        RECT 71.635 181.965 71.965 182.465 ;
        RECT 72.135 182.465 73.320 182.635 ;
        RECT 72.135 181.965 72.520 182.465 ;
        RECT 72.690 181.795 72.900 182.295 ;
        RECT 71.255 181.625 72.900 181.795 ;
        RECT 73.070 181.795 73.320 182.465 ;
        RECT 73.490 182.465 73.895 182.635 ;
        RECT 73.490 181.965 73.740 182.465 ;
        RECT 73.910 181.795 74.155 182.295 ;
        RECT 73.070 181.625 74.155 181.795 ;
        RECT 74.325 182.055 74.495 182.845 ;
        RECT 74.665 182.805 75.295 183.015 ;
        RECT 75.045 182.135 75.295 182.805 ;
        RECT 75.465 182.295 75.635 183.265 ;
        RECT 75.805 182.475 76.155 183.095 ;
        RECT 76.325 182.475 76.645 183.095 ;
        RECT 76.815 182.475 77.145 183.095 ;
        RECT 77.315 182.475 77.615 183.095 ;
        RECT 77.855 182.295 78.075 183.095 ;
        RECT 75.465 182.085 78.075 182.295 ;
        RECT 74.325 181.640 74.680 182.055 ;
        RECT 74.850 181.455 75.100 181.955 ;
        RECT 76.175 181.455 76.505 181.905 ;
        RECT 78.255 181.640 78.515 183.265 ;
        RECT 79.610 183.295 79.865 183.825 ;
        RECT 80.035 183.545 80.340 184.005 ;
        RECT 80.585 183.625 81.655 183.795 ;
        RECT 79.610 182.645 79.820 183.295 ;
        RECT 80.585 183.270 80.905 183.625 ;
        RECT 80.580 183.095 80.905 183.270 ;
        RECT 79.990 182.795 80.905 183.095 ;
        RECT 81.075 183.055 81.315 183.455 ;
        RECT 81.485 183.395 81.655 183.625 ;
        RECT 81.825 183.565 82.015 184.005 ;
        RECT 82.185 183.555 83.135 183.835 ;
        RECT 83.355 183.645 83.705 183.815 ;
        RECT 81.485 183.225 82.015 183.395 ;
        RECT 79.990 182.765 80.730 182.795 ;
        RECT 79.610 181.765 79.865 182.645 ;
        RECT 80.035 181.455 80.340 182.595 ;
        RECT 80.560 182.175 80.730 182.765 ;
        RECT 81.075 182.685 81.615 183.055 ;
        RECT 81.795 182.945 82.015 183.225 ;
        RECT 82.185 182.775 82.355 183.555 ;
        RECT 81.950 182.605 82.355 182.775 ;
        RECT 82.525 182.765 82.875 183.385 ;
        RECT 81.950 182.515 82.120 182.605 ;
        RECT 83.045 182.595 83.255 183.385 ;
        RECT 80.900 182.345 82.120 182.515 ;
        RECT 82.580 182.435 83.255 182.595 ;
        RECT 80.560 182.005 81.360 182.175 ;
        RECT 80.680 181.455 81.010 181.835 ;
        RECT 81.190 181.715 81.360 182.005 ;
        RECT 81.950 181.965 82.120 182.345 ;
        RECT 82.290 182.425 83.255 182.435 ;
        RECT 83.445 183.255 83.705 183.645 ;
        RECT 83.915 183.545 84.245 184.005 ;
        RECT 85.120 183.615 85.975 183.785 ;
        RECT 86.180 183.615 86.675 183.785 ;
        RECT 86.845 183.645 87.175 184.005 ;
        RECT 83.445 182.565 83.615 183.255 ;
        RECT 83.785 182.905 83.955 183.085 ;
        RECT 84.125 183.075 84.915 183.325 ;
        RECT 85.120 182.905 85.290 183.615 ;
        RECT 85.460 183.105 85.815 183.325 ;
        RECT 83.785 182.735 85.475 182.905 ;
        RECT 82.290 182.135 82.750 182.425 ;
        RECT 83.445 182.395 84.945 182.565 ;
        RECT 83.445 182.255 83.615 182.395 ;
        RECT 83.055 182.085 83.615 182.255 ;
        RECT 81.530 181.455 81.780 181.915 ;
        RECT 81.950 181.625 82.820 181.965 ;
        RECT 83.055 181.625 83.225 182.085 ;
        RECT 84.060 182.055 85.135 182.225 ;
        RECT 83.395 181.455 83.765 181.915 ;
        RECT 84.060 181.715 84.230 182.055 ;
        RECT 84.400 181.455 84.730 181.885 ;
        RECT 84.965 181.715 85.135 182.055 ;
        RECT 85.305 181.955 85.475 182.735 ;
        RECT 85.645 182.515 85.815 183.105 ;
        RECT 85.985 182.705 86.335 183.325 ;
        RECT 85.645 182.125 86.110 182.515 ;
        RECT 86.505 182.255 86.675 183.615 ;
        RECT 86.845 182.425 87.305 183.475 ;
        RECT 86.280 182.085 86.675 182.255 ;
        RECT 86.280 181.955 86.450 182.085 ;
        RECT 85.305 181.625 85.985 181.955 ;
        RECT 86.200 181.625 86.450 181.955 ;
        RECT 86.620 181.455 86.870 181.915 ;
        RECT 87.040 181.640 87.365 182.425 ;
        RECT 87.535 181.625 87.705 183.745 ;
        RECT 87.875 183.625 88.205 184.005 ;
        RECT 88.375 183.455 88.630 183.745 ;
        RECT 87.880 183.285 88.630 183.455 ;
        RECT 87.880 182.295 88.110 183.285 ;
        RECT 88.805 183.280 89.095 184.005 ;
        RECT 89.325 183.185 89.535 184.005 ;
        RECT 89.705 183.205 90.035 183.835 ;
        RECT 88.280 182.465 88.630 183.115 ;
        RECT 87.880 182.125 88.630 182.295 ;
        RECT 87.875 181.455 88.205 181.955 ;
        RECT 88.375 181.625 88.630 182.125 ;
        RECT 88.805 181.455 89.095 182.620 ;
        RECT 89.705 182.605 89.955 183.205 ;
        RECT 90.205 183.185 90.435 184.005 ;
        RECT 90.645 183.255 91.855 184.005 ;
        RECT 90.125 182.765 90.455 183.015 ;
        RECT 89.325 181.455 89.535 182.595 ;
        RECT 89.705 181.625 90.035 182.605 ;
        RECT 90.205 181.455 90.435 182.595 ;
        RECT 90.645 182.545 91.165 183.085 ;
        RECT 91.335 182.715 91.855 183.255 ;
        RECT 92.025 183.235 95.535 184.005 ;
        RECT 92.025 182.545 93.715 183.065 ;
        RECT 93.885 182.715 95.535 183.235 ;
        RECT 95.980 183.195 96.225 183.800 ;
        RECT 96.445 183.470 96.955 184.005 ;
        RECT 95.705 183.025 96.935 183.195 ;
        RECT 90.645 181.455 91.855 182.545 ;
        RECT 92.025 181.455 95.535 182.545 ;
        RECT 95.705 182.215 96.045 183.025 ;
        RECT 96.215 182.460 96.965 182.650 ;
        RECT 95.705 181.805 96.220 182.215 ;
        RECT 96.455 181.455 96.625 182.215 ;
        RECT 96.795 181.795 96.965 182.460 ;
        RECT 97.135 182.475 97.325 183.835 ;
        RECT 97.495 183.665 97.770 183.835 ;
        RECT 97.495 183.495 97.775 183.665 ;
        RECT 97.495 182.675 97.770 183.495 ;
        RECT 97.960 183.470 98.490 183.835 ;
        RECT 98.915 183.605 99.245 184.005 ;
        RECT 98.315 183.435 98.490 183.470 ;
        RECT 97.975 182.475 98.145 183.275 ;
        RECT 97.135 182.305 98.145 182.475 ;
        RECT 98.315 183.265 99.245 183.435 ;
        RECT 99.415 183.265 99.670 183.835 ;
        RECT 98.315 182.135 98.485 183.265 ;
        RECT 99.075 183.095 99.245 183.265 ;
        RECT 97.360 181.965 98.485 182.135 ;
        RECT 98.655 182.765 98.850 183.095 ;
        RECT 99.075 182.765 99.330 183.095 ;
        RECT 98.655 181.795 98.825 182.765 ;
        RECT 99.500 182.595 99.670 183.265 ;
        RECT 99.845 183.235 102.435 184.005 ;
        RECT 96.795 181.625 98.825 181.795 ;
        RECT 98.995 181.455 99.165 182.595 ;
        RECT 99.335 181.625 99.670 182.595 ;
        RECT 99.845 182.545 101.055 183.065 ;
        RECT 101.225 182.715 102.435 183.235 ;
        RECT 102.880 183.195 103.125 183.800 ;
        RECT 103.345 183.470 103.855 184.005 ;
        RECT 102.605 183.025 103.835 183.195 ;
        RECT 99.845 181.455 102.435 182.545 ;
        RECT 102.605 182.215 102.945 183.025 ;
        RECT 103.115 182.460 103.865 182.650 ;
        RECT 102.605 181.805 103.120 182.215 ;
        RECT 103.355 181.455 103.525 182.215 ;
        RECT 103.695 181.795 103.865 182.460 ;
        RECT 104.035 182.475 104.225 183.835 ;
        RECT 104.395 183.325 104.670 183.835 ;
        RECT 104.860 183.470 105.390 183.835 ;
        RECT 105.815 183.605 106.145 184.005 ;
        RECT 105.215 183.435 105.390 183.470 ;
        RECT 104.395 183.155 104.675 183.325 ;
        RECT 104.395 182.675 104.670 183.155 ;
        RECT 104.875 182.475 105.045 183.275 ;
        RECT 104.035 182.305 105.045 182.475 ;
        RECT 105.215 183.265 106.145 183.435 ;
        RECT 106.315 183.265 106.570 183.835 ;
        RECT 105.215 182.135 105.385 183.265 ;
        RECT 105.975 183.095 106.145 183.265 ;
        RECT 104.260 181.965 105.385 182.135 ;
        RECT 105.555 182.765 105.750 183.095 ;
        RECT 105.975 182.765 106.230 183.095 ;
        RECT 105.555 181.795 105.725 182.765 ;
        RECT 106.400 182.595 106.570 183.265 ;
        RECT 103.695 181.625 105.725 181.795 ;
        RECT 105.895 181.455 106.065 182.595 ;
        RECT 106.235 181.625 106.570 182.595 ;
        RECT 106.745 183.205 107.085 183.835 ;
        RECT 107.255 183.205 107.505 184.005 ;
        RECT 107.695 183.355 108.025 183.835 ;
        RECT 108.195 183.545 108.420 184.005 ;
        RECT 108.590 183.355 108.920 183.835 ;
        RECT 106.745 182.645 106.920 183.205 ;
        RECT 107.695 183.185 108.920 183.355 ;
        RECT 109.550 183.225 110.050 183.835 ;
        RECT 107.090 182.845 107.785 183.015 ;
        RECT 106.745 182.595 106.975 182.645 ;
        RECT 107.615 182.595 107.785 182.845 ;
        RECT 107.960 182.815 108.380 183.015 ;
        RECT 108.550 182.815 108.880 183.015 ;
        RECT 109.050 182.815 109.380 183.015 ;
        RECT 109.550 182.595 109.720 183.225 ;
        RECT 110.700 183.195 110.945 183.800 ;
        RECT 111.165 183.470 111.675 184.005 ;
        RECT 110.425 183.025 111.655 183.195 ;
        RECT 109.905 182.765 110.255 183.015 ;
        RECT 106.745 181.625 107.085 182.595 ;
        RECT 107.255 181.455 107.425 182.595 ;
        RECT 107.615 182.425 110.050 182.595 ;
        RECT 107.695 181.455 107.945 182.255 ;
        RECT 108.590 181.625 108.920 182.425 ;
        RECT 109.220 181.455 109.550 182.255 ;
        RECT 109.720 181.625 110.050 182.425 ;
        RECT 110.425 182.215 110.765 183.025 ;
        RECT 110.935 182.460 111.685 182.650 ;
        RECT 110.425 181.805 110.940 182.215 ;
        RECT 111.175 181.455 111.345 182.215 ;
        RECT 111.515 181.795 111.685 182.460 ;
        RECT 111.855 182.475 112.045 183.835 ;
        RECT 112.215 182.985 112.490 183.835 ;
        RECT 112.680 183.470 113.210 183.835 ;
        RECT 113.635 183.605 113.965 184.005 ;
        RECT 113.035 183.435 113.210 183.470 ;
        RECT 112.215 182.815 112.495 182.985 ;
        RECT 112.215 182.675 112.490 182.815 ;
        RECT 112.695 182.475 112.865 183.275 ;
        RECT 111.855 182.305 112.865 182.475 ;
        RECT 113.035 183.265 113.965 183.435 ;
        RECT 114.135 183.265 114.390 183.835 ;
        RECT 114.565 183.280 114.855 184.005 ;
        RECT 115.950 183.295 116.205 183.825 ;
        RECT 116.375 183.545 116.680 184.005 ;
        RECT 116.925 183.625 117.995 183.795 ;
        RECT 113.035 182.135 113.205 183.265 ;
        RECT 113.795 183.095 113.965 183.265 ;
        RECT 112.080 181.965 113.205 182.135 ;
        RECT 113.375 182.765 113.570 183.095 ;
        RECT 113.795 182.765 114.050 183.095 ;
        RECT 113.375 181.795 113.545 182.765 ;
        RECT 114.220 182.595 114.390 183.265 ;
        RECT 115.950 182.645 116.160 183.295 ;
        RECT 116.925 183.270 117.245 183.625 ;
        RECT 116.920 183.095 117.245 183.270 ;
        RECT 116.330 182.795 117.245 183.095 ;
        RECT 117.415 183.055 117.655 183.455 ;
        RECT 117.825 183.395 117.995 183.625 ;
        RECT 118.165 183.565 118.355 184.005 ;
        RECT 118.525 183.555 119.475 183.835 ;
        RECT 119.695 183.645 120.045 183.815 ;
        RECT 117.825 183.225 118.355 183.395 ;
        RECT 116.330 182.765 117.070 182.795 ;
        RECT 111.515 181.625 113.545 181.795 ;
        RECT 113.715 181.455 113.885 182.595 ;
        RECT 114.055 181.625 114.390 182.595 ;
        RECT 114.565 181.455 114.855 182.620 ;
        RECT 115.950 181.765 116.205 182.645 ;
        RECT 116.375 181.455 116.680 182.595 ;
        RECT 116.900 182.175 117.070 182.765 ;
        RECT 117.415 182.685 117.955 183.055 ;
        RECT 118.135 182.945 118.355 183.225 ;
        RECT 118.525 182.775 118.695 183.555 ;
        RECT 118.290 182.605 118.695 182.775 ;
        RECT 118.865 182.765 119.215 183.385 ;
        RECT 118.290 182.515 118.460 182.605 ;
        RECT 119.385 182.595 119.595 183.385 ;
        RECT 117.240 182.345 118.460 182.515 ;
        RECT 118.920 182.435 119.595 182.595 ;
        RECT 116.900 182.005 117.700 182.175 ;
        RECT 117.020 181.455 117.350 181.835 ;
        RECT 117.530 181.715 117.700 182.005 ;
        RECT 118.290 181.965 118.460 182.345 ;
        RECT 118.630 182.425 119.595 182.435 ;
        RECT 119.785 183.255 120.045 183.645 ;
        RECT 120.255 183.545 120.585 184.005 ;
        RECT 121.460 183.615 122.315 183.785 ;
        RECT 122.520 183.615 123.015 183.785 ;
        RECT 123.185 183.645 123.515 184.005 ;
        RECT 119.785 182.565 119.955 183.255 ;
        RECT 120.125 182.905 120.295 183.085 ;
        RECT 120.465 183.075 121.255 183.325 ;
        RECT 121.460 182.905 121.630 183.615 ;
        RECT 121.800 183.105 122.155 183.325 ;
        RECT 120.125 182.735 121.815 182.905 ;
        RECT 118.630 182.135 119.090 182.425 ;
        RECT 119.785 182.395 121.285 182.565 ;
        RECT 119.785 182.255 119.955 182.395 ;
        RECT 119.395 182.085 119.955 182.255 ;
        RECT 117.870 181.455 118.120 181.915 ;
        RECT 118.290 181.625 119.160 181.965 ;
        RECT 119.395 181.625 119.565 182.085 ;
        RECT 120.400 182.055 121.475 182.225 ;
        RECT 119.735 181.455 120.105 181.915 ;
        RECT 120.400 181.715 120.570 182.055 ;
        RECT 120.740 181.455 121.070 181.885 ;
        RECT 121.305 181.715 121.475 182.055 ;
        RECT 121.645 181.955 121.815 182.735 ;
        RECT 121.985 182.515 122.155 183.105 ;
        RECT 122.325 182.705 122.675 183.325 ;
        RECT 121.985 182.125 122.450 182.515 ;
        RECT 122.845 182.255 123.015 183.615 ;
        RECT 123.185 182.425 123.645 183.475 ;
        RECT 122.620 182.085 123.015 182.255 ;
        RECT 122.620 181.955 122.790 182.085 ;
        RECT 121.645 181.625 122.325 181.955 ;
        RECT 122.540 181.625 122.790 181.955 ;
        RECT 122.960 181.455 123.210 181.915 ;
        RECT 123.380 181.640 123.705 182.425 ;
        RECT 123.875 181.625 124.045 183.745 ;
        RECT 124.215 183.625 124.545 184.005 ;
        RECT 124.715 183.455 124.970 183.745 ;
        RECT 124.220 183.285 124.970 183.455 ;
        RECT 124.220 182.295 124.450 183.285 ;
        RECT 125.145 183.255 126.355 184.005 ;
        RECT 126.525 183.255 127.735 184.005 ;
        RECT 124.620 182.465 124.970 183.115 ;
        RECT 125.145 182.545 125.665 183.085 ;
        RECT 125.835 182.715 126.355 183.255 ;
        RECT 126.525 182.545 127.045 183.085 ;
        RECT 127.215 182.715 127.735 183.255 ;
        RECT 124.220 182.125 124.970 182.295 ;
        RECT 124.215 181.455 124.545 181.955 ;
        RECT 124.715 181.625 124.970 182.125 ;
        RECT 125.145 181.455 126.355 182.545 ;
        RECT 126.525 181.455 127.735 182.545 ;
        RECT 14.660 181.285 127.820 181.455 ;
        RECT 14.745 180.195 15.955 181.285 ;
        RECT 14.745 179.485 15.265 180.025 ;
        RECT 15.435 179.655 15.955 180.195 ;
        RECT 16.125 180.195 18.715 181.285 ;
        RECT 18.890 180.850 24.235 181.285 ;
        RECT 16.125 179.675 17.335 180.195 ;
        RECT 17.505 179.505 18.715 180.025 ;
        RECT 20.480 179.600 20.830 180.850 ;
        RECT 24.405 180.120 24.695 181.285 ;
        RECT 24.870 180.615 25.125 181.115 ;
        RECT 25.295 180.785 25.625 181.285 ;
        RECT 24.870 180.445 25.620 180.615 ;
        RECT 14.745 178.735 15.955 179.485 ;
        RECT 16.125 178.735 18.715 179.505 ;
        RECT 22.310 179.280 22.650 180.110 ;
        RECT 24.870 179.625 25.220 180.275 ;
        RECT 18.890 178.735 24.235 179.280 ;
        RECT 24.405 178.735 24.695 179.460 ;
        RECT 25.390 179.455 25.620 180.445 ;
        RECT 24.870 179.285 25.620 179.455 ;
        RECT 24.870 178.995 25.125 179.285 ;
        RECT 25.295 178.735 25.625 179.115 ;
        RECT 25.795 178.995 25.965 181.115 ;
        RECT 26.135 180.315 26.460 181.100 ;
        RECT 26.630 180.825 26.880 181.285 ;
        RECT 27.050 180.785 27.300 181.115 ;
        RECT 27.515 180.785 28.195 181.115 ;
        RECT 27.050 180.655 27.220 180.785 ;
        RECT 26.825 180.485 27.220 180.655 ;
        RECT 26.195 179.265 26.655 180.315 ;
        RECT 26.825 179.125 26.995 180.485 ;
        RECT 27.390 180.225 27.855 180.615 ;
        RECT 27.165 179.415 27.515 180.035 ;
        RECT 27.685 179.635 27.855 180.225 ;
        RECT 28.025 180.005 28.195 180.785 ;
        RECT 28.365 180.685 28.535 181.025 ;
        RECT 28.770 180.855 29.100 181.285 ;
        RECT 29.270 180.685 29.440 181.025 ;
        RECT 29.735 180.825 30.105 181.285 ;
        RECT 28.365 180.515 29.440 180.685 ;
        RECT 30.275 180.655 30.445 181.115 ;
        RECT 30.680 180.775 31.550 181.115 ;
        RECT 31.720 180.825 31.970 181.285 ;
        RECT 29.885 180.485 30.445 180.655 ;
        RECT 29.885 180.345 30.055 180.485 ;
        RECT 28.555 180.175 30.055 180.345 ;
        RECT 30.750 180.315 31.210 180.605 ;
        RECT 28.025 179.835 29.715 180.005 ;
        RECT 27.685 179.415 28.040 179.635 ;
        RECT 28.210 179.125 28.380 179.835 ;
        RECT 28.585 179.415 29.375 179.665 ;
        RECT 29.545 179.655 29.715 179.835 ;
        RECT 29.885 179.485 30.055 180.175 ;
        RECT 26.325 178.735 26.655 179.095 ;
        RECT 26.825 178.955 27.320 179.125 ;
        RECT 27.525 178.955 28.380 179.125 ;
        RECT 29.255 178.735 29.585 179.195 ;
        RECT 29.795 179.095 30.055 179.485 ;
        RECT 30.245 180.305 31.210 180.315 ;
        RECT 31.380 180.395 31.550 180.775 ;
        RECT 32.140 180.735 32.310 181.025 ;
        RECT 32.490 180.905 32.820 181.285 ;
        RECT 32.140 180.565 32.940 180.735 ;
        RECT 30.245 180.145 30.920 180.305 ;
        RECT 31.380 180.225 32.600 180.395 ;
        RECT 30.245 179.355 30.455 180.145 ;
        RECT 31.380 180.135 31.550 180.225 ;
        RECT 30.625 179.355 30.975 179.975 ;
        RECT 31.145 179.965 31.550 180.135 ;
        RECT 31.145 179.185 31.315 179.965 ;
        RECT 31.485 179.515 31.705 179.795 ;
        RECT 31.885 179.685 32.425 180.055 ;
        RECT 32.770 179.975 32.940 180.565 ;
        RECT 33.160 180.145 33.465 181.285 ;
        RECT 33.635 180.095 33.890 180.975 ;
        RECT 32.770 179.945 33.510 179.975 ;
        RECT 31.485 179.345 32.015 179.515 ;
        RECT 29.795 178.925 30.145 179.095 ;
        RECT 30.365 178.905 31.315 179.185 ;
        RECT 31.485 178.735 31.675 179.175 ;
        RECT 31.845 179.115 32.015 179.345 ;
        RECT 32.185 179.285 32.425 179.685 ;
        RECT 32.595 179.645 33.510 179.945 ;
        RECT 32.595 179.470 32.920 179.645 ;
        RECT 32.595 179.115 32.915 179.470 ;
        RECT 33.680 179.445 33.890 180.095 ;
        RECT 31.845 178.945 32.915 179.115 ;
        RECT 33.160 178.735 33.465 179.195 ;
        RECT 33.635 178.915 33.890 179.445 ;
        RECT 34.065 180.145 34.450 181.115 ;
        RECT 34.620 180.825 34.945 181.285 ;
        RECT 35.465 180.655 35.745 181.115 ;
        RECT 34.620 180.435 35.745 180.655 ;
        RECT 34.065 179.475 34.345 180.145 ;
        RECT 34.620 179.975 35.070 180.435 ;
        RECT 35.935 180.265 36.335 181.115 ;
        RECT 36.735 180.825 37.005 181.285 ;
        RECT 37.175 180.655 37.460 181.115 ;
        RECT 34.515 179.645 35.070 179.975 ;
        RECT 35.240 179.705 36.335 180.265 ;
        RECT 34.620 179.535 35.070 179.645 ;
        RECT 34.065 178.905 34.450 179.475 ;
        RECT 34.620 179.365 35.745 179.535 ;
        RECT 34.620 178.735 34.945 179.195 ;
        RECT 35.465 178.905 35.745 179.365 ;
        RECT 35.935 178.905 36.335 179.705 ;
        RECT 36.505 180.435 37.460 180.655 ;
        RECT 36.505 179.535 36.715 180.435 ;
        RECT 36.885 179.705 37.575 180.265 ;
        RECT 38.205 180.145 38.545 181.115 ;
        RECT 38.715 180.145 38.885 181.285 ;
        RECT 39.155 180.485 39.405 181.285 ;
        RECT 40.050 180.315 40.380 181.115 ;
        RECT 40.680 180.485 41.010 181.285 ;
        RECT 41.180 180.315 41.510 181.115 ;
        RECT 39.075 180.145 41.510 180.315 ;
        RECT 42.345 180.145 42.685 181.115 ;
        RECT 42.855 180.145 43.025 181.285 ;
        RECT 43.295 180.485 43.545 181.285 ;
        RECT 44.190 180.315 44.520 181.115 ;
        RECT 44.820 180.485 45.150 181.285 ;
        RECT 45.320 180.315 45.650 181.115 ;
        RECT 43.215 180.145 45.650 180.315 ;
        RECT 46.025 180.525 46.540 180.935 ;
        RECT 46.775 180.525 46.945 181.285 ;
        RECT 47.115 180.945 49.145 181.115 ;
        RECT 38.205 179.585 38.380 180.145 ;
        RECT 39.075 179.895 39.245 180.145 ;
        RECT 38.550 179.725 39.245 179.895 ;
        RECT 39.420 179.725 39.840 179.925 ;
        RECT 40.010 179.725 40.340 179.925 ;
        RECT 40.510 179.725 40.840 179.925 ;
        RECT 38.205 179.535 38.435 179.585 ;
        RECT 36.505 179.365 37.460 179.535 ;
        RECT 36.735 178.735 37.005 179.195 ;
        RECT 37.175 178.905 37.460 179.365 ;
        RECT 38.205 178.905 38.545 179.535 ;
        RECT 38.715 178.735 38.965 179.535 ;
        RECT 39.155 179.385 40.380 179.555 ;
        RECT 39.155 178.905 39.485 179.385 ;
        RECT 39.655 178.735 39.880 179.195 ;
        RECT 40.050 178.905 40.380 179.385 ;
        RECT 41.010 179.515 41.180 180.145 ;
        RECT 41.365 179.725 41.715 179.975 ;
        RECT 42.345 179.535 42.520 180.145 ;
        RECT 43.215 179.895 43.385 180.145 ;
        RECT 42.690 179.725 43.385 179.895 ;
        RECT 43.560 179.725 43.980 179.925 ;
        RECT 44.150 179.725 44.480 179.925 ;
        RECT 44.650 179.725 44.980 179.925 ;
        RECT 41.010 178.905 41.510 179.515 ;
        RECT 42.345 178.905 42.685 179.535 ;
        RECT 42.855 178.735 43.105 179.535 ;
        RECT 43.295 179.385 44.520 179.555 ;
        RECT 43.295 178.905 43.625 179.385 ;
        RECT 43.795 178.735 44.020 179.195 ;
        RECT 44.190 178.905 44.520 179.385 ;
        RECT 45.150 179.515 45.320 180.145 ;
        RECT 45.505 179.725 45.855 179.975 ;
        RECT 46.025 179.715 46.365 180.525 ;
        RECT 47.115 180.280 47.285 180.945 ;
        RECT 47.680 180.605 48.805 180.775 ;
        RECT 46.535 180.090 47.285 180.280 ;
        RECT 47.455 180.265 48.465 180.435 ;
        RECT 46.025 179.545 47.255 179.715 ;
        RECT 45.150 178.905 45.650 179.515 ;
        RECT 46.300 178.940 46.545 179.545 ;
        RECT 46.765 178.735 47.275 179.270 ;
        RECT 47.455 178.905 47.645 180.265 ;
        RECT 47.815 179.245 48.090 180.065 ;
        RECT 48.295 179.465 48.465 180.265 ;
        RECT 48.635 179.475 48.805 180.605 ;
        RECT 48.975 179.975 49.145 180.945 ;
        RECT 49.315 180.145 49.485 181.285 ;
        RECT 49.655 180.145 49.990 181.115 ;
        RECT 48.975 179.645 49.170 179.975 ;
        RECT 49.395 179.645 49.650 179.975 ;
        RECT 49.395 179.475 49.565 179.645 ;
        RECT 49.820 179.475 49.990 180.145 ;
        RECT 50.165 180.120 50.455 181.285 ;
        RECT 50.740 180.655 51.025 181.115 ;
        RECT 51.195 180.825 51.465 181.285 ;
        RECT 50.740 180.435 51.695 180.655 ;
        RECT 50.625 179.705 51.315 180.265 ;
        RECT 51.485 179.535 51.695 180.435 ;
        RECT 48.635 179.305 49.565 179.475 ;
        RECT 48.635 179.270 48.810 179.305 ;
        RECT 47.815 179.075 48.095 179.245 ;
        RECT 47.815 178.905 48.090 179.075 ;
        RECT 48.280 178.905 48.810 179.270 ;
        RECT 49.235 178.735 49.565 179.135 ;
        RECT 49.735 178.905 49.990 179.475 ;
        RECT 50.165 178.735 50.455 179.460 ;
        RECT 50.740 179.365 51.695 179.535 ;
        RECT 51.865 180.265 52.265 181.115 ;
        RECT 52.455 180.655 52.735 181.115 ;
        RECT 53.255 180.825 53.580 181.285 ;
        RECT 52.455 180.435 53.580 180.655 ;
        RECT 51.865 179.705 52.960 180.265 ;
        RECT 53.130 179.975 53.580 180.435 ;
        RECT 53.750 180.145 54.135 181.115 ;
        RECT 50.740 178.905 51.025 179.365 ;
        RECT 51.195 178.735 51.465 179.195 ;
        RECT 51.865 178.905 52.265 179.705 ;
        RECT 53.130 179.645 53.685 179.975 ;
        RECT 53.130 179.535 53.580 179.645 ;
        RECT 52.455 179.365 53.580 179.535 ;
        RECT 53.855 179.475 54.135 180.145 ;
        RECT 54.305 180.195 55.975 181.285 ;
        RECT 54.305 179.675 55.055 180.195 ;
        RECT 56.150 180.145 56.485 181.115 ;
        RECT 56.655 180.145 56.825 181.285 ;
        RECT 56.995 180.945 59.025 181.115 ;
        RECT 55.225 179.505 55.975 180.025 ;
        RECT 52.455 178.905 52.735 179.365 ;
        RECT 53.255 178.735 53.580 179.195 ;
        RECT 53.750 178.905 54.135 179.475 ;
        RECT 54.305 178.735 55.975 179.505 ;
        RECT 56.150 179.475 56.320 180.145 ;
        RECT 56.995 179.975 57.165 180.945 ;
        RECT 56.490 179.645 56.745 179.975 ;
        RECT 56.970 179.645 57.165 179.975 ;
        RECT 57.335 180.605 58.460 180.775 ;
        RECT 56.575 179.475 56.745 179.645 ;
        RECT 57.335 179.475 57.505 180.605 ;
        RECT 56.150 178.905 56.405 179.475 ;
        RECT 56.575 179.305 57.505 179.475 ;
        RECT 57.675 180.265 58.685 180.435 ;
        RECT 57.675 179.465 57.845 180.265 ;
        RECT 57.330 179.270 57.505 179.305 ;
        RECT 56.575 178.735 56.905 179.135 ;
        RECT 57.330 178.905 57.860 179.270 ;
        RECT 58.050 179.245 58.325 180.065 ;
        RECT 58.045 179.075 58.325 179.245 ;
        RECT 58.050 178.905 58.325 179.075 ;
        RECT 58.495 178.905 58.685 180.265 ;
        RECT 58.855 180.280 59.025 180.945 ;
        RECT 59.195 180.525 59.365 181.285 ;
        RECT 59.600 180.525 60.115 180.935 ;
        RECT 58.855 180.090 59.605 180.280 ;
        RECT 59.775 179.715 60.115 180.525 ;
        RECT 60.340 180.415 60.625 181.285 ;
        RECT 60.795 180.655 61.055 181.115 ;
        RECT 61.230 180.825 61.485 181.285 ;
        RECT 61.655 180.655 61.915 181.115 ;
        RECT 60.795 180.485 61.915 180.655 ;
        RECT 62.085 180.485 62.395 181.285 ;
        RECT 60.795 180.235 61.055 180.485 ;
        RECT 62.565 180.315 62.875 181.115 ;
        RECT 58.885 179.545 60.115 179.715 ;
        RECT 60.300 180.065 61.055 180.235 ;
        RECT 61.845 180.145 62.875 180.315 ;
        RECT 60.300 179.555 60.705 180.065 ;
        RECT 61.845 179.895 62.015 180.145 ;
        RECT 60.875 179.725 62.015 179.895 ;
        RECT 58.865 178.735 59.375 179.270 ;
        RECT 59.595 178.940 59.840 179.545 ;
        RECT 60.300 179.385 61.950 179.555 ;
        RECT 62.185 179.405 62.535 179.975 ;
        RECT 60.345 178.735 60.625 179.215 ;
        RECT 60.795 178.995 61.055 179.385 ;
        RECT 61.230 178.735 61.485 179.215 ;
        RECT 61.655 178.995 61.950 179.385 ;
        RECT 62.705 179.235 62.875 180.145 ;
        RECT 63.045 180.195 65.635 181.285 ;
        RECT 63.045 179.675 64.255 180.195 ;
        RECT 65.845 180.145 66.075 181.285 ;
        RECT 66.245 180.135 66.575 181.115 ;
        RECT 66.745 180.145 66.955 181.285 ;
        RECT 67.190 180.135 67.450 181.285 ;
        RECT 67.625 180.210 67.880 181.115 ;
        RECT 68.050 180.525 68.380 181.285 ;
        RECT 68.595 180.355 68.765 181.115 ;
        RECT 64.425 179.505 65.635 180.025 ;
        RECT 65.825 179.725 66.155 179.975 ;
        RECT 62.130 178.735 62.405 179.215 ;
        RECT 62.575 178.905 62.875 179.235 ;
        RECT 63.045 178.735 65.635 179.505 ;
        RECT 65.845 178.735 66.075 179.555 ;
        RECT 66.325 179.535 66.575 180.135 ;
        RECT 66.245 178.905 66.575 179.535 ;
        RECT 66.745 178.735 66.955 179.555 ;
        RECT 67.190 178.735 67.450 179.575 ;
        RECT 67.625 179.480 67.795 180.210 ;
        RECT 68.050 180.185 68.765 180.355 ;
        RECT 69.025 180.315 69.335 181.115 ;
        RECT 69.505 180.485 69.815 181.285 ;
        RECT 69.985 180.655 70.245 181.115 ;
        RECT 70.415 180.825 70.670 181.285 ;
        RECT 70.845 180.655 71.105 181.115 ;
        RECT 69.985 180.485 71.105 180.655 ;
        RECT 68.050 179.975 68.220 180.185 ;
        RECT 69.025 180.145 70.055 180.315 ;
        RECT 67.965 179.645 68.220 179.975 ;
        RECT 67.625 178.905 67.880 179.480 ;
        RECT 68.050 179.455 68.220 179.645 ;
        RECT 68.500 179.635 68.855 180.005 ;
        RECT 68.050 179.285 68.765 179.455 ;
        RECT 68.050 178.735 68.380 179.115 ;
        RECT 68.595 178.905 68.765 179.285 ;
        RECT 69.025 179.235 69.195 180.145 ;
        RECT 69.365 179.405 69.715 179.975 ;
        RECT 69.885 179.895 70.055 180.145 ;
        RECT 70.845 180.235 71.105 180.485 ;
        RECT 71.275 180.415 71.560 181.285 ;
        RECT 70.845 180.065 71.600 180.235 ;
        RECT 69.885 179.725 71.025 179.895 ;
        RECT 71.195 179.555 71.600 180.065 ;
        RECT 69.950 179.385 71.600 179.555 ;
        RECT 71.785 179.475 72.045 181.100 ;
        RECT 73.795 180.835 74.125 181.285 ;
        RECT 72.225 180.445 74.835 180.655 ;
        RECT 72.225 179.645 72.445 180.445 ;
        RECT 72.685 179.645 72.985 180.265 ;
        RECT 73.155 179.645 73.485 180.265 ;
        RECT 73.655 179.645 73.975 180.265 ;
        RECT 74.145 179.645 74.495 180.265 ;
        RECT 74.665 179.475 74.835 180.445 ;
        RECT 75.925 180.120 76.215 181.285 ;
        RECT 76.500 180.655 76.785 181.115 ;
        RECT 76.955 180.825 77.225 181.285 ;
        RECT 76.500 180.435 77.455 180.655 ;
        RECT 76.385 179.705 77.075 180.265 ;
        RECT 77.245 179.535 77.455 180.435 ;
        RECT 69.025 178.905 69.325 179.235 ;
        RECT 69.495 178.735 69.770 179.215 ;
        RECT 69.950 178.995 70.245 179.385 ;
        RECT 70.415 178.735 70.670 179.215 ;
        RECT 70.845 178.995 71.105 179.385 ;
        RECT 71.785 179.305 73.625 179.475 ;
        RECT 71.275 178.735 71.555 179.215 ;
        RECT 72.055 178.735 72.385 179.130 ;
        RECT 72.555 178.950 72.755 179.305 ;
        RECT 72.925 178.735 73.255 179.135 ;
        RECT 73.425 178.960 73.625 179.305 ;
        RECT 73.795 178.735 74.125 179.475 ;
        RECT 74.360 179.305 74.835 179.475 ;
        RECT 74.360 179.055 74.530 179.305 ;
        RECT 75.925 178.735 76.215 179.460 ;
        RECT 76.500 179.365 77.455 179.535 ;
        RECT 77.625 180.265 78.025 181.115 ;
        RECT 78.215 180.655 78.495 181.115 ;
        RECT 79.015 180.825 79.340 181.285 ;
        RECT 78.215 180.435 79.340 180.655 ;
        RECT 77.625 179.705 78.720 180.265 ;
        RECT 78.890 179.975 79.340 180.435 ;
        RECT 79.510 180.145 79.895 181.115 ;
        RECT 80.270 180.315 80.600 181.115 ;
        RECT 80.770 180.485 81.100 181.285 ;
        RECT 81.400 180.315 81.730 181.115 ;
        RECT 82.375 180.485 82.625 181.285 ;
        RECT 80.270 180.145 82.705 180.315 ;
        RECT 82.895 180.145 83.065 181.285 ;
        RECT 83.235 180.145 83.575 181.115 ;
        RECT 76.500 178.905 76.785 179.365 ;
        RECT 76.955 178.735 77.225 179.195 ;
        RECT 77.625 178.905 78.025 179.705 ;
        RECT 78.890 179.645 79.445 179.975 ;
        RECT 78.890 179.535 79.340 179.645 ;
        RECT 78.215 179.365 79.340 179.535 ;
        RECT 79.615 179.475 79.895 180.145 ;
        RECT 80.065 179.725 80.415 179.975 ;
        RECT 80.600 179.515 80.770 180.145 ;
        RECT 80.940 179.725 81.270 179.925 ;
        RECT 81.440 179.725 81.770 179.925 ;
        RECT 81.940 179.725 82.360 179.925 ;
        RECT 82.535 179.895 82.705 180.145 ;
        RECT 82.535 179.725 83.230 179.895 ;
        RECT 78.215 178.905 78.495 179.365 ;
        RECT 79.015 178.735 79.340 179.195 ;
        RECT 79.510 178.905 79.895 179.475 ;
        RECT 80.270 178.905 80.770 179.515 ;
        RECT 81.400 179.385 82.625 179.555 ;
        RECT 83.400 179.535 83.575 180.145 ;
        RECT 83.745 180.195 85.415 181.285 ;
        RECT 85.585 180.525 86.100 180.935 ;
        RECT 86.335 180.525 86.505 181.285 ;
        RECT 86.675 180.945 88.705 181.115 ;
        RECT 83.745 179.675 84.495 180.195 ;
        RECT 81.400 178.905 81.730 179.385 ;
        RECT 81.900 178.735 82.125 179.195 ;
        RECT 82.295 178.905 82.625 179.385 ;
        RECT 82.815 178.735 83.065 179.535 ;
        RECT 83.235 178.905 83.575 179.535 ;
        RECT 84.665 179.505 85.415 180.025 ;
        RECT 85.585 179.715 85.925 180.525 ;
        RECT 86.675 180.280 86.845 180.945 ;
        RECT 87.240 180.605 88.365 180.775 ;
        RECT 86.095 180.090 86.845 180.280 ;
        RECT 87.015 180.265 88.025 180.435 ;
        RECT 85.585 179.545 86.815 179.715 ;
        RECT 83.745 178.735 85.415 179.505 ;
        RECT 85.860 178.940 86.105 179.545 ;
        RECT 86.325 178.735 86.835 179.270 ;
        RECT 87.015 178.905 87.205 180.265 ;
        RECT 87.375 179.245 87.650 180.065 ;
        RECT 87.855 179.465 88.025 180.265 ;
        RECT 88.195 179.475 88.365 180.605 ;
        RECT 88.535 179.975 88.705 180.945 ;
        RECT 88.875 180.145 89.045 181.285 ;
        RECT 89.215 180.145 89.550 181.115 ;
        RECT 88.535 179.645 88.730 179.975 ;
        RECT 88.955 179.645 89.210 179.975 ;
        RECT 88.955 179.475 89.125 179.645 ;
        RECT 89.380 179.475 89.550 180.145 ;
        RECT 88.195 179.305 89.125 179.475 ;
        RECT 88.195 179.270 88.370 179.305 ;
        RECT 87.375 179.075 87.655 179.245 ;
        RECT 87.375 178.905 87.650 179.075 ;
        RECT 87.840 178.905 88.370 179.270 ;
        RECT 88.795 178.735 89.125 179.135 ;
        RECT 89.295 178.905 89.550 179.475 ;
        RECT 89.725 180.210 89.995 181.115 ;
        RECT 90.165 180.525 90.495 181.285 ;
        RECT 90.675 180.355 90.845 181.115 ;
        RECT 89.725 179.410 89.895 180.210 ;
        RECT 90.180 180.185 90.845 180.355 ;
        RECT 90.180 180.040 90.350 180.185 ;
        RECT 91.145 180.145 91.375 181.285 ;
        RECT 91.545 180.135 91.875 181.115 ;
        RECT 92.045 180.145 92.255 181.285 ;
        RECT 90.065 179.710 90.350 180.040 ;
        RECT 90.180 179.455 90.350 179.710 ;
        RECT 90.585 179.635 90.915 180.005 ;
        RECT 91.125 179.725 91.455 179.975 ;
        RECT 89.725 178.905 89.985 179.410 ;
        RECT 90.180 179.285 90.845 179.455 ;
        RECT 90.165 178.735 90.495 179.115 ;
        RECT 90.675 178.905 90.845 179.285 ;
        RECT 91.145 178.735 91.375 179.555 ;
        RECT 91.625 179.535 91.875 180.135 ;
        RECT 92.490 180.095 92.745 180.975 ;
        RECT 92.915 180.145 93.220 181.285 ;
        RECT 93.560 180.905 93.890 181.285 ;
        RECT 94.070 180.735 94.240 181.025 ;
        RECT 94.410 180.825 94.660 181.285 ;
        RECT 93.440 180.565 94.240 180.735 ;
        RECT 94.830 180.775 95.700 181.115 ;
        RECT 91.545 178.905 91.875 179.535 ;
        RECT 92.045 178.735 92.255 179.555 ;
        RECT 92.490 179.445 92.700 180.095 ;
        RECT 93.440 179.975 93.610 180.565 ;
        RECT 94.830 180.395 95.000 180.775 ;
        RECT 95.935 180.655 96.105 181.115 ;
        RECT 96.275 180.825 96.645 181.285 ;
        RECT 96.940 180.685 97.110 181.025 ;
        RECT 97.280 180.855 97.610 181.285 ;
        RECT 97.845 180.685 98.015 181.025 ;
        RECT 93.780 180.225 95.000 180.395 ;
        RECT 95.170 180.315 95.630 180.605 ;
        RECT 95.935 180.485 96.495 180.655 ;
        RECT 96.940 180.515 98.015 180.685 ;
        RECT 98.185 180.785 98.865 181.115 ;
        RECT 99.080 180.785 99.330 181.115 ;
        RECT 99.500 180.825 99.750 181.285 ;
        RECT 96.325 180.345 96.495 180.485 ;
        RECT 95.170 180.305 96.135 180.315 ;
        RECT 94.830 180.135 95.000 180.225 ;
        RECT 95.460 180.145 96.135 180.305 ;
        RECT 92.870 179.945 93.610 179.975 ;
        RECT 92.870 179.645 93.785 179.945 ;
        RECT 93.460 179.470 93.785 179.645 ;
        RECT 92.490 178.915 92.745 179.445 ;
        RECT 92.915 178.735 93.220 179.195 ;
        RECT 93.465 179.115 93.785 179.470 ;
        RECT 93.955 179.685 94.495 180.055 ;
        RECT 94.830 179.965 95.235 180.135 ;
        RECT 93.955 179.285 94.195 179.685 ;
        RECT 94.675 179.515 94.895 179.795 ;
        RECT 94.365 179.345 94.895 179.515 ;
        RECT 94.365 179.115 94.535 179.345 ;
        RECT 95.065 179.185 95.235 179.965 ;
        RECT 95.405 179.355 95.755 179.975 ;
        RECT 95.925 179.355 96.135 180.145 ;
        RECT 96.325 180.175 97.825 180.345 ;
        RECT 96.325 179.485 96.495 180.175 ;
        RECT 98.185 180.005 98.355 180.785 ;
        RECT 99.160 180.655 99.330 180.785 ;
        RECT 96.665 179.835 98.355 180.005 ;
        RECT 98.525 180.225 98.990 180.615 ;
        RECT 99.160 180.485 99.555 180.655 ;
        RECT 96.665 179.655 96.835 179.835 ;
        RECT 93.465 178.945 94.535 179.115 ;
        RECT 94.705 178.735 94.895 179.175 ;
        RECT 95.065 178.905 96.015 179.185 ;
        RECT 96.325 179.095 96.585 179.485 ;
        RECT 97.005 179.415 97.795 179.665 ;
        RECT 96.235 178.925 96.585 179.095 ;
        RECT 96.795 178.735 97.125 179.195 ;
        RECT 98.000 179.125 98.170 179.835 ;
        RECT 98.525 179.635 98.695 180.225 ;
        RECT 98.340 179.415 98.695 179.635 ;
        RECT 98.865 179.415 99.215 180.035 ;
        RECT 99.385 179.125 99.555 180.485 ;
        RECT 99.920 180.315 100.245 181.100 ;
        RECT 99.725 179.265 100.185 180.315 ;
        RECT 98.000 178.955 98.855 179.125 ;
        RECT 99.060 178.955 99.555 179.125 ;
        RECT 99.725 178.735 100.055 179.095 ;
        RECT 100.415 178.995 100.585 181.115 ;
        RECT 100.755 180.785 101.085 181.285 ;
        RECT 101.255 180.615 101.510 181.115 ;
        RECT 100.760 180.445 101.510 180.615 ;
        RECT 100.760 179.455 100.990 180.445 ;
        RECT 101.160 179.625 101.510 180.275 ;
        RECT 101.685 180.120 101.975 181.285 ;
        RECT 102.145 180.145 102.530 181.115 ;
        RECT 102.700 180.825 103.025 181.285 ;
        RECT 103.545 180.655 103.825 181.115 ;
        RECT 102.700 180.435 103.825 180.655 ;
        RECT 102.145 179.475 102.425 180.145 ;
        RECT 102.700 179.975 103.150 180.435 ;
        RECT 104.015 180.265 104.415 181.115 ;
        RECT 104.815 180.825 105.085 181.285 ;
        RECT 105.255 180.655 105.540 181.115 ;
        RECT 102.595 179.645 103.150 179.975 ;
        RECT 103.320 179.705 104.415 180.265 ;
        RECT 102.700 179.535 103.150 179.645 ;
        RECT 100.760 179.285 101.510 179.455 ;
        RECT 100.755 178.735 101.085 179.115 ;
        RECT 101.255 178.995 101.510 179.285 ;
        RECT 101.685 178.735 101.975 179.460 ;
        RECT 102.145 178.905 102.530 179.475 ;
        RECT 102.700 179.365 103.825 179.535 ;
        RECT 102.700 178.735 103.025 179.195 ;
        RECT 103.545 178.905 103.825 179.365 ;
        RECT 104.015 178.905 104.415 179.705 ;
        RECT 104.585 180.435 105.540 180.655 ;
        RECT 104.585 179.535 104.795 180.435 ;
        RECT 104.965 179.705 105.655 180.265 ;
        RECT 105.825 180.145 106.210 181.115 ;
        RECT 106.380 180.825 106.705 181.285 ;
        RECT 107.225 180.655 107.505 181.115 ;
        RECT 106.380 180.435 107.505 180.655 ;
        RECT 104.585 179.365 105.540 179.535 ;
        RECT 104.815 178.735 105.085 179.195 ;
        RECT 105.255 178.905 105.540 179.365 ;
        RECT 105.825 179.475 106.105 180.145 ;
        RECT 106.380 179.975 106.830 180.435 ;
        RECT 107.695 180.265 108.095 181.115 ;
        RECT 108.495 180.825 108.765 181.285 ;
        RECT 108.935 180.655 109.220 181.115 ;
        RECT 106.275 179.645 106.830 179.975 ;
        RECT 107.000 179.705 108.095 180.265 ;
        RECT 106.380 179.535 106.830 179.645 ;
        RECT 105.825 178.905 106.210 179.475 ;
        RECT 106.380 179.365 107.505 179.535 ;
        RECT 106.380 178.735 106.705 179.195 ;
        RECT 107.225 178.905 107.505 179.365 ;
        RECT 107.695 178.905 108.095 179.705 ;
        RECT 108.265 180.435 109.220 180.655 ;
        RECT 108.265 179.535 108.475 180.435 ;
        RECT 108.645 179.705 109.335 180.265 ;
        RECT 110.005 180.145 110.235 181.285 ;
        RECT 110.405 180.135 110.735 181.115 ;
        RECT 110.905 180.145 111.115 181.285 ;
        RECT 109.985 179.725 110.315 179.975 ;
        RECT 108.265 179.365 109.220 179.535 ;
        RECT 108.495 178.735 108.765 179.195 ;
        RECT 108.935 178.905 109.220 179.365 ;
        RECT 110.005 178.735 110.235 179.555 ;
        RECT 110.485 179.535 110.735 180.135 ;
        RECT 111.350 180.095 111.605 180.975 ;
        RECT 111.775 180.145 112.080 181.285 ;
        RECT 112.420 180.905 112.750 181.285 ;
        RECT 112.930 180.735 113.100 181.025 ;
        RECT 113.270 180.825 113.520 181.285 ;
        RECT 112.300 180.565 113.100 180.735 ;
        RECT 113.690 180.775 114.560 181.115 ;
        RECT 110.405 178.905 110.735 179.535 ;
        RECT 110.905 178.735 111.115 179.555 ;
        RECT 111.350 179.445 111.560 180.095 ;
        RECT 112.300 179.975 112.470 180.565 ;
        RECT 113.690 180.395 113.860 180.775 ;
        RECT 114.795 180.655 114.965 181.115 ;
        RECT 115.135 180.825 115.505 181.285 ;
        RECT 115.800 180.685 115.970 181.025 ;
        RECT 116.140 180.855 116.470 181.285 ;
        RECT 116.705 180.685 116.875 181.025 ;
        RECT 112.640 180.225 113.860 180.395 ;
        RECT 114.030 180.315 114.490 180.605 ;
        RECT 114.795 180.485 115.355 180.655 ;
        RECT 115.800 180.515 116.875 180.685 ;
        RECT 117.045 180.785 117.725 181.115 ;
        RECT 117.940 180.785 118.190 181.115 ;
        RECT 118.360 180.825 118.610 181.285 ;
        RECT 115.185 180.345 115.355 180.485 ;
        RECT 114.030 180.305 114.995 180.315 ;
        RECT 113.690 180.135 113.860 180.225 ;
        RECT 114.320 180.145 114.995 180.305 ;
        RECT 111.730 179.945 112.470 179.975 ;
        RECT 111.730 179.645 112.645 179.945 ;
        RECT 112.320 179.470 112.645 179.645 ;
        RECT 111.350 178.915 111.605 179.445 ;
        RECT 111.775 178.735 112.080 179.195 ;
        RECT 112.325 179.115 112.645 179.470 ;
        RECT 112.815 179.685 113.355 180.055 ;
        RECT 113.690 179.965 114.095 180.135 ;
        RECT 112.815 179.285 113.055 179.685 ;
        RECT 113.535 179.515 113.755 179.795 ;
        RECT 113.225 179.345 113.755 179.515 ;
        RECT 113.225 179.115 113.395 179.345 ;
        RECT 113.925 179.185 114.095 179.965 ;
        RECT 114.265 179.355 114.615 179.975 ;
        RECT 114.785 179.355 114.995 180.145 ;
        RECT 115.185 180.175 116.685 180.345 ;
        RECT 115.185 179.485 115.355 180.175 ;
        RECT 117.045 180.005 117.215 180.785 ;
        RECT 118.020 180.655 118.190 180.785 ;
        RECT 115.525 179.835 117.215 180.005 ;
        RECT 117.385 180.225 117.850 180.615 ;
        RECT 118.020 180.485 118.415 180.655 ;
        RECT 115.525 179.655 115.695 179.835 ;
        RECT 112.325 178.945 113.395 179.115 ;
        RECT 113.565 178.735 113.755 179.175 ;
        RECT 113.925 178.905 114.875 179.185 ;
        RECT 115.185 179.095 115.445 179.485 ;
        RECT 115.865 179.415 116.655 179.665 ;
        RECT 115.095 178.925 115.445 179.095 ;
        RECT 115.655 178.735 115.985 179.195 ;
        RECT 116.860 179.125 117.030 179.835 ;
        RECT 117.385 179.635 117.555 180.225 ;
        RECT 117.200 179.415 117.555 179.635 ;
        RECT 117.725 179.415 118.075 180.035 ;
        RECT 118.245 179.125 118.415 180.485 ;
        RECT 118.780 180.315 119.105 181.100 ;
        RECT 118.585 179.265 119.045 180.315 ;
        RECT 116.860 178.955 117.715 179.125 ;
        RECT 117.920 178.955 118.415 179.125 ;
        RECT 118.585 178.735 118.915 179.095 ;
        RECT 119.275 178.995 119.445 181.115 ;
        RECT 119.615 180.785 119.945 181.285 ;
        RECT 120.115 180.615 120.370 181.115 ;
        RECT 119.620 180.445 120.370 180.615 ;
        RECT 119.620 179.455 119.850 180.445 ;
        RECT 120.020 179.625 120.370 180.275 ;
        RECT 120.585 180.145 120.815 181.285 ;
        RECT 120.985 180.135 121.315 181.115 ;
        RECT 121.485 180.145 121.695 181.285 ;
        RECT 122.015 180.355 122.185 181.115 ;
        RECT 122.365 180.525 122.695 181.285 ;
        RECT 122.015 180.185 122.680 180.355 ;
        RECT 122.865 180.210 123.135 181.115 ;
        RECT 120.565 179.725 120.895 179.975 ;
        RECT 119.620 179.285 120.370 179.455 ;
        RECT 119.615 178.735 119.945 179.115 ;
        RECT 120.115 178.995 120.370 179.285 ;
        RECT 120.585 178.735 120.815 179.555 ;
        RECT 121.065 179.535 121.315 180.135 ;
        RECT 122.510 180.040 122.680 180.185 ;
        RECT 121.945 179.635 122.275 180.005 ;
        RECT 122.510 179.710 122.795 180.040 ;
        RECT 120.985 178.905 121.315 179.535 ;
        RECT 121.485 178.735 121.695 179.555 ;
        RECT 122.510 179.455 122.680 179.710 ;
        RECT 122.015 179.285 122.680 179.455 ;
        RECT 122.965 179.410 123.135 180.210 ;
        RECT 123.765 180.195 126.355 181.285 ;
        RECT 126.525 180.195 127.735 181.285 ;
        RECT 123.765 179.675 124.975 180.195 ;
        RECT 125.145 179.505 126.355 180.025 ;
        RECT 126.525 179.655 127.045 180.195 ;
        RECT 122.015 178.905 122.185 179.285 ;
        RECT 122.365 178.735 122.695 179.115 ;
        RECT 122.875 178.905 123.135 179.410 ;
        RECT 123.765 178.735 126.355 179.505 ;
        RECT 127.215 179.485 127.735 180.025 ;
        RECT 126.525 178.735 127.735 179.485 ;
        RECT 14.660 178.565 127.820 178.735 ;
        RECT 14.745 177.815 15.955 178.565 ;
        RECT 14.745 177.275 15.265 177.815 ;
        RECT 16.125 177.795 19.635 178.565 ;
        RECT 19.810 178.020 25.155 178.565 ;
        RECT 15.435 177.105 15.955 177.645 ;
        RECT 14.745 176.015 15.955 177.105 ;
        RECT 16.125 177.105 17.815 177.625 ;
        RECT 17.985 177.275 19.635 177.795 ;
        RECT 16.125 176.015 19.635 177.105 ;
        RECT 21.400 176.450 21.750 177.700 ;
        RECT 23.230 177.190 23.570 178.020 ;
        RECT 25.385 177.745 25.595 178.565 ;
        RECT 25.765 177.765 26.095 178.395 ;
        RECT 25.765 177.165 26.015 177.765 ;
        RECT 26.265 177.745 26.495 178.565 ;
        RECT 26.745 177.745 26.975 178.565 ;
        RECT 27.145 177.765 27.475 178.395 ;
        RECT 26.185 177.325 26.515 177.575 ;
        RECT 26.725 177.325 27.055 177.575 ;
        RECT 27.225 177.165 27.475 177.765 ;
        RECT 27.645 177.745 27.855 178.565 ;
        RECT 28.090 177.855 28.345 178.385 ;
        RECT 28.515 178.105 28.820 178.565 ;
        RECT 29.065 178.185 30.135 178.355 ;
        RECT 19.810 176.015 25.155 176.450 ;
        RECT 25.385 176.015 25.595 177.155 ;
        RECT 25.765 176.185 26.095 177.165 ;
        RECT 26.265 176.015 26.495 177.155 ;
        RECT 26.745 176.015 26.975 177.155 ;
        RECT 27.145 176.185 27.475 177.165 ;
        RECT 28.090 177.205 28.300 177.855 ;
        RECT 29.065 177.830 29.385 178.185 ;
        RECT 29.060 177.655 29.385 177.830 ;
        RECT 28.470 177.355 29.385 177.655 ;
        RECT 29.555 177.615 29.795 178.015 ;
        RECT 29.965 177.955 30.135 178.185 ;
        RECT 30.305 178.125 30.495 178.565 ;
        RECT 30.665 178.115 31.615 178.395 ;
        RECT 31.835 178.205 32.185 178.375 ;
        RECT 29.965 177.785 30.495 177.955 ;
        RECT 28.470 177.325 29.210 177.355 ;
        RECT 27.645 176.015 27.855 177.155 ;
        RECT 28.090 176.325 28.345 177.205 ;
        RECT 28.515 176.015 28.820 177.155 ;
        RECT 29.040 176.735 29.210 177.325 ;
        RECT 29.555 177.245 30.095 177.615 ;
        RECT 30.275 177.505 30.495 177.785 ;
        RECT 30.665 177.335 30.835 178.115 ;
        RECT 30.430 177.165 30.835 177.335 ;
        RECT 31.005 177.325 31.355 177.945 ;
        RECT 30.430 177.075 30.600 177.165 ;
        RECT 31.525 177.155 31.735 177.945 ;
        RECT 29.380 176.905 30.600 177.075 ;
        RECT 31.060 176.995 31.735 177.155 ;
        RECT 29.040 176.565 29.840 176.735 ;
        RECT 29.160 176.015 29.490 176.395 ;
        RECT 29.670 176.275 29.840 176.565 ;
        RECT 30.430 176.525 30.600 176.905 ;
        RECT 30.770 176.985 31.735 176.995 ;
        RECT 31.925 177.815 32.185 178.205 ;
        RECT 32.395 178.105 32.725 178.565 ;
        RECT 33.600 178.175 34.455 178.345 ;
        RECT 34.660 178.175 35.155 178.345 ;
        RECT 35.325 178.205 35.655 178.565 ;
        RECT 31.925 177.125 32.095 177.815 ;
        RECT 32.265 177.465 32.435 177.645 ;
        RECT 32.605 177.635 33.395 177.885 ;
        RECT 33.600 177.465 33.770 178.175 ;
        RECT 33.940 177.665 34.295 177.885 ;
        RECT 32.265 177.295 33.955 177.465 ;
        RECT 30.770 176.695 31.230 176.985 ;
        RECT 31.925 176.955 33.425 177.125 ;
        RECT 31.925 176.815 32.095 176.955 ;
        RECT 31.535 176.645 32.095 176.815 ;
        RECT 30.010 176.015 30.260 176.475 ;
        RECT 30.430 176.185 31.300 176.525 ;
        RECT 31.535 176.185 31.705 176.645 ;
        RECT 32.540 176.615 33.615 176.785 ;
        RECT 31.875 176.015 32.245 176.475 ;
        RECT 32.540 176.275 32.710 176.615 ;
        RECT 32.880 176.015 33.210 176.445 ;
        RECT 33.445 176.275 33.615 176.615 ;
        RECT 33.785 176.515 33.955 177.295 ;
        RECT 34.125 177.075 34.295 177.665 ;
        RECT 34.465 177.265 34.815 177.885 ;
        RECT 34.125 176.685 34.590 177.075 ;
        RECT 34.985 176.815 35.155 178.175 ;
        RECT 35.325 176.985 35.785 178.035 ;
        RECT 34.760 176.645 35.155 176.815 ;
        RECT 34.760 176.515 34.930 176.645 ;
        RECT 33.785 176.185 34.465 176.515 ;
        RECT 34.680 176.185 34.930 176.515 ;
        RECT 35.100 176.015 35.350 176.475 ;
        RECT 35.520 176.200 35.845 176.985 ;
        RECT 36.015 176.185 36.185 178.305 ;
        RECT 36.355 178.185 36.685 178.565 ;
        RECT 36.855 178.015 37.110 178.305 ;
        RECT 36.360 177.845 37.110 178.015 ;
        RECT 36.360 176.855 36.590 177.845 ;
        RECT 37.285 177.840 37.575 178.565 ;
        RECT 38.020 177.755 38.265 178.360 ;
        RECT 38.485 178.030 38.995 178.565 ;
        RECT 36.760 177.025 37.110 177.675 ;
        RECT 37.745 177.585 38.975 177.755 ;
        RECT 36.360 176.685 37.110 176.855 ;
        RECT 36.355 176.015 36.685 176.515 ;
        RECT 36.855 176.185 37.110 176.685 ;
        RECT 37.285 176.015 37.575 177.180 ;
        RECT 37.745 176.775 38.085 177.585 ;
        RECT 38.255 177.020 39.005 177.210 ;
        RECT 37.745 176.365 38.260 176.775 ;
        RECT 38.495 176.015 38.665 176.775 ;
        RECT 38.835 176.355 39.005 177.020 ;
        RECT 39.175 177.035 39.365 178.395 ;
        RECT 39.535 178.225 39.810 178.395 ;
        RECT 39.535 178.055 39.815 178.225 ;
        RECT 39.535 177.235 39.810 178.055 ;
        RECT 40.000 178.030 40.530 178.395 ;
        RECT 40.955 178.165 41.285 178.565 ;
        RECT 40.355 177.995 40.530 178.030 ;
        RECT 40.015 177.035 40.185 177.835 ;
        RECT 39.175 176.865 40.185 177.035 ;
        RECT 40.355 177.825 41.285 177.995 ;
        RECT 41.455 177.825 41.710 178.395 ;
        RECT 40.355 176.695 40.525 177.825 ;
        RECT 41.115 177.655 41.285 177.825 ;
        RECT 39.400 176.525 40.525 176.695 ;
        RECT 40.695 177.325 40.890 177.655 ;
        RECT 41.115 177.325 41.370 177.655 ;
        RECT 40.695 176.355 40.865 177.325 ;
        RECT 41.540 177.155 41.710 177.825 ;
        RECT 42.920 177.935 43.205 178.395 ;
        RECT 43.375 178.105 43.645 178.565 ;
        RECT 42.920 177.765 43.875 177.935 ;
        RECT 38.835 176.185 40.865 176.355 ;
        RECT 41.035 176.015 41.205 177.155 ;
        RECT 41.375 176.185 41.710 177.155 ;
        RECT 42.805 177.035 43.495 177.595 ;
        RECT 43.665 176.865 43.875 177.765 ;
        RECT 42.920 176.645 43.875 176.865 ;
        RECT 44.045 177.595 44.445 178.395 ;
        RECT 44.635 177.935 44.915 178.395 ;
        RECT 45.435 178.105 45.760 178.565 ;
        RECT 44.635 177.765 45.760 177.935 ;
        RECT 45.930 177.825 46.315 178.395 ;
        RECT 45.310 177.655 45.760 177.765 ;
        RECT 44.045 177.035 45.140 177.595 ;
        RECT 45.310 177.325 45.865 177.655 ;
        RECT 42.920 176.185 43.205 176.645 ;
        RECT 43.375 176.015 43.645 176.475 ;
        RECT 44.045 176.185 44.445 177.035 ;
        RECT 45.310 176.865 45.760 177.325 ;
        RECT 46.035 177.155 46.315 177.825 ;
        RECT 46.690 177.785 47.190 178.395 ;
        RECT 46.485 177.325 46.835 177.575 ;
        RECT 47.020 177.155 47.190 177.785 ;
        RECT 47.820 177.915 48.150 178.395 ;
        RECT 48.320 178.105 48.545 178.565 ;
        RECT 48.715 177.915 49.045 178.395 ;
        RECT 47.820 177.745 49.045 177.915 ;
        RECT 49.235 177.765 49.485 178.565 ;
        RECT 49.655 177.765 49.995 178.395 ;
        RECT 50.280 177.935 50.565 178.395 ;
        RECT 50.735 178.105 51.005 178.565 ;
        RECT 50.280 177.765 51.235 177.935 ;
        RECT 47.360 177.375 47.690 177.575 ;
        RECT 47.860 177.375 48.190 177.575 ;
        RECT 48.360 177.375 48.780 177.575 ;
        RECT 48.955 177.405 49.650 177.575 ;
        RECT 48.955 177.155 49.125 177.405 ;
        RECT 49.820 177.155 49.995 177.765 ;
        RECT 44.635 176.645 45.760 176.865 ;
        RECT 44.635 176.185 44.915 176.645 ;
        RECT 45.435 176.015 45.760 176.475 ;
        RECT 45.930 176.185 46.315 177.155 ;
        RECT 46.690 176.985 49.125 177.155 ;
        RECT 46.690 176.185 47.020 176.985 ;
        RECT 47.190 176.015 47.520 176.815 ;
        RECT 47.820 176.185 48.150 176.985 ;
        RECT 48.795 176.015 49.045 176.815 ;
        RECT 49.315 176.015 49.485 177.155 ;
        RECT 49.655 176.185 49.995 177.155 ;
        RECT 50.165 177.035 50.855 177.595 ;
        RECT 51.025 176.865 51.235 177.765 ;
        RECT 50.280 176.645 51.235 176.865 ;
        RECT 51.405 177.595 51.805 178.395 ;
        RECT 51.995 177.935 52.275 178.395 ;
        RECT 52.795 178.105 53.120 178.565 ;
        RECT 51.995 177.765 53.120 177.935 ;
        RECT 53.290 177.825 53.675 178.395 ;
        RECT 52.670 177.655 53.120 177.765 ;
        RECT 51.405 177.035 52.500 177.595 ;
        RECT 52.670 177.325 53.225 177.655 ;
        RECT 50.280 176.185 50.565 176.645 ;
        RECT 50.735 176.015 51.005 176.475 ;
        RECT 51.405 176.185 51.805 177.035 ;
        RECT 52.670 176.865 53.120 177.325 ;
        RECT 53.395 177.155 53.675 177.825 ;
        RECT 51.995 176.645 53.120 176.865 ;
        RECT 51.995 176.185 52.275 176.645 ;
        RECT 52.795 176.015 53.120 176.475 ;
        RECT 53.290 176.185 53.675 177.155 ;
        RECT 53.850 177.855 54.105 178.385 ;
        RECT 54.275 178.105 54.580 178.565 ;
        RECT 54.825 178.185 55.895 178.355 ;
        RECT 53.850 177.205 54.060 177.855 ;
        RECT 54.825 177.830 55.145 178.185 ;
        RECT 54.820 177.655 55.145 177.830 ;
        RECT 54.230 177.355 55.145 177.655 ;
        RECT 55.315 177.615 55.555 178.015 ;
        RECT 55.725 177.955 55.895 178.185 ;
        RECT 56.065 178.125 56.255 178.565 ;
        RECT 56.425 178.115 57.375 178.395 ;
        RECT 57.595 178.205 57.945 178.375 ;
        RECT 55.725 177.785 56.255 177.955 ;
        RECT 54.230 177.325 54.970 177.355 ;
        RECT 53.850 176.325 54.105 177.205 ;
        RECT 54.275 176.015 54.580 177.155 ;
        RECT 54.800 176.735 54.970 177.325 ;
        RECT 55.315 177.245 55.855 177.615 ;
        RECT 56.035 177.505 56.255 177.785 ;
        RECT 56.425 177.335 56.595 178.115 ;
        RECT 56.190 177.165 56.595 177.335 ;
        RECT 56.765 177.325 57.115 177.945 ;
        RECT 56.190 177.075 56.360 177.165 ;
        RECT 57.285 177.155 57.495 177.945 ;
        RECT 55.140 176.905 56.360 177.075 ;
        RECT 56.820 176.995 57.495 177.155 ;
        RECT 54.800 176.565 55.600 176.735 ;
        RECT 54.920 176.015 55.250 176.395 ;
        RECT 55.430 176.275 55.600 176.565 ;
        RECT 56.190 176.525 56.360 176.905 ;
        RECT 56.530 176.985 57.495 176.995 ;
        RECT 57.685 177.815 57.945 178.205 ;
        RECT 58.155 178.105 58.485 178.565 ;
        RECT 59.360 178.175 60.215 178.345 ;
        RECT 60.420 178.175 60.915 178.345 ;
        RECT 61.085 178.205 61.415 178.565 ;
        RECT 57.685 177.125 57.855 177.815 ;
        RECT 58.025 177.465 58.195 177.645 ;
        RECT 58.365 177.635 59.155 177.885 ;
        RECT 59.360 177.465 59.530 178.175 ;
        RECT 59.700 177.665 60.055 177.885 ;
        RECT 58.025 177.295 59.715 177.465 ;
        RECT 56.530 176.695 56.990 176.985 ;
        RECT 57.685 176.955 59.185 177.125 ;
        RECT 57.685 176.815 57.855 176.955 ;
        RECT 57.295 176.645 57.855 176.815 ;
        RECT 55.770 176.015 56.020 176.475 ;
        RECT 56.190 176.185 57.060 176.525 ;
        RECT 57.295 176.185 57.465 176.645 ;
        RECT 58.300 176.615 59.375 176.785 ;
        RECT 57.635 176.015 58.005 176.475 ;
        RECT 58.300 176.275 58.470 176.615 ;
        RECT 58.640 176.015 58.970 176.445 ;
        RECT 59.205 176.275 59.375 176.615 ;
        RECT 59.545 176.515 59.715 177.295 ;
        RECT 59.885 177.075 60.055 177.665 ;
        RECT 60.225 177.265 60.575 177.885 ;
        RECT 59.885 176.685 60.350 177.075 ;
        RECT 60.745 176.815 60.915 178.175 ;
        RECT 61.085 176.985 61.545 178.035 ;
        RECT 60.520 176.645 60.915 176.815 ;
        RECT 60.520 176.515 60.690 176.645 ;
        RECT 59.545 176.185 60.225 176.515 ;
        RECT 60.440 176.185 60.690 176.515 ;
        RECT 60.860 176.015 61.110 176.475 ;
        RECT 61.280 176.200 61.605 176.985 ;
        RECT 61.775 176.185 61.945 178.305 ;
        RECT 62.115 178.185 62.445 178.565 ;
        RECT 62.615 178.015 62.870 178.305 ;
        RECT 62.120 177.845 62.870 178.015 ;
        RECT 62.120 176.855 62.350 177.845 ;
        RECT 63.045 177.840 63.335 178.565 ;
        RECT 63.505 177.890 63.765 178.395 ;
        RECT 63.945 178.185 64.275 178.565 ;
        RECT 64.455 178.015 64.625 178.395 ;
        RECT 62.520 177.025 62.870 177.675 ;
        RECT 62.120 176.685 62.870 176.855 ;
        RECT 62.115 176.015 62.445 176.515 ;
        RECT 62.615 176.185 62.870 176.685 ;
        RECT 63.045 176.015 63.335 177.180 ;
        RECT 63.505 177.090 63.675 177.890 ;
        RECT 63.960 177.845 64.625 178.015 ;
        RECT 63.960 177.590 64.130 177.845 ;
        RECT 64.885 177.795 67.475 178.565 ;
        RECT 63.845 177.260 64.130 177.590 ;
        RECT 64.365 177.295 64.695 177.665 ;
        RECT 63.960 177.115 64.130 177.260 ;
        RECT 63.505 176.185 63.775 177.090 ;
        RECT 63.960 176.945 64.625 177.115 ;
        RECT 63.945 176.015 64.275 176.775 ;
        RECT 64.455 176.185 64.625 176.945 ;
        RECT 64.885 177.105 66.095 177.625 ;
        RECT 66.265 177.275 67.475 177.795 ;
        RECT 67.650 177.725 67.910 178.565 ;
        RECT 68.085 177.820 68.340 178.395 ;
        RECT 68.510 178.185 68.840 178.565 ;
        RECT 69.055 178.015 69.225 178.395 ;
        RECT 68.510 177.845 69.225 178.015 ;
        RECT 69.575 178.015 69.745 178.395 ;
        RECT 69.960 178.185 70.290 178.565 ;
        RECT 69.575 177.845 70.290 178.015 ;
        RECT 64.885 176.015 67.475 177.105 ;
        RECT 67.650 176.015 67.910 177.165 ;
        RECT 68.085 177.090 68.255 177.820 ;
        RECT 68.510 177.655 68.680 177.845 ;
        RECT 68.425 177.325 68.680 177.655 ;
        RECT 68.510 177.115 68.680 177.325 ;
        RECT 68.960 177.295 69.315 177.665 ;
        RECT 69.485 177.295 69.840 177.665 ;
        RECT 70.120 177.655 70.290 177.845 ;
        RECT 70.460 177.820 70.715 178.395 ;
        RECT 70.120 177.325 70.375 177.655 ;
        RECT 70.120 177.115 70.290 177.325 ;
        RECT 68.085 176.185 68.340 177.090 ;
        RECT 68.510 176.945 69.225 177.115 ;
        RECT 68.510 176.015 68.840 176.775 ;
        RECT 69.055 176.185 69.225 176.945 ;
        RECT 69.575 176.945 70.290 177.115 ;
        RECT 70.545 177.090 70.715 177.820 ;
        RECT 70.890 177.725 71.150 178.565 ;
        RECT 71.415 178.015 71.585 178.395 ;
        RECT 71.800 178.185 72.130 178.565 ;
        RECT 71.415 177.845 72.130 178.015 ;
        RECT 71.325 177.295 71.680 177.665 ;
        RECT 71.960 177.655 72.130 177.845 ;
        RECT 72.300 177.820 72.555 178.395 ;
        RECT 71.960 177.325 72.215 177.655 ;
        RECT 69.575 176.185 69.745 176.945 ;
        RECT 69.960 176.015 70.290 176.775 ;
        RECT 70.460 176.185 70.715 177.090 ;
        RECT 70.890 176.015 71.150 177.165 ;
        RECT 71.960 177.115 72.130 177.325 ;
        RECT 71.415 176.945 72.130 177.115 ;
        RECT 72.385 177.090 72.555 177.820 ;
        RECT 72.730 177.725 72.990 178.565 ;
        RECT 73.165 177.805 73.875 178.395 ;
        RECT 74.385 178.035 74.715 178.395 ;
        RECT 74.915 178.205 75.245 178.565 ;
        RECT 75.415 178.035 75.745 178.395 ;
        RECT 74.385 177.825 75.745 178.035 ;
        RECT 71.415 176.185 71.585 176.945 ;
        RECT 71.800 176.015 72.130 176.775 ;
        RECT 72.300 176.185 72.555 177.090 ;
        RECT 72.730 176.015 72.990 177.165 ;
        RECT 73.165 176.835 73.370 177.805 ;
        RECT 76.590 177.785 77.090 178.395 ;
        RECT 73.540 177.035 73.870 177.575 ;
        RECT 74.045 177.325 74.540 177.655 ;
        RECT 74.860 177.325 75.235 177.655 ;
        RECT 75.445 177.325 75.755 177.655 ;
        RECT 76.385 177.325 76.735 177.575 ;
        RECT 74.045 177.035 74.370 177.325 ;
        RECT 74.565 176.835 74.895 177.055 ;
        RECT 73.165 176.605 74.895 176.835 ;
        RECT 73.165 176.185 73.865 176.605 ;
        RECT 74.065 176.015 74.395 176.375 ;
        RECT 74.565 176.205 74.895 176.605 ;
        RECT 75.065 176.400 75.235 177.325 ;
        RECT 76.920 177.155 77.090 177.785 ;
        RECT 77.720 177.915 78.050 178.395 ;
        RECT 78.220 178.105 78.445 178.565 ;
        RECT 78.615 177.915 78.945 178.395 ;
        RECT 77.720 177.745 78.945 177.915 ;
        RECT 79.135 177.765 79.385 178.565 ;
        RECT 79.555 177.765 79.895 178.395 ;
        RECT 77.260 177.375 77.590 177.575 ;
        RECT 77.760 177.375 78.090 177.575 ;
        RECT 78.260 177.375 78.680 177.575 ;
        RECT 78.855 177.405 79.550 177.575 ;
        RECT 78.855 177.155 79.025 177.405 ;
        RECT 79.720 177.205 79.895 177.765 ;
        RECT 79.665 177.155 79.895 177.205 ;
        RECT 75.415 176.015 75.745 177.075 ;
        RECT 76.590 176.985 79.025 177.155 ;
        RECT 76.590 176.185 76.920 176.985 ;
        RECT 77.090 176.015 77.420 176.815 ;
        RECT 77.720 176.185 78.050 176.985 ;
        RECT 78.695 176.015 78.945 176.815 ;
        RECT 79.215 176.015 79.385 177.155 ;
        RECT 79.555 176.185 79.895 177.155 ;
        RECT 80.065 177.765 80.405 178.395 ;
        RECT 80.575 177.765 80.825 178.565 ;
        RECT 81.015 177.915 81.345 178.395 ;
        RECT 81.515 178.105 81.740 178.565 ;
        RECT 81.910 177.915 82.240 178.395 ;
        RECT 80.065 177.715 80.295 177.765 ;
        RECT 81.015 177.745 82.240 177.915 ;
        RECT 82.870 177.785 83.370 178.395 ;
        RECT 83.745 177.815 84.955 178.565 ;
        RECT 80.065 177.155 80.240 177.715 ;
        RECT 80.410 177.405 81.105 177.575 ;
        RECT 80.935 177.155 81.105 177.405 ;
        RECT 81.280 177.375 81.700 177.575 ;
        RECT 81.870 177.375 82.200 177.575 ;
        RECT 82.370 177.375 82.700 177.575 ;
        RECT 82.870 177.155 83.040 177.785 ;
        RECT 83.225 177.325 83.575 177.575 ;
        RECT 80.065 176.185 80.405 177.155 ;
        RECT 80.575 176.015 80.745 177.155 ;
        RECT 80.935 176.985 83.370 177.155 ;
        RECT 81.015 176.015 81.265 176.815 ;
        RECT 81.910 176.185 82.240 176.985 ;
        RECT 82.540 176.015 82.870 176.815 ;
        RECT 83.040 176.185 83.370 176.985 ;
        RECT 83.745 177.105 84.265 177.645 ;
        RECT 84.435 177.275 84.955 177.815 ;
        RECT 85.240 177.935 85.525 178.395 ;
        RECT 85.695 178.105 85.965 178.565 ;
        RECT 85.240 177.765 86.195 177.935 ;
        RECT 83.745 176.015 84.955 177.105 ;
        RECT 85.125 177.035 85.815 177.595 ;
        RECT 85.985 176.865 86.195 177.765 ;
        RECT 85.240 176.645 86.195 176.865 ;
        RECT 86.365 177.595 86.765 178.395 ;
        RECT 86.955 177.935 87.235 178.395 ;
        RECT 87.755 178.105 88.080 178.565 ;
        RECT 86.955 177.765 88.080 177.935 ;
        RECT 88.250 177.825 88.635 178.395 ;
        RECT 88.805 177.840 89.095 178.565 ;
        RECT 87.630 177.655 88.080 177.765 ;
        RECT 86.365 177.035 87.460 177.595 ;
        RECT 87.630 177.325 88.185 177.655 ;
        RECT 85.240 176.185 85.525 176.645 ;
        RECT 85.695 176.015 85.965 176.475 ;
        RECT 86.365 176.185 86.765 177.035 ;
        RECT 87.630 176.865 88.080 177.325 ;
        RECT 88.355 177.155 88.635 177.825 ;
        RECT 89.265 177.795 92.775 178.565 ;
        RECT 92.950 178.020 98.295 178.565 ;
        RECT 86.955 176.645 88.080 176.865 ;
        RECT 86.955 176.185 87.235 176.645 ;
        RECT 87.755 176.015 88.080 176.475 ;
        RECT 88.250 176.185 88.635 177.155 ;
        RECT 88.805 176.015 89.095 177.180 ;
        RECT 89.265 177.105 90.955 177.625 ;
        RECT 91.125 177.275 92.775 177.795 ;
        RECT 89.265 176.015 92.775 177.105 ;
        RECT 94.540 176.450 94.890 177.700 ;
        RECT 96.370 177.190 96.710 178.020 ;
        RECT 98.670 177.785 99.170 178.395 ;
        RECT 98.465 177.325 98.815 177.575 ;
        RECT 99.000 177.155 99.170 177.785 ;
        RECT 99.800 177.915 100.130 178.395 ;
        RECT 100.300 178.105 100.525 178.565 ;
        RECT 100.695 177.915 101.025 178.395 ;
        RECT 99.800 177.745 101.025 177.915 ;
        RECT 101.215 177.765 101.465 178.565 ;
        RECT 101.635 177.765 101.975 178.395 ;
        RECT 99.340 177.375 99.670 177.575 ;
        RECT 99.840 177.375 100.170 177.575 ;
        RECT 100.340 177.375 100.760 177.575 ;
        RECT 100.935 177.405 101.630 177.575 ;
        RECT 100.935 177.155 101.105 177.405 ;
        RECT 101.800 177.155 101.975 177.765 ;
        RECT 98.670 176.985 101.105 177.155 ;
        RECT 92.950 176.015 98.295 176.450 ;
        RECT 98.670 176.185 99.000 176.985 ;
        RECT 99.170 176.015 99.500 176.815 ;
        RECT 99.800 176.185 100.130 176.985 ;
        RECT 100.775 176.015 101.025 176.815 ;
        RECT 101.295 176.015 101.465 177.155 ;
        RECT 101.635 176.185 101.975 177.155 ;
        RECT 102.145 177.890 102.405 178.395 ;
        RECT 102.585 178.185 102.915 178.565 ;
        RECT 103.095 178.015 103.265 178.395 ;
        RECT 102.145 177.090 102.315 177.890 ;
        RECT 102.600 177.845 103.265 178.015 ;
        RECT 102.600 177.590 102.770 177.845 ;
        RECT 103.525 177.815 104.735 178.565 ;
        RECT 102.485 177.260 102.770 177.590 ;
        RECT 103.005 177.295 103.335 177.665 ;
        RECT 102.600 177.115 102.770 177.260 ;
        RECT 102.145 176.185 102.415 177.090 ;
        RECT 102.600 176.945 103.265 177.115 ;
        RECT 102.585 176.015 102.915 176.775 ;
        RECT 103.095 176.185 103.265 176.945 ;
        RECT 103.525 177.105 104.045 177.645 ;
        RECT 104.215 177.275 104.735 177.815 ;
        RECT 104.905 177.765 105.245 178.395 ;
        RECT 105.415 177.765 105.665 178.565 ;
        RECT 105.855 177.915 106.185 178.395 ;
        RECT 106.355 178.105 106.580 178.565 ;
        RECT 106.750 177.915 107.080 178.395 ;
        RECT 104.905 177.155 105.080 177.765 ;
        RECT 105.855 177.745 107.080 177.915 ;
        RECT 107.710 177.785 108.210 178.395 ;
        RECT 108.585 177.795 110.255 178.565 ;
        RECT 105.250 177.405 105.945 177.575 ;
        RECT 105.775 177.155 105.945 177.405 ;
        RECT 106.120 177.375 106.540 177.575 ;
        RECT 106.710 177.375 107.040 177.575 ;
        RECT 107.210 177.375 107.540 177.575 ;
        RECT 107.710 177.155 107.880 177.785 ;
        RECT 108.065 177.325 108.415 177.575 ;
        RECT 103.525 176.015 104.735 177.105 ;
        RECT 104.905 176.185 105.245 177.155 ;
        RECT 105.415 176.015 105.585 177.155 ;
        RECT 105.775 176.985 108.210 177.155 ;
        RECT 105.855 176.015 106.105 176.815 ;
        RECT 106.750 176.185 107.080 176.985 ;
        RECT 107.380 176.015 107.710 176.815 ;
        RECT 107.880 176.185 108.210 176.985 ;
        RECT 108.585 177.105 109.335 177.625 ;
        RECT 109.505 177.275 110.255 177.795 ;
        RECT 110.700 177.755 110.945 178.360 ;
        RECT 111.165 178.030 111.675 178.565 ;
        RECT 110.425 177.585 111.655 177.755 ;
        RECT 108.585 176.015 110.255 177.105 ;
        RECT 110.425 176.775 110.765 177.585 ;
        RECT 110.935 177.020 111.685 177.210 ;
        RECT 110.425 176.365 110.940 176.775 ;
        RECT 111.175 176.015 111.345 176.775 ;
        RECT 111.515 176.355 111.685 177.020 ;
        RECT 111.855 177.035 112.045 178.395 ;
        RECT 112.215 178.225 112.490 178.395 ;
        RECT 112.215 178.055 112.495 178.225 ;
        RECT 112.215 177.235 112.490 178.055 ;
        RECT 112.680 178.030 113.210 178.395 ;
        RECT 113.635 178.165 113.965 178.565 ;
        RECT 113.035 177.995 113.210 178.030 ;
        RECT 112.695 177.035 112.865 177.835 ;
        RECT 111.855 176.865 112.865 177.035 ;
        RECT 113.035 177.825 113.965 177.995 ;
        RECT 114.135 177.825 114.390 178.395 ;
        RECT 114.565 177.840 114.855 178.565 ;
        RECT 113.035 176.695 113.205 177.825 ;
        RECT 113.795 177.655 113.965 177.825 ;
        RECT 112.080 176.525 113.205 176.695 ;
        RECT 113.375 177.325 113.570 177.655 ;
        RECT 113.795 177.325 114.050 177.655 ;
        RECT 113.375 176.355 113.545 177.325 ;
        RECT 114.220 177.155 114.390 177.825 ;
        RECT 115.025 177.795 116.695 178.565 ;
        RECT 116.955 178.015 117.125 178.395 ;
        RECT 117.305 178.185 117.635 178.565 ;
        RECT 116.955 177.845 117.620 178.015 ;
        RECT 117.815 177.890 118.075 178.395 ;
        RECT 111.515 176.185 113.545 176.355 ;
        RECT 113.715 176.015 113.885 177.155 ;
        RECT 114.055 176.185 114.390 177.155 ;
        RECT 114.565 176.015 114.855 177.180 ;
        RECT 115.025 177.105 115.775 177.625 ;
        RECT 115.945 177.275 116.695 177.795 ;
        RECT 116.885 177.295 117.215 177.665 ;
        RECT 117.450 177.590 117.620 177.845 ;
        RECT 117.450 177.260 117.735 177.590 ;
        RECT 117.450 177.115 117.620 177.260 ;
        RECT 115.025 176.015 116.695 177.105 ;
        RECT 116.955 176.945 117.620 177.115 ;
        RECT 117.905 177.090 118.075 177.890 ;
        RECT 118.245 177.795 120.835 178.565 ;
        RECT 121.010 178.020 126.355 178.565 ;
        RECT 116.955 176.185 117.125 176.945 ;
        RECT 117.305 176.015 117.635 176.775 ;
        RECT 117.805 176.185 118.075 177.090 ;
        RECT 118.245 177.105 119.455 177.625 ;
        RECT 119.625 177.275 120.835 177.795 ;
        RECT 118.245 176.015 120.835 177.105 ;
        RECT 122.600 176.450 122.950 177.700 ;
        RECT 124.430 177.190 124.770 178.020 ;
        RECT 126.525 177.815 127.735 178.565 ;
        RECT 126.525 177.105 127.045 177.645 ;
        RECT 127.215 177.275 127.735 177.815 ;
        RECT 121.010 176.015 126.355 176.450 ;
        RECT 126.525 176.015 127.735 177.105 ;
        RECT 14.660 175.845 127.820 176.015 ;
        RECT 14.745 174.755 15.955 175.845 ;
        RECT 14.745 174.045 15.265 174.585 ;
        RECT 15.435 174.215 15.955 174.755 ;
        RECT 16.125 174.755 18.715 175.845 ;
        RECT 18.890 175.410 24.235 175.845 ;
        RECT 16.125 174.235 17.335 174.755 ;
        RECT 17.505 174.065 18.715 174.585 ;
        RECT 20.480 174.160 20.830 175.410 ;
        RECT 24.405 174.680 24.695 175.845 ;
        RECT 25.785 174.770 26.055 175.675 ;
        RECT 26.225 175.085 26.555 175.845 ;
        RECT 26.735 174.915 26.905 175.675 ;
        RECT 27.280 175.215 27.565 175.675 ;
        RECT 27.735 175.385 28.005 175.845 ;
        RECT 27.280 174.995 28.235 175.215 ;
        RECT 14.745 173.295 15.955 174.045 ;
        RECT 16.125 173.295 18.715 174.065 ;
        RECT 22.310 173.840 22.650 174.670 ;
        RECT 18.890 173.295 24.235 173.840 ;
        RECT 24.405 173.295 24.695 174.020 ;
        RECT 25.785 173.970 25.955 174.770 ;
        RECT 26.240 174.745 26.905 174.915 ;
        RECT 26.240 174.600 26.410 174.745 ;
        RECT 26.125 174.270 26.410 174.600 ;
        RECT 26.240 174.015 26.410 174.270 ;
        RECT 26.645 174.195 26.975 174.565 ;
        RECT 27.165 174.265 27.855 174.825 ;
        RECT 28.025 174.095 28.235 174.995 ;
        RECT 25.785 173.465 26.045 173.970 ;
        RECT 26.240 173.845 26.905 174.015 ;
        RECT 26.225 173.295 26.555 173.675 ;
        RECT 26.735 173.465 26.905 173.845 ;
        RECT 27.280 173.925 28.235 174.095 ;
        RECT 28.405 174.825 28.805 175.675 ;
        RECT 28.995 175.215 29.275 175.675 ;
        RECT 29.795 175.385 30.120 175.845 ;
        RECT 28.995 174.995 30.120 175.215 ;
        RECT 28.405 174.265 29.500 174.825 ;
        RECT 29.670 174.535 30.120 174.995 ;
        RECT 30.290 174.705 30.675 175.675 ;
        RECT 27.280 173.465 27.565 173.925 ;
        RECT 27.735 173.295 28.005 173.755 ;
        RECT 28.405 173.465 28.805 174.265 ;
        RECT 29.670 174.205 30.225 174.535 ;
        RECT 29.670 174.095 30.120 174.205 ;
        RECT 28.995 173.925 30.120 174.095 ;
        RECT 30.395 174.035 30.675 174.705 ;
        RECT 28.995 173.465 29.275 173.925 ;
        RECT 29.795 173.295 30.120 173.755 ;
        RECT 30.290 173.465 30.675 174.035 ;
        RECT 30.850 174.705 31.185 175.675 ;
        RECT 31.355 174.705 31.525 175.845 ;
        RECT 31.695 175.505 33.725 175.675 ;
        RECT 30.850 174.035 31.020 174.705 ;
        RECT 31.695 174.535 31.865 175.505 ;
        RECT 31.190 174.205 31.445 174.535 ;
        RECT 31.670 174.205 31.865 174.535 ;
        RECT 32.035 175.165 33.160 175.335 ;
        RECT 31.275 174.035 31.445 174.205 ;
        RECT 32.035 174.035 32.205 175.165 ;
        RECT 30.850 173.465 31.105 174.035 ;
        RECT 31.275 173.865 32.205 174.035 ;
        RECT 32.375 174.825 33.385 174.995 ;
        RECT 32.375 174.025 32.545 174.825 ;
        RECT 32.750 174.485 33.025 174.625 ;
        RECT 32.745 174.315 33.025 174.485 ;
        RECT 32.030 173.830 32.205 173.865 ;
        RECT 31.275 173.295 31.605 173.695 ;
        RECT 32.030 173.465 32.560 173.830 ;
        RECT 32.750 173.465 33.025 174.315 ;
        RECT 33.195 173.465 33.385 174.825 ;
        RECT 33.555 174.840 33.725 175.505 ;
        RECT 33.895 175.085 34.065 175.845 ;
        RECT 34.300 175.085 34.815 175.495 ;
        RECT 33.555 174.650 34.305 174.840 ;
        RECT 34.475 174.275 34.815 175.085 ;
        RECT 35.650 174.875 35.980 175.675 ;
        RECT 36.150 175.045 36.480 175.845 ;
        RECT 36.780 174.875 37.110 175.675 ;
        RECT 37.755 175.045 38.005 175.845 ;
        RECT 35.650 174.705 38.085 174.875 ;
        RECT 38.275 174.705 38.445 175.845 ;
        RECT 38.615 174.705 38.955 175.675 ;
        RECT 35.445 174.285 35.795 174.535 ;
        RECT 33.585 174.105 34.815 174.275 ;
        RECT 33.565 173.295 34.075 173.830 ;
        RECT 34.295 173.500 34.540 174.105 ;
        RECT 35.980 174.075 36.150 174.705 ;
        RECT 36.320 174.285 36.650 174.485 ;
        RECT 36.820 174.285 37.150 174.485 ;
        RECT 37.320 174.285 37.740 174.485 ;
        RECT 37.915 174.455 38.085 174.705 ;
        RECT 37.915 174.285 38.610 174.455 ;
        RECT 38.780 174.145 38.955 174.705 ;
        RECT 35.650 173.465 36.150 174.075 ;
        RECT 36.780 173.945 38.005 174.115 ;
        RECT 38.725 174.095 38.955 174.145 ;
        RECT 36.780 173.465 37.110 173.945 ;
        RECT 37.280 173.295 37.505 173.755 ;
        RECT 37.675 173.465 38.005 173.945 ;
        RECT 38.195 173.295 38.445 174.095 ;
        RECT 38.615 173.465 38.955 174.095 ;
        RECT 39.125 174.705 39.465 175.675 ;
        RECT 39.635 174.705 39.805 175.845 ;
        RECT 40.075 175.045 40.325 175.845 ;
        RECT 40.970 174.875 41.300 175.675 ;
        RECT 41.600 175.045 41.930 175.845 ;
        RECT 42.100 174.875 42.430 175.675 ;
        RECT 39.995 174.705 42.430 174.875 ;
        RECT 43.010 174.875 43.340 175.675 ;
        RECT 43.510 175.045 43.840 175.845 ;
        RECT 44.140 174.875 44.470 175.675 ;
        RECT 45.115 175.045 45.365 175.845 ;
        RECT 43.010 174.705 45.445 174.875 ;
        RECT 45.635 174.705 45.805 175.845 ;
        RECT 45.975 174.705 46.315 175.675 ;
        RECT 46.600 175.215 46.885 175.675 ;
        RECT 47.055 175.385 47.325 175.845 ;
        RECT 46.600 174.995 47.555 175.215 ;
        RECT 39.125 174.095 39.300 174.705 ;
        RECT 39.995 174.455 40.165 174.705 ;
        RECT 39.470 174.285 40.165 174.455 ;
        RECT 40.340 174.285 40.760 174.485 ;
        RECT 40.930 174.285 41.260 174.485 ;
        RECT 41.430 174.285 41.760 174.485 ;
        RECT 39.125 173.465 39.465 174.095 ;
        RECT 39.635 173.295 39.885 174.095 ;
        RECT 40.075 173.945 41.300 174.115 ;
        RECT 40.075 173.465 40.405 173.945 ;
        RECT 40.575 173.295 40.800 173.755 ;
        RECT 40.970 173.465 41.300 173.945 ;
        RECT 41.930 174.075 42.100 174.705 ;
        RECT 42.285 174.285 42.635 174.535 ;
        RECT 42.805 174.285 43.155 174.535 ;
        RECT 43.340 174.075 43.510 174.705 ;
        RECT 43.680 174.285 44.010 174.485 ;
        RECT 44.180 174.285 44.510 174.485 ;
        RECT 44.680 174.285 45.100 174.485 ;
        RECT 45.275 174.455 45.445 174.705 ;
        RECT 45.275 174.285 45.970 174.455 ;
        RECT 46.140 174.145 46.315 174.705 ;
        RECT 46.485 174.265 47.175 174.825 ;
        RECT 41.930 173.465 42.430 174.075 ;
        RECT 43.010 173.465 43.510 174.075 ;
        RECT 44.140 173.945 45.365 174.115 ;
        RECT 46.085 174.095 46.315 174.145 ;
        RECT 47.345 174.095 47.555 174.995 ;
        RECT 44.140 173.465 44.470 173.945 ;
        RECT 44.640 173.295 44.865 173.755 ;
        RECT 45.035 173.465 45.365 173.945 ;
        RECT 45.555 173.295 45.805 174.095 ;
        RECT 45.975 173.465 46.315 174.095 ;
        RECT 46.600 173.925 47.555 174.095 ;
        RECT 47.725 174.825 48.125 175.675 ;
        RECT 48.315 175.215 48.595 175.675 ;
        RECT 49.115 175.385 49.440 175.845 ;
        RECT 48.315 174.995 49.440 175.215 ;
        RECT 47.725 174.265 48.820 174.825 ;
        RECT 48.990 174.535 49.440 174.995 ;
        RECT 49.610 174.705 49.995 175.675 ;
        RECT 46.600 173.465 46.885 173.925 ;
        RECT 47.055 173.295 47.325 173.755 ;
        RECT 47.725 173.465 48.125 174.265 ;
        RECT 48.990 174.205 49.545 174.535 ;
        RECT 48.990 174.095 49.440 174.205 ;
        RECT 48.315 173.925 49.440 174.095 ;
        RECT 49.715 174.035 49.995 174.705 ;
        RECT 50.165 174.680 50.455 175.845 ;
        RECT 50.625 174.755 53.215 175.845 ;
        RECT 53.385 175.085 53.900 175.495 ;
        RECT 54.135 175.085 54.305 175.845 ;
        RECT 54.475 175.505 56.505 175.675 ;
        RECT 50.625 174.235 51.835 174.755 ;
        RECT 52.005 174.065 53.215 174.585 ;
        RECT 53.385 174.275 53.725 175.085 ;
        RECT 54.475 174.840 54.645 175.505 ;
        RECT 55.040 175.165 56.165 175.335 ;
        RECT 53.895 174.650 54.645 174.840 ;
        RECT 54.815 174.825 55.825 174.995 ;
        RECT 53.385 174.105 54.615 174.275 ;
        RECT 48.315 173.465 48.595 173.925 ;
        RECT 49.115 173.295 49.440 173.755 ;
        RECT 49.610 173.465 49.995 174.035 ;
        RECT 50.165 173.295 50.455 174.020 ;
        RECT 50.625 173.295 53.215 174.065 ;
        RECT 53.660 173.500 53.905 174.105 ;
        RECT 54.125 173.295 54.635 173.830 ;
        RECT 54.815 173.465 55.005 174.825 ;
        RECT 55.175 174.485 55.450 174.625 ;
        RECT 55.175 174.315 55.455 174.485 ;
        RECT 55.175 173.465 55.450 174.315 ;
        RECT 55.655 174.025 55.825 174.825 ;
        RECT 55.995 174.035 56.165 175.165 ;
        RECT 56.335 174.535 56.505 175.505 ;
        RECT 56.675 174.705 56.845 175.845 ;
        RECT 57.015 174.705 57.350 175.675 ;
        RECT 56.335 174.205 56.530 174.535 ;
        RECT 56.755 174.205 57.010 174.535 ;
        RECT 56.755 174.035 56.925 174.205 ;
        RECT 57.180 174.035 57.350 174.705 ;
        RECT 55.995 173.865 56.925 174.035 ;
        RECT 55.995 173.830 56.170 173.865 ;
        RECT 55.640 173.465 56.170 173.830 ;
        RECT 56.595 173.295 56.925 173.695 ;
        RECT 57.095 173.465 57.350 174.035 ;
        RECT 57.530 174.655 57.785 175.535 ;
        RECT 57.955 174.705 58.260 175.845 ;
        RECT 58.600 175.465 58.930 175.845 ;
        RECT 59.110 175.295 59.280 175.585 ;
        RECT 59.450 175.385 59.700 175.845 ;
        RECT 58.480 175.125 59.280 175.295 ;
        RECT 59.870 175.335 60.740 175.675 ;
        RECT 57.530 174.005 57.740 174.655 ;
        RECT 58.480 174.535 58.650 175.125 ;
        RECT 59.870 174.955 60.040 175.335 ;
        RECT 60.975 175.215 61.145 175.675 ;
        RECT 61.315 175.385 61.685 175.845 ;
        RECT 61.980 175.245 62.150 175.585 ;
        RECT 62.320 175.415 62.650 175.845 ;
        RECT 62.885 175.245 63.055 175.585 ;
        RECT 58.820 174.785 60.040 174.955 ;
        RECT 60.210 174.875 60.670 175.165 ;
        RECT 60.975 175.045 61.535 175.215 ;
        RECT 61.980 175.075 63.055 175.245 ;
        RECT 63.225 175.345 63.905 175.675 ;
        RECT 64.120 175.345 64.370 175.675 ;
        RECT 64.540 175.385 64.790 175.845 ;
        RECT 61.365 174.905 61.535 175.045 ;
        RECT 60.210 174.865 61.175 174.875 ;
        RECT 59.870 174.695 60.040 174.785 ;
        RECT 60.500 174.705 61.175 174.865 ;
        RECT 57.910 174.505 58.650 174.535 ;
        RECT 57.910 174.205 58.825 174.505 ;
        RECT 58.500 174.030 58.825 174.205 ;
        RECT 57.530 173.475 57.785 174.005 ;
        RECT 57.955 173.295 58.260 173.755 ;
        RECT 58.505 173.675 58.825 174.030 ;
        RECT 58.995 174.245 59.535 174.615 ;
        RECT 59.870 174.525 60.275 174.695 ;
        RECT 58.995 173.845 59.235 174.245 ;
        RECT 59.715 174.075 59.935 174.355 ;
        RECT 59.405 173.905 59.935 174.075 ;
        RECT 59.405 173.675 59.575 173.905 ;
        RECT 60.105 173.745 60.275 174.525 ;
        RECT 60.445 173.915 60.795 174.535 ;
        RECT 60.965 173.915 61.175 174.705 ;
        RECT 61.365 174.735 62.865 174.905 ;
        RECT 61.365 174.045 61.535 174.735 ;
        RECT 63.225 174.565 63.395 175.345 ;
        RECT 64.200 175.215 64.370 175.345 ;
        RECT 61.705 174.395 63.395 174.565 ;
        RECT 63.565 174.785 64.030 175.175 ;
        RECT 64.200 175.045 64.595 175.215 ;
        RECT 61.705 174.215 61.875 174.395 ;
        RECT 58.505 173.505 59.575 173.675 ;
        RECT 59.745 173.295 59.935 173.735 ;
        RECT 60.105 173.465 61.055 173.745 ;
        RECT 61.365 173.655 61.625 174.045 ;
        RECT 62.045 173.975 62.835 174.225 ;
        RECT 61.275 173.485 61.625 173.655 ;
        RECT 61.835 173.295 62.165 173.755 ;
        RECT 63.040 173.685 63.210 174.395 ;
        RECT 63.565 174.195 63.735 174.785 ;
        RECT 63.380 173.975 63.735 174.195 ;
        RECT 63.905 173.975 64.255 174.595 ;
        RECT 64.425 173.685 64.595 175.045 ;
        RECT 64.960 174.875 65.285 175.660 ;
        RECT 64.765 173.825 65.225 174.875 ;
        RECT 63.040 173.515 63.895 173.685 ;
        RECT 64.100 173.515 64.595 173.685 ;
        RECT 64.765 173.295 65.095 173.655 ;
        RECT 65.455 173.555 65.625 175.675 ;
        RECT 65.795 175.345 66.125 175.845 ;
        RECT 66.295 175.175 66.550 175.675 ;
        RECT 65.800 175.005 66.550 175.175 ;
        RECT 65.800 174.015 66.030 175.005 ;
        RECT 66.200 174.185 66.550 174.835 ;
        RECT 66.725 174.755 68.395 175.845 ;
        RECT 68.575 174.865 68.905 175.675 ;
        RECT 69.075 175.045 69.315 175.845 ;
        RECT 66.725 174.235 67.475 174.755 ;
        RECT 68.575 174.695 69.290 174.865 ;
        RECT 67.645 174.065 68.395 174.585 ;
        RECT 68.570 174.285 68.950 174.525 ;
        RECT 69.120 174.455 69.290 174.695 ;
        RECT 69.495 174.825 69.665 175.675 ;
        RECT 69.835 175.045 70.165 175.845 ;
        RECT 70.335 174.825 70.505 175.675 ;
        RECT 69.495 174.655 70.505 174.825 ;
        RECT 70.675 174.695 71.005 175.845 ;
        RECT 71.330 174.695 71.590 175.845 ;
        RECT 71.765 174.770 72.020 175.675 ;
        RECT 72.190 175.085 72.520 175.845 ;
        RECT 72.735 174.915 72.905 175.675 ;
        RECT 69.120 174.285 69.620 174.455 ;
        RECT 69.120 174.115 69.290 174.285 ;
        RECT 70.010 174.115 70.505 174.655 ;
        RECT 65.800 173.845 66.550 174.015 ;
        RECT 65.795 173.295 66.125 173.675 ;
        RECT 66.295 173.555 66.550 173.845 ;
        RECT 66.725 173.295 68.395 174.065 ;
        RECT 68.655 173.945 69.290 174.115 ;
        RECT 69.495 173.945 70.505 174.115 ;
        RECT 68.655 173.465 68.825 173.945 ;
        RECT 69.005 173.295 69.245 173.775 ;
        RECT 69.495 173.465 69.665 173.945 ;
        RECT 69.835 173.295 70.165 173.775 ;
        RECT 70.335 173.465 70.505 173.945 ;
        RECT 70.675 173.295 71.005 174.095 ;
        RECT 71.330 173.295 71.590 174.135 ;
        RECT 71.765 174.040 71.935 174.770 ;
        RECT 72.190 174.745 72.905 174.915 ;
        RECT 73.165 174.755 75.755 175.845 ;
        RECT 72.190 174.535 72.360 174.745 ;
        RECT 72.105 174.205 72.360 174.535 ;
        RECT 71.765 173.465 72.020 174.040 ;
        RECT 72.190 174.015 72.360 174.205 ;
        RECT 72.640 174.195 72.995 174.565 ;
        RECT 73.165 174.235 74.375 174.755 ;
        RECT 75.925 174.680 76.215 175.845 ;
        RECT 77.305 174.755 80.815 175.845 ;
        RECT 74.545 174.065 75.755 174.585 ;
        RECT 77.305 174.235 78.995 174.755 ;
        RECT 80.985 174.705 81.325 175.675 ;
        RECT 81.495 174.705 81.665 175.845 ;
        RECT 81.935 175.045 82.185 175.845 ;
        RECT 82.830 174.875 83.160 175.675 ;
        RECT 83.460 175.045 83.790 175.845 ;
        RECT 83.960 174.875 84.290 175.675 ;
        RECT 85.130 175.410 90.475 175.845 ;
        RECT 90.650 175.410 95.995 175.845 ;
        RECT 96.170 175.410 101.515 175.845 ;
        RECT 81.855 174.705 84.290 174.875 ;
        RECT 79.165 174.065 80.815 174.585 ;
        RECT 72.190 173.845 72.905 174.015 ;
        RECT 72.190 173.295 72.520 173.675 ;
        RECT 72.735 173.465 72.905 173.845 ;
        RECT 73.165 173.295 75.755 174.065 ;
        RECT 75.925 173.295 76.215 174.020 ;
        RECT 77.305 173.295 80.815 174.065 ;
        RECT 80.985 174.145 81.160 174.705 ;
        RECT 81.855 174.455 82.025 174.705 ;
        RECT 81.330 174.285 82.025 174.455 ;
        RECT 82.200 174.285 82.620 174.485 ;
        RECT 82.790 174.285 83.120 174.485 ;
        RECT 83.290 174.285 83.620 174.485 ;
        RECT 80.985 174.095 81.215 174.145 ;
        RECT 80.985 173.465 81.325 174.095 ;
        RECT 81.495 173.295 81.745 174.095 ;
        RECT 81.935 173.945 83.160 174.115 ;
        RECT 81.935 173.465 82.265 173.945 ;
        RECT 82.435 173.295 82.660 173.755 ;
        RECT 82.830 173.465 83.160 173.945 ;
        RECT 83.790 174.075 83.960 174.705 ;
        RECT 84.145 174.285 84.495 174.535 ;
        RECT 86.720 174.160 87.070 175.410 ;
        RECT 83.790 173.465 84.290 174.075 ;
        RECT 88.550 173.840 88.890 174.670 ;
        RECT 92.240 174.160 92.590 175.410 ;
        RECT 94.070 173.840 94.410 174.670 ;
        RECT 97.760 174.160 98.110 175.410 ;
        RECT 101.685 174.680 101.975 175.845 ;
        RECT 102.145 174.755 103.815 175.845 ;
        RECT 104.190 174.875 104.520 175.675 ;
        RECT 104.690 175.045 105.020 175.845 ;
        RECT 105.320 174.875 105.650 175.675 ;
        RECT 106.295 175.045 106.545 175.845 ;
        RECT 99.590 173.840 99.930 174.670 ;
        RECT 102.145 174.235 102.895 174.755 ;
        RECT 104.190 174.705 106.625 174.875 ;
        RECT 106.815 174.705 106.985 175.845 ;
        RECT 107.155 174.705 107.495 175.675 ;
        RECT 103.065 174.065 103.815 174.585 ;
        RECT 103.985 174.285 104.335 174.535 ;
        RECT 104.520 174.075 104.690 174.705 ;
        RECT 104.860 174.285 105.190 174.485 ;
        RECT 105.360 174.285 105.690 174.485 ;
        RECT 105.860 174.285 106.280 174.485 ;
        RECT 106.455 174.455 106.625 174.705 ;
        RECT 106.455 174.285 107.150 174.455 ;
        RECT 85.130 173.295 90.475 173.840 ;
        RECT 90.650 173.295 95.995 173.840 ;
        RECT 96.170 173.295 101.515 173.840 ;
        RECT 101.685 173.295 101.975 174.020 ;
        RECT 102.145 173.295 103.815 174.065 ;
        RECT 104.190 173.465 104.690 174.075 ;
        RECT 105.320 173.945 106.545 174.115 ;
        RECT 107.320 174.095 107.495 174.705 ;
        RECT 105.320 173.465 105.650 173.945 ;
        RECT 105.820 173.295 106.045 173.755 ;
        RECT 106.215 173.465 106.545 173.945 ;
        RECT 106.735 173.295 106.985 174.095 ;
        RECT 107.155 173.465 107.495 174.095 ;
        RECT 107.665 174.705 108.005 175.675 ;
        RECT 108.175 174.705 108.345 175.845 ;
        RECT 108.615 175.045 108.865 175.845 ;
        RECT 109.510 174.875 109.840 175.675 ;
        RECT 110.140 175.045 110.470 175.845 ;
        RECT 110.640 174.875 110.970 175.675 ;
        RECT 108.535 174.705 110.970 174.875 ;
        RECT 111.345 174.755 112.555 175.845 ;
        RECT 112.730 175.410 118.075 175.845 ;
        RECT 107.665 174.145 107.840 174.705 ;
        RECT 108.535 174.455 108.705 174.705 ;
        RECT 108.010 174.285 108.705 174.455 ;
        RECT 108.880 174.285 109.300 174.485 ;
        RECT 109.470 174.285 109.800 174.485 ;
        RECT 109.970 174.285 110.300 174.485 ;
        RECT 107.665 174.095 107.895 174.145 ;
        RECT 107.665 173.465 108.005 174.095 ;
        RECT 108.175 173.295 108.425 174.095 ;
        RECT 108.615 173.945 109.840 174.115 ;
        RECT 108.615 173.465 108.945 173.945 ;
        RECT 109.115 173.295 109.340 173.755 ;
        RECT 109.510 173.465 109.840 173.945 ;
        RECT 110.470 174.075 110.640 174.705 ;
        RECT 110.825 174.285 111.175 174.535 ;
        RECT 111.345 174.215 111.865 174.755 ;
        RECT 110.470 173.465 110.970 174.075 ;
        RECT 112.035 174.045 112.555 174.585 ;
        RECT 114.320 174.160 114.670 175.410 ;
        RECT 118.285 174.705 118.515 175.845 ;
        RECT 118.685 174.695 119.015 175.675 ;
        RECT 119.185 174.705 119.395 175.845 ;
        RECT 119.625 174.755 120.835 175.845 ;
        RECT 121.010 175.410 126.355 175.845 ;
        RECT 111.345 173.295 112.555 174.045 ;
        RECT 116.150 173.840 116.490 174.670 ;
        RECT 118.265 174.285 118.595 174.535 ;
        RECT 112.730 173.295 118.075 173.840 ;
        RECT 118.285 173.295 118.515 174.115 ;
        RECT 118.765 174.095 119.015 174.695 ;
        RECT 119.625 174.215 120.145 174.755 ;
        RECT 118.685 173.465 119.015 174.095 ;
        RECT 119.185 173.295 119.395 174.115 ;
        RECT 120.315 174.045 120.835 174.585 ;
        RECT 122.600 174.160 122.950 175.410 ;
        RECT 126.525 174.755 127.735 175.845 ;
        RECT 119.625 173.295 120.835 174.045 ;
        RECT 124.430 173.840 124.770 174.670 ;
        RECT 126.525 174.215 127.045 174.755 ;
        RECT 127.215 174.045 127.735 174.585 ;
        RECT 121.010 173.295 126.355 173.840 ;
        RECT 126.525 173.295 127.735 174.045 ;
        RECT 14.660 173.125 127.820 173.295 ;
        RECT 14.745 172.375 15.955 173.125 ;
        RECT 14.745 171.835 15.265 172.375 ;
        RECT 17.045 172.355 20.555 173.125 ;
        RECT 20.730 172.580 26.075 173.125 ;
        RECT 26.250 172.580 31.595 173.125 ;
        RECT 31.770 172.580 37.115 173.125 ;
        RECT 15.435 171.665 15.955 172.205 ;
        RECT 14.745 170.575 15.955 171.665 ;
        RECT 17.045 171.665 18.735 172.185 ;
        RECT 18.905 171.835 20.555 172.355 ;
        RECT 17.045 170.575 20.555 171.665 ;
        RECT 22.320 171.010 22.670 172.260 ;
        RECT 24.150 171.750 24.490 172.580 ;
        RECT 27.840 171.010 28.190 172.260 ;
        RECT 29.670 171.750 30.010 172.580 ;
        RECT 33.360 171.010 33.710 172.260 ;
        RECT 35.190 171.750 35.530 172.580 ;
        RECT 37.285 172.400 37.575 173.125 ;
        RECT 37.745 172.325 38.085 172.955 ;
        RECT 38.255 172.325 38.505 173.125 ;
        RECT 38.695 172.475 39.025 172.955 ;
        RECT 39.195 172.665 39.420 173.125 ;
        RECT 39.590 172.475 39.920 172.955 ;
        RECT 20.730 170.575 26.075 171.010 ;
        RECT 26.250 170.575 31.595 171.010 ;
        RECT 31.770 170.575 37.115 171.010 ;
        RECT 37.285 170.575 37.575 171.740 ;
        RECT 37.745 171.715 37.920 172.325 ;
        RECT 38.695 172.305 39.920 172.475 ;
        RECT 40.550 172.345 41.050 172.955 ;
        RECT 41.885 172.450 42.145 172.955 ;
        RECT 42.325 172.745 42.655 173.125 ;
        RECT 42.835 172.575 43.005 172.955 ;
        RECT 38.090 171.965 38.785 172.135 ;
        RECT 38.615 171.715 38.785 171.965 ;
        RECT 38.960 171.935 39.380 172.135 ;
        RECT 39.550 171.935 39.880 172.135 ;
        RECT 40.050 171.935 40.380 172.135 ;
        RECT 40.550 171.715 40.720 172.345 ;
        RECT 40.905 171.885 41.255 172.135 ;
        RECT 37.745 170.745 38.085 171.715 ;
        RECT 38.255 170.575 38.425 171.715 ;
        RECT 38.615 171.545 41.050 171.715 ;
        RECT 38.695 170.575 38.945 171.375 ;
        RECT 39.590 170.745 39.920 171.545 ;
        RECT 40.220 170.575 40.550 171.375 ;
        RECT 40.720 170.745 41.050 171.545 ;
        RECT 41.885 171.650 42.055 172.450 ;
        RECT 42.340 172.405 43.005 172.575 ;
        RECT 42.340 172.150 42.510 172.405 ;
        RECT 44.185 172.325 44.525 172.955 ;
        RECT 44.695 172.325 44.945 173.125 ;
        RECT 45.135 172.475 45.465 172.955 ;
        RECT 45.635 172.665 45.860 173.125 ;
        RECT 46.030 172.475 46.360 172.955 ;
        RECT 42.225 171.820 42.510 172.150 ;
        RECT 42.745 171.855 43.075 172.225 ;
        RECT 42.340 171.675 42.510 171.820 ;
        RECT 44.185 171.715 44.360 172.325 ;
        RECT 45.135 172.305 46.360 172.475 ;
        RECT 46.990 172.345 47.490 172.955 ;
        RECT 44.530 171.965 45.225 172.135 ;
        RECT 45.055 171.715 45.225 171.965 ;
        RECT 45.400 171.935 45.820 172.135 ;
        RECT 45.990 171.935 46.320 172.135 ;
        RECT 46.490 171.935 46.820 172.135 ;
        RECT 46.990 171.715 47.160 172.345 ;
        RECT 47.865 172.325 48.205 172.955 ;
        RECT 48.375 172.325 48.625 173.125 ;
        RECT 48.815 172.475 49.145 172.955 ;
        RECT 49.315 172.665 49.540 173.125 ;
        RECT 49.710 172.475 50.040 172.955 ;
        RECT 47.345 171.885 47.695 172.135 ;
        RECT 47.865 171.715 48.040 172.325 ;
        RECT 48.815 172.305 50.040 172.475 ;
        RECT 50.670 172.345 51.170 172.955 ;
        RECT 48.210 171.965 48.905 172.135 ;
        RECT 48.735 171.715 48.905 171.965 ;
        RECT 49.080 171.935 49.500 172.135 ;
        RECT 49.670 171.935 50.000 172.135 ;
        RECT 50.170 171.935 50.500 172.135 ;
        RECT 50.670 171.715 50.840 172.345 ;
        RECT 51.545 172.325 51.885 172.955 ;
        RECT 52.055 172.325 52.305 173.125 ;
        RECT 52.495 172.475 52.825 172.955 ;
        RECT 52.995 172.665 53.220 173.125 ;
        RECT 53.390 172.475 53.720 172.955 ;
        RECT 51.025 171.885 51.375 172.135 ;
        RECT 51.545 171.715 51.720 172.325 ;
        RECT 52.495 172.305 53.720 172.475 ;
        RECT 54.350 172.345 54.850 172.955 ;
        RECT 55.225 172.375 56.435 173.125 ;
        RECT 51.890 171.965 52.585 172.135 ;
        RECT 52.415 171.715 52.585 171.965 ;
        RECT 52.760 171.935 53.180 172.135 ;
        RECT 53.350 171.935 53.680 172.135 ;
        RECT 53.850 171.935 54.180 172.135 ;
        RECT 54.350 171.715 54.520 172.345 ;
        RECT 54.705 171.885 55.055 172.135 ;
        RECT 41.885 170.745 42.155 171.650 ;
        RECT 42.340 171.505 43.005 171.675 ;
        RECT 42.325 170.575 42.655 171.335 ;
        RECT 42.835 170.745 43.005 171.505 ;
        RECT 44.185 170.745 44.525 171.715 ;
        RECT 44.695 170.575 44.865 171.715 ;
        RECT 45.055 171.545 47.490 171.715 ;
        RECT 45.135 170.575 45.385 171.375 ;
        RECT 46.030 170.745 46.360 171.545 ;
        RECT 46.660 170.575 46.990 171.375 ;
        RECT 47.160 170.745 47.490 171.545 ;
        RECT 47.865 170.745 48.205 171.715 ;
        RECT 48.375 170.575 48.545 171.715 ;
        RECT 48.735 171.545 51.170 171.715 ;
        RECT 48.815 170.575 49.065 171.375 ;
        RECT 49.710 170.745 50.040 171.545 ;
        RECT 50.340 170.575 50.670 171.375 ;
        RECT 50.840 170.745 51.170 171.545 ;
        RECT 51.545 170.745 51.885 171.715 ;
        RECT 52.055 170.575 52.225 171.715 ;
        RECT 52.415 171.545 54.850 171.715 ;
        RECT 52.495 170.575 52.745 171.375 ;
        RECT 53.390 170.745 53.720 171.545 ;
        RECT 54.020 170.575 54.350 171.375 ;
        RECT 54.520 170.745 54.850 171.545 ;
        RECT 55.225 171.665 55.745 172.205 ;
        RECT 55.915 171.835 56.435 172.375 ;
        RECT 56.605 172.355 60.115 173.125 ;
        RECT 56.605 171.665 58.295 172.185 ;
        RECT 58.465 171.835 60.115 172.355 ;
        RECT 60.345 172.305 60.555 173.125 ;
        RECT 60.725 172.325 61.055 172.955 ;
        RECT 60.725 171.725 60.975 172.325 ;
        RECT 61.225 172.305 61.455 173.125 ;
        RECT 61.755 172.575 61.925 172.955 ;
        RECT 62.105 172.745 62.435 173.125 ;
        RECT 61.755 172.405 62.420 172.575 ;
        RECT 62.615 172.450 62.875 172.955 ;
        RECT 61.145 171.885 61.475 172.135 ;
        RECT 61.685 171.855 62.015 172.225 ;
        RECT 62.250 172.150 62.420 172.405 ;
        RECT 62.250 171.820 62.535 172.150 ;
        RECT 55.225 170.575 56.435 171.665 ;
        RECT 56.605 170.575 60.115 171.665 ;
        RECT 60.345 170.575 60.555 171.715 ;
        RECT 60.725 170.745 61.055 171.725 ;
        RECT 61.225 170.575 61.455 171.715 ;
        RECT 62.250 171.675 62.420 171.820 ;
        RECT 61.755 171.505 62.420 171.675 ;
        RECT 62.705 171.650 62.875 172.450 ;
        RECT 63.045 172.400 63.335 173.125 ;
        RECT 63.965 172.355 65.635 173.125 ;
        RECT 65.810 172.580 71.155 173.125 ;
        RECT 71.330 172.580 76.675 173.125 ;
        RECT 76.850 172.580 82.195 173.125 ;
        RECT 61.755 170.745 61.925 171.505 ;
        RECT 62.105 170.575 62.435 171.335 ;
        RECT 62.605 170.745 62.875 171.650 ;
        RECT 63.045 170.575 63.335 171.740 ;
        RECT 63.965 171.665 64.715 172.185 ;
        RECT 64.885 171.835 65.635 172.355 ;
        RECT 63.965 170.575 65.635 171.665 ;
        RECT 67.400 171.010 67.750 172.260 ;
        RECT 69.230 171.750 69.570 172.580 ;
        RECT 72.920 171.010 73.270 172.260 ;
        RECT 74.750 171.750 75.090 172.580 ;
        RECT 78.440 171.010 78.790 172.260 ;
        RECT 80.270 171.750 80.610 172.580 ;
        RECT 82.455 172.475 82.625 172.955 ;
        RECT 82.805 172.645 83.045 173.125 ;
        RECT 83.295 172.475 83.465 172.955 ;
        RECT 83.635 172.645 83.965 173.125 ;
        RECT 84.135 172.475 84.305 172.955 ;
        RECT 82.455 172.305 83.090 172.475 ;
        RECT 83.295 172.305 84.305 172.475 ;
        RECT 84.475 172.325 84.805 173.125 ;
        RECT 85.240 172.495 85.525 172.955 ;
        RECT 85.695 172.665 85.965 173.125 ;
        RECT 85.240 172.325 86.195 172.495 ;
        RECT 82.920 172.135 83.090 172.305 ;
        RECT 83.805 172.275 84.305 172.305 ;
        RECT 82.370 171.895 82.750 172.135 ;
        RECT 82.920 171.965 83.420 172.135 ;
        RECT 82.920 171.725 83.090 171.965 ;
        RECT 83.810 171.765 84.305 172.275 ;
        RECT 82.375 171.555 83.090 171.725 ;
        RECT 83.295 171.595 84.305 171.765 ;
        RECT 65.810 170.575 71.155 171.010 ;
        RECT 71.330 170.575 76.675 171.010 ;
        RECT 76.850 170.575 82.195 171.010 ;
        RECT 82.375 170.745 82.705 171.555 ;
        RECT 82.875 170.575 83.115 171.375 ;
        RECT 83.295 170.745 83.465 171.595 ;
        RECT 83.635 170.575 83.965 171.375 ;
        RECT 84.135 170.745 84.305 171.595 ;
        RECT 84.475 170.575 84.805 171.725 ;
        RECT 85.125 171.595 85.815 172.155 ;
        RECT 85.985 171.425 86.195 172.325 ;
        RECT 85.240 171.205 86.195 171.425 ;
        RECT 86.365 172.155 86.765 172.955 ;
        RECT 86.955 172.495 87.235 172.955 ;
        RECT 87.755 172.665 88.080 173.125 ;
        RECT 86.955 172.325 88.080 172.495 ;
        RECT 88.250 172.385 88.635 172.955 ;
        RECT 88.805 172.400 89.095 173.125 ;
        RECT 87.630 172.215 88.080 172.325 ;
        RECT 86.365 171.595 87.460 172.155 ;
        RECT 87.630 171.885 88.185 172.215 ;
        RECT 85.240 170.745 85.525 171.205 ;
        RECT 85.695 170.575 85.965 171.035 ;
        RECT 86.365 170.745 86.765 171.595 ;
        RECT 87.630 171.425 88.080 171.885 ;
        RECT 88.355 171.715 88.635 172.385 ;
        RECT 89.765 172.305 89.995 173.125 ;
        RECT 90.165 172.325 90.495 172.955 ;
        RECT 89.745 171.885 90.075 172.135 ;
        RECT 86.955 171.205 88.080 171.425 ;
        RECT 86.955 170.745 87.235 171.205 ;
        RECT 87.755 170.575 88.080 171.035 ;
        RECT 88.250 170.745 88.635 171.715 ;
        RECT 88.805 170.575 89.095 171.740 ;
        RECT 90.245 171.725 90.495 172.325 ;
        RECT 90.665 172.305 90.875 173.125 ;
        RECT 91.110 172.415 91.365 172.945 ;
        RECT 91.535 172.665 91.840 173.125 ;
        RECT 92.085 172.745 93.155 172.915 ;
        RECT 89.765 170.575 89.995 171.715 ;
        RECT 90.165 170.745 90.495 171.725 ;
        RECT 91.110 171.765 91.320 172.415 ;
        RECT 92.085 172.390 92.405 172.745 ;
        RECT 92.080 172.215 92.405 172.390 ;
        RECT 91.490 171.915 92.405 172.215 ;
        RECT 92.575 172.175 92.815 172.575 ;
        RECT 92.985 172.515 93.155 172.745 ;
        RECT 93.325 172.685 93.515 173.125 ;
        RECT 93.685 172.675 94.635 172.955 ;
        RECT 94.855 172.765 95.205 172.935 ;
        RECT 92.985 172.345 93.515 172.515 ;
        RECT 91.490 171.885 92.230 171.915 ;
        RECT 90.665 170.575 90.875 171.715 ;
        RECT 91.110 170.885 91.365 171.765 ;
        RECT 91.535 170.575 91.840 171.715 ;
        RECT 92.060 171.295 92.230 171.885 ;
        RECT 92.575 171.805 93.115 172.175 ;
        RECT 93.295 172.065 93.515 172.345 ;
        RECT 93.685 171.895 93.855 172.675 ;
        RECT 93.450 171.725 93.855 171.895 ;
        RECT 94.025 171.885 94.375 172.505 ;
        RECT 93.450 171.635 93.620 171.725 ;
        RECT 94.545 171.715 94.755 172.505 ;
        RECT 92.400 171.465 93.620 171.635 ;
        RECT 94.080 171.555 94.755 171.715 ;
        RECT 92.060 171.125 92.860 171.295 ;
        RECT 92.180 170.575 92.510 170.955 ;
        RECT 92.690 170.835 92.860 171.125 ;
        RECT 93.450 171.085 93.620 171.465 ;
        RECT 93.790 171.545 94.755 171.555 ;
        RECT 94.945 172.375 95.205 172.765 ;
        RECT 95.415 172.665 95.745 173.125 ;
        RECT 96.620 172.735 97.475 172.905 ;
        RECT 97.680 172.735 98.175 172.905 ;
        RECT 98.345 172.765 98.675 173.125 ;
        RECT 94.945 171.685 95.115 172.375 ;
        RECT 95.285 172.025 95.455 172.205 ;
        RECT 95.625 172.195 96.415 172.445 ;
        RECT 96.620 172.025 96.790 172.735 ;
        RECT 96.960 172.225 97.315 172.445 ;
        RECT 95.285 171.855 96.975 172.025 ;
        RECT 93.790 171.255 94.250 171.545 ;
        RECT 94.945 171.515 96.445 171.685 ;
        RECT 94.945 171.375 95.115 171.515 ;
        RECT 94.555 171.205 95.115 171.375 ;
        RECT 93.030 170.575 93.280 171.035 ;
        RECT 93.450 170.745 94.320 171.085 ;
        RECT 94.555 170.745 94.725 171.205 ;
        RECT 95.560 171.175 96.635 171.345 ;
        RECT 94.895 170.575 95.265 171.035 ;
        RECT 95.560 170.835 95.730 171.175 ;
        RECT 95.900 170.575 96.230 171.005 ;
        RECT 96.465 170.835 96.635 171.175 ;
        RECT 96.805 171.075 96.975 171.855 ;
        RECT 97.145 171.635 97.315 172.225 ;
        RECT 97.485 171.825 97.835 172.445 ;
        RECT 97.145 171.245 97.610 171.635 ;
        RECT 98.005 171.375 98.175 172.735 ;
        RECT 98.345 171.545 98.805 172.595 ;
        RECT 97.780 171.205 98.175 171.375 ;
        RECT 97.780 171.075 97.950 171.205 ;
        RECT 96.805 170.745 97.485 171.075 ;
        RECT 97.700 170.745 97.950 171.075 ;
        RECT 98.120 170.575 98.370 171.035 ;
        RECT 98.540 170.760 98.865 171.545 ;
        RECT 99.035 170.745 99.205 172.865 ;
        RECT 99.375 172.745 99.705 173.125 ;
        RECT 99.875 172.575 100.130 172.865 ;
        RECT 101.230 172.580 106.575 173.125 ;
        RECT 99.380 172.405 100.130 172.575 ;
        RECT 99.380 171.415 99.610 172.405 ;
        RECT 99.780 171.585 100.130 172.235 ;
        RECT 99.380 171.245 100.130 171.415 ;
        RECT 99.375 170.575 99.705 171.075 ;
        RECT 99.875 170.745 100.130 171.245 ;
        RECT 102.820 171.010 103.170 172.260 ;
        RECT 104.650 171.750 104.990 172.580 ;
        RECT 106.805 172.305 107.015 173.125 ;
        RECT 107.185 172.325 107.515 172.955 ;
        RECT 107.185 171.725 107.435 172.325 ;
        RECT 107.685 172.305 107.915 173.125 ;
        RECT 108.330 172.345 108.830 172.955 ;
        RECT 107.605 171.885 107.935 172.135 ;
        RECT 108.125 171.885 108.475 172.135 ;
        RECT 101.230 170.575 106.575 171.010 ;
        RECT 106.805 170.575 107.015 171.715 ;
        RECT 107.185 170.745 107.515 171.725 ;
        RECT 108.660 171.715 108.830 172.345 ;
        RECT 109.460 172.475 109.790 172.955 ;
        RECT 109.960 172.665 110.185 173.125 ;
        RECT 110.355 172.475 110.685 172.955 ;
        RECT 109.460 172.305 110.685 172.475 ;
        RECT 110.875 172.325 111.125 173.125 ;
        RECT 111.295 172.325 111.635 172.955 ;
        RECT 111.805 172.375 113.015 173.125 ;
        RECT 109.000 171.935 109.330 172.135 ;
        RECT 109.500 171.935 109.830 172.135 ;
        RECT 110.000 171.935 110.420 172.135 ;
        RECT 110.595 171.965 111.290 172.135 ;
        RECT 110.595 171.715 110.765 171.965 ;
        RECT 111.460 171.715 111.635 172.325 ;
        RECT 107.685 170.575 107.915 171.715 ;
        RECT 108.330 171.545 110.765 171.715 ;
        RECT 108.330 170.745 108.660 171.545 ;
        RECT 108.830 170.575 109.160 171.375 ;
        RECT 109.460 170.745 109.790 171.545 ;
        RECT 110.435 170.575 110.685 171.375 ;
        RECT 110.955 170.575 111.125 171.715 ;
        RECT 111.295 170.745 111.635 171.715 ;
        RECT 111.805 171.665 112.325 172.205 ;
        RECT 112.495 171.835 113.015 172.375 ;
        RECT 113.225 172.305 113.455 173.125 ;
        RECT 113.625 172.325 113.955 172.955 ;
        RECT 113.205 171.885 113.535 172.135 ;
        RECT 113.705 171.725 113.955 172.325 ;
        RECT 114.125 172.305 114.335 173.125 ;
        RECT 114.565 172.400 114.855 173.125 ;
        RECT 115.950 172.415 116.205 172.945 ;
        RECT 116.375 172.665 116.680 173.125 ;
        RECT 116.925 172.745 117.995 172.915 ;
        RECT 115.950 171.765 116.160 172.415 ;
        RECT 116.925 172.390 117.245 172.745 ;
        RECT 116.920 172.215 117.245 172.390 ;
        RECT 116.330 171.915 117.245 172.215 ;
        RECT 117.415 172.175 117.655 172.575 ;
        RECT 117.825 172.515 117.995 172.745 ;
        RECT 118.165 172.685 118.355 173.125 ;
        RECT 118.525 172.675 119.475 172.955 ;
        RECT 119.695 172.765 120.045 172.935 ;
        RECT 117.825 172.345 118.355 172.515 ;
        RECT 116.330 171.885 117.070 171.915 ;
        RECT 111.805 170.575 113.015 171.665 ;
        RECT 113.225 170.575 113.455 171.715 ;
        RECT 113.625 170.745 113.955 171.725 ;
        RECT 114.125 170.575 114.335 171.715 ;
        RECT 114.565 170.575 114.855 171.740 ;
        RECT 115.950 170.885 116.205 171.765 ;
        RECT 116.375 170.575 116.680 171.715 ;
        RECT 116.900 171.295 117.070 171.885 ;
        RECT 117.415 171.805 117.955 172.175 ;
        RECT 118.135 172.065 118.355 172.345 ;
        RECT 118.525 171.895 118.695 172.675 ;
        RECT 118.290 171.725 118.695 171.895 ;
        RECT 118.865 171.885 119.215 172.505 ;
        RECT 118.290 171.635 118.460 171.725 ;
        RECT 119.385 171.715 119.595 172.505 ;
        RECT 117.240 171.465 118.460 171.635 ;
        RECT 118.920 171.555 119.595 171.715 ;
        RECT 116.900 171.125 117.700 171.295 ;
        RECT 117.020 170.575 117.350 170.955 ;
        RECT 117.530 170.835 117.700 171.125 ;
        RECT 118.290 171.085 118.460 171.465 ;
        RECT 118.630 171.545 119.595 171.555 ;
        RECT 119.785 172.375 120.045 172.765 ;
        RECT 120.255 172.665 120.585 173.125 ;
        RECT 121.460 172.735 122.315 172.905 ;
        RECT 122.520 172.735 123.015 172.905 ;
        RECT 123.185 172.765 123.515 173.125 ;
        RECT 119.785 171.685 119.955 172.375 ;
        RECT 120.125 172.025 120.295 172.205 ;
        RECT 120.465 172.195 121.255 172.445 ;
        RECT 121.460 172.025 121.630 172.735 ;
        RECT 121.800 172.225 122.155 172.445 ;
        RECT 120.125 171.855 121.815 172.025 ;
        RECT 118.630 171.255 119.090 171.545 ;
        RECT 119.785 171.515 121.285 171.685 ;
        RECT 119.785 171.375 119.955 171.515 ;
        RECT 119.395 171.205 119.955 171.375 ;
        RECT 117.870 170.575 118.120 171.035 ;
        RECT 118.290 170.745 119.160 171.085 ;
        RECT 119.395 170.745 119.565 171.205 ;
        RECT 120.400 171.175 121.475 171.345 ;
        RECT 119.735 170.575 120.105 171.035 ;
        RECT 120.400 170.835 120.570 171.175 ;
        RECT 120.740 170.575 121.070 171.005 ;
        RECT 121.305 170.835 121.475 171.175 ;
        RECT 121.645 171.075 121.815 171.855 ;
        RECT 121.985 171.635 122.155 172.225 ;
        RECT 122.325 171.825 122.675 172.445 ;
        RECT 121.985 171.245 122.450 171.635 ;
        RECT 122.845 171.375 123.015 172.735 ;
        RECT 123.185 171.545 123.645 172.595 ;
        RECT 122.620 171.205 123.015 171.375 ;
        RECT 122.620 171.075 122.790 171.205 ;
        RECT 121.645 170.745 122.325 171.075 ;
        RECT 122.540 170.745 122.790 171.075 ;
        RECT 122.960 170.575 123.210 171.035 ;
        RECT 123.380 170.760 123.705 171.545 ;
        RECT 123.875 170.745 124.045 172.865 ;
        RECT 124.215 172.745 124.545 173.125 ;
        RECT 124.715 172.575 124.970 172.865 ;
        RECT 124.220 172.405 124.970 172.575 ;
        RECT 124.220 171.415 124.450 172.405 ;
        RECT 125.145 172.375 126.355 173.125 ;
        RECT 126.525 172.375 127.735 173.125 ;
        RECT 124.620 171.585 124.970 172.235 ;
        RECT 125.145 171.665 125.665 172.205 ;
        RECT 125.835 171.835 126.355 172.375 ;
        RECT 126.525 171.665 127.045 172.205 ;
        RECT 127.215 171.835 127.735 172.375 ;
        RECT 124.220 171.245 124.970 171.415 ;
        RECT 124.215 170.575 124.545 171.075 ;
        RECT 124.715 170.745 124.970 171.245 ;
        RECT 125.145 170.575 126.355 171.665 ;
        RECT 126.525 170.575 127.735 171.665 ;
        RECT 14.660 170.405 127.820 170.575 ;
        RECT 14.745 169.315 15.955 170.405 ;
        RECT 14.745 168.605 15.265 169.145 ;
        RECT 15.435 168.775 15.955 169.315 ;
        RECT 16.125 169.315 18.715 170.405 ;
        RECT 18.890 169.970 24.235 170.405 ;
        RECT 16.125 168.795 17.335 169.315 ;
        RECT 17.505 168.625 18.715 169.145 ;
        RECT 20.480 168.720 20.830 169.970 ;
        RECT 24.405 169.240 24.695 170.405 ;
        RECT 25.325 169.315 26.995 170.405 ;
        RECT 14.745 167.855 15.955 168.605 ;
        RECT 16.125 167.855 18.715 168.625 ;
        RECT 22.310 168.400 22.650 169.230 ;
        RECT 25.325 168.795 26.075 169.315 ;
        RECT 27.205 169.265 27.435 170.405 ;
        RECT 27.605 169.255 27.935 170.235 ;
        RECT 28.105 169.265 28.315 170.405 ;
        RECT 29.005 169.315 32.515 170.405 ;
        RECT 26.245 168.625 26.995 169.145 ;
        RECT 27.185 168.845 27.515 169.095 ;
        RECT 18.890 167.855 24.235 168.400 ;
        RECT 24.405 167.855 24.695 168.580 ;
        RECT 25.325 167.855 26.995 168.625 ;
        RECT 27.205 167.855 27.435 168.675 ;
        RECT 27.685 168.655 27.935 169.255 ;
        RECT 29.005 168.795 30.695 169.315 ;
        RECT 32.745 169.265 32.955 170.405 ;
        RECT 33.125 169.255 33.455 170.235 ;
        RECT 33.625 169.265 33.855 170.405 ;
        RECT 34.065 169.315 35.275 170.405 ;
        RECT 35.535 169.660 35.805 170.405 ;
        RECT 36.435 170.400 42.710 170.405 ;
        RECT 35.975 169.490 36.265 170.230 ;
        RECT 36.435 169.675 36.690 170.400 ;
        RECT 36.875 169.505 37.135 170.230 ;
        RECT 37.305 169.675 37.550 170.400 ;
        RECT 37.735 169.505 37.995 170.230 ;
        RECT 38.165 169.675 38.410 170.400 ;
        RECT 38.595 169.505 38.855 170.230 ;
        RECT 39.025 169.675 39.270 170.400 ;
        RECT 39.440 169.505 39.700 170.230 ;
        RECT 39.870 169.675 40.130 170.400 ;
        RECT 40.300 169.505 40.560 170.230 ;
        RECT 40.730 169.675 40.990 170.400 ;
        RECT 41.160 169.505 41.420 170.230 ;
        RECT 41.590 169.675 41.850 170.400 ;
        RECT 42.020 169.505 42.280 170.230 ;
        RECT 42.450 169.605 42.710 170.400 ;
        RECT 36.875 169.490 42.280 169.505 ;
        RECT 27.605 168.025 27.935 168.655 ;
        RECT 28.105 167.855 28.315 168.675 ;
        RECT 30.865 168.625 32.515 169.145 ;
        RECT 29.005 167.855 32.515 168.625 ;
        RECT 32.745 167.855 32.955 168.675 ;
        RECT 33.125 168.655 33.375 169.255 ;
        RECT 33.545 168.845 33.875 169.095 ;
        RECT 34.065 168.775 34.585 169.315 ;
        RECT 35.535 169.265 42.280 169.490 ;
        RECT 33.125 168.025 33.455 168.655 ;
        RECT 33.625 167.855 33.855 168.675 ;
        RECT 34.755 168.605 35.275 169.145 ;
        RECT 34.065 167.855 35.275 168.605 ;
        RECT 35.535 168.675 36.700 169.265 ;
        RECT 42.880 169.095 43.130 170.230 ;
        RECT 43.310 169.595 43.570 170.405 ;
        RECT 43.745 169.095 43.990 170.235 ;
        RECT 44.170 169.595 44.465 170.405 ;
        RECT 44.650 169.970 49.995 170.405 ;
        RECT 36.870 168.845 43.990 169.095 ;
        RECT 35.535 168.505 42.280 168.675 ;
        RECT 35.535 167.855 35.835 168.335 ;
        RECT 36.005 168.050 36.265 168.505 ;
        RECT 36.435 167.855 36.695 168.335 ;
        RECT 36.875 168.050 37.135 168.505 ;
        RECT 37.305 167.855 37.555 168.335 ;
        RECT 37.735 168.050 37.995 168.505 ;
        RECT 38.165 167.855 38.415 168.335 ;
        RECT 38.595 168.050 38.855 168.505 ;
        RECT 39.025 167.855 39.270 168.335 ;
        RECT 39.440 168.050 39.715 168.505 ;
        RECT 39.885 167.855 40.130 168.335 ;
        RECT 40.300 168.050 40.560 168.505 ;
        RECT 40.730 167.855 40.990 168.335 ;
        RECT 41.160 168.050 41.420 168.505 ;
        RECT 41.590 167.855 41.850 168.335 ;
        RECT 42.020 168.050 42.280 168.505 ;
        RECT 42.450 167.855 42.710 168.415 ;
        RECT 42.880 168.035 43.130 168.845 ;
        RECT 43.310 167.855 43.570 168.380 ;
        RECT 43.740 168.035 43.990 168.845 ;
        RECT 44.160 168.535 44.475 169.095 ;
        RECT 46.240 168.720 46.590 169.970 ;
        RECT 50.165 169.240 50.455 170.405 ;
        RECT 50.625 169.315 51.835 170.405 ;
        RECT 52.010 169.970 57.355 170.405 ;
        RECT 57.530 169.970 62.875 170.405 ;
        RECT 63.050 169.970 68.395 170.405 ;
        RECT 48.070 168.400 48.410 169.230 ;
        RECT 50.625 168.775 51.145 169.315 ;
        RECT 51.315 168.605 51.835 169.145 ;
        RECT 53.600 168.720 53.950 169.970 ;
        RECT 44.170 167.855 44.475 168.365 ;
        RECT 44.650 167.855 49.995 168.400 ;
        RECT 50.165 167.855 50.455 168.580 ;
        RECT 50.625 167.855 51.835 168.605 ;
        RECT 55.430 168.400 55.770 169.230 ;
        RECT 59.120 168.720 59.470 169.970 ;
        RECT 60.950 168.400 61.290 169.230 ;
        RECT 64.640 168.720 64.990 169.970 ;
        RECT 68.570 169.255 68.830 170.405 ;
        RECT 69.005 169.330 69.260 170.235 ;
        RECT 69.430 169.645 69.760 170.405 ;
        RECT 69.975 169.475 70.145 170.235 ;
        RECT 66.470 168.400 66.810 169.230 ;
        RECT 52.010 167.855 57.355 168.400 ;
        RECT 57.530 167.855 62.875 168.400 ;
        RECT 63.050 167.855 68.395 168.400 ;
        RECT 68.570 167.855 68.830 168.695 ;
        RECT 69.005 168.600 69.175 169.330 ;
        RECT 69.430 169.305 70.145 169.475 ;
        RECT 69.430 169.095 69.600 169.305 ;
        RECT 70.410 169.255 70.670 170.405 ;
        RECT 70.845 169.330 71.100 170.235 ;
        RECT 71.270 169.645 71.600 170.405 ;
        RECT 71.815 169.475 71.985 170.235 ;
        RECT 69.345 168.765 69.600 169.095 ;
        RECT 69.005 168.025 69.260 168.600 ;
        RECT 69.430 168.575 69.600 168.765 ;
        RECT 69.880 168.755 70.235 169.125 ;
        RECT 69.430 168.405 70.145 168.575 ;
        RECT 69.430 167.855 69.760 168.235 ;
        RECT 69.975 168.025 70.145 168.405 ;
        RECT 70.410 167.855 70.670 168.695 ;
        RECT 70.845 168.600 71.015 169.330 ;
        RECT 71.270 169.305 71.985 169.475 ;
        RECT 72.245 169.315 75.755 170.405 ;
        RECT 71.270 169.095 71.440 169.305 ;
        RECT 71.185 168.765 71.440 169.095 ;
        RECT 70.845 168.025 71.100 168.600 ;
        RECT 71.270 168.575 71.440 168.765 ;
        RECT 71.720 168.755 72.075 169.125 ;
        RECT 72.245 168.795 73.935 169.315 ;
        RECT 75.925 169.240 76.215 170.405 ;
        RECT 76.385 169.645 76.900 170.055 ;
        RECT 77.135 169.645 77.305 170.405 ;
        RECT 77.475 170.065 79.505 170.235 ;
        RECT 74.105 168.625 75.755 169.145 ;
        RECT 76.385 168.835 76.725 169.645 ;
        RECT 77.475 169.400 77.645 170.065 ;
        RECT 78.040 169.725 79.165 169.895 ;
        RECT 76.895 169.210 77.645 169.400 ;
        RECT 77.815 169.385 78.825 169.555 ;
        RECT 76.385 168.665 77.615 168.835 ;
        RECT 71.270 168.405 71.985 168.575 ;
        RECT 71.270 167.855 71.600 168.235 ;
        RECT 71.815 168.025 71.985 168.405 ;
        RECT 72.245 167.855 75.755 168.625 ;
        RECT 75.925 167.855 76.215 168.580 ;
        RECT 76.660 168.060 76.905 168.665 ;
        RECT 77.125 167.855 77.635 168.390 ;
        RECT 77.815 168.025 78.005 169.385 ;
        RECT 78.175 168.365 78.450 169.185 ;
        RECT 78.655 168.585 78.825 169.385 ;
        RECT 78.995 168.595 79.165 169.725 ;
        RECT 79.335 169.095 79.505 170.065 ;
        RECT 79.675 169.265 79.845 170.405 ;
        RECT 80.015 169.265 80.350 170.235 ;
        RECT 79.335 168.765 79.530 169.095 ;
        RECT 79.755 168.765 80.010 169.095 ;
        RECT 79.755 168.595 79.925 168.765 ;
        RECT 80.180 168.595 80.350 169.265 ;
        RECT 80.900 169.425 81.155 170.095 ;
        RECT 81.335 169.605 81.620 170.405 ;
        RECT 81.800 169.685 82.130 170.195 ;
        RECT 80.900 168.705 81.080 169.425 ;
        RECT 81.800 169.095 82.050 169.685 ;
        RECT 82.400 169.535 82.570 170.145 ;
        RECT 82.740 169.715 83.070 170.405 ;
        RECT 83.300 169.855 83.540 170.145 ;
        RECT 83.740 170.025 84.160 170.405 ;
        RECT 84.340 169.935 84.970 170.185 ;
        RECT 85.440 170.025 85.770 170.405 ;
        RECT 84.340 169.855 84.510 169.935 ;
        RECT 85.940 169.855 86.110 170.145 ;
        RECT 86.290 170.025 86.670 170.405 ;
        RECT 86.910 170.020 87.740 170.190 ;
        RECT 83.300 169.685 84.510 169.855 ;
        RECT 81.250 168.765 82.050 169.095 ;
        RECT 78.995 168.425 79.925 168.595 ;
        RECT 78.995 168.390 79.170 168.425 ;
        RECT 78.175 168.195 78.455 168.365 ;
        RECT 78.175 168.025 78.450 168.195 ;
        RECT 78.640 168.025 79.170 168.390 ;
        RECT 79.595 167.855 79.925 168.255 ;
        RECT 80.095 168.025 80.350 168.595 ;
        RECT 80.815 168.565 81.080 168.705 ;
        RECT 80.815 168.535 81.155 168.565 ;
        RECT 80.900 168.035 81.155 168.535 ;
        RECT 81.335 167.855 81.620 168.315 ;
        RECT 81.800 168.115 82.050 168.765 ;
        RECT 82.250 169.515 82.570 169.535 ;
        RECT 82.250 169.345 84.170 169.515 ;
        RECT 82.250 168.450 82.440 169.345 ;
        RECT 84.340 169.175 84.510 169.685 ;
        RECT 84.680 169.425 85.200 169.735 ;
        RECT 82.610 169.005 84.510 169.175 ;
        RECT 82.610 168.945 82.940 169.005 ;
        RECT 83.090 168.775 83.420 168.835 ;
        RECT 82.760 168.505 83.420 168.775 ;
        RECT 82.250 168.120 82.570 168.450 ;
        RECT 82.750 167.855 83.410 168.335 ;
        RECT 83.610 168.245 83.780 169.005 ;
        RECT 84.680 168.835 84.860 169.245 ;
        RECT 83.950 168.665 84.280 168.785 ;
        RECT 85.030 168.665 85.200 169.425 ;
        RECT 83.950 168.495 85.200 168.665 ;
        RECT 85.370 169.605 86.740 169.855 ;
        RECT 85.370 168.835 85.560 169.605 ;
        RECT 86.490 169.345 86.740 169.605 ;
        RECT 85.730 169.175 85.980 169.335 ;
        RECT 86.910 169.175 87.080 170.020 ;
        RECT 87.975 169.735 88.145 170.235 ;
        RECT 88.315 169.905 88.645 170.405 ;
        RECT 87.250 169.345 87.750 169.725 ;
        RECT 87.975 169.565 88.670 169.735 ;
        RECT 85.730 169.005 87.080 169.175 ;
        RECT 86.660 168.965 87.080 169.005 ;
        RECT 85.370 168.495 85.790 168.835 ;
        RECT 86.080 168.505 86.490 168.835 ;
        RECT 83.610 168.075 84.460 168.245 ;
        RECT 85.020 167.855 85.340 168.315 ;
        RECT 85.540 168.065 85.790 168.495 ;
        RECT 86.080 167.855 86.490 168.295 ;
        RECT 86.660 168.235 86.830 168.965 ;
        RECT 87.000 168.415 87.350 168.785 ;
        RECT 87.530 168.475 87.750 169.345 ;
        RECT 87.920 168.775 88.330 169.395 ;
        RECT 88.500 168.595 88.670 169.565 ;
        RECT 87.975 168.405 88.670 168.595 ;
        RECT 86.660 168.035 87.675 168.235 ;
        RECT 87.975 168.075 88.145 168.405 ;
        RECT 88.315 167.855 88.645 168.235 ;
        RECT 88.860 168.115 89.085 170.235 ;
        RECT 89.255 169.905 89.585 170.405 ;
        RECT 89.755 169.735 89.925 170.235 ;
        RECT 89.260 169.565 89.925 169.735 ;
        RECT 89.260 168.575 89.490 169.565 ;
        RECT 89.660 168.745 90.010 169.395 ;
        RECT 90.185 169.315 91.395 170.405 ;
        RECT 91.565 169.645 92.080 170.055 ;
        RECT 92.315 169.645 92.485 170.405 ;
        RECT 92.655 170.065 94.685 170.235 ;
        RECT 90.185 168.775 90.705 169.315 ;
        RECT 90.875 168.605 91.395 169.145 ;
        RECT 91.565 168.835 91.905 169.645 ;
        RECT 92.655 169.400 92.825 170.065 ;
        RECT 93.220 169.725 94.345 169.895 ;
        RECT 92.075 169.210 92.825 169.400 ;
        RECT 92.995 169.385 94.005 169.555 ;
        RECT 91.565 168.665 92.795 168.835 ;
        RECT 89.260 168.405 89.925 168.575 ;
        RECT 89.255 167.855 89.585 168.235 ;
        RECT 89.755 168.115 89.925 168.405 ;
        RECT 90.185 167.855 91.395 168.605 ;
        RECT 91.840 168.060 92.085 168.665 ;
        RECT 92.305 167.855 92.815 168.390 ;
        RECT 92.995 168.025 93.185 169.385 ;
        RECT 93.355 169.045 93.630 169.185 ;
        RECT 93.355 168.875 93.635 169.045 ;
        RECT 93.355 168.025 93.630 168.875 ;
        RECT 93.835 168.585 94.005 169.385 ;
        RECT 94.175 168.595 94.345 169.725 ;
        RECT 94.515 169.095 94.685 170.065 ;
        RECT 94.855 169.265 95.025 170.405 ;
        RECT 95.195 169.265 95.530 170.235 ;
        RECT 96.255 169.475 96.425 170.235 ;
        RECT 96.605 169.645 96.935 170.405 ;
        RECT 96.255 169.305 96.920 169.475 ;
        RECT 97.105 169.330 97.375 170.235 ;
        RECT 94.515 168.765 94.710 169.095 ;
        RECT 94.935 168.765 95.190 169.095 ;
        RECT 94.935 168.595 95.105 168.765 ;
        RECT 95.360 168.595 95.530 169.265 ;
        RECT 96.750 169.160 96.920 169.305 ;
        RECT 96.185 168.755 96.515 169.125 ;
        RECT 96.750 168.830 97.035 169.160 ;
        RECT 94.175 168.425 95.105 168.595 ;
        RECT 94.175 168.390 94.350 168.425 ;
        RECT 93.820 168.025 94.350 168.390 ;
        RECT 94.775 167.855 95.105 168.255 ;
        RECT 95.275 168.025 95.530 168.595 ;
        RECT 96.750 168.575 96.920 168.830 ;
        RECT 96.255 168.405 96.920 168.575 ;
        RECT 97.205 168.530 97.375 169.330 ;
        RECT 98.005 169.315 101.515 170.405 ;
        RECT 98.005 168.795 99.695 169.315 ;
        RECT 101.685 169.240 101.975 170.405 ;
        RECT 103.070 169.215 103.325 170.095 ;
        RECT 103.495 169.265 103.800 170.405 ;
        RECT 104.140 170.025 104.470 170.405 ;
        RECT 104.650 169.855 104.820 170.145 ;
        RECT 104.990 169.945 105.240 170.405 ;
        RECT 104.020 169.685 104.820 169.855 ;
        RECT 105.410 169.895 106.280 170.235 ;
        RECT 99.865 168.625 101.515 169.145 ;
        RECT 96.255 168.025 96.425 168.405 ;
        RECT 96.605 167.855 96.935 168.235 ;
        RECT 97.115 168.025 97.375 168.530 ;
        RECT 98.005 167.855 101.515 168.625 ;
        RECT 101.685 167.855 101.975 168.580 ;
        RECT 103.070 168.565 103.280 169.215 ;
        RECT 104.020 169.095 104.190 169.685 ;
        RECT 105.410 169.515 105.580 169.895 ;
        RECT 106.515 169.775 106.685 170.235 ;
        RECT 106.855 169.945 107.225 170.405 ;
        RECT 107.520 169.805 107.690 170.145 ;
        RECT 107.860 169.975 108.190 170.405 ;
        RECT 108.425 169.805 108.595 170.145 ;
        RECT 104.360 169.345 105.580 169.515 ;
        RECT 105.750 169.435 106.210 169.725 ;
        RECT 106.515 169.605 107.075 169.775 ;
        RECT 107.520 169.635 108.595 169.805 ;
        RECT 108.765 169.905 109.445 170.235 ;
        RECT 109.660 169.905 109.910 170.235 ;
        RECT 110.080 169.945 110.330 170.405 ;
        RECT 106.905 169.465 107.075 169.605 ;
        RECT 105.750 169.425 106.715 169.435 ;
        RECT 105.410 169.255 105.580 169.345 ;
        RECT 106.040 169.265 106.715 169.425 ;
        RECT 103.450 169.065 104.190 169.095 ;
        RECT 103.450 168.765 104.365 169.065 ;
        RECT 104.040 168.590 104.365 168.765 ;
        RECT 103.070 168.035 103.325 168.565 ;
        RECT 103.495 167.855 103.800 168.315 ;
        RECT 104.045 168.235 104.365 168.590 ;
        RECT 104.535 168.805 105.075 169.175 ;
        RECT 105.410 169.085 105.815 169.255 ;
        RECT 104.535 168.405 104.775 168.805 ;
        RECT 105.255 168.635 105.475 168.915 ;
        RECT 104.945 168.465 105.475 168.635 ;
        RECT 104.945 168.235 105.115 168.465 ;
        RECT 105.645 168.305 105.815 169.085 ;
        RECT 105.985 168.475 106.335 169.095 ;
        RECT 106.505 168.475 106.715 169.265 ;
        RECT 106.905 169.295 108.405 169.465 ;
        RECT 106.905 168.605 107.075 169.295 ;
        RECT 108.765 169.125 108.935 169.905 ;
        RECT 109.740 169.775 109.910 169.905 ;
        RECT 107.245 168.955 108.935 169.125 ;
        RECT 109.105 169.345 109.570 169.735 ;
        RECT 109.740 169.605 110.135 169.775 ;
        RECT 107.245 168.775 107.415 168.955 ;
        RECT 104.045 168.065 105.115 168.235 ;
        RECT 105.285 167.855 105.475 168.295 ;
        RECT 105.645 168.025 106.595 168.305 ;
        RECT 106.905 168.215 107.165 168.605 ;
        RECT 107.585 168.535 108.375 168.785 ;
        RECT 106.815 168.045 107.165 168.215 ;
        RECT 107.375 167.855 107.705 168.315 ;
        RECT 108.580 168.245 108.750 168.955 ;
        RECT 109.105 168.755 109.275 169.345 ;
        RECT 108.920 168.535 109.275 168.755 ;
        RECT 109.445 168.535 109.795 169.155 ;
        RECT 109.965 168.245 110.135 169.605 ;
        RECT 110.500 169.435 110.825 170.220 ;
        RECT 110.305 168.385 110.765 169.435 ;
        RECT 108.580 168.075 109.435 168.245 ;
        RECT 109.640 168.075 110.135 168.245 ;
        RECT 110.305 167.855 110.635 168.215 ;
        RECT 110.995 168.115 111.165 170.235 ;
        RECT 111.335 169.905 111.665 170.405 ;
        RECT 111.835 169.735 112.090 170.235 ;
        RECT 111.340 169.565 112.090 169.735 ;
        RECT 111.340 168.575 111.570 169.565 ;
        RECT 111.740 168.745 112.090 169.395 ;
        RECT 112.730 169.265 113.065 170.235 ;
        RECT 113.235 169.265 113.405 170.405 ;
        RECT 113.575 170.065 115.605 170.235 ;
        RECT 112.730 168.595 112.900 169.265 ;
        RECT 113.575 169.095 113.745 170.065 ;
        RECT 113.070 168.765 113.325 169.095 ;
        RECT 113.550 168.765 113.745 169.095 ;
        RECT 113.915 169.725 115.040 169.895 ;
        RECT 113.155 168.595 113.325 168.765 ;
        RECT 113.915 168.595 114.085 169.725 ;
        RECT 111.340 168.405 112.090 168.575 ;
        RECT 111.335 167.855 111.665 168.235 ;
        RECT 111.835 168.115 112.090 168.405 ;
        RECT 112.730 168.025 112.985 168.595 ;
        RECT 113.155 168.425 114.085 168.595 ;
        RECT 114.255 169.385 115.265 169.555 ;
        RECT 114.255 168.585 114.425 169.385 ;
        RECT 114.630 169.045 114.905 169.185 ;
        RECT 114.625 168.875 114.905 169.045 ;
        RECT 113.910 168.390 114.085 168.425 ;
        RECT 113.155 167.855 113.485 168.255 ;
        RECT 113.910 168.025 114.440 168.390 ;
        RECT 114.630 168.025 114.905 168.875 ;
        RECT 115.075 168.025 115.265 169.385 ;
        RECT 115.435 169.400 115.605 170.065 ;
        RECT 115.775 169.645 115.945 170.405 ;
        RECT 116.180 169.645 116.695 170.055 ;
        RECT 115.435 169.210 116.185 169.400 ;
        RECT 116.355 168.835 116.695 169.645 ;
        RECT 115.465 168.665 116.695 168.835 ;
        RECT 116.865 169.265 117.250 170.235 ;
        RECT 117.420 169.945 117.745 170.405 ;
        RECT 118.265 169.775 118.545 170.235 ;
        RECT 117.420 169.555 118.545 169.775 ;
        RECT 115.445 167.855 115.955 168.390 ;
        RECT 116.175 168.060 116.420 168.665 ;
        RECT 116.865 168.595 117.145 169.265 ;
        RECT 117.420 169.095 117.870 169.555 ;
        RECT 118.735 169.385 119.135 170.235 ;
        RECT 119.535 169.945 119.805 170.405 ;
        RECT 119.975 169.775 120.260 170.235 ;
        RECT 117.315 168.765 117.870 169.095 ;
        RECT 118.040 168.825 119.135 169.385 ;
        RECT 117.420 168.655 117.870 168.765 ;
        RECT 116.865 168.025 117.250 168.595 ;
        RECT 117.420 168.485 118.545 168.655 ;
        RECT 117.420 167.855 117.745 168.315 ;
        RECT 118.265 168.025 118.545 168.485 ;
        RECT 118.735 168.025 119.135 168.825 ;
        RECT 119.305 169.555 120.260 169.775 ;
        RECT 119.305 168.655 119.515 169.555 ;
        RECT 120.635 169.475 120.805 170.235 ;
        RECT 120.985 169.645 121.315 170.405 ;
        RECT 119.685 168.825 120.375 169.385 ;
        RECT 120.635 169.305 121.300 169.475 ;
        RECT 121.485 169.330 121.755 170.235 ;
        RECT 121.930 169.980 122.265 170.405 ;
        RECT 122.435 169.800 122.620 170.205 ;
        RECT 121.130 169.160 121.300 169.305 ;
        RECT 120.565 168.755 120.895 169.125 ;
        RECT 121.130 168.830 121.415 169.160 ;
        RECT 119.305 168.485 120.260 168.655 ;
        RECT 121.130 168.575 121.300 168.830 ;
        RECT 119.535 167.855 119.805 168.315 ;
        RECT 119.975 168.025 120.260 168.485 ;
        RECT 120.635 168.405 121.300 168.575 ;
        RECT 121.585 168.530 121.755 169.330 ;
        RECT 120.635 168.025 120.805 168.405 ;
        RECT 120.985 167.855 121.315 168.235 ;
        RECT 121.495 168.025 121.755 168.530 ;
        RECT 121.955 169.625 122.620 169.800 ;
        RECT 122.825 169.625 123.155 170.405 ;
        RECT 121.955 168.595 122.295 169.625 ;
        RECT 123.325 169.435 123.595 170.205 ;
        RECT 122.465 169.265 123.595 169.435 ;
        RECT 122.465 168.765 122.715 169.265 ;
        RECT 121.955 168.425 122.640 168.595 ;
        RECT 122.895 168.515 123.255 169.095 ;
        RECT 121.930 167.855 122.265 168.255 ;
        RECT 122.435 168.025 122.640 168.425 ;
        RECT 123.425 168.355 123.595 169.265 ;
        RECT 123.765 169.315 126.355 170.405 ;
        RECT 126.525 169.315 127.735 170.405 ;
        RECT 123.765 168.795 124.975 169.315 ;
        RECT 125.145 168.625 126.355 169.145 ;
        RECT 126.525 168.775 127.045 169.315 ;
        RECT 122.850 167.855 123.125 168.335 ;
        RECT 123.335 168.025 123.595 168.355 ;
        RECT 123.765 167.855 126.355 168.625 ;
        RECT 127.215 168.605 127.735 169.145 ;
        RECT 126.525 167.855 127.735 168.605 ;
        RECT 14.660 167.685 127.820 167.855 ;
        RECT 14.745 166.935 15.955 167.685 ;
        RECT 14.745 166.395 15.265 166.935 ;
        RECT 16.125 166.915 17.795 167.685 ;
        RECT 17.970 167.140 23.315 167.685 ;
        RECT 15.435 166.225 15.955 166.765 ;
        RECT 14.745 165.135 15.955 166.225 ;
        RECT 16.125 166.225 16.875 166.745 ;
        RECT 17.045 166.395 17.795 166.915 ;
        RECT 16.125 165.135 17.795 166.225 ;
        RECT 19.560 165.570 19.910 166.820 ;
        RECT 21.390 166.310 21.730 167.140 ;
        RECT 23.490 167.135 23.745 167.425 ;
        RECT 23.915 167.305 24.245 167.685 ;
        RECT 23.490 166.965 24.240 167.135 ;
        RECT 23.490 166.145 23.840 166.795 ;
        RECT 24.010 165.975 24.240 166.965 ;
        RECT 23.490 165.805 24.240 165.975 ;
        RECT 17.970 165.135 23.315 165.570 ;
        RECT 23.490 165.305 23.745 165.805 ;
        RECT 23.915 165.135 24.245 165.635 ;
        RECT 24.415 165.305 24.585 167.425 ;
        RECT 24.945 167.325 25.275 167.685 ;
        RECT 25.445 167.295 25.940 167.465 ;
        RECT 26.145 167.295 27.000 167.465 ;
        RECT 24.815 166.105 25.275 167.155 ;
        RECT 24.755 165.320 25.080 166.105 ;
        RECT 25.445 165.935 25.615 167.295 ;
        RECT 25.785 166.385 26.135 167.005 ;
        RECT 26.305 166.785 26.660 167.005 ;
        RECT 26.305 166.195 26.475 166.785 ;
        RECT 26.830 166.585 27.000 167.295 ;
        RECT 27.875 167.225 28.205 167.685 ;
        RECT 28.415 167.325 28.765 167.495 ;
        RECT 27.205 166.755 27.995 167.005 ;
        RECT 28.415 166.935 28.675 167.325 ;
        RECT 28.985 167.235 29.935 167.515 ;
        RECT 30.105 167.245 30.295 167.685 ;
        RECT 30.465 167.305 31.535 167.475 ;
        RECT 28.165 166.585 28.335 166.765 ;
        RECT 25.445 165.765 25.840 165.935 ;
        RECT 26.010 165.805 26.475 166.195 ;
        RECT 26.645 166.415 28.335 166.585 ;
        RECT 25.670 165.635 25.840 165.765 ;
        RECT 26.645 165.635 26.815 166.415 ;
        RECT 28.505 166.245 28.675 166.935 ;
        RECT 27.175 166.075 28.675 166.245 ;
        RECT 28.865 166.275 29.075 167.065 ;
        RECT 29.245 166.445 29.595 167.065 ;
        RECT 29.765 166.455 29.935 167.235 ;
        RECT 30.465 167.075 30.635 167.305 ;
        RECT 30.105 166.905 30.635 167.075 ;
        RECT 30.105 166.625 30.325 166.905 ;
        RECT 30.805 166.735 31.045 167.135 ;
        RECT 29.765 166.285 30.170 166.455 ;
        RECT 30.505 166.365 31.045 166.735 ;
        RECT 31.215 166.950 31.535 167.305 ;
        RECT 31.780 167.225 32.085 167.685 ;
        RECT 32.255 166.975 32.510 167.505 ;
        RECT 31.215 166.775 31.540 166.950 ;
        RECT 31.215 166.475 32.130 166.775 ;
        RECT 31.390 166.445 32.130 166.475 ;
        RECT 28.865 166.115 29.540 166.275 ;
        RECT 30.000 166.195 30.170 166.285 ;
        RECT 28.865 166.105 29.830 166.115 ;
        RECT 28.505 165.935 28.675 166.075 ;
        RECT 25.250 165.135 25.500 165.595 ;
        RECT 25.670 165.305 25.920 165.635 ;
        RECT 26.135 165.305 26.815 165.635 ;
        RECT 26.985 165.735 28.060 165.905 ;
        RECT 28.505 165.765 29.065 165.935 ;
        RECT 29.370 165.815 29.830 166.105 ;
        RECT 30.000 166.025 31.220 166.195 ;
        RECT 26.985 165.395 27.155 165.735 ;
        RECT 27.390 165.135 27.720 165.565 ;
        RECT 27.890 165.395 28.060 165.735 ;
        RECT 28.355 165.135 28.725 165.595 ;
        RECT 28.895 165.305 29.065 165.765 ;
        RECT 30.000 165.645 30.170 166.025 ;
        RECT 31.390 165.855 31.560 166.445 ;
        RECT 32.300 166.325 32.510 166.975 ;
        RECT 29.300 165.305 30.170 165.645 ;
        RECT 30.760 165.685 31.560 165.855 ;
        RECT 30.340 165.135 30.590 165.595 ;
        RECT 30.760 165.395 30.930 165.685 ;
        RECT 31.110 165.135 31.440 165.515 ;
        RECT 31.780 165.135 32.085 166.275 ;
        RECT 32.255 165.445 32.510 166.325 ;
        RECT 32.685 167.010 32.945 167.515 ;
        RECT 33.125 167.305 33.455 167.685 ;
        RECT 33.635 167.135 33.805 167.515 ;
        RECT 34.165 167.220 34.415 167.685 ;
        RECT 32.685 166.210 32.855 167.010 ;
        RECT 33.140 166.965 33.805 167.135 ;
        RECT 34.585 167.045 34.755 167.515 ;
        RECT 35.005 167.225 35.175 167.685 ;
        RECT 35.425 167.045 35.595 167.515 ;
        RECT 35.845 167.225 36.015 167.685 ;
        RECT 36.265 167.045 36.435 167.515 ;
        RECT 36.805 167.225 37.070 167.685 ;
        RECT 33.140 166.710 33.310 166.965 ;
        RECT 34.065 166.865 36.435 167.045 ;
        RECT 37.285 166.960 37.575 167.685 ;
        RECT 37.785 166.865 38.015 167.685 ;
        RECT 38.185 166.885 38.515 167.515 ;
        RECT 33.025 166.380 33.310 166.710 ;
        RECT 33.545 166.415 33.875 166.785 ;
        RECT 33.140 166.235 33.310 166.380 ;
        RECT 34.065 166.275 34.415 166.865 ;
        RECT 34.585 166.445 37.095 166.695 ;
        RECT 37.765 166.445 38.095 166.695 ;
        RECT 32.685 165.305 32.955 166.210 ;
        RECT 33.140 166.065 33.805 166.235 ;
        RECT 34.065 166.105 36.515 166.275 ;
        RECT 34.065 166.085 34.835 166.105 ;
        RECT 33.125 165.135 33.455 165.895 ;
        RECT 33.635 165.305 33.805 166.065 ;
        RECT 34.165 165.135 34.335 165.595 ;
        RECT 34.505 165.305 34.835 166.085 ;
        RECT 35.005 165.135 35.175 165.935 ;
        RECT 35.345 165.305 35.675 166.105 ;
        RECT 35.845 165.135 36.015 165.935 ;
        RECT 36.185 165.305 36.515 166.105 ;
        RECT 36.775 165.135 37.070 166.275 ;
        RECT 37.285 165.135 37.575 166.300 ;
        RECT 38.265 166.285 38.515 166.885 ;
        RECT 38.685 166.865 38.895 167.685 ;
        RECT 39.240 167.055 39.525 167.515 ;
        RECT 39.695 167.225 39.965 167.685 ;
        RECT 39.240 166.885 40.195 167.055 ;
        RECT 37.785 165.135 38.015 166.275 ;
        RECT 38.185 165.305 38.515 166.285 ;
        RECT 38.685 165.135 38.895 166.275 ;
        RECT 39.125 166.155 39.815 166.715 ;
        RECT 39.985 165.985 40.195 166.885 ;
        RECT 39.240 165.765 40.195 165.985 ;
        RECT 40.365 166.715 40.765 167.515 ;
        RECT 40.955 167.055 41.235 167.515 ;
        RECT 41.755 167.225 42.080 167.685 ;
        RECT 40.955 166.885 42.080 167.055 ;
        RECT 42.250 166.945 42.635 167.515 ;
        RECT 41.630 166.775 42.080 166.885 ;
        RECT 40.365 166.155 41.460 166.715 ;
        RECT 41.630 166.445 42.185 166.775 ;
        RECT 39.240 165.305 39.525 165.765 ;
        RECT 39.695 165.135 39.965 165.595 ;
        RECT 40.365 165.305 40.765 166.155 ;
        RECT 41.630 165.985 42.080 166.445 ;
        RECT 42.355 166.275 42.635 166.945 ;
        RECT 40.955 165.765 42.080 165.985 ;
        RECT 40.955 165.305 41.235 165.765 ;
        RECT 41.755 165.135 42.080 165.595 ;
        RECT 42.250 165.305 42.635 166.275 ;
        RECT 42.805 166.945 43.190 167.515 ;
        RECT 43.360 167.225 43.685 167.685 ;
        RECT 44.205 167.055 44.485 167.515 ;
        RECT 42.805 166.275 43.085 166.945 ;
        RECT 43.360 166.885 44.485 167.055 ;
        RECT 43.360 166.775 43.810 166.885 ;
        RECT 43.255 166.445 43.810 166.775 ;
        RECT 44.675 166.715 45.075 167.515 ;
        RECT 45.475 167.225 45.745 167.685 ;
        RECT 45.915 167.055 46.200 167.515 ;
        RECT 42.805 165.305 43.190 166.275 ;
        RECT 43.360 165.985 43.810 166.445 ;
        RECT 43.980 166.155 45.075 166.715 ;
        RECT 43.360 165.765 44.485 165.985 ;
        RECT 43.360 165.135 43.685 165.595 ;
        RECT 44.205 165.305 44.485 165.765 ;
        RECT 44.675 165.305 45.075 166.155 ;
        RECT 45.245 166.885 46.200 167.055 ;
        RECT 47.410 166.975 47.665 167.505 ;
        RECT 47.835 167.225 48.140 167.685 ;
        RECT 48.385 167.305 49.455 167.475 ;
        RECT 45.245 165.985 45.455 166.885 ;
        RECT 45.625 166.155 46.315 166.715 ;
        RECT 47.410 166.325 47.620 166.975 ;
        RECT 48.385 166.950 48.705 167.305 ;
        RECT 48.380 166.775 48.705 166.950 ;
        RECT 47.790 166.475 48.705 166.775 ;
        RECT 48.875 166.735 49.115 167.135 ;
        RECT 49.285 167.075 49.455 167.305 ;
        RECT 49.625 167.245 49.815 167.685 ;
        RECT 49.985 167.235 50.935 167.515 ;
        RECT 51.155 167.325 51.505 167.495 ;
        RECT 49.285 166.905 49.815 167.075 ;
        RECT 47.790 166.445 48.530 166.475 ;
        RECT 45.245 165.765 46.200 165.985 ;
        RECT 45.475 165.135 45.745 165.595 ;
        RECT 45.915 165.305 46.200 165.765 ;
        RECT 47.410 165.445 47.665 166.325 ;
        RECT 47.835 165.135 48.140 166.275 ;
        RECT 48.360 165.855 48.530 166.445 ;
        RECT 48.875 166.365 49.415 166.735 ;
        RECT 49.595 166.625 49.815 166.905 ;
        RECT 49.985 166.455 50.155 167.235 ;
        RECT 49.750 166.285 50.155 166.455 ;
        RECT 50.325 166.445 50.675 167.065 ;
        RECT 49.750 166.195 49.920 166.285 ;
        RECT 50.845 166.275 51.055 167.065 ;
        RECT 48.700 166.025 49.920 166.195 ;
        RECT 50.380 166.115 51.055 166.275 ;
        RECT 48.360 165.685 49.160 165.855 ;
        RECT 48.480 165.135 48.810 165.515 ;
        RECT 48.990 165.395 49.160 165.685 ;
        RECT 49.750 165.645 49.920 166.025 ;
        RECT 50.090 166.105 51.055 166.115 ;
        RECT 51.245 166.935 51.505 167.325 ;
        RECT 51.715 167.225 52.045 167.685 ;
        RECT 52.920 167.295 53.775 167.465 ;
        RECT 53.980 167.295 54.475 167.465 ;
        RECT 54.645 167.325 54.975 167.685 ;
        RECT 51.245 166.245 51.415 166.935 ;
        RECT 51.585 166.585 51.755 166.765 ;
        RECT 51.925 166.755 52.715 167.005 ;
        RECT 52.920 166.585 53.090 167.295 ;
        RECT 53.260 166.785 53.615 167.005 ;
        RECT 51.585 166.415 53.275 166.585 ;
        RECT 50.090 165.815 50.550 166.105 ;
        RECT 51.245 166.075 52.745 166.245 ;
        RECT 51.245 165.935 51.415 166.075 ;
        RECT 50.855 165.765 51.415 165.935 ;
        RECT 49.330 165.135 49.580 165.595 ;
        RECT 49.750 165.305 50.620 165.645 ;
        RECT 50.855 165.305 51.025 165.765 ;
        RECT 51.860 165.735 52.935 165.905 ;
        RECT 51.195 165.135 51.565 165.595 ;
        RECT 51.860 165.395 52.030 165.735 ;
        RECT 52.200 165.135 52.530 165.565 ;
        RECT 52.765 165.395 52.935 165.735 ;
        RECT 53.105 165.635 53.275 166.415 ;
        RECT 53.445 166.195 53.615 166.785 ;
        RECT 53.785 166.385 54.135 167.005 ;
        RECT 53.445 165.805 53.910 166.195 ;
        RECT 54.305 165.935 54.475 167.295 ;
        RECT 54.645 166.105 55.105 167.155 ;
        RECT 54.080 165.765 54.475 165.935 ;
        RECT 54.080 165.635 54.250 165.765 ;
        RECT 53.105 165.305 53.785 165.635 ;
        RECT 54.000 165.305 54.250 165.635 ;
        RECT 54.420 165.135 54.670 165.595 ;
        RECT 54.840 165.320 55.165 166.105 ;
        RECT 55.335 165.305 55.505 167.425 ;
        RECT 55.675 167.305 56.005 167.685 ;
        RECT 56.175 167.135 56.430 167.425 ;
        RECT 55.680 166.965 56.430 167.135 ;
        RECT 55.680 165.975 55.910 166.965 ;
        RECT 56.605 166.915 58.275 167.685 ;
        RECT 56.080 166.145 56.430 166.795 ;
        RECT 56.605 166.225 57.355 166.745 ;
        RECT 57.525 166.395 58.275 166.915 ;
        RECT 58.505 166.865 58.715 167.685 ;
        RECT 58.885 166.885 59.215 167.515 ;
        RECT 58.885 166.285 59.135 166.885 ;
        RECT 59.385 166.865 59.615 167.685 ;
        RECT 60.435 166.885 60.765 167.685 ;
        RECT 60.935 167.035 61.105 167.515 ;
        RECT 61.275 167.205 61.605 167.685 ;
        RECT 61.775 167.035 61.945 167.515 ;
        RECT 62.195 167.205 62.435 167.685 ;
        RECT 62.615 167.035 62.785 167.515 ;
        RECT 60.935 166.865 61.945 167.035 ;
        RECT 62.150 166.865 62.785 167.035 ;
        RECT 63.045 166.960 63.335 167.685 ;
        RECT 63.505 166.915 65.175 167.685 ;
        RECT 65.405 167.205 65.685 167.685 ;
        RECT 65.855 167.035 66.115 167.425 ;
        RECT 66.290 167.205 66.545 167.685 ;
        RECT 66.715 167.035 67.010 167.425 ;
        RECT 67.190 167.205 67.465 167.685 ;
        RECT 67.635 167.185 67.935 167.515 ;
        RECT 59.305 166.445 59.635 166.695 ;
        RECT 60.935 166.665 61.430 166.865 ;
        RECT 62.150 166.695 62.320 166.865 ;
        RECT 60.935 166.495 61.435 166.665 ;
        RECT 61.820 166.525 62.320 166.695 ;
        RECT 60.935 166.325 61.430 166.495 ;
        RECT 55.680 165.805 56.430 165.975 ;
        RECT 55.675 165.135 56.005 165.635 ;
        RECT 56.175 165.305 56.430 165.805 ;
        RECT 56.605 165.135 58.275 166.225 ;
        RECT 58.505 165.135 58.715 166.275 ;
        RECT 58.885 165.305 59.215 166.285 ;
        RECT 59.385 165.135 59.615 166.275 ;
        RECT 60.435 165.135 60.765 166.285 ;
        RECT 60.935 166.155 61.945 166.325 ;
        RECT 60.935 165.305 61.105 166.155 ;
        RECT 61.275 165.135 61.605 165.935 ;
        RECT 61.775 165.305 61.945 166.155 ;
        RECT 62.150 166.285 62.320 166.525 ;
        RECT 62.490 166.455 62.870 166.695 ;
        RECT 62.150 166.115 62.865 166.285 ;
        RECT 62.125 165.135 62.365 165.935 ;
        RECT 62.535 165.305 62.865 166.115 ;
        RECT 63.045 165.135 63.335 166.300 ;
        RECT 63.505 166.225 64.255 166.745 ;
        RECT 64.425 166.395 65.175 166.915 ;
        RECT 65.360 166.865 67.010 167.035 ;
        RECT 65.360 166.355 65.765 166.865 ;
        RECT 65.935 166.525 67.075 166.695 ;
        RECT 63.505 165.135 65.175 166.225 ;
        RECT 65.360 166.185 66.115 166.355 ;
        RECT 65.400 165.135 65.685 166.005 ;
        RECT 65.855 165.935 66.115 166.185 ;
        RECT 66.905 166.275 67.075 166.525 ;
        RECT 67.245 166.445 67.595 167.015 ;
        RECT 67.765 166.275 67.935 167.185 ;
        RECT 66.905 166.105 67.935 166.275 ;
        RECT 65.855 165.765 66.975 165.935 ;
        RECT 65.855 165.305 66.115 165.765 ;
        RECT 66.290 165.135 66.545 165.595 ;
        RECT 66.715 165.305 66.975 165.765 ;
        RECT 67.145 165.135 67.455 165.935 ;
        RECT 67.625 165.305 67.935 166.105 ;
        RECT 68.105 167.185 68.405 167.515 ;
        RECT 68.575 167.205 68.850 167.685 ;
        RECT 68.105 166.275 68.275 167.185 ;
        RECT 69.030 167.035 69.325 167.425 ;
        RECT 69.495 167.205 69.750 167.685 ;
        RECT 69.925 167.035 70.185 167.425 ;
        RECT 70.355 167.205 70.635 167.685 ;
        RECT 70.875 167.155 71.205 167.515 ;
        RECT 71.375 167.325 71.705 167.685 ;
        RECT 71.905 167.155 72.235 167.515 ;
        RECT 68.445 166.445 68.795 167.015 ;
        RECT 69.030 166.865 70.680 167.035 ;
        RECT 70.875 166.945 72.235 167.155 ;
        RECT 72.745 166.925 73.455 167.515 ;
        RECT 68.965 166.525 70.105 166.695 ;
        RECT 68.965 166.275 69.135 166.525 ;
        RECT 70.275 166.355 70.680 166.865 ;
        RECT 73.225 166.835 73.455 166.925 ;
        RECT 73.625 166.915 75.295 167.685 ;
        RECT 70.865 166.445 71.175 166.775 ;
        RECT 71.385 166.445 71.760 166.775 ;
        RECT 72.080 166.445 72.575 166.775 ;
        RECT 68.105 166.105 69.135 166.275 ;
        RECT 69.925 166.185 70.680 166.355 ;
        RECT 68.105 165.305 68.415 166.105 ;
        RECT 69.925 165.935 70.185 166.185 ;
        RECT 68.585 165.135 68.895 165.935 ;
        RECT 69.065 165.765 70.185 165.935 ;
        RECT 69.065 165.305 69.325 165.765 ;
        RECT 69.495 165.135 69.750 165.595 ;
        RECT 69.925 165.305 70.185 165.765 ;
        RECT 70.355 165.135 70.640 166.005 ;
        RECT 70.875 165.135 71.205 166.195 ;
        RECT 71.385 165.520 71.555 166.445 ;
        RECT 71.725 165.955 72.055 166.175 ;
        RECT 72.250 166.155 72.575 166.445 ;
        RECT 72.750 166.155 73.080 166.695 ;
        RECT 73.250 165.955 73.455 166.835 ;
        RECT 71.725 165.725 73.455 165.955 ;
        RECT 71.725 165.325 72.055 165.725 ;
        RECT 72.225 165.135 72.555 165.495 ;
        RECT 72.755 165.305 73.455 165.725 ;
        RECT 73.625 166.225 74.375 166.745 ;
        RECT 74.545 166.395 75.295 166.915 ;
        RECT 75.840 166.975 76.095 167.505 ;
        RECT 76.275 167.225 76.560 167.685 ;
        RECT 73.625 165.135 75.295 166.225 ;
        RECT 75.840 166.115 76.020 166.975 ;
        RECT 76.740 166.775 76.990 167.425 ;
        RECT 76.190 166.445 76.990 166.775 ;
        RECT 75.840 165.645 76.095 166.115 ;
        RECT 75.755 165.475 76.095 165.645 ;
        RECT 75.840 165.445 76.095 165.475 ;
        RECT 76.275 165.135 76.560 165.935 ;
        RECT 76.740 165.855 76.990 166.445 ;
        RECT 77.190 167.090 77.510 167.420 ;
        RECT 77.690 167.205 78.350 167.685 ;
        RECT 78.550 167.295 79.400 167.465 ;
        RECT 77.190 166.195 77.380 167.090 ;
        RECT 77.700 166.765 78.360 167.035 ;
        RECT 78.030 166.705 78.360 166.765 ;
        RECT 77.550 166.535 77.880 166.595 ;
        RECT 78.550 166.535 78.720 167.295 ;
        RECT 79.960 167.225 80.280 167.685 ;
        RECT 80.480 167.045 80.730 167.475 ;
        RECT 81.020 167.245 81.430 167.685 ;
        RECT 81.600 167.305 82.615 167.505 ;
        RECT 78.890 166.875 80.140 167.045 ;
        RECT 78.890 166.755 79.220 166.875 ;
        RECT 77.550 166.365 79.450 166.535 ;
        RECT 77.190 166.025 79.110 166.195 ;
        RECT 77.190 166.005 77.510 166.025 ;
        RECT 76.740 165.345 77.070 165.855 ;
        RECT 77.340 165.395 77.510 166.005 ;
        RECT 79.280 165.855 79.450 166.365 ;
        RECT 79.620 166.295 79.800 166.705 ;
        RECT 79.970 166.115 80.140 166.875 ;
        RECT 77.680 165.135 78.010 165.825 ;
        RECT 78.240 165.685 79.450 165.855 ;
        RECT 79.620 165.805 80.140 166.115 ;
        RECT 80.310 166.705 80.730 167.045 ;
        RECT 81.020 166.705 81.430 167.035 ;
        RECT 80.310 165.935 80.500 166.705 ;
        RECT 81.600 166.575 81.770 167.305 ;
        RECT 82.915 167.135 83.085 167.465 ;
        RECT 83.255 167.305 83.585 167.685 ;
        RECT 81.940 166.755 82.290 167.125 ;
        RECT 81.600 166.535 82.020 166.575 ;
        RECT 80.670 166.365 82.020 166.535 ;
        RECT 80.670 166.205 80.920 166.365 ;
        RECT 81.430 165.935 81.680 166.195 ;
        RECT 80.310 165.685 81.680 165.935 ;
        RECT 78.240 165.395 78.480 165.685 ;
        RECT 79.280 165.605 79.450 165.685 ;
        RECT 78.680 165.135 79.100 165.515 ;
        RECT 79.280 165.355 79.910 165.605 ;
        RECT 80.380 165.135 80.710 165.515 ;
        RECT 80.880 165.395 81.050 165.685 ;
        RECT 81.850 165.520 82.020 166.365 ;
        RECT 82.470 166.195 82.690 167.065 ;
        RECT 82.915 166.945 83.610 167.135 ;
        RECT 82.190 165.815 82.690 166.195 ;
        RECT 82.860 166.145 83.270 166.765 ;
        RECT 83.440 165.975 83.610 166.945 ;
        RECT 82.915 165.805 83.610 165.975 ;
        RECT 81.230 165.135 81.610 165.515 ;
        RECT 81.850 165.350 82.680 165.520 ;
        RECT 82.915 165.305 83.085 165.805 ;
        RECT 83.255 165.135 83.585 165.635 ;
        RECT 83.800 165.305 84.025 167.425 ;
        RECT 84.195 167.305 84.525 167.685 ;
        RECT 84.695 167.135 84.865 167.425 ;
        RECT 84.200 166.965 84.865 167.135 ;
        RECT 84.200 165.975 84.430 166.965 ;
        RECT 85.185 166.865 85.395 167.685 ;
        RECT 85.565 166.885 85.895 167.515 ;
        RECT 84.600 166.145 84.950 166.795 ;
        RECT 85.565 166.285 85.815 166.885 ;
        RECT 86.065 166.865 86.295 167.685 ;
        RECT 86.565 166.865 86.775 167.685 ;
        RECT 86.945 166.885 87.275 167.515 ;
        RECT 85.985 166.445 86.315 166.695 ;
        RECT 86.945 166.285 87.195 166.885 ;
        RECT 87.445 166.865 87.675 167.685 ;
        RECT 88.805 166.960 89.095 167.685 ;
        RECT 89.725 166.915 93.235 167.685 ;
        RECT 87.365 166.445 87.695 166.695 ;
        RECT 84.200 165.805 84.865 165.975 ;
        RECT 84.195 165.135 84.525 165.635 ;
        RECT 84.695 165.305 84.865 165.805 ;
        RECT 85.185 165.135 85.395 166.275 ;
        RECT 85.565 165.305 85.895 166.285 ;
        RECT 86.065 165.135 86.295 166.275 ;
        RECT 86.565 165.135 86.775 166.275 ;
        RECT 86.945 165.305 87.275 166.285 ;
        RECT 87.445 165.135 87.675 166.275 ;
        RECT 88.805 165.135 89.095 166.300 ;
        RECT 89.725 166.225 91.415 166.745 ;
        RECT 91.585 166.395 93.235 166.915 ;
        RECT 93.680 166.875 93.925 167.480 ;
        RECT 94.145 167.150 94.655 167.685 ;
        RECT 93.405 166.705 94.635 166.875 ;
        RECT 89.725 165.135 93.235 166.225 ;
        RECT 93.405 165.895 93.745 166.705 ;
        RECT 93.915 166.140 94.665 166.330 ;
        RECT 93.405 165.485 93.920 165.895 ;
        RECT 94.155 165.135 94.325 165.895 ;
        RECT 94.495 165.475 94.665 166.140 ;
        RECT 94.835 166.155 95.025 167.515 ;
        RECT 95.195 166.665 95.470 167.515 ;
        RECT 95.660 167.150 96.190 167.515 ;
        RECT 96.615 167.285 96.945 167.685 ;
        RECT 96.015 167.115 96.190 167.150 ;
        RECT 95.195 166.495 95.475 166.665 ;
        RECT 95.195 166.355 95.470 166.495 ;
        RECT 95.675 166.155 95.845 166.955 ;
        RECT 94.835 165.985 95.845 166.155 ;
        RECT 96.015 166.945 96.945 167.115 ;
        RECT 97.115 166.945 97.370 167.515 ;
        RECT 96.015 165.815 96.185 166.945 ;
        RECT 96.775 166.775 96.945 166.945 ;
        RECT 95.060 165.645 96.185 165.815 ;
        RECT 96.355 166.445 96.550 166.775 ;
        RECT 96.775 166.445 97.030 166.775 ;
        RECT 96.355 165.475 96.525 166.445 ;
        RECT 97.200 166.275 97.370 166.945 ;
        RECT 97.920 166.975 98.175 167.505 ;
        RECT 98.355 167.225 98.640 167.685 ;
        RECT 97.920 166.325 98.100 166.975 ;
        RECT 98.820 166.775 99.070 167.425 ;
        RECT 98.270 166.445 99.070 166.775 ;
        RECT 94.495 165.305 96.525 165.475 ;
        RECT 96.695 165.135 96.865 166.275 ;
        RECT 97.035 165.305 97.370 166.275 ;
        RECT 97.835 166.155 98.100 166.325 ;
        RECT 97.920 166.115 98.100 166.155 ;
        RECT 97.920 165.445 98.175 166.115 ;
        RECT 98.355 165.135 98.640 165.935 ;
        RECT 98.820 165.855 99.070 166.445 ;
        RECT 99.270 167.090 99.590 167.420 ;
        RECT 99.770 167.205 100.430 167.685 ;
        RECT 100.630 167.295 101.480 167.465 ;
        RECT 99.270 166.195 99.460 167.090 ;
        RECT 99.780 166.765 100.440 167.035 ;
        RECT 100.110 166.705 100.440 166.765 ;
        RECT 99.630 166.535 99.960 166.595 ;
        RECT 100.630 166.535 100.800 167.295 ;
        RECT 102.040 167.225 102.360 167.685 ;
        RECT 102.560 167.045 102.810 167.475 ;
        RECT 103.100 167.245 103.510 167.685 ;
        RECT 103.680 167.305 104.695 167.505 ;
        RECT 100.970 166.875 102.220 167.045 ;
        RECT 100.970 166.755 101.300 166.875 ;
        RECT 99.630 166.365 101.530 166.535 ;
        RECT 99.270 166.025 101.190 166.195 ;
        RECT 99.270 166.005 99.590 166.025 ;
        RECT 98.820 165.345 99.150 165.855 ;
        RECT 99.420 165.395 99.590 166.005 ;
        RECT 101.360 165.855 101.530 166.365 ;
        RECT 101.700 166.295 101.880 166.705 ;
        RECT 102.050 166.115 102.220 166.875 ;
        RECT 99.760 165.135 100.090 165.825 ;
        RECT 100.320 165.685 101.530 165.855 ;
        RECT 101.700 165.805 102.220 166.115 ;
        RECT 102.390 166.705 102.810 167.045 ;
        RECT 103.100 166.705 103.510 167.035 ;
        RECT 102.390 165.935 102.580 166.705 ;
        RECT 103.680 166.575 103.850 167.305 ;
        RECT 104.995 167.135 105.165 167.465 ;
        RECT 105.335 167.305 105.665 167.685 ;
        RECT 104.020 166.755 104.370 167.125 ;
        RECT 103.680 166.535 104.100 166.575 ;
        RECT 102.750 166.365 104.100 166.535 ;
        RECT 102.750 166.205 103.000 166.365 ;
        RECT 103.510 165.935 103.760 166.195 ;
        RECT 102.390 165.685 103.760 165.935 ;
        RECT 100.320 165.395 100.560 165.685 ;
        RECT 101.360 165.605 101.530 165.685 ;
        RECT 100.760 165.135 101.180 165.515 ;
        RECT 101.360 165.355 101.990 165.605 ;
        RECT 102.460 165.135 102.790 165.515 ;
        RECT 102.960 165.395 103.130 165.685 ;
        RECT 103.930 165.520 104.100 166.365 ;
        RECT 104.550 166.195 104.770 167.065 ;
        RECT 104.995 166.945 105.690 167.135 ;
        RECT 104.270 165.815 104.770 166.195 ;
        RECT 104.940 166.145 105.350 166.765 ;
        RECT 105.520 165.975 105.690 166.945 ;
        RECT 104.995 165.805 105.690 165.975 ;
        RECT 103.310 165.135 103.690 165.515 ;
        RECT 103.930 165.350 104.760 165.520 ;
        RECT 104.995 165.305 105.165 165.805 ;
        RECT 105.335 165.135 105.665 165.635 ;
        RECT 105.880 165.305 106.105 167.425 ;
        RECT 106.275 167.305 106.605 167.685 ;
        RECT 106.775 167.135 106.945 167.425 ;
        RECT 106.280 166.965 106.945 167.135 ;
        RECT 107.320 167.055 107.605 167.515 ;
        RECT 107.775 167.225 108.045 167.685 ;
        RECT 106.280 165.975 106.510 166.965 ;
        RECT 107.320 166.885 108.275 167.055 ;
        RECT 106.680 166.145 107.030 166.795 ;
        RECT 107.205 166.155 107.895 166.715 ;
        RECT 108.065 165.985 108.275 166.885 ;
        RECT 106.280 165.805 106.945 165.975 ;
        RECT 106.275 165.135 106.605 165.635 ;
        RECT 106.775 165.305 106.945 165.805 ;
        RECT 107.320 165.765 108.275 165.985 ;
        RECT 108.445 166.715 108.845 167.515 ;
        RECT 109.035 167.055 109.315 167.515 ;
        RECT 109.835 167.225 110.160 167.685 ;
        RECT 109.035 166.885 110.160 167.055 ;
        RECT 110.330 166.945 110.715 167.515 ;
        RECT 109.710 166.775 110.160 166.885 ;
        RECT 108.445 166.155 109.540 166.715 ;
        RECT 109.710 166.445 110.265 166.775 ;
        RECT 107.320 165.305 107.605 165.765 ;
        RECT 107.775 165.135 108.045 165.595 ;
        RECT 108.445 165.305 108.845 166.155 ;
        RECT 109.710 165.985 110.160 166.445 ;
        RECT 110.435 166.275 110.715 166.945 ;
        RECT 111.000 167.055 111.285 167.515 ;
        RECT 111.455 167.225 111.725 167.685 ;
        RECT 111.000 166.885 111.955 167.055 ;
        RECT 109.035 165.765 110.160 165.985 ;
        RECT 109.035 165.305 109.315 165.765 ;
        RECT 109.835 165.135 110.160 165.595 ;
        RECT 110.330 165.305 110.715 166.275 ;
        RECT 110.885 166.155 111.575 166.715 ;
        RECT 111.745 165.985 111.955 166.885 ;
        RECT 111.000 165.765 111.955 165.985 ;
        RECT 112.125 166.715 112.525 167.515 ;
        RECT 112.715 167.055 112.995 167.515 ;
        RECT 113.515 167.225 113.840 167.685 ;
        RECT 112.715 166.885 113.840 167.055 ;
        RECT 114.010 166.945 114.395 167.515 ;
        RECT 114.565 166.960 114.855 167.685 ;
        RECT 115.950 166.975 116.205 167.505 ;
        RECT 116.375 167.225 116.680 167.685 ;
        RECT 116.925 167.305 117.995 167.475 ;
        RECT 113.390 166.775 113.840 166.885 ;
        RECT 112.125 166.155 113.220 166.715 ;
        RECT 113.390 166.445 113.945 166.775 ;
        RECT 111.000 165.305 111.285 165.765 ;
        RECT 111.455 165.135 111.725 165.595 ;
        RECT 112.125 165.305 112.525 166.155 ;
        RECT 113.390 165.985 113.840 166.445 ;
        RECT 114.115 166.275 114.395 166.945 ;
        RECT 115.950 166.325 116.160 166.975 ;
        RECT 116.925 166.950 117.245 167.305 ;
        RECT 116.920 166.775 117.245 166.950 ;
        RECT 116.330 166.475 117.245 166.775 ;
        RECT 117.415 166.735 117.655 167.135 ;
        RECT 117.825 167.075 117.995 167.305 ;
        RECT 118.165 167.245 118.355 167.685 ;
        RECT 118.525 167.235 119.475 167.515 ;
        RECT 119.695 167.325 120.045 167.495 ;
        RECT 117.825 166.905 118.355 167.075 ;
        RECT 116.330 166.445 117.070 166.475 ;
        RECT 112.715 165.765 113.840 165.985 ;
        RECT 112.715 165.305 112.995 165.765 ;
        RECT 113.515 165.135 113.840 165.595 ;
        RECT 114.010 165.305 114.395 166.275 ;
        RECT 114.565 165.135 114.855 166.300 ;
        RECT 115.950 165.445 116.205 166.325 ;
        RECT 116.375 165.135 116.680 166.275 ;
        RECT 116.900 165.855 117.070 166.445 ;
        RECT 117.415 166.365 117.955 166.735 ;
        RECT 118.135 166.625 118.355 166.905 ;
        RECT 118.525 166.455 118.695 167.235 ;
        RECT 118.290 166.285 118.695 166.455 ;
        RECT 118.865 166.445 119.215 167.065 ;
        RECT 118.290 166.195 118.460 166.285 ;
        RECT 119.385 166.275 119.595 167.065 ;
        RECT 117.240 166.025 118.460 166.195 ;
        RECT 118.920 166.115 119.595 166.275 ;
        RECT 116.900 165.685 117.700 165.855 ;
        RECT 117.020 165.135 117.350 165.515 ;
        RECT 117.530 165.395 117.700 165.685 ;
        RECT 118.290 165.645 118.460 166.025 ;
        RECT 118.630 166.105 119.595 166.115 ;
        RECT 119.785 166.935 120.045 167.325 ;
        RECT 120.255 167.225 120.585 167.685 ;
        RECT 121.460 167.295 122.315 167.465 ;
        RECT 122.520 167.295 123.015 167.465 ;
        RECT 123.185 167.325 123.515 167.685 ;
        RECT 119.785 166.245 119.955 166.935 ;
        RECT 120.125 166.585 120.295 166.765 ;
        RECT 120.465 166.755 121.255 167.005 ;
        RECT 121.460 166.585 121.630 167.295 ;
        RECT 121.800 166.785 122.155 167.005 ;
        RECT 120.125 166.415 121.815 166.585 ;
        RECT 118.630 165.815 119.090 166.105 ;
        RECT 119.785 166.075 121.285 166.245 ;
        RECT 119.785 165.935 119.955 166.075 ;
        RECT 119.395 165.765 119.955 165.935 ;
        RECT 117.870 165.135 118.120 165.595 ;
        RECT 118.290 165.305 119.160 165.645 ;
        RECT 119.395 165.305 119.565 165.765 ;
        RECT 120.400 165.735 121.475 165.905 ;
        RECT 119.735 165.135 120.105 165.595 ;
        RECT 120.400 165.395 120.570 165.735 ;
        RECT 120.740 165.135 121.070 165.565 ;
        RECT 121.305 165.395 121.475 165.735 ;
        RECT 121.645 165.635 121.815 166.415 ;
        RECT 121.985 166.195 122.155 166.785 ;
        RECT 122.325 166.385 122.675 167.005 ;
        RECT 121.985 165.805 122.450 166.195 ;
        RECT 122.845 165.935 123.015 167.295 ;
        RECT 123.185 166.105 123.645 167.155 ;
        RECT 122.620 165.765 123.015 165.935 ;
        RECT 122.620 165.635 122.790 165.765 ;
        RECT 121.645 165.305 122.325 165.635 ;
        RECT 122.540 165.305 122.790 165.635 ;
        RECT 122.960 165.135 123.210 165.595 ;
        RECT 123.380 165.320 123.705 166.105 ;
        RECT 123.875 165.305 124.045 167.425 ;
        RECT 124.215 167.305 124.545 167.685 ;
        RECT 124.715 167.135 124.970 167.425 ;
        RECT 124.220 166.965 124.970 167.135 ;
        RECT 124.220 165.975 124.450 166.965 ;
        RECT 125.145 166.935 126.355 167.685 ;
        RECT 126.525 166.935 127.735 167.685 ;
        RECT 124.620 166.145 124.970 166.795 ;
        RECT 125.145 166.225 125.665 166.765 ;
        RECT 125.835 166.395 126.355 166.935 ;
        RECT 126.525 166.225 127.045 166.765 ;
        RECT 127.215 166.395 127.735 166.935 ;
        RECT 124.220 165.805 124.970 165.975 ;
        RECT 124.215 165.135 124.545 165.635 ;
        RECT 124.715 165.305 124.970 165.805 ;
        RECT 125.145 165.135 126.355 166.225 ;
        RECT 126.525 165.135 127.735 166.225 ;
        RECT 14.660 164.965 127.820 165.135 ;
        RECT 14.745 163.875 15.955 164.965 ;
        RECT 14.745 163.165 15.265 163.705 ;
        RECT 15.435 163.335 15.955 163.875 ;
        RECT 16.125 163.875 18.715 164.965 ;
        RECT 18.890 164.530 24.235 164.965 ;
        RECT 16.125 163.355 17.335 163.875 ;
        RECT 17.505 163.185 18.715 163.705 ;
        RECT 20.480 163.280 20.830 164.530 ;
        RECT 24.405 163.800 24.695 164.965 ;
        RECT 25.785 163.890 26.055 164.795 ;
        RECT 26.225 164.205 26.555 164.965 ;
        RECT 26.735 164.035 26.905 164.795 ;
        RECT 27.170 164.295 27.425 164.795 ;
        RECT 27.595 164.465 27.925 164.965 ;
        RECT 27.170 164.125 27.920 164.295 ;
        RECT 14.745 162.415 15.955 163.165 ;
        RECT 16.125 162.415 18.715 163.185 ;
        RECT 22.310 162.960 22.650 163.790 ;
        RECT 18.890 162.415 24.235 162.960 ;
        RECT 24.405 162.415 24.695 163.140 ;
        RECT 25.785 163.090 25.955 163.890 ;
        RECT 26.240 163.865 26.905 164.035 ;
        RECT 26.240 163.720 26.410 163.865 ;
        RECT 26.125 163.390 26.410 163.720 ;
        RECT 26.240 163.135 26.410 163.390 ;
        RECT 26.645 163.315 26.975 163.685 ;
        RECT 27.170 163.305 27.520 163.955 ;
        RECT 27.690 163.135 27.920 164.125 ;
        RECT 25.785 162.585 26.045 163.090 ;
        RECT 26.240 162.965 26.905 163.135 ;
        RECT 26.225 162.415 26.555 162.795 ;
        RECT 26.735 162.585 26.905 162.965 ;
        RECT 27.170 162.965 27.920 163.135 ;
        RECT 27.170 162.675 27.425 162.965 ;
        RECT 27.595 162.415 27.925 162.795 ;
        RECT 28.095 162.675 28.265 164.795 ;
        RECT 28.435 163.995 28.760 164.780 ;
        RECT 28.930 164.505 29.180 164.965 ;
        RECT 29.350 164.465 29.600 164.795 ;
        RECT 29.815 164.465 30.495 164.795 ;
        RECT 29.350 164.335 29.520 164.465 ;
        RECT 29.125 164.165 29.520 164.335 ;
        RECT 28.495 162.945 28.955 163.995 ;
        RECT 29.125 162.805 29.295 164.165 ;
        RECT 29.690 163.905 30.155 164.295 ;
        RECT 29.465 163.095 29.815 163.715 ;
        RECT 29.985 163.315 30.155 163.905 ;
        RECT 30.325 163.685 30.495 164.465 ;
        RECT 30.665 164.365 30.835 164.705 ;
        RECT 31.070 164.535 31.400 164.965 ;
        RECT 31.570 164.365 31.740 164.705 ;
        RECT 32.035 164.505 32.405 164.965 ;
        RECT 30.665 164.195 31.740 164.365 ;
        RECT 32.575 164.335 32.745 164.795 ;
        RECT 32.980 164.455 33.850 164.795 ;
        RECT 34.020 164.505 34.270 164.965 ;
        RECT 32.185 164.165 32.745 164.335 ;
        RECT 32.185 164.025 32.355 164.165 ;
        RECT 30.855 163.855 32.355 164.025 ;
        RECT 33.050 163.995 33.510 164.285 ;
        RECT 30.325 163.515 32.015 163.685 ;
        RECT 29.985 163.095 30.340 163.315 ;
        RECT 30.510 162.805 30.680 163.515 ;
        RECT 30.885 163.095 31.675 163.345 ;
        RECT 31.845 163.335 32.015 163.515 ;
        RECT 32.185 163.165 32.355 163.855 ;
        RECT 28.625 162.415 28.955 162.775 ;
        RECT 29.125 162.635 29.620 162.805 ;
        RECT 29.825 162.635 30.680 162.805 ;
        RECT 31.555 162.415 31.885 162.875 ;
        RECT 32.095 162.775 32.355 163.165 ;
        RECT 32.545 163.985 33.510 163.995 ;
        RECT 33.680 164.075 33.850 164.455 ;
        RECT 34.440 164.415 34.610 164.705 ;
        RECT 34.790 164.585 35.120 164.965 ;
        RECT 34.440 164.245 35.240 164.415 ;
        RECT 32.545 163.825 33.220 163.985 ;
        RECT 33.680 163.905 34.900 164.075 ;
        RECT 32.545 163.035 32.755 163.825 ;
        RECT 33.680 163.815 33.850 163.905 ;
        RECT 32.925 163.035 33.275 163.655 ;
        RECT 33.445 163.645 33.850 163.815 ;
        RECT 33.445 162.865 33.615 163.645 ;
        RECT 33.785 163.195 34.005 163.475 ;
        RECT 34.185 163.365 34.725 163.735 ;
        RECT 35.070 163.655 35.240 164.245 ;
        RECT 35.460 163.825 35.765 164.965 ;
        RECT 35.935 163.775 36.190 164.655 ;
        RECT 35.070 163.625 35.810 163.655 ;
        RECT 33.785 163.025 34.315 163.195 ;
        RECT 32.095 162.605 32.445 162.775 ;
        RECT 32.665 162.585 33.615 162.865 ;
        RECT 33.785 162.415 33.975 162.855 ;
        RECT 34.145 162.795 34.315 163.025 ;
        RECT 34.485 162.965 34.725 163.365 ;
        RECT 34.895 163.325 35.810 163.625 ;
        RECT 34.895 163.150 35.220 163.325 ;
        RECT 34.895 162.795 35.215 163.150 ;
        RECT 35.980 163.125 36.190 163.775 ;
        RECT 34.145 162.625 35.215 162.795 ;
        RECT 35.460 162.415 35.765 162.875 ;
        RECT 35.935 162.595 36.190 163.125 ;
        RECT 36.370 163.775 36.625 164.655 ;
        RECT 36.795 163.825 37.100 164.965 ;
        RECT 37.440 164.585 37.770 164.965 ;
        RECT 37.950 164.415 38.120 164.705 ;
        RECT 38.290 164.505 38.540 164.965 ;
        RECT 37.320 164.245 38.120 164.415 ;
        RECT 38.710 164.455 39.580 164.795 ;
        RECT 36.370 163.125 36.580 163.775 ;
        RECT 37.320 163.655 37.490 164.245 ;
        RECT 38.710 164.075 38.880 164.455 ;
        RECT 39.815 164.335 39.985 164.795 ;
        RECT 40.155 164.505 40.525 164.965 ;
        RECT 40.820 164.365 40.990 164.705 ;
        RECT 41.160 164.535 41.490 164.965 ;
        RECT 41.725 164.365 41.895 164.705 ;
        RECT 37.660 163.905 38.880 164.075 ;
        RECT 39.050 163.995 39.510 164.285 ;
        RECT 39.815 164.165 40.375 164.335 ;
        RECT 40.820 164.195 41.895 164.365 ;
        RECT 42.065 164.465 42.745 164.795 ;
        RECT 42.960 164.465 43.210 164.795 ;
        RECT 43.380 164.505 43.630 164.965 ;
        RECT 40.205 164.025 40.375 164.165 ;
        RECT 39.050 163.985 40.015 163.995 ;
        RECT 38.710 163.815 38.880 163.905 ;
        RECT 39.340 163.825 40.015 163.985 ;
        RECT 36.750 163.625 37.490 163.655 ;
        RECT 36.750 163.325 37.665 163.625 ;
        RECT 37.340 163.150 37.665 163.325 ;
        RECT 36.370 162.595 36.625 163.125 ;
        RECT 36.795 162.415 37.100 162.875 ;
        RECT 37.345 162.795 37.665 163.150 ;
        RECT 37.835 163.365 38.375 163.735 ;
        RECT 38.710 163.645 39.115 163.815 ;
        RECT 37.835 162.965 38.075 163.365 ;
        RECT 38.555 163.195 38.775 163.475 ;
        RECT 38.245 163.025 38.775 163.195 ;
        RECT 38.245 162.795 38.415 163.025 ;
        RECT 38.945 162.865 39.115 163.645 ;
        RECT 39.285 163.035 39.635 163.655 ;
        RECT 39.805 163.035 40.015 163.825 ;
        RECT 40.205 163.855 41.705 164.025 ;
        RECT 40.205 163.165 40.375 163.855 ;
        RECT 42.065 163.685 42.235 164.465 ;
        RECT 43.040 164.335 43.210 164.465 ;
        RECT 40.545 163.515 42.235 163.685 ;
        RECT 42.405 163.905 42.870 164.295 ;
        RECT 43.040 164.165 43.435 164.335 ;
        RECT 40.545 163.335 40.715 163.515 ;
        RECT 37.345 162.625 38.415 162.795 ;
        RECT 38.585 162.415 38.775 162.855 ;
        RECT 38.945 162.585 39.895 162.865 ;
        RECT 40.205 162.775 40.465 163.165 ;
        RECT 40.885 163.095 41.675 163.345 ;
        RECT 40.115 162.605 40.465 162.775 ;
        RECT 40.675 162.415 41.005 162.875 ;
        RECT 41.880 162.805 42.050 163.515 ;
        RECT 42.405 163.315 42.575 163.905 ;
        RECT 42.220 163.095 42.575 163.315 ;
        RECT 42.745 163.095 43.095 163.715 ;
        RECT 43.265 162.805 43.435 164.165 ;
        RECT 43.800 163.995 44.125 164.780 ;
        RECT 43.605 162.945 44.065 163.995 ;
        RECT 41.880 162.635 42.735 162.805 ;
        RECT 42.940 162.635 43.435 162.805 ;
        RECT 43.605 162.415 43.935 162.775 ;
        RECT 44.295 162.675 44.465 164.795 ;
        RECT 44.635 164.465 44.965 164.965 ;
        RECT 45.135 164.295 45.390 164.795 ;
        RECT 44.640 164.125 45.390 164.295 ;
        RECT 46.600 164.335 46.885 164.795 ;
        RECT 47.055 164.505 47.325 164.965 ;
        RECT 44.640 163.135 44.870 164.125 ;
        RECT 46.600 164.115 47.555 164.335 ;
        RECT 45.040 163.305 45.390 163.955 ;
        RECT 46.485 163.385 47.175 163.945 ;
        RECT 47.345 163.215 47.555 164.115 ;
        RECT 44.640 162.965 45.390 163.135 ;
        RECT 44.635 162.415 44.965 162.795 ;
        RECT 45.135 162.675 45.390 162.965 ;
        RECT 46.600 163.045 47.555 163.215 ;
        RECT 47.725 163.945 48.125 164.795 ;
        RECT 48.315 164.335 48.595 164.795 ;
        RECT 49.115 164.505 49.440 164.965 ;
        RECT 48.315 164.115 49.440 164.335 ;
        RECT 47.725 163.385 48.820 163.945 ;
        RECT 48.990 163.655 49.440 164.115 ;
        RECT 49.610 163.825 49.995 164.795 ;
        RECT 46.600 162.585 46.885 163.045 ;
        RECT 47.055 162.415 47.325 162.875 ;
        RECT 47.725 162.585 48.125 163.385 ;
        RECT 48.990 163.325 49.545 163.655 ;
        RECT 48.990 163.215 49.440 163.325 ;
        RECT 48.315 163.045 49.440 163.215 ;
        RECT 49.715 163.155 49.995 163.825 ;
        RECT 50.165 163.800 50.455 164.965 ;
        RECT 50.685 163.825 50.895 164.965 ;
        RECT 51.065 163.815 51.395 164.795 ;
        RECT 51.565 163.825 51.795 164.965 ;
        RECT 52.005 163.875 53.675 164.965 ;
        RECT 53.935 164.035 54.105 164.795 ;
        RECT 54.285 164.205 54.615 164.965 ;
        RECT 48.315 162.585 48.595 163.045 ;
        RECT 49.115 162.415 49.440 162.875 ;
        RECT 49.610 162.585 49.995 163.155 ;
        RECT 50.165 162.415 50.455 163.140 ;
        RECT 50.685 162.415 50.895 163.235 ;
        RECT 51.065 163.215 51.315 163.815 ;
        RECT 51.485 163.405 51.815 163.655 ;
        RECT 52.005 163.355 52.755 163.875 ;
        RECT 53.935 163.865 54.600 164.035 ;
        RECT 54.785 163.890 55.055 164.795 ;
        RECT 54.430 163.720 54.600 163.865 ;
        RECT 51.065 162.585 51.395 163.215 ;
        RECT 51.565 162.415 51.795 163.235 ;
        RECT 52.925 163.185 53.675 163.705 ;
        RECT 53.865 163.315 54.195 163.685 ;
        RECT 54.430 163.390 54.715 163.720 ;
        RECT 52.005 162.415 53.675 163.185 ;
        RECT 54.430 163.135 54.600 163.390 ;
        RECT 53.935 162.965 54.600 163.135 ;
        RECT 54.885 163.090 55.055 163.890 ;
        RECT 53.935 162.585 54.105 162.965 ;
        RECT 54.285 162.415 54.615 162.795 ;
        RECT 54.795 162.585 55.055 163.090 ;
        RECT 55.230 163.775 55.485 164.655 ;
        RECT 55.655 163.825 55.960 164.965 ;
        RECT 56.300 164.585 56.630 164.965 ;
        RECT 56.810 164.415 56.980 164.705 ;
        RECT 57.150 164.505 57.400 164.965 ;
        RECT 56.180 164.245 56.980 164.415 ;
        RECT 57.570 164.455 58.440 164.795 ;
        RECT 55.230 163.125 55.440 163.775 ;
        RECT 56.180 163.655 56.350 164.245 ;
        RECT 57.570 164.075 57.740 164.455 ;
        RECT 58.675 164.335 58.845 164.795 ;
        RECT 59.015 164.505 59.385 164.965 ;
        RECT 59.680 164.365 59.850 164.705 ;
        RECT 60.020 164.535 60.350 164.965 ;
        RECT 60.585 164.365 60.755 164.705 ;
        RECT 56.520 163.905 57.740 164.075 ;
        RECT 57.910 163.995 58.370 164.285 ;
        RECT 58.675 164.165 59.235 164.335 ;
        RECT 59.680 164.195 60.755 164.365 ;
        RECT 60.925 164.465 61.605 164.795 ;
        RECT 61.820 164.465 62.070 164.795 ;
        RECT 62.240 164.505 62.490 164.965 ;
        RECT 59.065 164.025 59.235 164.165 ;
        RECT 57.910 163.985 58.875 163.995 ;
        RECT 57.570 163.815 57.740 163.905 ;
        RECT 58.200 163.825 58.875 163.985 ;
        RECT 55.610 163.625 56.350 163.655 ;
        RECT 55.610 163.325 56.525 163.625 ;
        RECT 56.200 163.150 56.525 163.325 ;
        RECT 55.230 162.595 55.485 163.125 ;
        RECT 55.655 162.415 55.960 162.875 ;
        RECT 56.205 162.795 56.525 163.150 ;
        RECT 56.695 163.365 57.235 163.735 ;
        RECT 57.570 163.645 57.975 163.815 ;
        RECT 56.695 162.965 56.935 163.365 ;
        RECT 57.415 163.195 57.635 163.475 ;
        RECT 57.105 163.025 57.635 163.195 ;
        RECT 57.105 162.795 57.275 163.025 ;
        RECT 57.805 162.865 57.975 163.645 ;
        RECT 58.145 163.035 58.495 163.655 ;
        RECT 58.665 163.035 58.875 163.825 ;
        RECT 59.065 163.855 60.565 164.025 ;
        RECT 59.065 163.165 59.235 163.855 ;
        RECT 60.925 163.685 61.095 164.465 ;
        RECT 61.900 164.335 62.070 164.465 ;
        RECT 59.405 163.515 61.095 163.685 ;
        RECT 61.265 163.905 61.730 164.295 ;
        RECT 61.900 164.165 62.295 164.335 ;
        RECT 59.405 163.335 59.575 163.515 ;
        RECT 56.205 162.625 57.275 162.795 ;
        RECT 57.445 162.415 57.635 162.855 ;
        RECT 57.805 162.585 58.755 162.865 ;
        RECT 59.065 162.775 59.325 163.165 ;
        RECT 59.745 163.095 60.535 163.345 ;
        RECT 58.975 162.605 59.325 162.775 ;
        RECT 59.535 162.415 59.865 162.875 ;
        RECT 60.740 162.805 60.910 163.515 ;
        RECT 61.265 163.315 61.435 163.905 ;
        RECT 61.080 163.095 61.435 163.315 ;
        RECT 61.605 163.095 61.955 163.715 ;
        RECT 62.125 162.805 62.295 164.165 ;
        RECT 62.660 163.995 62.985 164.780 ;
        RECT 62.465 162.945 62.925 163.995 ;
        RECT 60.740 162.635 61.595 162.805 ;
        RECT 61.800 162.635 62.295 162.805 ;
        RECT 62.465 162.415 62.795 162.775 ;
        RECT 63.155 162.675 63.325 164.795 ;
        RECT 63.495 164.465 63.825 164.965 ;
        RECT 63.995 164.295 64.250 164.795 ;
        RECT 63.500 164.125 64.250 164.295 ;
        RECT 63.500 163.135 63.730 164.125 ;
        RECT 63.900 163.305 64.250 163.955 ;
        RECT 64.575 163.815 64.905 164.965 ;
        RECT 65.075 163.945 65.245 164.795 ;
        RECT 65.415 164.165 65.745 164.965 ;
        RECT 65.915 163.945 66.085 164.795 ;
        RECT 66.265 164.165 66.505 164.965 ;
        RECT 66.675 163.985 67.005 164.795 ;
        RECT 67.240 164.095 67.525 164.965 ;
        RECT 67.695 164.335 67.955 164.795 ;
        RECT 68.130 164.505 68.385 164.965 ;
        RECT 68.555 164.335 68.815 164.795 ;
        RECT 67.695 164.165 68.815 164.335 ;
        RECT 68.985 164.165 69.295 164.965 ;
        RECT 65.075 163.775 66.085 163.945 ;
        RECT 66.290 163.815 67.005 163.985 ;
        RECT 67.695 163.915 67.955 164.165 ;
        RECT 69.465 163.995 69.775 164.795 ;
        RECT 70.410 164.530 75.755 164.965 ;
        RECT 65.075 163.265 65.570 163.775 ;
        RECT 66.290 163.575 66.460 163.815 ;
        RECT 67.200 163.745 67.955 163.915 ;
        RECT 68.745 163.825 69.775 163.995 ;
        RECT 65.960 163.405 66.460 163.575 ;
        RECT 66.630 163.405 67.010 163.645 ;
        RECT 65.075 163.235 65.575 163.265 ;
        RECT 66.290 163.235 66.460 163.405 ;
        RECT 67.200 163.235 67.605 163.745 ;
        RECT 68.745 163.575 68.915 163.825 ;
        RECT 67.775 163.405 68.915 163.575 ;
        RECT 63.500 162.965 64.250 163.135 ;
        RECT 63.495 162.415 63.825 162.795 ;
        RECT 63.995 162.675 64.250 162.965 ;
        RECT 64.575 162.415 64.905 163.215 ;
        RECT 65.075 163.065 66.085 163.235 ;
        RECT 66.290 163.065 66.925 163.235 ;
        RECT 67.200 163.065 68.850 163.235 ;
        RECT 69.085 163.085 69.435 163.655 ;
        RECT 65.075 162.585 65.245 163.065 ;
        RECT 65.415 162.415 65.745 162.895 ;
        RECT 65.915 162.585 66.085 163.065 ;
        RECT 66.335 162.415 66.575 162.895 ;
        RECT 66.755 162.585 66.925 163.065 ;
        RECT 67.245 162.415 67.525 162.895 ;
        RECT 67.695 162.675 67.955 163.065 ;
        RECT 68.130 162.415 68.385 162.895 ;
        RECT 68.555 162.675 68.850 163.065 ;
        RECT 69.605 162.915 69.775 163.825 ;
        RECT 72.000 163.280 72.350 164.530 ;
        RECT 75.925 163.800 76.215 164.965 ;
        RECT 76.385 163.875 78.055 164.965 ;
        RECT 78.225 164.205 78.740 164.615 ;
        RECT 78.975 164.205 79.145 164.965 ;
        RECT 79.315 164.625 81.345 164.795 ;
        RECT 73.830 162.960 74.170 163.790 ;
        RECT 76.385 163.355 77.135 163.875 ;
        RECT 77.305 163.185 78.055 163.705 ;
        RECT 78.225 163.395 78.565 164.205 ;
        RECT 79.315 163.960 79.485 164.625 ;
        RECT 79.880 164.285 81.005 164.455 ;
        RECT 78.735 163.770 79.485 163.960 ;
        RECT 79.655 163.945 80.665 164.115 ;
        RECT 78.225 163.225 79.455 163.395 ;
        RECT 69.030 162.415 69.305 162.895 ;
        RECT 69.475 162.585 69.775 162.915 ;
        RECT 70.410 162.415 75.755 162.960 ;
        RECT 75.925 162.415 76.215 163.140 ;
        RECT 76.385 162.415 78.055 163.185 ;
        RECT 78.500 162.620 78.745 163.225 ;
        RECT 78.965 162.415 79.475 162.950 ;
        RECT 79.655 162.585 79.845 163.945 ;
        RECT 80.015 162.925 80.290 163.745 ;
        RECT 80.495 163.145 80.665 163.945 ;
        RECT 80.835 163.155 81.005 164.285 ;
        RECT 81.175 163.655 81.345 164.625 ;
        RECT 81.515 163.825 81.685 164.965 ;
        RECT 81.855 163.825 82.190 164.795 ;
        RECT 82.455 164.035 82.625 164.795 ;
        RECT 82.805 164.205 83.135 164.965 ;
        RECT 82.455 163.865 83.120 164.035 ;
        RECT 83.305 163.890 83.575 164.795 ;
        RECT 81.175 163.325 81.370 163.655 ;
        RECT 81.595 163.325 81.850 163.655 ;
        RECT 81.595 163.155 81.765 163.325 ;
        RECT 82.020 163.155 82.190 163.825 ;
        RECT 82.950 163.720 83.120 163.865 ;
        RECT 82.385 163.315 82.715 163.685 ;
        RECT 82.950 163.390 83.235 163.720 ;
        RECT 80.835 162.985 81.765 163.155 ;
        RECT 80.835 162.950 81.010 162.985 ;
        RECT 80.015 162.755 80.295 162.925 ;
        RECT 80.015 162.585 80.290 162.755 ;
        RECT 80.480 162.585 81.010 162.950 ;
        RECT 81.435 162.415 81.765 162.815 ;
        RECT 81.935 162.585 82.190 163.155 ;
        RECT 82.950 163.135 83.120 163.390 ;
        RECT 82.455 162.965 83.120 163.135 ;
        RECT 83.405 163.090 83.575 163.890 ;
        RECT 83.745 163.875 85.415 164.965 ;
        RECT 85.675 164.035 85.845 164.795 ;
        RECT 86.025 164.205 86.355 164.965 ;
        RECT 83.745 163.355 84.495 163.875 ;
        RECT 85.675 163.865 86.340 164.035 ;
        RECT 86.525 163.890 86.795 164.795 ;
        RECT 86.970 164.530 92.315 164.965 ;
        RECT 86.170 163.720 86.340 163.865 ;
        RECT 84.665 163.185 85.415 163.705 ;
        RECT 85.605 163.315 85.935 163.685 ;
        RECT 86.170 163.390 86.455 163.720 ;
        RECT 82.455 162.585 82.625 162.965 ;
        RECT 82.805 162.415 83.135 162.795 ;
        RECT 83.315 162.585 83.575 163.090 ;
        RECT 83.745 162.415 85.415 163.185 ;
        RECT 86.170 163.135 86.340 163.390 ;
        RECT 85.675 162.965 86.340 163.135 ;
        RECT 86.625 163.090 86.795 163.890 ;
        RECT 88.560 163.280 88.910 164.530 ;
        RECT 92.575 164.220 92.845 164.965 ;
        RECT 93.475 164.960 99.750 164.965 ;
        RECT 93.015 164.050 93.305 164.790 ;
        RECT 93.475 164.235 93.730 164.960 ;
        RECT 93.915 164.065 94.175 164.790 ;
        RECT 94.345 164.235 94.590 164.960 ;
        RECT 94.775 164.065 95.035 164.790 ;
        RECT 95.205 164.235 95.450 164.960 ;
        RECT 95.635 164.065 95.895 164.790 ;
        RECT 96.065 164.235 96.310 164.960 ;
        RECT 96.480 164.065 96.740 164.790 ;
        RECT 96.910 164.235 97.170 164.960 ;
        RECT 97.340 164.065 97.600 164.790 ;
        RECT 97.770 164.235 98.030 164.960 ;
        RECT 98.200 164.065 98.460 164.790 ;
        RECT 98.630 164.235 98.890 164.960 ;
        RECT 99.060 164.065 99.320 164.790 ;
        RECT 99.490 164.165 99.750 164.960 ;
        RECT 93.915 164.050 99.320 164.065 ;
        RECT 92.575 163.825 99.320 164.050 ;
        RECT 85.675 162.585 85.845 162.965 ;
        RECT 86.025 162.415 86.355 162.795 ;
        RECT 86.535 162.585 86.795 163.090 ;
        RECT 90.390 162.960 90.730 163.790 ;
        RECT 92.575 163.235 93.740 163.825 ;
        RECT 99.920 163.655 100.170 164.790 ;
        RECT 100.350 164.155 100.610 164.965 ;
        RECT 100.785 163.655 101.030 164.795 ;
        RECT 101.210 164.155 101.505 164.965 ;
        RECT 101.685 163.800 101.975 164.965 ;
        RECT 102.145 164.205 102.660 164.615 ;
        RECT 102.895 164.205 103.065 164.965 ;
        RECT 103.235 164.625 105.265 164.795 ;
        RECT 93.910 163.405 101.030 163.655 ;
        RECT 92.575 163.065 99.320 163.235 ;
        RECT 86.970 162.415 92.315 162.960 ;
        RECT 92.575 162.415 92.875 162.895 ;
        RECT 93.045 162.610 93.305 163.065 ;
        RECT 93.475 162.415 93.735 162.895 ;
        RECT 93.915 162.610 94.175 163.065 ;
        RECT 94.345 162.415 94.595 162.895 ;
        RECT 94.775 162.610 95.035 163.065 ;
        RECT 95.205 162.415 95.455 162.895 ;
        RECT 95.635 162.610 95.895 163.065 ;
        RECT 96.065 162.415 96.310 162.895 ;
        RECT 96.480 162.610 96.755 163.065 ;
        RECT 96.925 162.415 97.170 162.895 ;
        RECT 97.340 162.610 97.600 163.065 ;
        RECT 97.770 162.415 98.030 162.895 ;
        RECT 98.200 162.610 98.460 163.065 ;
        RECT 98.630 162.415 98.890 162.895 ;
        RECT 99.060 162.610 99.320 163.065 ;
        RECT 99.490 162.415 99.750 162.975 ;
        RECT 99.920 162.595 100.170 163.405 ;
        RECT 100.350 162.415 100.610 162.940 ;
        RECT 100.780 162.595 101.030 163.405 ;
        RECT 101.200 163.095 101.515 163.655 ;
        RECT 102.145 163.395 102.485 164.205 ;
        RECT 103.235 163.960 103.405 164.625 ;
        RECT 103.800 164.285 104.925 164.455 ;
        RECT 102.655 163.770 103.405 163.960 ;
        RECT 103.575 163.945 104.585 164.115 ;
        RECT 102.145 163.225 103.375 163.395 ;
        RECT 101.210 162.415 101.515 162.925 ;
        RECT 101.685 162.415 101.975 163.140 ;
        RECT 102.420 162.620 102.665 163.225 ;
        RECT 102.885 162.415 103.395 162.950 ;
        RECT 103.575 162.585 103.765 163.945 ;
        RECT 103.935 163.265 104.210 163.745 ;
        RECT 103.935 163.095 104.215 163.265 ;
        RECT 104.415 163.145 104.585 163.945 ;
        RECT 104.755 163.155 104.925 164.285 ;
        RECT 105.095 163.655 105.265 164.625 ;
        RECT 105.435 163.825 105.605 164.965 ;
        RECT 105.775 163.825 106.110 164.795 ;
        RECT 105.095 163.325 105.290 163.655 ;
        RECT 105.515 163.325 105.770 163.655 ;
        RECT 105.515 163.155 105.685 163.325 ;
        RECT 105.940 163.155 106.110 163.825 ;
        RECT 103.935 162.585 104.210 163.095 ;
        RECT 104.755 162.985 105.685 163.155 ;
        RECT 104.755 162.950 104.930 162.985 ;
        RECT 104.400 162.585 104.930 162.950 ;
        RECT 105.355 162.415 105.685 162.815 ;
        RECT 105.855 162.585 106.110 163.155 ;
        RECT 106.750 163.825 107.085 164.795 ;
        RECT 107.255 163.825 107.425 164.965 ;
        RECT 107.595 164.625 109.625 164.795 ;
        RECT 106.750 163.155 106.920 163.825 ;
        RECT 107.595 163.655 107.765 164.625 ;
        RECT 107.090 163.325 107.345 163.655 ;
        RECT 107.570 163.325 107.765 163.655 ;
        RECT 107.935 164.285 109.060 164.455 ;
        RECT 107.175 163.155 107.345 163.325 ;
        RECT 107.935 163.155 108.105 164.285 ;
        RECT 106.750 162.585 107.005 163.155 ;
        RECT 107.175 162.985 108.105 163.155 ;
        RECT 108.275 163.945 109.285 164.115 ;
        RECT 108.275 163.145 108.445 163.945 ;
        RECT 107.930 162.950 108.105 162.985 ;
        RECT 107.175 162.415 107.505 162.815 ;
        RECT 107.930 162.585 108.460 162.950 ;
        RECT 108.650 162.925 108.925 163.745 ;
        RECT 108.645 162.755 108.925 162.925 ;
        RECT 108.650 162.585 108.925 162.755 ;
        RECT 109.095 162.585 109.285 163.945 ;
        RECT 109.455 163.960 109.625 164.625 ;
        RECT 109.795 164.205 109.965 164.965 ;
        RECT 110.200 164.205 110.715 164.615 ;
        RECT 109.455 163.770 110.205 163.960 ;
        RECT 110.375 163.395 110.715 164.205 ;
        RECT 111.035 163.815 111.365 164.965 ;
        RECT 111.535 163.945 111.705 164.795 ;
        RECT 111.875 164.165 112.205 164.965 ;
        RECT 112.375 163.945 112.545 164.795 ;
        RECT 112.725 164.165 112.965 164.965 ;
        RECT 113.135 163.985 113.465 164.795 ;
        RECT 109.485 163.225 110.715 163.395 ;
        RECT 111.535 163.775 112.545 163.945 ;
        RECT 112.750 163.815 113.465 163.985 ;
        RECT 111.535 163.265 112.030 163.775 ;
        RECT 112.750 163.575 112.920 163.815 ;
        RECT 113.650 163.775 113.905 164.655 ;
        RECT 114.075 163.825 114.380 164.965 ;
        RECT 114.720 164.585 115.050 164.965 ;
        RECT 115.230 164.415 115.400 164.705 ;
        RECT 115.570 164.505 115.820 164.965 ;
        RECT 114.600 164.245 115.400 164.415 ;
        RECT 115.990 164.455 116.860 164.795 ;
        RECT 112.420 163.405 112.920 163.575 ;
        RECT 113.090 163.405 113.470 163.645 ;
        RECT 111.535 163.235 112.035 163.265 ;
        RECT 112.750 163.235 112.920 163.405 ;
        RECT 109.465 162.415 109.975 162.950 ;
        RECT 110.195 162.620 110.440 163.225 ;
        RECT 111.035 162.415 111.365 163.215 ;
        RECT 111.535 163.065 112.545 163.235 ;
        RECT 112.750 163.065 113.385 163.235 ;
        RECT 111.535 162.585 111.705 163.065 ;
        RECT 111.875 162.415 112.205 162.895 ;
        RECT 112.375 162.585 112.545 163.065 ;
        RECT 112.795 162.415 113.035 162.895 ;
        RECT 113.215 162.585 113.385 163.065 ;
        RECT 113.650 163.125 113.860 163.775 ;
        RECT 114.600 163.655 114.770 164.245 ;
        RECT 115.990 164.075 116.160 164.455 ;
        RECT 117.095 164.335 117.265 164.795 ;
        RECT 117.435 164.505 117.805 164.965 ;
        RECT 118.100 164.365 118.270 164.705 ;
        RECT 118.440 164.535 118.770 164.965 ;
        RECT 119.005 164.365 119.175 164.705 ;
        RECT 114.940 163.905 116.160 164.075 ;
        RECT 116.330 163.995 116.790 164.285 ;
        RECT 117.095 164.165 117.655 164.335 ;
        RECT 118.100 164.195 119.175 164.365 ;
        RECT 119.345 164.465 120.025 164.795 ;
        RECT 120.240 164.465 120.490 164.795 ;
        RECT 120.660 164.505 120.910 164.965 ;
        RECT 117.485 164.025 117.655 164.165 ;
        RECT 116.330 163.985 117.295 163.995 ;
        RECT 115.990 163.815 116.160 163.905 ;
        RECT 116.620 163.825 117.295 163.985 ;
        RECT 114.030 163.625 114.770 163.655 ;
        RECT 114.030 163.325 114.945 163.625 ;
        RECT 114.620 163.150 114.945 163.325 ;
        RECT 113.650 162.595 113.905 163.125 ;
        RECT 114.075 162.415 114.380 162.875 ;
        RECT 114.625 162.795 114.945 163.150 ;
        RECT 115.115 163.365 115.655 163.735 ;
        RECT 115.990 163.645 116.395 163.815 ;
        RECT 115.115 162.965 115.355 163.365 ;
        RECT 115.835 163.195 116.055 163.475 ;
        RECT 115.525 163.025 116.055 163.195 ;
        RECT 115.525 162.795 115.695 163.025 ;
        RECT 116.225 162.865 116.395 163.645 ;
        RECT 116.565 163.035 116.915 163.655 ;
        RECT 117.085 163.035 117.295 163.825 ;
        RECT 117.485 163.855 118.985 164.025 ;
        RECT 117.485 163.165 117.655 163.855 ;
        RECT 119.345 163.685 119.515 164.465 ;
        RECT 120.320 164.335 120.490 164.465 ;
        RECT 117.825 163.515 119.515 163.685 ;
        RECT 119.685 163.905 120.150 164.295 ;
        RECT 120.320 164.165 120.715 164.335 ;
        RECT 117.825 163.335 117.995 163.515 ;
        RECT 114.625 162.625 115.695 162.795 ;
        RECT 115.865 162.415 116.055 162.855 ;
        RECT 116.225 162.585 117.175 162.865 ;
        RECT 117.485 162.775 117.745 163.165 ;
        RECT 118.165 163.095 118.955 163.345 ;
        RECT 117.395 162.605 117.745 162.775 ;
        RECT 117.955 162.415 118.285 162.875 ;
        RECT 119.160 162.805 119.330 163.515 ;
        RECT 119.685 163.315 119.855 163.905 ;
        RECT 119.500 163.095 119.855 163.315 ;
        RECT 120.025 163.095 120.375 163.715 ;
        RECT 120.545 162.805 120.715 164.165 ;
        RECT 121.080 163.995 121.405 164.780 ;
        RECT 120.885 162.945 121.345 163.995 ;
        RECT 119.160 162.635 120.015 162.805 ;
        RECT 120.220 162.635 120.715 162.805 ;
        RECT 120.885 162.415 121.215 162.775 ;
        RECT 121.575 162.675 121.745 164.795 ;
        RECT 121.915 164.465 122.245 164.965 ;
        RECT 122.415 164.295 122.670 164.795 ;
        RECT 121.920 164.125 122.670 164.295 ;
        RECT 121.920 163.135 122.150 164.125 ;
        RECT 122.320 163.305 122.670 163.955 ;
        RECT 122.845 163.890 123.115 164.795 ;
        RECT 123.285 164.205 123.615 164.965 ;
        RECT 123.795 164.035 123.965 164.795 ;
        RECT 121.920 162.965 122.670 163.135 ;
        RECT 121.915 162.415 122.245 162.795 ;
        RECT 122.415 162.675 122.670 162.965 ;
        RECT 122.845 163.090 123.015 163.890 ;
        RECT 123.300 163.865 123.965 164.035 ;
        RECT 124.685 163.875 126.355 164.965 ;
        RECT 126.525 163.875 127.735 164.965 ;
        RECT 123.300 163.720 123.470 163.865 ;
        RECT 123.185 163.390 123.470 163.720 ;
        RECT 123.300 163.135 123.470 163.390 ;
        RECT 123.705 163.315 124.035 163.685 ;
        RECT 124.685 163.355 125.435 163.875 ;
        RECT 125.605 163.185 126.355 163.705 ;
        RECT 126.525 163.335 127.045 163.875 ;
        RECT 122.845 162.585 123.105 163.090 ;
        RECT 123.300 162.965 123.965 163.135 ;
        RECT 123.285 162.415 123.615 162.795 ;
        RECT 123.795 162.585 123.965 162.965 ;
        RECT 124.685 162.415 126.355 163.185 ;
        RECT 127.215 163.165 127.735 163.705 ;
        RECT 126.525 162.415 127.735 163.165 ;
        RECT 14.660 162.245 127.820 162.415 ;
        RECT 14.745 161.495 15.955 162.245 ;
        RECT 14.745 160.955 15.265 161.495 ;
        RECT 16.125 161.475 17.795 162.245 ;
        RECT 15.435 160.785 15.955 161.325 ;
        RECT 14.745 159.695 15.955 160.785 ;
        RECT 16.125 160.785 16.875 161.305 ;
        RECT 17.045 160.955 17.795 161.475 ;
        RECT 18.340 161.535 18.595 162.065 ;
        RECT 18.775 161.785 19.060 162.245 ;
        RECT 16.125 159.695 17.795 160.785 ;
        RECT 18.340 160.675 18.520 161.535 ;
        RECT 19.240 161.335 19.490 161.985 ;
        RECT 18.690 161.005 19.490 161.335 ;
        RECT 18.340 160.205 18.595 160.675 ;
        RECT 18.255 160.035 18.595 160.205 ;
        RECT 18.340 160.005 18.595 160.035 ;
        RECT 18.775 159.695 19.060 160.495 ;
        RECT 19.240 160.415 19.490 161.005 ;
        RECT 19.690 161.650 20.010 161.980 ;
        RECT 20.190 161.765 20.850 162.245 ;
        RECT 21.050 161.855 21.900 162.025 ;
        RECT 19.690 160.755 19.880 161.650 ;
        RECT 20.200 161.325 20.860 161.595 ;
        RECT 20.530 161.265 20.860 161.325 ;
        RECT 20.050 161.095 20.380 161.155 ;
        RECT 21.050 161.095 21.220 161.855 ;
        RECT 22.460 161.785 22.780 162.245 ;
        RECT 22.980 161.605 23.230 162.035 ;
        RECT 23.520 161.805 23.930 162.245 ;
        RECT 24.100 161.865 25.115 162.065 ;
        RECT 21.390 161.435 22.640 161.605 ;
        RECT 21.390 161.315 21.720 161.435 ;
        RECT 20.050 160.925 21.950 161.095 ;
        RECT 19.690 160.585 21.610 160.755 ;
        RECT 19.690 160.565 20.010 160.585 ;
        RECT 19.240 159.905 19.570 160.415 ;
        RECT 19.840 159.955 20.010 160.565 ;
        RECT 21.780 160.415 21.950 160.925 ;
        RECT 22.120 160.855 22.300 161.265 ;
        RECT 22.470 160.675 22.640 161.435 ;
        RECT 20.180 159.695 20.510 160.385 ;
        RECT 20.740 160.245 21.950 160.415 ;
        RECT 22.120 160.365 22.640 160.675 ;
        RECT 22.810 161.265 23.230 161.605 ;
        RECT 23.520 161.265 23.930 161.595 ;
        RECT 22.810 160.495 23.000 161.265 ;
        RECT 24.100 161.135 24.270 161.865 ;
        RECT 25.415 161.695 25.585 162.025 ;
        RECT 25.755 161.865 26.085 162.245 ;
        RECT 24.440 161.315 24.790 161.685 ;
        RECT 24.100 161.095 24.520 161.135 ;
        RECT 23.170 160.925 24.520 161.095 ;
        RECT 23.170 160.765 23.420 160.925 ;
        RECT 23.930 160.495 24.180 160.755 ;
        RECT 22.810 160.245 24.180 160.495 ;
        RECT 20.740 159.955 20.980 160.245 ;
        RECT 21.780 160.165 21.950 160.245 ;
        RECT 21.180 159.695 21.600 160.075 ;
        RECT 21.780 159.915 22.410 160.165 ;
        RECT 22.880 159.695 23.210 160.075 ;
        RECT 23.380 159.955 23.550 160.245 ;
        RECT 24.350 160.080 24.520 160.925 ;
        RECT 24.970 160.755 25.190 161.625 ;
        RECT 25.415 161.505 26.110 161.695 ;
        RECT 24.690 160.375 25.190 160.755 ;
        RECT 25.360 160.705 25.770 161.325 ;
        RECT 25.940 160.535 26.110 161.505 ;
        RECT 25.415 160.365 26.110 160.535 ;
        RECT 23.730 159.695 24.110 160.075 ;
        RECT 24.350 159.910 25.180 160.080 ;
        RECT 25.415 159.865 25.585 160.365 ;
        RECT 25.755 159.695 26.085 160.195 ;
        RECT 26.300 159.865 26.525 161.985 ;
        RECT 26.695 161.865 27.025 162.245 ;
        RECT 27.195 161.695 27.365 161.985 ;
        RECT 26.700 161.525 27.365 161.695 ;
        RECT 26.700 160.535 26.930 161.525 ;
        RECT 27.630 161.505 27.885 162.075 ;
        RECT 28.055 161.845 28.385 162.245 ;
        RECT 28.810 161.710 29.340 162.075 ;
        RECT 28.810 161.675 28.985 161.710 ;
        RECT 28.055 161.505 28.985 161.675 ;
        RECT 29.530 161.565 29.805 162.075 ;
        RECT 27.100 160.705 27.450 161.355 ;
        RECT 27.630 160.835 27.800 161.505 ;
        RECT 28.055 161.335 28.225 161.505 ;
        RECT 27.970 161.005 28.225 161.335 ;
        RECT 28.450 161.005 28.645 161.335 ;
        RECT 26.700 160.365 27.365 160.535 ;
        RECT 26.695 159.695 27.025 160.195 ;
        RECT 27.195 159.865 27.365 160.365 ;
        RECT 27.630 159.865 27.965 160.835 ;
        RECT 28.135 159.695 28.305 160.835 ;
        RECT 28.475 160.035 28.645 161.005 ;
        RECT 28.815 160.375 28.985 161.505 ;
        RECT 29.155 160.715 29.325 161.515 ;
        RECT 29.525 161.395 29.805 161.565 ;
        RECT 29.530 160.915 29.805 161.395 ;
        RECT 29.975 160.715 30.165 162.075 ;
        RECT 30.345 161.710 30.855 162.245 ;
        RECT 31.075 161.435 31.320 162.040 ;
        RECT 31.765 161.495 32.975 162.245 ;
        RECT 30.365 161.265 31.595 161.435 ;
        RECT 29.155 160.545 30.165 160.715 ;
        RECT 30.335 160.700 31.085 160.890 ;
        RECT 28.815 160.205 29.940 160.375 ;
        RECT 30.335 160.035 30.505 160.700 ;
        RECT 31.255 160.455 31.595 161.265 ;
        RECT 28.475 159.865 30.505 160.035 ;
        RECT 30.675 159.695 30.845 160.455 ;
        RECT 31.080 160.045 31.595 160.455 ;
        RECT 31.765 160.785 32.285 161.325 ;
        RECT 32.455 160.955 32.975 161.495 ;
        RECT 33.150 161.505 33.405 162.075 ;
        RECT 33.575 161.845 33.905 162.245 ;
        RECT 34.330 161.710 34.860 162.075 ;
        RECT 34.330 161.675 34.505 161.710 ;
        RECT 33.575 161.505 34.505 161.675 ;
        RECT 35.050 161.565 35.325 162.075 ;
        RECT 33.150 160.835 33.320 161.505 ;
        RECT 33.575 161.335 33.745 161.505 ;
        RECT 33.490 161.005 33.745 161.335 ;
        RECT 33.970 161.005 34.165 161.335 ;
        RECT 31.765 159.695 32.975 160.785 ;
        RECT 33.150 159.865 33.485 160.835 ;
        RECT 33.655 159.695 33.825 160.835 ;
        RECT 33.995 160.035 34.165 161.005 ;
        RECT 34.335 160.375 34.505 161.505 ;
        RECT 34.675 160.715 34.845 161.515 ;
        RECT 35.045 161.395 35.325 161.565 ;
        RECT 35.050 160.915 35.325 161.395 ;
        RECT 35.495 160.715 35.685 162.075 ;
        RECT 35.865 161.710 36.375 162.245 ;
        RECT 36.595 161.435 36.840 162.040 ;
        RECT 37.285 161.520 37.575 162.245 ;
        RECT 38.205 161.475 39.875 162.245 ;
        RECT 35.885 161.265 37.115 161.435 ;
        RECT 34.675 160.545 35.685 160.715 ;
        RECT 35.855 160.700 36.605 160.890 ;
        RECT 34.335 160.205 35.460 160.375 ;
        RECT 35.855 160.035 36.025 160.700 ;
        RECT 36.775 160.455 37.115 161.265 ;
        RECT 33.995 159.865 36.025 160.035 ;
        RECT 36.195 159.695 36.365 160.455 ;
        RECT 36.600 160.045 37.115 160.455 ;
        RECT 37.285 159.695 37.575 160.860 ;
        RECT 38.205 160.785 38.955 161.305 ;
        RECT 39.125 160.955 39.875 161.475 ;
        RECT 40.160 161.615 40.445 162.075 ;
        RECT 40.615 161.785 40.885 162.245 ;
        RECT 40.160 161.445 41.115 161.615 ;
        RECT 38.205 159.695 39.875 160.785 ;
        RECT 40.045 160.715 40.735 161.275 ;
        RECT 40.905 160.545 41.115 161.445 ;
        RECT 40.160 160.325 41.115 160.545 ;
        RECT 41.285 161.275 41.685 162.075 ;
        RECT 41.875 161.615 42.155 162.075 ;
        RECT 42.675 161.785 43.000 162.245 ;
        RECT 41.875 161.445 43.000 161.615 ;
        RECT 43.170 161.505 43.555 162.075 ;
        RECT 42.550 161.335 43.000 161.445 ;
        RECT 41.285 160.715 42.380 161.275 ;
        RECT 42.550 161.005 43.105 161.335 ;
        RECT 40.160 159.865 40.445 160.325 ;
        RECT 40.615 159.695 40.885 160.155 ;
        RECT 41.285 159.865 41.685 160.715 ;
        RECT 42.550 160.545 43.000 161.005 ;
        RECT 43.275 160.835 43.555 161.505 ;
        RECT 41.875 160.325 43.000 160.545 ;
        RECT 41.875 159.865 42.155 160.325 ;
        RECT 42.675 159.695 43.000 160.155 ;
        RECT 43.170 159.865 43.555 160.835 ;
        RECT 43.730 161.505 43.985 162.075 ;
        RECT 44.155 161.845 44.485 162.245 ;
        RECT 44.910 161.710 45.440 162.075 ;
        RECT 45.630 161.905 45.905 162.075 ;
        RECT 45.625 161.735 45.905 161.905 ;
        RECT 44.910 161.675 45.085 161.710 ;
        RECT 44.155 161.505 45.085 161.675 ;
        RECT 43.730 160.835 43.900 161.505 ;
        RECT 44.155 161.335 44.325 161.505 ;
        RECT 44.070 161.005 44.325 161.335 ;
        RECT 44.550 161.005 44.745 161.335 ;
        RECT 43.730 159.865 44.065 160.835 ;
        RECT 44.235 159.695 44.405 160.835 ;
        RECT 44.575 160.035 44.745 161.005 ;
        RECT 44.915 160.375 45.085 161.505 ;
        RECT 45.255 160.715 45.425 161.515 ;
        RECT 45.630 160.915 45.905 161.735 ;
        RECT 46.075 160.715 46.265 162.075 ;
        RECT 46.445 161.710 46.955 162.245 ;
        RECT 47.175 161.435 47.420 162.040 ;
        RECT 47.865 161.570 48.125 162.075 ;
        RECT 48.305 161.865 48.635 162.245 ;
        RECT 48.815 161.695 48.985 162.075 ;
        RECT 46.465 161.265 47.695 161.435 ;
        RECT 45.255 160.545 46.265 160.715 ;
        RECT 46.435 160.700 47.185 160.890 ;
        RECT 44.915 160.205 46.040 160.375 ;
        RECT 46.435 160.035 46.605 160.700 ;
        RECT 47.355 160.455 47.695 161.265 ;
        RECT 44.575 159.865 46.605 160.035 ;
        RECT 46.775 159.695 46.945 160.455 ;
        RECT 47.180 160.045 47.695 160.455 ;
        RECT 47.865 160.770 48.035 161.570 ;
        RECT 48.320 161.525 48.985 161.695 ;
        RECT 48.320 161.270 48.490 161.525 ;
        RECT 49.250 161.505 49.505 162.075 ;
        RECT 49.675 161.845 50.005 162.245 ;
        RECT 50.430 161.710 50.960 162.075 ;
        RECT 50.430 161.675 50.605 161.710 ;
        RECT 49.675 161.505 50.605 161.675 ;
        RECT 48.205 160.940 48.490 161.270 ;
        RECT 48.725 160.975 49.055 161.345 ;
        RECT 48.320 160.795 48.490 160.940 ;
        RECT 49.250 160.835 49.420 161.505 ;
        RECT 49.675 161.335 49.845 161.505 ;
        RECT 49.590 161.005 49.845 161.335 ;
        RECT 50.070 161.005 50.265 161.335 ;
        RECT 47.865 159.865 48.135 160.770 ;
        RECT 48.320 160.625 48.985 160.795 ;
        RECT 48.305 159.695 48.635 160.455 ;
        RECT 48.815 159.865 48.985 160.625 ;
        RECT 49.250 159.865 49.585 160.835 ;
        RECT 49.755 159.695 49.925 160.835 ;
        RECT 50.095 160.035 50.265 161.005 ;
        RECT 50.435 160.375 50.605 161.505 ;
        RECT 50.775 160.715 50.945 161.515 ;
        RECT 51.150 161.225 51.425 162.075 ;
        RECT 51.145 161.055 51.425 161.225 ;
        RECT 51.150 160.915 51.425 161.055 ;
        RECT 51.595 160.715 51.785 162.075 ;
        RECT 51.965 161.710 52.475 162.245 ;
        RECT 52.695 161.435 52.940 162.040 ;
        RECT 53.660 161.435 53.905 162.040 ;
        RECT 54.125 161.710 54.635 162.245 ;
        RECT 51.985 161.265 53.215 161.435 ;
        RECT 50.775 160.545 51.785 160.715 ;
        RECT 51.955 160.700 52.705 160.890 ;
        RECT 50.435 160.205 51.560 160.375 ;
        RECT 51.955 160.035 52.125 160.700 ;
        RECT 52.875 160.455 53.215 161.265 ;
        RECT 50.095 159.865 52.125 160.035 ;
        RECT 52.295 159.695 52.465 160.455 ;
        RECT 52.700 160.045 53.215 160.455 ;
        RECT 53.385 161.265 54.615 161.435 ;
        RECT 53.385 160.455 53.725 161.265 ;
        RECT 53.895 160.700 54.645 160.890 ;
        RECT 53.385 160.045 53.900 160.455 ;
        RECT 54.135 159.695 54.305 160.455 ;
        RECT 54.475 160.035 54.645 160.700 ;
        RECT 54.815 160.715 55.005 162.075 ;
        RECT 55.175 161.905 55.450 162.075 ;
        RECT 55.175 161.735 55.455 161.905 ;
        RECT 55.175 160.915 55.450 161.735 ;
        RECT 55.640 161.710 56.170 162.075 ;
        RECT 56.595 161.845 56.925 162.245 ;
        RECT 55.995 161.675 56.170 161.710 ;
        RECT 55.655 160.715 55.825 161.515 ;
        RECT 54.815 160.545 55.825 160.715 ;
        RECT 55.995 161.505 56.925 161.675 ;
        RECT 57.095 161.505 57.350 162.075 ;
        RECT 55.995 160.375 56.165 161.505 ;
        RECT 56.755 161.335 56.925 161.505 ;
        RECT 55.040 160.205 56.165 160.375 ;
        RECT 56.335 161.005 56.530 161.335 ;
        RECT 56.755 161.005 57.010 161.335 ;
        RECT 56.335 160.035 56.505 161.005 ;
        RECT 57.180 160.835 57.350 161.505 ;
        RECT 57.985 161.475 59.655 162.245 ;
        RECT 59.915 161.695 60.085 162.075 ;
        RECT 60.265 161.865 60.595 162.245 ;
        RECT 59.915 161.525 60.580 161.695 ;
        RECT 60.775 161.570 61.035 162.075 ;
        RECT 54.475 159.865 56.505 160.035 ;
        RECT 56.675 159.695 56.845 160.835 ;
        RECT 57.015 159.865 57.350 160.835 ;
        RECT 57.985 160.785 58.735 161.305 ;
        RECT 58.905 160.955 59.655 161.475 ;
        RECT 59.845 160.975 60.175 161.345 ;
        RECT 60.410 161.270 60.580 161.525 ;
        RECT 60.410 160.940 60.695 161.270 ;
        RECT 60.410 160.795 60.580 160.940 ;
        RECT 57.985 159.695 59.655 160.785 ;
        RECT 59.915 160.625 60.580 160.795 ;
        RECT 60.865 160.770 61.035 161.570 ;
        RECT 61.205 161.475 62.875 162.245 ;
        RECT 63.045 161.520 63.335 162.245 ;
        RECT 63.505 161.495 64.715 162.245 ;
        RECT 59.915 159.865 60.085 160.625 ;
        RECT 60.265 159.695 60.595 160.455 ;
        RECT 60.765 159.865 61.035 160.770 ;
        RECT 61.205 160.785 61.955 161.305 ;
        RECT 62.125 160.955 62.875 161.475 ;
        RECT 61.205 159.695 62.875 160.785 ;
        RECT 63.045 159.695 63.335 160.860 ;
        RECT 63.505 160.785 64.025 161.325 ;
        RECT 64.195 160.955 64.715 161.495 ;
        RECT 64.890 161.405 65.150 162.245 ;
        RECT 65.325 161.500 65.580 162.075 ;
        RECT 65.750 161.865 66.080 162.245 ;
        RECT 66.295 161.695 66.465 162.075 ;
        RECT 65.750 161.525 66.465 161.695 ;
        RECT 63.505 159.695 64.715 160.785 ;
        RECT 64.890 159.695 65.150 160.845 ;
        RECT 65.325 160.770 65.495 161.500 ;
        RECT 65.750 161.335 65.920 161.525 ;
        RECT 66.730 161.405 66.990 162.245 ;
        RECT 67.165 161.500 67.420 162.075 ;
        RECT 67.590 161.865 67.920 162.245 ;
        RECT 68.135 161.695 68.305 162.075 ;
        RECT 67.590 161.525 68.305 161.695 ;
        RECT 68.655 161.695 68.825 162.075 ;
        RECT 69.040 161.865 69.370 162.245 ;
        RECT 68.655 161.525 69.370 161.695 ;
        RECT 65.665 161.005 65.920 161.335 ;
        RECT 65.750 160.795 65.920 161.005 ;
        RECT 66.200 160.975 66.555 161.345 ;
        RECT 65.325 159.865 65.580 160.770 ;
        RECT 65.750 160.625 66.465 160.795 ;
        RECT 65.750 159.695 66.080 160.455 ;
        RECT 66.295 159.865 66.465 160.625 ;
        RECT 66.730 159.695 66.990 160.845 ;
        RECT 67.165 160.770 67.335 161.500 ;
        RECT 67.590 161.335 67.760 161.525 ;
        RECT 67.505 161.005 67.760 161.335 ;
        RECT 67.590 160.795 67.760 161.005 ;
        RECT 68.040 160.975 68.395 161.345 ;
        RECT 68.565 160.975 68.920 161.345 ;
        RECT 69.200 161.335 69.370 161.525 ;
        RECT 69.540 161.500 69.795 162.075 ;
        RECT 69.200 161.005 69.455 161.335 ;
        RECT 69.200 160.795 69.370 161.005 ;
        RECT 67.165 159.865 67.420 160.770 ;
        RECT 67.590 160.625 68.305 160.795 ;
        RECT 67.590 159.695 67.920 160.455 ;
        RECT 68.135 159.865 68.305 160.625 ;
        RECT 68.655 160.625 69.370 160.795 ;
        RECT 69.625 160.770 69.795 161.500 ;
        RECT 69.970 161.405 70.230 162.245 ;
        RECT 70.495 161.695 70.665 162.075 ;
        RECT 70.880 161.865 71.210 162.245 ;
        RECT 70.495 161.525 71.210 161.695 ;
        RECT 70.405 160.975 70.760 161.345 ;
        RECT 71.040 161.335 71.210 161.525 ;
        RECT 71.380 161.500 71.635 162.075 ;
        RECT 71.040 161.005 71.295 161.335 ;
        RECT 68.655 159.865 68.825 160.625 ;
        RECT 69.040 159.695 69.370 160.455 ;
        RECT 69.540 159.865 69.795 160.770 ;
        RECT 69.970 159.695 70.230 160.845 ;
        RECT 71.040 160.795 71.210 161.005 ;
        RECT 70.495 160.625 71.210 160.795 ;
        RECT 71.465 160.770 71.635 161.500 ;
        RECT 71.810 161.405 72.070 162.245 ;
        RECT 72.705 161.475 75.295 162.245 ;
        RECT 75.470 161.700 80.815 162.245 ;
        RECT 70.495 159.865 70.665 160.625 ;
        RECT 70.880 159.695 71.210 160.455 ;
        RECT 71.380 159.865 71.635 160.770 ;
        RECT 71.810 159.695 72.070 160.845 ;
        RECT 72.705 160.785 73.915 161.305 ;
        RECT 74.085 160.955 75.295 161.475 ;
        RECT 72.705 159.695 75.295 160.785 ;
        RECT 77.060 160.130 77.410 161.380 ;
        RECT 78.890 160.870 79.230 161.700 ;
        RECT 81.045 161.425 81.255 162.245 ;
        RECT 81.425 161.445 81.755 162.075 ;
        RECT 81.425 160.845 81.675 161.445 ;
        RECT 81.925 161.425 82.155 162.245 ;
        RECT 82.640 161.435 82.885 162.040 ;
        RECT 83.105 161.710 83.615 162.245 ;
        RECT 82.365 161.265 83.595 161.435 ;
        RECT 81.845 161.005 82.175 161.255 ;
        RECT 75.470 159.695 80.815 160.130 ;
        RECT 81.045 159.695 81.255 160.835 ;
        RECT 81.425 159.865 81.755 160.845 ;
        RECT 81.925 159.695 82.155 160.835 ;
        RECT 82.365 160.455 82.705 161.265 ;
        RECT 82.875 160.700 83.625 160.890 ;
        RECT 82.365 160.045 82.880 160.455 ;
        RECT 83.115 159.695 83.285 160.455 ;
        RECT 83.455 160.035 83.625 160.700 ;
        RECT 83.795 160.715 83.985 162.075 ;
        RECT 84.155 161.565 84.430 162.075 ;
        RECT 84.620 161.710 85.150 162.075 ;
        RECT 85.575 161.845 85.905 162.245 ;
        RECT 84.975 161.675 85.150 161.710 ;
        RECT 84.155 161.395 84.435 161.565 ;
        RECT 84.155 160.915 84.430 161.395 ;
        RECT 84.635 160.715 84.805 161.515 ;
        RECT 83.795 160.545 84.805 160.715 ;
        RECT 84.975 161.505 85.905 161.675 ;
        RECT 86.075 161.505 86.330 162.075 ;
        RECT 86.595 161.695 86.765 162.075 ;
        RECT 86.945 161.865 87.275 162.245 ;
        RECT 86.595 161.525 87.260 161.695 ;
        RECT 87.455 161.570 87.715 162.075 ;
        RECT 84.975 160.375 85.145 161.505 ;
        RECT 85.735 161.335 85.905 161.505 ;
        RECT 84.020 160.205 85.145 160.375 ;
        RECT 85.315 161.005 85.510 161.335 ;
        RECT 85.735 161.005 85.990 161.335 ;
        RECT 85.315 160.035 85.485 161.005 ;
        RECT 86.160 160.835 86.330 161.505 ;
        RECT 86.525 160.975 86.855 161.345 ;
        RECT 87.090 161.270 87.260 161.525 ;
        RECT 83.455 159.865 85.485 160.035 ;
        RECT 85.655 159.695 85.825 160.835 ;
        RECT 85.995 159.865 86.330 160.835 ;
        RECT 87.090 160.940 87.375 161.270 ;
        RECT 87.090 160.795 87.260 160.940 ;
        RECT 86.595 160.625 87.260 160.795 ;
        RECT 87.545 160.770 87.715 161.570 ;
        RECT 88.805 161.520 89.095 162.245 ;
        RECT 90.100 161.905 90.355 162.065 ;
        RECT 90.015 161.735 90.355 161.905 ;
        RECT 90.535 161.785 90.820 162.245 ;
        RECT 90.100 161.535 90.355 161.735 ;
        RECT 86.595 159.865 86.765 160.625 ;
        RECT 86.945 159.695 87.275 160.455 ;
        RECT 87.445 159.865 87.715 160.770 ;
        RECT 88.805 159.695 89.095 160.860 ;
        RECT 90.100 160.675 90.280 161.535 ;
        RECT 91.000 161.335 91.250 161.985 ;
        RECT 90.450 161.005 91.250 161.335 ;
        RECT 90.100 160.005 90.355 160.675 ;
        RECT 90.535 159.695 90.820 160.495 ;
        RECT 91.000 160.415 91.250 161.005 ;
        RECT 91.450 161.650 91.770 161.980 ;
        RECT 91.950 161.765 92.610 162.245 ;
        RECT 92.810 161.855 93.660 162.025 ;
        RECT 91.450 160.755 91.640 161.650 ;
        RECT 91.960 161.325 92.620 161.595 ;
        RECT 92.290 161.265 92.620 161.325 ;
        RECT 91.810 161.095 92.140 161.155 ;
        RECT 92.810 161.095 92.980 161.855 ;
        RECT 94.220 161.785 94.540 162.245 ;
        RECT 94.740 161.605 94.990 162.035 ;
        RECT 95.280 161.805 95.690 162.245 ;
        RECT 95.860 161.865 96.875 162.065 ;
        RECT 93.150 161.435 94.400 161.605 ;
        RECT 93.150 161.315 93.480 161.435 ;
        RECT 91.810 160.925 93.710 161.095 ;
        RECT 91.450 160.585 93.370 160.755 ;
        RECT 91.450 160.565 91.770 160.585 ;
        RECT 91.000 159.905 91.330 160.415 ;
        RECT 91.600 159.955 91.770 160.565 ;
        RECT 93.540 160.415 93.710 160.925 ;
        RECT 93.880 160.855 94.060 161.265 ;
        RECT 94.230 160.675 94.400 161.435 ;
        RECT 91.940 159.695 92.270 160.385 ;
        RECT 92.500 160.245 93.710 160.415 ;
        RECT 93.880 160.365 94.400 160.675 ;
        RECT 94.570 161.265 94.990 161.605 ;
        RECT 95.280 161.265 95.690 161.595 ;
        RECT 94.570 160.495 94.760 161.265 ;
        RECT 95.860 161.135 96.030 161.865 ;
        RECT 97.175 161.695 97.345 162.025 ;
        RECT 97.515 161.865 97.845 162.245 ;
        RECT 96.200 161.315 96.550 161.685 ;
        RECT 95.860 161.095 96.280 161.135 ;
        RECT 94.930 160.925 96.280 161.095 ;
        RECT 94.930 160.765 95.180 160.925 ;
        RECT 95.690 160.495 95.940 160.755 ;
        RECT 94.570 160.245 95.940 160.495 ;
        RECT 92.500 159.955 92.740 160.245 ;
        RECT 93.540 160.165 93.710 160.245 ;
        RECT 92.940 159.695 93.360 160.075 ;
        RECT 93.540 159.915 94.170 160.165 ;
        RECT 94.640 159.695 94.970 160.075 ;
        RECT 95.140 159.955 95.310 160.245 ;
        RECT 96.110 160.080 96.280 160.925 ;
        RECT 96.730 160.755 96.950 161.625 ;
        RECT 97.175 161.505 97.870 161.695 ;
        RECT 96.450 160.375 96.950 160.755 ;
        RECT 97.120 160.705 97.530 161.325 ;
        RECT 97.700 160.535 97.870 161.505 ;
        RECT 97.175 160.365 97.870 160.535 ;
        RECT 95.490 159.695 95.870 160.075 ;
        RECT 96.110 159.910 96.940 160.080 ;
        RECT 97.175 159.865 97.345 160.365 ;
        RECT 97.515 159.695 97.845 160.195 ;
        RECT 98.060 159.865 98.285 161.985 ;
        RECT 98.455 161.865 98.785 162.245 ;
        RECT 98.955 161.695 99.125 161.985 ;
        RECT 99.485 161.780 99.735 162.245 ;
        RECT 98.460 161.525 99.125 161.695 ;
        RECT 99.905 161.605 100.075 162.075 ;
        RECT 100.325 161.785 100.495 162.245 ;
        RECT 100.745 161.605 100.915 162.075 ;
        RECT 101.165 161.785 101.335 162.245 ;
        RECT 101.585 161.605 101.755 162.075 ;
        RECT 102.125 161.785 102.390 162.245 ;
        RECT 98.460 160.535 98.690 161.525 ;
        RECT 99.385 161.425 101.755 161.605 ;
        RECT 102.720 161.615 103.005 162.075 ;
        RECT 103.175 161.785 103.445 162.245 ;
        RECT 102.720 161.445 103.675 161.615 ;
        RECT 98.860 160.705 99.210 161.355 ;
        RECT 99.385 160.835 99.735 161.425 ;
        RECT 99.905 161.005 102.415 161.255 ;
        RECT 99.385 160.665 101.835 160.835 ;
        RECT 99.385 160.645 100.155 160.665 ;
        RECT 98.460 160.365 99.125 160.535 ;
        RECT 98.455 159.695 98.785 160.195 ;
        RECT 98.955 159.865 99.125 160.365 ;
        RECT 99.485 159.695 99.655 160.155 ;
        RECT 99.825 159.865 100.155 160.645 ;
        RECT 100.325 159.695 100.495 160.495 ;
        RECT 100.665 159.865 100.995 160.665 ;
        RECT 101.165 159.695 101.335 160.495 ;
        RECT 101.505 159.865 101.835 160.665 ;
        RECT 102.095 159.695 102.390 160.835 ;
        RECT 102.605 160.715 103.295 161.275 ;
        RECT 103.465 160.545 103.675 161.445 ;
        RECT 102.720 160.325 103.675 160.545 ;
        RECT 103.845 161.275 104.245 162.075 ;
        RECT 104.435 161.615 104.715 162.075 ;
        RECT 105.235 161.785 105.560 162.245 ;
        RECT 104.435 161.445 105.560 161.615 ;
        RECT 105.730 161.505 106.115 162.075 ;
        RECT 105.110 161.335 105.560 161.445 ;
        RECT 103.845 160.715 104.940 161.275 ;
        RECT 105.110 161.005 105.665 161.335 ;
        RECT 102.720 159.865 103.005 160.325 ;
        RECT 103.175 159.695 103.445 160.155 ;
        RECT 103.845 159.865 104.245 160.715 ;
        RECT 105.110 160.545 105.560 161.005 ;
        RECT 105.835 160.835 106.115 161.505 ;
        RECT 106.860 161.615 107.145 162.075 ;
        RECT 107.315 161.785 107.585 162.245 ;
        RECT 106.860 161.445 107.815 161.615 ;
        RECT 104.435 160.325 105.560 160.545 ;
        RECT 104.435 159.865 104.715 160.325 ;
        RECT 105.235 159.695 105.560 160.155 ;
        RECT 105.730 159.865 106.115 160.835 ;
        RECT 106.745 160.715 107.435 161.275 ;
        RECT 107.605 160.545 107.815 161.445 ;
        RECT 106.860 160.325 107.815 160.545 ;
        RECT 107.985 161.275 108.385 162.075 ;
        RECT 108.575 161.615 108.855 162.075 ;
        RECT 109.375 161.785 109.700 162.245 ;
        RECT 108.575 161.445 109.700 161.615 ;
        RECT 109.870 161.505 110.255 162.075 ;
        RECT 109.250 161.335 109.700 161.445 ;
        RECT 107.985 160.715 109.080 161.275 ;
        RECT 109.250 161.005 109.805 161.335 ;
        RECT 106.860 159.865 107.145 160.325 ;
        RECT 107.315 159.695 107.585 160.155 ;
        RECT 107.985 159.865 108.385 160.715 ;
        RECT 109.250 160.545 109.700 161.005 ;
        RECT 109.975 160.835 110.255 161.505 ;
        RECT 110.700 161.435 110.945 162.040 ;
        RECT 111.165 161.710 111.675 162.245 ;
        RECT 108.575 160.325 109.700 160.545 ;
        RECT 108.575 159.865 108.855 160.325 ;
        RECT 109.375 159.695 109.700 160.155 ;
        RECT 109.870 159.865 110.255 160.835 ;
        RECT 110.425 161.265 111.655 161.435 ;
        RECT 110.425 160.455 110.765 161.265 ;
        RECT 110.935 160.700 111.685 160.890 ;
        RECT 110.425 160.045 110.940 160.455 ;
        RECT 111.175 159.695 111.345 160.455 ;
        RECT 111.515 160.035 111.685 160.700 ;
        RECT 111.855 160.715 112.045 162.075 ;
        RECT 112.215 161.225 112.490 162.075 ;
        RECT 112.680 161.710 113.210 162.075 ;
        RECT 113.635 161.845 113.965 162.245 ;
        RECT 113.035 161.675 113.210 161.710 ;
        RECT 112.215 161.055 112.495 161.225 ;
        RECT 112.215 160.915 112.490 161.055 ;
        RECT 112.695 160.715 112.865 161.515 ;
        RECT 111.855 160.545 112.865 160.715 ;
        RECT 113.035 161.505 113.965 161.675 ;
        RECT 114.135 161.505 114.390 162.075 ;
        RECT 114.565 161.520 114.855 162.245 ;
        RECT 113.035 160.375 113.205 161.505 ;
        RECT 113.795 161.335 113.965 161.505 ;
        RECT 112.080 160.205 113.205 160.375 ;
        RECT 113.375 161.005 113.570 161.335 ;
        RECT 113.795 161.005 114.050 161.335 ;
        RECT 113.375 160.035 113.545 161.005 ;
        RECT 114.220 160.835 114.390 161.505 ;
        RECT 115.300 161.435 115.545 162.040 ;
        RECT 115.765 161.710 116.275 162.245 ;
        RECT 115.025 161.265 116.255 161.435 ;
        RECT 111.515 159.865 113.545 160.035 ;
        RECT 113.715 159.695 113.885 160.835 ;
        RECT 114.055 159.865 114.390 160.835 ;
        RECT 114.565 159.695 114.855 160.860 ;
        RECT 115.025 160.455 115.365 161.265 ;
        RECT 115.535 160.700 116.285 160.890 ;
        RECT 115.025 160.045 115.540 160.455 ;
        RECT 115.775 159.695 115.945 160.455 ;
        RECT 116.115 160.035 116.285 160.700 ;
        RECT 116.455 160.715 116.645 162.075 ;
        RECT 116.815 161.905 117.090 162.075 ;
        RECT 116.815 161.735 117.095 161.905 ;
        RECT 116.815 160.915 117.090 161.735 ;
        RECT 117.280 161.710 117.810 162.075 ;
        RECT 118.235 161.845 118.565 162.245 ;
        RECT 117.635 161.675 117.810 161.710 ;
        RECT 117.295 160.715 117.465 161.515 ;
        RECT 116.455 160.545 117.465 160.715 ;
        RECT 117.635 161.505 118.565 161.675 ;
        RECT 118.735 161.505 118.990 162.075 ;
        RECT 117.635 160.375 117.805 161.505 ;
        RECT 118.395 161.335 118.565 161.505 ;
        RECT 116.680 160.205 117.805 160.375 ;
        RECT 117.975 161.005 118.170 161.335 ;
        RECT 118.395 161.005 118.650 161.335 ;
        RECT 117.975 160.035 118.145 161.005 ;
        RECT 118.820 160.835 118.990 161.505 ;
        RECT 119.205 161.425 119.435 162.245 ;
        RECT 119.605 161.445 119.935 162.075 ;
        RECT 119.185 161.005 119.515 161.255 ;
        RECT 119.685 160.845 119.935 161.445 ;
        RECT 120.105 161.425 120.315 162.245 ;
        RECT 121.095 161.695 121.265 162.075 ;
        RECT 121.445 161.865 121.775 162.245 ;
        RECT 121.095 161.525 121.760 161.695 ;
        RECT 121.955 161.570 122.215 162.075 ;
        RECT 121.025 160.975 121.355 161.345 ;
        RECT 121.590 161.270 121.760 161.525 ;
        RECT 116.115 159.865 118.145 160.035 ;
        RECT 118.315 159.695 118.485 160.835 ;
        RECT 118.655 159.865 118.990 160.835 ;
        RECT 119.205 159.695 119.435 160.835 ;
        RECT 119.605 159.865 119.935 160.845 ;
        RECT 121.590 160.940 121.875 161.270 ;
        RECT 120.105 159.695 120.315 160.835 ;
        RECT 121.590 160.795 121.760 160.940 ;
        RECT 121.095 160.625 121.760 160.795 ;
        RECT 122.045 160.770 122.215 161.570 ;
        RECT 122.845 161.475 126.355 162.245 ;
        RECT 126.525 161.495 127.735 162.245 ;
        RECT 121.095 159.865 121.265 160.625 ;
        RECT 121.445 159.695 121.775 160.455 ;
        RECT 121.945 159.865 122.215 160.770 ;
        RECT 122.845 160.785 124.535 161.305 ;
        RECT 124.705 160.955 126.355 161.475 ;
        RECT 126.525 160.785 127.045 161.325 ;
        RECT 127.215 160.955 127.735 161.495 ;
        RECT 122.845 159.695 126.355 160.785 ;
        RECT 126.525 159.695 127.735 160.785 ;
        RECT 14.660 159.525 127.820 159.695 ;
        RECT 14.745 158.435 15.955 159.525 ;
        RECT 14.745 157.725 15.265 158.265 ;
        RECT 15.435 157.895 15.955 158.435 ;
        RECT 16.125 158.435 17.335 159.525 ;
        RECT 16.125 157.895 16.645 158.435 ;
        RECT 17.565 158.385 17.775 159.525 ;
        RECT 17.945 158.375 18.275 159.355 ;
        RECT 18.445 158.385 18.675 159.525 ;
        RECT 18.925 158.385 19.155 159.525 ;
        RECT 19.325 158.375 19.655 159.355 ;
        RECT 19.825 158.385 20.035 159.525 ;
        RECT 20.265 158.765 20.780 159.175 ;
        RECT 21.015 158.765 21.185 159.525 ;
        RECT 21.355 159.185 23.385 159.355 ;
        RECT 16.815 157.725 17.335 158.265 ;
        RECT 14.745 156.975 15.955 157.725 ;
        RECT 16.125 156.975 17.335 157.725 ;
        RECT 17.565 156.975 17.775 157.795 ;
        RECT 17.945 157.775 18.195 158.375 ;
        RECT 18.365 157.965 18.695 158.215 ;
        RECT 18.905 157.965 19.235 158.215 ;
        RECT 17.945 157.145 18.275 157.775 ;
        RECT 18.445 156.975 18.675 157.795 ;
        RECT 18.925 156.975 19.155 157.795 ;
        RECT 19.405 157.775 19.655 158.375 ;
        RECT 20.265 157.955 20.605 158.765 ;
        RECT 21.355 158.520 21.525 159.185 ;
        RECT 21.920 158.845 23.045 159.015 ;
        RECT 20.775 158.330 21.525 158.520 ;
        RECT 21.695 158.505 22.705 158.675 ;
        RECT 19.325 157.145 19.655 157.775 ;
        RECT 19.825 156.975 20.035 157.795 ;
        RECT 20.265 157.785 21.495 157.955 ;
        RECT 20.540 157.180 20.785 157.785 ;
        RECT 21.005 156.975 21.515 157.510 ;
        RECT 21.695 157.145 21.885 158.505 ;
        RECT 22.055 157.485 22.330 158.305 ;
        RECT 22.535 157.705 22.705 158.505 ;
        RECT 22.875 157.715 23.045 158.845 ;
        RECT 23.215 158.215 23.385 159.185 ;
        RECT 23.555 158.385 23.725 159.525 ;
        RECT 23.895 158.385 24.230 159.355 ;
        RECT 23.215 157.885 23.410 158.215 ;
        RECT 23.635 157.885 23.890 158.215 ;
        RECT 23.635 157.715 23.805 157.885 ;
        RECT 24.060 157.715 24.230 158.385 ;
        RECT 24.405 158.360 24.695 159.525 ;
        RECT 24.955 158.595 25.125 159.355 ;
        RECT 25.305 158.765 25.635 159.525 ;
        RECT 24.955 158.425 25.620 158.595 ;
        RECT 25.805 158.450 26.075 159.355 ;
        RECT 25.450 158.280 25.620 158.425 ;
        RECT 24.885 157.875 25.215 158.245 ;
        RECT 25.450 157.950 25.735 158.280 ;
        RECT 22.875 157.545 23.805 157.715 ;
        RECT 22.875 157.510 23.050 157.545 ;
        RECT 22.055 157.315 22.335 157.485 ;
        RECT 22.055 157.145 22.330 157.315 ;
        RECT 22.520 157.145 23.050 157.510 ;
        RECT 23.475 156.975 23.805 157.375 ;
        RECT 23.975 157.145 24.230 157.715 ;
        RECT 24.405 156.975 24.695 157.700 ;
        RECT 25.450 157.695 25.620 157.950 ;
        RECT 24.955 157.525 25.620 157.695 ;
        RECT 25.905 157.650 26.075 158.450 ;
        RECT 26.245 158.435 27.915 159.525 ;
        RECT 28.200 158.895 28.485 159.355 ;
        RECT 28.655 159.065 28.925 159.525 ;
        RECT 28.200 158.675 29.155 158.895 ;
        RECT 26.245 157.915 26.995 158.435 ;
        RECT 27.165 157.745 27.915 158.265 ;
        RECT 28.085 157.945 28.775 158.505 ;
        RECT 28.945 157.775 29.155 158.675 ;
        RECT 24.955 157.145 25.125 157.525 ;
        RECT 25.305 156.975 25.635 157.355 ;
        RECT 25.815 157.145 26.075 157.650 ;
        RECT 26.245 156.975 27.915 157.745 ;
        RECT 28.200 157.605 29.155 157.775 ;
        RECT 29.325 158.505 29.725 159.355 ;
        RECT 29.915 158.895 30.195 159.355 ;
        RECT 30.715 159.065 31.040 159.525 ;
        RECT 29.915 158.675 31.040 158.895 ;
        RECT 29.325 157.945 30.420 158.505 ;
        RECT 30.590 158.215 31.040 158.675 ;
        RECT 31.210 158.385 31.595 159.355 ;
        RECT 31.880 158.895 32.165 159.355 ;
        RECT 32.335 159.065 32.605 159.525 ;
        RECT 31.880 158.675 32.835 158.895 ;
        RECT 28.200 157.145 28.485 157.605 ;
        RECT 28.655 156.975 28.925 157.435 ;
        RECT 29.325 157.145 29.725 157.945 ;
        RECT 30.590 157.885 31.145 158.215 ;
        RECT 30.590 157.775 31.040 157.885 ;
        RECT 29.915 157.605 31.040 157.775 ;
        RECT 31.315 157.715 31.595 158.385 ;
        RECT 31.765 157.945 32.455 158.505 ;
        RECT 32.625 157.775 32.835 158.675 ;
        RECT 29.915 157.145 30.195 157.605 ;
        RECT 30.715 156.975 31.040 157.435 ;
        RECT 31.210 157.145 31.595 157.715 ;
        RECT 31.880 157.605 32.835 157.775 ;
        RECT 33.005 158.505 33.405 159.355 ;
        RECT 33.595 158.895 33.875 159.355 ;
        RECT 34.395 159.065 34.720 159.525 ;
        RECT 33.595 158.675 34.720 158.895 ;
        RECT 33.005 157.945 34.100 158.505 ;
        RECT 34.270 158.215 34.720 158.675 ;
        RECT 34.890 158.385 35.275 159.355 ;
        RECT 31.880 157.145 32.165 157.605 ;
        RECT 32.335 156.975 32.605 157.435 ;
        RECT 33.005 157.145 33.405 157.945 ;
        RECT 34.270 157.885 34.825 158.215 ;
        RECT 34.270 157.775 34.720 157.885 ;
        RECT 33.595 157.605 34.720 157.775 ;
        RECT 34.995 157.715 35.275 158.385 ;
        RECT 35.445 158.435 38.955 159.525 ;
        RECT 39.330 158.555 39.660 159.355 ;
        RECT 39.830 158.725 40.160 159.525 ;
        RECT 40.460 158.555 40.790 159.355 ;
        RECT 41.435 158.725 41.685 159.525 ;
        RECT 35.445 157.915 37.135 158.435 ;
        RECT 39.330 158.385 41.765 158.555 ;
        RECT 41.955 158.385 42.125 159.525 ;
        RECT 42.295 158.385 42.635 159.355 ;
        RECT 43.010 158.555 43.340 159.355 ;
        RECT 43.510 158.725 43.840 159.525 ;
        RECT 44.140 158.555 44.470 159.355 ;
        RECT 45.115 158.725 45.365 159.525 ;
        RECT 43.010 158.385 45.445 158.555 ;
        RECT 45.635 158.385 45.805 159.525 ;
        RECT 45.975 158.385 46.315 159.355 ;
        RECT 46.600 158.895 46.885 159.355 ;
        RECT 47.055 159.065 47.325 159.525 ;
        RECT 46.600 158.675 47.555 158.895 ;
        RECT 37.305 157.745 38.955 158.265 ;
        RECT 39.125 157.965 39.475 158.215 ;
        RECT 39.660 157.755 39.830 158.385 ;
        RECT 40.000 157.965 40.330 158.165 ;
        RECT 40.500 157.965 40.830 158.165 ;
        RECT 41.000 157.965 41.420 158.165 ;
        RECT 41.595 158.135 41.765 158.385 ;
        RECT 41.595 157.965 42.290 158.135 ;
        RECT 33.595 157.145 33.875 157.605 ;
        RECT 34.395 156.975 34.720 157.435 ;
        RECT 34.890 157.145 35.275 157.715 ;
        RECT 35.445 156.975 38.955 157.745 ;
        RECT 39.330 157.145 39.830 157.755 ;
        RECT 40.460 157.625 41.685 157.795 ;
        RECT 42.460 157.775 42.635 158.385 ;
        RECT 42.805 157.965 43.155 158.215 ;
        RECT 40.460 157.145 40.790 157.625 ;
        RECT 40.960 156.975 41.185 157.435 ;
        RECT 41.355 157.145 41.685 157.625 ;
        RECT 41.875 156.975 42.125 157.775 ;
        RECT 42.295 157.145 42.635 157.775 ;
        RECT 43.340 157.755 43.510 158.385 ;
        RECT 43.680 157.965 44.010 158.165 ;
        RECT 44.180 157.965 44.510 158.165 ;
        RECT 44.680 157.965 45.100 158.165 ;
        RECT 45.275 158.135 45.445 158.385 ;
        RECT 45.275 157.965 45.970 158.135 ;
        RECT 43.010 157.145 43.510 157.755 ;
        RECT 44.140 157.625 45.365 157.795 ;
        RECT 46.140 157.775 46.315 158.385 ;
        RECT 46.485 157.945 47.175 158.505 ;
        RECT 47.345 157.775 47.555 158.675 ;
        RECT 44.140 157.145 44.470 157.625 ;
        RECT 44.640 156.975 44.865 157.435 ;
        RECT 45.035 157.145 45.365 157.625 ;
        RECT 45.555 156.975 45.805 157.775 ;
        RECT 45.975 157.145 46.315 157.775 ;
        RECT 46.600 157.605 47.555 157.775 ;
        RECT 47.725 158.505 48.125 159.355 ;
        RECT 48.315 158.895 48.595 159.355 ;
        RECT 49.115 159.065 49.440 159.525 ;
        RECT 48.315 158.675 49.440 158.895 ;
        RECT 47.725 157.945 48.820 158.505 ;
        RECT 48.990 158.215 49.440 158.675 ;
        RECT 49.610 158.385 49.995 159.355 ;
        RECT 46.600 157.145 46.885 157.605 ;
        RECT 47.055 156.975 47.325 157.435 ;
        RECT 47.725 157.145 48.125 157.945 ;
        RECT 48.990 157.885 49.545 158.215 ;
        RECT 48.990 157.775 49.440 157.885 ;
        RECT 48.315 157.605 49.440 157.775 ;
        RECT 49.715 157.715 49.995 158.385 ;
        RECT 50.165 158.360 50.455 159.525 ;
        RECT 50.625 158.385 50.965 159.355 ;
        RECT 51.135 158.385 51.305 159.525 ;
        RECT 51.575 158.725 51.825 159.525 ;
        RECT 52.470 158.555 52.800 159.355 ;
        RECT 53.100 158.725 53.430 159.525 ;
        RECT 53.600 158.555 53.930 159.355 ;
        RECT 54.770 159.090 60.115 159.525 ;
        RECT 51.495 158.385 53.930 158.555 ;
        RECT 48.315 157.145 48.595 157.605 ;
        RECT 49.115 156.975 49.440 157.435 ;
        RECT 49.610 157.145 49.995 157.715 ;
        RECT 50.625 157.775 50.800 158.385 ;
        RECT 51.495 158.135 51.665 158.385 ;
        RECT 50.970 157.965 51.665 158.135 ;
        RECT 51.840 157.965 52.260 158.165 ;
        RECT 52.430 157.965 52.760 158.165 ;
        RECT 52.930 157.965 53.260 158.165 ;
        RECT 50.165 156.975 50.455 157.700 ;
        RECT 50.625 157.145 50.965 157.775 ;
        RECT 51.135 156.975 51.385 157.775 ;
        RECT 51.575 157.625 52.800 157.795 ;
        RECT 51.575 157.145 51.905 157.625 ;
        RECT 52.075 156.975 52.300 157.435 ;
        RECT 52.470 157.145 52.800 157.625 ;
        RECT 53.430 157.755 53.600 158.385 ;
        RECT 53.785 157.965 54.135 158.215 ;
        RECT 56.360 157.840 56.710 159.090 ;
        RECT 60.345 158.385 60.555 159.525 ;
        RECT 60.725 158.375 61.055 159.355 ;
        RECT 61.225 158.385 61.455 159.525 ;
        RECT 61.815 158.375 62.145 159.525 ;
        RECT 62.315 158.505 62.485 159.355 ;
        RECT 62.655 158.725 62.985 159.525 ;
        RECT 63.155 158.505 63.325 159.355 ;
        RECT 63.505 158.725 63.745 159.525 ;
        RECT 63.915 158.545 64.245 159.355 ;
        RECT 53.430 157.145 53.930 157.755 ;
        RECT 58.190 157.520 58.530 158.350 ;
        RECT 54.770 156.975 60.115 157.520 ;
        RECT 60.345 156.975 60.555 157.795 ;
        RECT 60.725 157.775 60.975 158.375 ;
        RECT 62.315 158.335 63.325 158.505 ;
        RECT 63.530 158.375 64.245 158.545 ;
        RECT 64.885 158.435 68.395 159.525 ;
        RECT 68.655 158.595 68.825 159.355 ;
        RECT 69.040 158.765 69.370 159.525 ;
        RECT 61.145 157.965 61.475 158.215 ;
        RECT 62.315 158.165 62.810 158.335 ;
        RECT 62.315 157.995 62.815 158.165 ;
        RECT 63.530 158.135 63.700 158.375 ;
        RECT 62.315 157.795 62.810 157.995 ;
        RECT 63.200 157.965 63.700 158.135 ;
        RECT 63.870 157.965 64.250 158.205 ;
        RECT 63.530 157.795 63.700 157.965 ;
        RECT 64.885 157.915 66.575 158.435 ;
        RECT 68.655 158.425 69.370 158.595 ;
        RECT 69.540 158.450 69.795 159.355 ;
        RECT 60.725 157.145 61.055 157.775 ;
        RECT 61.225 156.975 61.455 157.795 ;
        RECT 61.815 156.975 62.145 157.775 ;
        RECT 62.315 157.625 63.325 157.795 ;
        RECT 63.530 157.625 64.165 157.795 ;
        RECT 66.745 157.745 68.395 158.265 ;
        RECT 68.565 157.875 68.920 158.245 ;
        RECT 69.200 158.215 69.370 158.425 ;
        RECT 69.200 157.885 69.455 158.215 ;
        RECT 62.315 157.145 62.485 157.625 ;
        RECT 62.655 156.975 62.985 157.455 ;
        RECT 63.155 157.145 63.325 157.625 ;
        RECT 63.575 156.975 63.815 157.455 ;
        RECT 63.995 157.145 64.165 157.625 ;
        RECT 64.885 156.975 68.395 157.745 ;
        RECT 69.200 157.695 69.370 157.885 ;
        RECT 69.625 157.720 69.795 158.450 ;
        RECT 69.970 158.375 70.230 159.525 ;
        RECT 70.495 158.595 70.665 159.355 ;
        RECT 70.880 158.765 71.210 159.525 ;
        RECT 70.495 158.425 71.210 158.595 ;
        RECT 71.380 158.450 71.635 159.355 ;
        RECT 70.405 157.875 70.760 158.245 ;
        RECT 71.040 158.215 71.210 158.425 ;
        RECT 71.040 157.885 71.295 158.215 ;
        RECT 68.655 157.525 69.370 157.695 ;
        RECT 68.655 157.145 68.825 157.525 ;
        RECT 69.040 156.975 69.370 157.355 ;
        RECT 69.540 157.145 69.795 157.720 ;
        RECT 69.970 156.975 70.230 157.815 ;
        RECT 71.040 157.695 71.210 157.885 ;
        RECT 71.465 157.720 71.635 158.450 ;
        RECT 71.810 158.375 72.070 159.525 ;
        RECT 72.450 158.555 72.780 159.355 ;
        RECT 72.950 158.725 73.280 159.525 ;
        RECT 73.580 158.555 73.910 159.355 ;
        RECT 74.555 158.725 74.805 159.525 ;
        RECT 72.450 158.385 74.885 158.555 ;
        RECT 75.075 158.385 75.245 159.525 ;
        RECT 75.415 158.385 75.755 159.355 ;
        RECT 72.245 157.965 72.595 158.215 ;
        RECT 70.495 157.525 71.210 157.695 ;
        RECT 70.495 157.145 70.665 157.525 ;
        RECT 70.880 156.975 71.210 157.355 ;
        RECT 71.380 157.145 71.635 157.720 ;
        RECT 71.810 156.975 72.070 157.815 ;
        RECT 72.780 157.755 72.950 158.385 ;
        RECT 73.120 157.965 73.450 158.165 ;
        RECT 73.620 157.965 73.950 158.165 ;
        RECT 74.120 157.965 74.540 158.165 ;
        RECT 74.715 158.135 74.885 158.385 ;
        RECT 74.715 157.965 75.410 158.135 ;
        RECT 72.450 157.145 72.950 157.755 ;
        RECT 73.580 157.625 74.805 157.795 ;
        RECT 75.580 157.775 75.755 158.385 ;
        RECT 75.925 158.360 76.215 159.525 ;
        RECT 77.050 158.555 77.380 159.355 ;
        RECT 77.550 158.725 77.880 159.525 ;
        RECT 78.180 158.555 78.510 159.355 ;
        RECT 79.155 158.725 79.405 159.525 ;
        RECT 77.050 158.385 79.485 158.555 ;
        RECT 79.675 158.385 79.845 159.525 ;
        RECT 80.015 158.385 80.355 159.355 ;
        RECT 81.360 159.185 81.615 159.215 ;
        RECT 81.275 159.015 81.615 159.185 ;
        RECT 76.845 157.965 77.195 158.215 ;
        RECT 73.580 157.145 73.910 157.625 ;
        RECT 74.080 156.975 74.305 157.435 ;
        RECT 74.475 157.145 74.805 157.625 ;
        RECT 74.995 156.975 75.245 157.775 ;
        RECT 75.415 157.145 75.755 157.775 ;
        RECT 77.380 157.755 77.550 158.385 ;
        RECT 77.720 157.965 78.050 158.165 ;
        RECT 78.220 157.965 78.550 158.165 ;
        RECT 78.720 157.965 79.140 158.165 ;
        RECT 79.315 158.135 79.485 158.385 ;
        RECT 79.315 157.965 80.010 158.135 ;
        RECT 75.925 156.975 76.215 157.700 ;
        RECT 77.050 157.145 77.550 157.755 ;
        RECT 78.180 157.625 79.405 157.795 ;
        RECT 80.180 157.775 80.355 158.385 ;
        RECT 78.180 157.145 78.510 157.625 ;
        RECT 78.680 156.975 78.905 157.435 ;
        RECT 79.075 157.145 79.405 157.625 ;
        RECT 79.595 156.975 79.845 157.775 ;
        RECT 80.015 157.145 80.355 157.775 ;
        RECT 81.360 158.545 81.615 159.015 ;
        RECT 81.795 158.725 82.080 159.525 ;
        RECT 82.260 158.805 82.590 159.315 ;
        RECT 81.360 157.685 81.540 158.545 ;
        RECT 82.260 158.215 82.510 158.805 ;
        RECT 82.860 158.655 83.030 159.265 ;
        RECT 83.200 158.835 83.530 159.525 ;
        RECT 83.760 158.975 84.000 159.265 ;
        RECT 84.200 159.145 84.620 159.525 ;
        RECT 84.800 159.055 85.430 159.305 ;
        RECT 85.900 159.145 86.230 159.525 ;
        RECT 84.800 158.975 84.970 159.055 ;
        RECT 86.400 158.975 86.570 159.265 ;
        RECT 86.750 159.145 87.130 159.525 ;
        RECT 87.370 159.140 88.200 159.310 ;
        RECT 83.760 158.805 84.970 158.975 ;
        RECT 81.710 157.885 82.510 158.215 ;
        RECT 81.360 157.155 81.615 157.685 ;
        RECT 81.795 156.975 82.080 157.435 ;
        RECT 82.260 157.235 82.510 157.885 ;
        RECT 82.710 158.635 83.030 158.655 ;
        RECT 82.710 158.465 84.630 158.635 ;
        RECT 82.710 157.570 82.900 158.465 ;
        RECT 84.800 158.295 84.970 158.805 ;
        RECT 85.140 158.545 85.660 158.855 ;
        RECT 83.070 158.125 84.970 158.295 ;
        RECT 83.070 158.065 83.400 158.125 ;
        RECT 83.550 157.895 83.880 157.955 ;
        RECT 83.220 157.625 83.880 157.895 ;
        RECT 82.710 157.240 83.030 157.570 ;
        RECT 83.210 156.975 83.870 157.455 ;
        RECT 84.070 157.365 84.240 158.125 ;
        RECT 85.140 157.955 85.320 158.365 ;
        RECT 84.410 157.785 84.740 157.905 ;
        RECT 85.490 157.785 85.660 158.545 ;
        RECT 84.410 157.615 85.660 157.785 ;
        RECT 85.830 158.725 87.200 158.975 ;
        RECT 85.830 157.955 86.020 158.725 ;
        RECT 86.950 158.465 87.200 158.725 ;
        RECT 86.190 158.295 86.440 158.455 ;
        RECT 87.370 158.295 87.540 159.140 ;
        RECT 88.435 158.855 88.605 159.355 ;
        RECT 88.775 159.025 89.105 159.525 ;
        RECT 87.710 158.465 88.210 158.845 ;
        RECT 88.435 158.685 89.130 158.855 ;
        RECT 86.190 158.125 87.540 158.295 ;
        RECT 87.120 158.085 87.540 158.125 ;
        RECT 85.830 157.615 86.250 157.955 ;
        RECT 86.540 157.625 86.950 157.955 ;
        RECT 84.070 157.195 84.920 157.365 ;
        RECT 85.480 156.975 85.800 157.435 ;
        RECT 86.000 157.185 86.250 157.615 ;
        RECT 86.540 156.975 86.950 157.415 ;
        RECT 87.120 157.355 87.290 158.085 ;
        RECT 87.460 157.535 87.810 157.905 ;
        RECT 87.990 157.595 88.210 158.465 ;
        RECT 88.380 157.895 88.790 158.515 ;
        RECT 88.960 157.715 89.130 158.685 ;
        RECT 88.435 157.525 89.130 157.715 ;
        RECT 87.120 157.155 88.135 157.355 ;
        RECT 88.435 157.195 88.605 157.525 ;
        RECT 88.775 156.975 89.105 157.355 ;
        RECT 89.320 157.235 89.545 159.355 ;
        RECT 89.715 159.025 90.045 159.525 ;
        RECT 90.215 158.855 90.385 159.355 ;
        RECT 89.720 158.685 90.385 158.855 ;
        RECT 89.720 157.695 89.950 158.685 ;
        RECT 90.120 157.865 90.470 158.515 ;
        RECT 91.105 158.435 92.775 159.525 ;
        RECT 91.105 157.915 91.855 158.435 ;
        RECT 92.985 158.385 93.215 159.525 ;
        RECT 93.385 158.375 93.715 159.355 ;
        RECT 93.885 158.385 94.095 159.525 ;
        RECT 94.785 158.435 96.455 159.525 ;
        RECT 96.715 158.595 96.885 159.355 ;
        RECT 97.065 158.765 97.395 159.525 ;
        RECT 92.025 157.745 92.775 158.265 ;
        RECT 92.965 157.965 93.295 158.215 ;
        RECT 89.720 157.525 90.385 157.695 ;
        RECT 89.715 156.975 90.045 157.355 ;
        RECT 90.215 157.235 90.385 157.525 ;
        RECT 91.105 156.975 92.775 157.745 ;
        RECT 92.985 156.975 93.215 157.795 ;
        RECT 93.465 157.775 93.715 158.375 ;
        RECT 94.785 157.915 95.535 158.435 ;
        RECT 96.715 158.425 97.380 158.595 ;
        RECT 97.565 158.450 97.835 159.355 ;
        RECT 97.210 158.280 97.380 158.425 ;
        RECT 93.385 157.145 93.715 157.775 ;
        RECT 93.885 156.975 94.095 157.795 ;
        RECT 95.705 157.745 96.455 158.265 ;
        RECT 96.645 157.875 96.975 158.245 ;
        RECT 97.210 157.950 97.495 158.280 ;
        RECT 94.785 156.975 96.455 157.745 ;
        RECT 97.210 157.695 97.380 157.950 ;
        RECT 96.715 157.525 97.380 157.695 ;
        RECT 97.665 157.650 97.835 158.450 ;
        RECT 98.005 158.435 99.675 159.525 ;
        RECT 98.005 157.915 98.755 158.435 ;
        RECT 99.885 158.385 100.115 159.525 ;
        RECT 100.285 158.375 100.615 159.355 ;
        RECT 100.785 158.385 100.995 159.525 ;
        RECT 98.925 157.745 99.675 158.265 ;
        RECT 99.865 157.965 100.195 158.215 ;
        RECT 96.715 157.145 96.885 157.525 ;
        RECT 97.065 156.975 97.395 157.355 ;
        RECT 97.575 157.145 97.835 157.650 ;
        RECT 98.005 156.975 99.675 157.745 ;
        RECT 99.885 156.975 100.115 157.795 ;
        RECT 100.365 157.775 100.615 158.375 ;
        RECT 101.685 158.360 101.975 159.525 ;
        RECT 102.605 158.435 104.275 159.525 ;
        RECT 104.445 158.450 104.715 159.355 ;
        RECT 104.885 158.765 105.215 159.525 ;
        RECT 105.395 158.595 105.565 159.355 ;
        RECT 102.605 157.915 103.355 158.435 ;
        RECT 100.285 157.145 100.615 157.775 ;
        RECT 100.785 156.975 100.995 157.795 ;
        RECT 103.525 157.745 104.275 158.265 ;
        RECT 101.685 156.975 101.975 157.700 ;
        RECT 102.605 156.975 104.275 157.745 ;
        RECT 104.445 157.650 104.615 158.450 ;
        RECT 104.900 158.425 105.565 158.595 ;
        RECT 105.915 158.595 106.085 159.355 ;
        RECT 106.265 158.765 106.595 159.525 ;
        RECT 105.915 158.425 106.580 158.595 ;
        RECT 106.765 158.450 107.035 159.355 ;
        RECT 104.900 158.280 105.070 158.425 ;
        RECT 104.785 157.950 105.070 158.280 ;
        RECT 106.410 158.280 106.580 158.425 ;
        RECT 104.900 157.695 105.070 157.950 ;
        RECT 105.305 157.875 105.635 158.245 ;
        RECT 105.845 157.875 106.175 158.245 ;
        RECT 106.410 157.950 106.695 158.280 ;
        RECT 106.410 157.695 106.580 157.950 ;
        RECT 104.445 157.145 104.705 157.650 ;
        RECT 104.900 157.525 105.565 157.695 ;
        RECT 104.885 156.975 105.215 157.355 ;
        RECT 105.395 157.145 105.565 157.525 ;
        RECT 105.915 157.525 106.580 157.695 ;
        RECT 106.865 157.650 107.035 158.450 ;
        RECT 105.915 157.145 106.085 157.525 ;
        RECT 106.265 156.975 106.595 157.355 ;
        RECT 106.775 157.145 107.035 157.650 ;
        RECT 108.125 158.385 108.465 159.355 ;
        RECT 108.635 158.385 108.805 159.525 ;
        RECT 109.075 158.725 109.325 159.525 ;
        RECT 109.970 158.555 110.300 159.355 ;
        RECT 110.600 158.725 110.930 159.525 ;
        RECT 111.100 158.555 111.430 159.355 ;
        RECT 108.995 158.385 111.430 158.555 ;
        RECT 112.725 158.435 116.235 159.525 ;
        RECT 116.520 158.895 116.805 159.355 ;
        RECT 116.975 159.065 117.245 159.525 ;
        RECT 116.520 158.675 117.475 158.895 ;
        RECT 108.125 157.775 108.300 158.385 ;
        RECT 108.995 158.135 109.165 158.385 ;
        RECT 108.470 157.965 109.165 158.135 ;
        RECT 109.340 157.965 109.760 158.165 ;
        RECT 109.930 157.965 110.260 158.165 ;
        RECT 110.430 157.965 110.760 158.165 ;
        RECT 108.125 157.145 108.465 157.775 ;
        RECT 108.635 156.975 108.885 157.775 ;
        RECT 109.075 157.625 110.300 157.795 ;
        RECT 109.075 157.145 109.405 157.625 ;
        RECT 109.575 156.975 109.800 157.435 ;
        RECT 109.970 157.145 110.300 157.625 ;
        RECT 110.930 157.755 111.100 158.385 ;
        RECT 111.285 157.965 111.635 158.215 ;
        RECT 112.725 157.915 114.415 158.435 ;
        RECT 110.930 157.145 111.430 157.755 ;
        RECT 114.585 157.745 116.235 158.265 ;
        RECT 116.405 157.945 117.095 158.505 ;
        RECT 117.265 157.775 117.475 158.675 ;
        RECT 112.725 156.975 116.235 157.745 ;
        RECT 116.520 157.605 117.475 157.775 ;
        RECT 117.645 158.505 118.045 159.355 ;
        RECT 118.235 158.895 118.515 159.355 ;
        RECT 119.035 159.065 119.360 159.525 ;
        RECT 118.235 158.675 119.360 158.895 ;
        RECT 117.645 157.945 118.740 158.505 ;
        RECT 118.910 158.215 119.360 158.675 ;
        RECT 119.530 158.385 119.915 159.355 ;
        RECT 121.010 159.090 126.355 159.525 ;
        RECT 116.520 157.145 116.805 157.605 ;
        RECT 116.975 156.975 117.245 157.435 ;
        RECT 117.645 157.145 118.045 157.945 ;
        RECT 118.910 157.885 119.465 158.215 ;
        RECT 118.910 157.775 119.360 157.885 ;
        RECT 118.235 157.605 119.360 157.775 ;
        RECT 119.635 157.715 119.915 158.385 ;
        RECT 122.600 157.840 122.950 159.090 ;
        RECT 126.525 158.435 127.735 159.525 ;
        RECT 118.235 157.145 118.515 157.605 ;
        RECT 119.035 156.975 119.360 157.435 ;
        RECT 119.530 157.145 119.915 157.715 ;
        RECT 124.430 157.520 124.770 158.350 ;
        RECT 126.525 157.895 127.045 158.435 ;
        RECT 127.215 157.725 127.735 158.265 ;
        RECT 121.010 156.975 126.355 157.520 ;
        RECT 126.525 156.975 127.735 157.725 ;
        RECT 14.660 156.805 127.820 156.975 ;
        RECT 14.745 156.055 15.955 156.805 ;
        RECT 17.420 156.465 17.675 156.625 ;
        RECT 17.335 156.295 17.675 156.465 ;
        RECT 17.855 156.345 18.140 156.805 ;
        RECT 17.420 156.095 17.675 156.295 ;
        RECT 14.745 155.515 15.265 156.055 ;
        RECT 15.435 155.345 15.955 155.885 ;
        RECT 14.745 154.255 15.955 155.345 ;
        RECT 17.420 155.235 17.600 156.095 ;
        RECT 18.320 155.895 18.570 156.545 ;
        RECT 17.770 155.565 18.570 155.895 ;
        RECT 17.420 154.565 17.675 155.235 ;
        RECT 17.855 154.255 18.140 155.055 ;
        RECT 18.320 154.975 18.570 155.565 ;
        RECT 18.770 156.210 19.090 156.540 ;
        RECT 19.270 156.325 19.930 156.805 ;
        RECT 20.130 156.415 20.980 156.585 ;
        RECT 18.770 155.315 18.960 156.210 ;
        RECT 19.280 155.885 19.940 156.155 ;
        RECT 19.610 155.825 19.940 155.885 ;
        RECT 19.130 155.655 19.460 155.715 ;
        RECT 20.130 155.655 20.300 156.415 ;
        RECT 21.540 156.345 21.860 156.805 ;
        RECT 22.060 156.165 22.310 156.595 ;
        RECT 22.600 156.365 23.010 156.805 ;
        RECT 23.180 156.425 24.195 156.625 ;
        RECT 20.470 155.995 21.720 156.165 ;
        RECT 20.470 155.875 20.800 155.995 ;
        RECT 19.130 155.485 21.030 155.655 ;
        RECT 18.770 155.145 20.690 155.315 ;
        RECT 18.770 155.125 19.090 155.145 ;
        RECT 18.320 154.465 18.650 154.975 ;
        RECT 18.920 154.515 19.090 155.125 ;
        RECT 20.860 154.975 21.030 155.485 ;
        RECT 21.200 155.415 21.380 155.825 ;
        RECT 21.550 155.235 21.720 155.995 ;
        RECT 19.260 154.255 19.590 154.945 ;
        RECT 19.820 154.805 21.030 154.975 ;
        RECT 21.200 154.925 21.720 155.235 ;
        RECT 21.890 155.825 22.310 156.165 ;
        RECT 22.600 155.825 23.010 156.155 ;
        RECT 21.890 155.055 22.080 155.825 ;
        RECT 23.180 155.695 23.350 156.425 ;
        RECT 24.495 156.255 24.665 156.585 ;
        RECT 24.835 156.425 25.165 156.805 ;
        RECT 23.520 155.875 23.870 156.245 ;
        RECT 23.180 155.655 23.600 155.695 ;
        RECT 22.250 155.485 23.600 155.655 ;
        RECT 22.250 155.325 22.500 155.485 ;
        RECT 23.010 155.055 23.260 155.315 ;
        RECT 21.890 154.805 23.260 155.055 ;
        RECT 19.820 154.515 20.060 154.805 ;
        RECT 20.860 154.725 21.030 154.805 ;
        RECT 20.260 154.255 20.680 154.635 ;
        RECT 20.860 154.475 21.490 154.725 ;
        RECT 21.960 154.255 22.290 154.635 ;
        RECT 22.460 154.515 22.630 154.805 ;
        RECT 23.430 154.640 23.600 155.485 ;
        RECT 24.050 155.315 24.270 156.185 ;
        RECT 24.495 156.065 25.190 156.255 ;
        RECT 23.770 154.935 24.270 155.315 ;
        RECT 24.440 155.265 24.850 155.885 ;
        RECT 25.020 155.095 25.190 156.065 ;
        RECT 24.495 154.925 25.190 155.095 ;
        RECT 22.810 154.255 23.190 154.635 ;
        RECT 23.430 154.470 24.260 154.640 ;
        RECT 24.495 154.425 24.665 154.925 ;
        RECT 24.835 154.255 25.165 154.755 ;
        RECT 25.380 154.425 25.605 156.545 ;
        RECT 25.775 156.425 26.105 156.805 ;
        RECT 26.275 156.255 26.445 156.545 ;
        RECT 25.780 156.085 26.445 156.255 ;
        RECT 26.705 156.130 26.965 156.635 ;
        RECT 27.145 156.425 27.475 156.805 ;
        RECT 27.655 156.255 27.825 156.635 ;
        RECT 25.780 155.095 26.010 156.085 ;
        RECT 26.180 155.265 26.530 155.915 ;
        RECT 26.705 155.330 26.875 156.130 ;
        RECT 27.160 156.085 27.825 156.255 ;
        RECT 27.160 155.830 27.330 156.085 ;
        RECT 28.085 156.055 29.295 156.805 ;
        RECT 27.045 155.500 27.330 155.830 ;
        RECT 27.565 155.535 27.895 155.905 ;
        RECT 27.160 155.355 27.330 155.500 ;
        RECT 25.780 154.925 26.445 155.095 ;
        RECT 25.775 154.255 26.105 154.755 ;
        RECT 26.275 154.425 26.445 154.925 ;
        RECT 26.705 154.425 26.975 155.330 ;
        RECT 27.160 155.185 27.825 155.355 ;
        RECT 27.145 154.255 27.475 155.015 ;
        RECT 27.655 154.425 27.825 155.185 ;
        RECT 28.085 155.345 28.605 155.885 ;
        RECT 28.775 155.515 29.295 156.055 ;
        RECT 29.465 156.035 32.975 156.805 ;
        RECT 29.465 155.345 31.155 155.865 ;
        RECT 31.325 155.515 32.975 156.035 ;
        RECT 33.420 155.995 33.665 156.600 ;
        RECT 33.885 156.270 34.395 156.805 ;
        RECT 33.145 155.825 34.375 155.995 ;
        RECT 28.085 154.255 29.295 155.345 ;
        RECT 29.465 154.255 32.975 155.345 ;
        RECT 33.145 155.015 33.485 155.825 ;
        RECT 33.655 155.260 34.405 155.450 ;
        RECT 33.145 154.605 33.660 155.015 ;
        RECT 33.895 154.255 34.065 155.015 ;
        RECT 34.235 154.595 34.405 155.260 ;
        RECT 34.575 155.275 34.765 156.635 ;
        RECT 34.935 156.465 35.210 156.635 ;
        RECT 34.935 156.295 35.215 156.465 ;
        RECT 34.935 155.475 35.210 156.295 ;
        RECT 35.400 156.270 35.930 156.635 ;
        RECT 36.355 156.405 36.685 156.805 ;
        RECT 35.755 156.235 35.930 156.270 ;
        RECT 35.415 155.275 35.585 156.075 ;
        RECT 34.575 155.105 35.585 155.275 ;
        RECT 35.755 156.065 36.685 156.235 ;
        RECT 36.855 156.065 37.110 156.635 ;
        RECT 37.285 156.080 37.575 156.805 ;
        RECT 35.755 154.935 35.925 156.065 ;
        RECT 36.515 155.895 36.685 156.065 ;
        RECT 34.800 154.765 35.925 154.935 ;
        RECT 36.095 155.565 36.290 155.895 ;
        RECT 36.515 155.565 36.770 155.895 ;
        RECT 36.095 154.595 36.265 155.565 ;
        RECT 36.940 155.395 37.110 156.065 ;
        RECT 38.205 156.035 39.875 156.805 ;
        RECT 34.235 154.425 36.265 154.595 ;
        RECT 36.435 154.255 36.605 155.395 ;
        RECT 36.775 154.425 37.110 155.395 ;
        RECT 37.285 154.255 37.575 155.420 ;
        RECT 38.205 155.345 38.955 155.865 ;
        RECT 39.125 155.515 39.875 156.035 ;
        RECT 40.045 156.005 40.385 156.635 ;
        RECT 40.555 156.005 40.805 156.805 ;
        RECT 40.995 156.155 41.325 156.635 ;
        RECT 41.495 156.345 41.720 156.805 ;
        RECT 41.890 156.155 42.220 156.635 ;
        RECT 40.045 155.395 40.220 156.005 ;
        RECT 40.995 155.985 42.220 156.155 ;
        RECT 42.850 156.025 43.350 156.635 ;
        RECT 40.390 155.645 41.085 155.815 ;
        RECT 40.915 155.395 41.085 155.645 ;
        RECT 41.260 155.615 41.680 155.815 ;
        RECT 41.850 155.615 42.180 155.815 ;
        RECT 42.350 155.615 42.680 155.815 ;
        RECT 42.850 155.395 43.020 156.025 ;
        RECT 43.725 156.005 44.065 156.635 ;
        RECT 44.235 156.005 44.485 156.805 ;
        RECT 44.675 156.155 45.005 156.635 ;
        RECT 45.175 156.345 45.400 156.805 ;
        RECT 45.570 156.155 45.900 156.635 ;
        RECT 43.205 155.565 43.555 155.815 ;
        RECT 43.725 155.395 43.900 156.005 ;
        RECT 44.675 155.985 45.900 156.155 ;
        RECT 46.530 156.025 47.030 156.635 ;
        RECT 44.070 155.645 44.765 155.815 ;
        RECT 44.595 155.395 44.765 155.645 ;
        RECT 44.940 155.615 45.360 155.815 ;
        RECT 45.530 155.615 45.860 155.815 ;
        RECT 46.030 155.615 46.360 155.815 ;
        RECT 46.530 155.395 46.700 156.025 ;
        RECT 47.405 156.005 47.745 156.635 ;
        RECT 47.915 156.005 48.165 156.805 ;
        RECT 48.355 156.155 48.685 156.635 ;
        RECT 48.855 156.345 49.080 156.805 ;
        RECT 49.250 156.155 49.580 156.635 ;
        RECT 46.885 155.565 47.235 155.815 ;
        RECT 47.405 155.395 47.580 156.005 ;
        RECT 48.355 155.985 49.580 156.155 ;
        RECT 50.210 156.025 50.710 156.635 ;
        RECT 51.545 156.035 53.215 156.805 ;
        RECT 47.750 155.645 48.445 155.815 ;
        RECT 48.275 155.395 48.445 155.645 ;
        RECT 48.620 155.615 49.040 155.815 ;
        RECT 49.210 155.615 49.540 155.815 ;
        RECT 49.710 155.615 50.040 155.815 ;
        RECT 50.210 155.395 50.380 156.025 ;
        RECT 50.565 155.565 50.915 155.815 ;
        RECT 38.205 154.255 39.875 155.345 ;
        RECT 40.045 154.425 40.385 155.395 ;
        RECT 40.555 154.255 40.725 155.395 ;
        RECT 40.915 155.225 43.350 155.395 ;
        RECT 40.995 154.255 41.245 155.055 ;
        RECT 41.890 154.425 42.220 155.225 ;
        RECT 42.520 154.255 42.850 155.055 ;
        RECT 43.020 154.425 43.350 155.225 ;
        RECT 43.725 154.425 44.065 155.395 ;
        RECT 44.235 154.255 44.405 155.395 ;
        RECT 44.595 155.225 47.030 155.395 ;
        RECT 44.675 154.255 44.925 155.055 ;
        RECT 45.570 154.425 45.900 155.225 ;
        RECT 46.200 154.255 46.530 155.055 ;
        RECT 46.700 154.425 47.030 155.225 ;
        RECT 47.405 154.425 47.745 155.395 ;
        RECT 47.915 154.255 48.085 155.395 ;
        RECT 48.275 155.225 50.710 155.395 ;
        RECT 48.355 154.255 48.605 155.055 ;
        RECT 49.250 154.425 49.580 155.225 ;
        RECT 49.880 154.255 50.210 155.055 ;
        RECT 50.380 154.425 50.710 155.225 ;
        RECT 51.545 155.345 52.295 155.865 ;
        RECT 52.465 155.515 53.215 156.035 ;
        RECT 53.760 156.095 54.015 156.625 ;
        RECT 54.195 156.345 54.480 156.805 ;
        RECT 51.545 154.255 53.215 155.345 ;
        RECT 53.760 155.235 53.940 156.095 ;
        RECT 54.660 155.895 54.910 156.545 ;
        RECT 54.110 155.565 54.910 155.895 ;
        RECT 53.760 154.765 54.015 155.235 ;
        RECT 53.675 154.595 54.015 154.765 ;
        RECT 53.760 154.565 54.015 154.595 ;
        RECT 54.195 154.255 54.480 155.055 ;
        RECT 54.660 154.975 54.910 155.565 ;
        RECT 55.110 156.210 55.430 156.540 ;
        RECT 55.610 156.325 56.270 156.805 ;
        RECT 56.470 156.415 57.320 156.585 ;
        RECT 55.110 155.315 55.300 156.210 ;
        RECT 55.620 155.885 56.280 156.155 ;
        RECT 55.950 155.825 56.280 155.885 ;
        RECT 55.470 155.655 55.800 155.715 ;
        RECT 56.470 155.655 56.640 156.415 ;
        RECT 57.880 156.345 58.200 156.805 ;
        RECT 58.400 156.165 58.650 156.595 ;
        RECT 58.940 156.365 59.350 156.805 ;
        RECT 59.520 156.425 60.535 156.625 ;
        RECT 56.810 155.995 58.060 156.165 ;
        RECT 56.810 155.875 57.140 155.995 ;
        RECT 55.470 155.485 57.370 155.655 ;
        RECT 55.110 155.145 57.030 155.315 ;
        RECT 55.110 155.125 55.430 155.145 ;
        RECT 54.660 154.465 54.990 154.975 ;
        RECT 55.260 154.515 55.430 155.125 ;
        RECT 57.200 154.975 57.370 155.485 ;
        RECT 57.540 155.415 57.720 155.825 ;
        RECT 57.890 155.235 58.060 155.995 ;
        RECT 55.600 154.255 55.930 154.945 ;
        RECT 56.160 154.805 57.370 154.975 ;
        RECT 57.540 154.925 58.060 155.235 ;
        RECT 58.230 155.825 58.650 156.165 ;
        RECT 58.940 155.825 59.350 156.155 ;
        RECT 58.230 155.055 58.420 155.825 ;
        RECT 59.520 155.695 59.690 156.425 ;
        RECT 60.835 156.255 61.005 156.585 ;
        RECT 61.175 156.425 61.505 156.805 ;
        RECT 59.860 155.875 60.210 156.245 ;
        RECT 59.520 155.655 59.940 155.695 ;
        RECT 58.590 155.485 59.940 155.655 ;
        RECT 58.590 155.325 58.840 155.485 ;
        RECT 59.350 155.055 59.600 155.315 ;
        RECT 58.230 154.805 59.600 155.055 ;
        RECT 56.160 154.515 56.400 154.805 ;
        RECT 57.200 154.725 57.370 154.805 ;
        RECT 56.600 154.255 57.020 154.635 ;
        RECT 57.200 154.475 57.830 154.725 ;
        RECT 58.300 154.255 58.630 154.635 ;
        RECT 58.800 154.515 58.970 154.805 ;
        RECT 59.770 154.640 59.940 155.485 ;
        RECT 60.390 155.315 60.610 156.185 ;
        RECT 60.835 156.065 61.530 156.255 ;
        RECT 60.110 154.935 60.610 155.315 ;
        RECT 60.780 155.265 61.190 155.885 ;
        RECT 61.360 155.095 61.530 156.065 ;
        RECT 60.835 154.925 61.530 155.095 ;
        RECT 59.150 154.255 59.530 154.635 ;
        RECT 59.770 154.470 60.600 154.640 ;
        RECT 60.835 154.425 61.005 154.925 ;
        RECT 61.175 154.255 61.505 154.755 ;
        RECT 61.720 154.425 61.945 156.545 ;
        RECT 62.115 156.425 62.445 156.805 ;
        RECT 62.615 156.255 62.785 156.545 ;
        RECT 62.120 156.085 62.785 156.255 ;
        RECT 62.120 155.095 62.350 156.085 ;
        RECT 63.045 156.080 63.335 156.805 ;
        RECT 63.965 156.035 65.635 156.805 ;
        RECT 65.895 156.325 66.195 156.805 ;
        RECT 66.365 156.155 66.625 156.610 ;
        RECT 66.795 156.325 67.055 156.805 ;
        RECT 67.235 156.155 67.495 156.610 ;
        RECT 67.665 156.325 67.915 156.805 ;
        RECT 68.095 156.155 68.355 156.610 ;
        RECT 68.525 156.325 68.775 156.805 ;
        RECT 68.955 156.155 69.215 156.610 ;
        RECT 69.385 156.325 69.630 156.805 ;
        RECT 69.800 156.155 70.075 156.610 ;
        RECT 70.245 156.325 70.490 156.805 ;
        RECT 70.660 156.155 70.920 156.610 ;
        RECT 71.090 156.325 71.350 156.805 ;
        RECT 71.520 156.155 71.780 156.610 ;
        RECT 71.950 156.325 72.210 156.805 ;
        RECT 72.380 156.155 72.640 156.610 ;
        RECT 72.810 156.245 73.070 156.805 ;
        RECT 62.520 155.265 62.870 155.915 ;
        RECT 62.120 154.925 62.785 155.095 ;
        RECT 62.115 154.255 62.445 154.755 ;
        RECT 62.615 154.425 62.785 154.925 ;
        RECT 63.045 154.255 63.335 155.420 ;
        RECT 63.965 155.345 64.715 155.865 ;
        RECT 64.885 155.515 65.635 156.035 ;
        RECT 65.895 155.985 72.640 156.155 ;
        RECT 65.895 155.445 67.060 155.985 ;
        RECT 73.240 155.815 73.490 156.625 ;
        RECT 73.670 156.280 73.930 156.805 ;
        RECT 74.100 155.815 74.350 156.625 ;
        RECT 74.530 156.295 74.835 156.805 ;
        RECT 67.230 155.565 74.350 155.815 ;
        RECT 74.520 155.565 74.835 156.125 ;
        RECT 75.005 156.035 76.675 156.805 ;
        RECT 65.865 155.395 67.060 155.445 ;
        RECT 63.965 154.255 65.635 155.345 ;
        RECT 65.865 155.275 72.640 155.395 ;
        RECT 65.895 155.170 72.640 155.275 ;
        RECT 65.895 154.255 66.165 155.000 ;
        RECT 66.335 154.430 66.625 155.170 ;
        RECT 67.235 155.155 72.640 155.170 ;
        RECT 66.795 154.260 67.050 154.985 ;
        RECT 67.235 154.430 67.495 155.155 ;
        RECT 67.665 154.260 67.910 154.985 ;
        RECT 68.095 154.430 68.355 155.155 ;
        RECT 68.525 154.260 68.770 154.985 ;
        RECT 68.955 154.430 69.215 155.155 ;
        RECT 69.385 154.260 69.630 154.985 ;
        RECT 69.800 154.430 70.060 155.155 ;
        RECT 70.230 154.260 70.490 154.985 ;
        RECT 70.660 154.430 70.920 155.155 ;
        RECT 71.090 154.260 71.350 154.985 ;
        RECT 71.520 154.430 71.780 155.155 ;
        RECT 71.950 154.260 72.210 154.985 ;
        RECT 72.380 154.430 72.640 155.155 ;
        RECT 72.810 154.260 73.070 155.055 ;
        RECT 73.240 154.430 73.490 155.565 ;
        RECT 66.795 154.255 73.070 154.260 ;
        RECT 73.670 154.255 73.930 155.065 ;
        RECT 74.105 154.425 74.350 155.565 ;
        RECT 75.005 155.345 75.755 155.865 ;
        RECT 75.925 155.515 76.675 156.035 ;
        RECT 76.845 156.005 77.185 156.635 ;
        RECT 77.355 156.005 77.605 156.805 ;
        RECT 77.795 156.155 78.125 156.635 ;
        RECT 78.295 156.345 78.520 156.805 ;
        RECT 78.690 156.155 79.020 156.635 ;
        RECT 76.845 155.395 77.020 156.005 ;
        RECT 77.795 155.985 79.020 156.155 ;
        RECT 79.650 156.025 80.150 156.635 ;
        RECT 77.190 155.645 77.885 155.815 ;
        RECT 77.715 155.395 77.885 155.645 ;
        RECT 78.060 155.615 78.480 155.815 ;
        RECT 78.650 155.615 78.980 155.815 ;
        RECT 79.150 155.615 79.480 155.815 ;
        RECT 79.650 155.395 79.820 156.025 ;
        RECT 80.525 156.005 80.865 156.635 ;
        RECT 81.035 156.005 81.285 156.805 ;
        RECT 81.475 156.155 81.805 156.635 ;
        RECT 81.975 156.345 82.200 156.805 ;
        RECT 82.370 156.155 82.700 156.635 ;
        RECT 80.005 155.565 80.355 155.815 ;
        RECT 80.525 155.395 80.700 156.005 ;
        RECT 81.475 155.985 82.700 156.155 ;
        RECT 83.330 156.025 83.830 156.635 ;
        RECT 85.125 156.035 88.635 156.805 ;
        RECT 88.805 156.080 89.095 156.805 ;
        RECT 89.265 156.035 91.855 156.805 ;
        RECT 92.030 156.260 97.375 156.805 ;
        RECT 80.870 155.645 81.565 155.815 ;
        RECT 81.395 155.395 81.565 155.645 ;
        RECT 81.740 155.615 82.160 155.815 ;
        RECT 82.330 155.615 82.660 155.815 ;
        RECT 82.830 155.615 83.160 155.815 ;
        RECT 83.330 155.395 83.500 156.025 ;
        RECT 83.685 155.565 84.035 155.815 ;
        RECT 74.530 154.255 74.825 155.065 ;
        RECT 75.005 154.255 76.675 155.345 ;
        RECT 76.845 154.425 77.185 155.395 ;
        RECT 77.355 154.255 77.525 155.395 ;
        RECT 77.715 155.225 80.150 155.395 ;
        RECT 77.795 154.255 78.045 155.055 ;
        RECT 78.690 154.425 79.020 155.225 ;
        RECT 79.320 154.255 79.650 155.055 ;
        RECT 79.820 154.425 80.150 155.225 ;
        RECT 80.525 154.425 80.865 155.395 ;
        RECT 81.035 154.255 81.205 155.395 ;
        RECT 81.395 155.225 83.830 155.395 ;
        RECT 81.475 154.255 81.725 155.055 ;
        RECT 82.370 154.425 82.700 155.225 ;
        RECT 83.000 154.255 83.330 155.055 ;
        RECT 83.500 154.425 83.830 155.225 ;
        RECT 85.125 155.345 86.815 155.865 ;
        RECT 86.985 155.515 88.635 156.035 ;
        RECT 85.125 154.255 88.635 155.345 ;
        RECT 88.805 154.255 89.095 155.420 ;
        RECT 89.265 155.345 90.475 155.865 ;
        RECT 90.645 155.515 91.855 156.035 ;
        RECT 89.265 154.255 91.855 155.345 ;
        RECT 93.620 154.690 93.970 155.940 ;
        RECT 95.450 155.430 95.790 156.260 ;
        RECT 97.750 156.025 98.250 156.635 ;
        RECT 97.545 155.565 97.895 155.815 ;
        RECT 98.080 155.395 98.250 156.025 ;
        RECT 98.880 156.155 99.210 156.635 ;
        RECT 99.380 156.345 99.605 156.805 ;
        RECT 99.775 156.155 100.105 156.635 ;
        RECT 98.880 155.985 100.105 156.155 ;
        RECT 100.295 156.005 100.545 156.805 ;
        RECT 100.715 156.005 101.055 156.635 ;
        RECT 101.685 156.035 103.355 156.805 ;
        RECT 98.420 155.615 98.750 155.815 ;
        RECT 98.920 155.615 99.250 155.815 ;
        RECT 99.420 155.615 99.840 155.815 ;
        RECT 100.015 155.645 100.710 155.815 ;
        RECT 100.015 155.395 100.185 155.645 ;
        RECT 100.880 155.395 101.055 156.005 ;
        RECT 97.750 155.225 100.185 155.395 ;
        RECT 92.030 154.255 97.375 154.690 ;
        RECT 97.750 154.425 98.080 155.225 ;
        RECT 98.250 154.255 98.580 155.055 ;
        RECT 98.880 154.425 99.210 155.225 ;
        RECT 99.855 154.255 100.105 155.055 ;
        RECT 100.375 154.255 100.545 155.395 ;
        RECT 100.715 154.425 101.055 155.395 ;
        RECT 101.685 155.345 102.435 155.865 ;
        RECT 102.605 155.515 103.355 156.035 ;
        RECT 103.525 156.005 103.865 156.635 ;
        RECT 104.035 156.005 104.285 156.805 ;
        RECT 104.475 156.155 104.805 156.635 ;
        RECT 104.975 156.345 105.200 156.805 ;
        RECT 105.370 156.155 105.700 156.635 ;
        RECT 103.525 155.395 103.700 156.005 ;
        RECT 104.475 155.985 105.700 156.155 ;
        RECT 106.330 156.025 106.830 156.635 ;
        RECT 107.410 156.025 107.910 156.635 ;
        RECT 103.870 155.645 104.565 155.815 ;
        RECT 104.395 155.395 104.565 155.645 ;
        RECT 104.740 155.615 105.160 155.815 ;
        RECT 105.330 155.615 105.660 155.815 ;
        RECT 105.830 155.615 106.160 155.815 ;
        RECT 106.330 155.395 106.500 156.025 ;
        RECT 106.685 155.565 107.035 155.815 ;
        RECT 107.205 155.565 107.555 155.815 ;
        RECT 107.740 155.395 107.910 156.025 ;
        RECT 108.540 156.155 108.870 156.635 ;
        RECT 109.040 156.345 109.265 156.805 ;
        RECT 109.435 156.155 109.765 156.635 ;
        RECT 108.540 155.985 109.765 156.155 ;
        RECT 109.955 156.005 110.205 156.805 ;
        RECT 110.375 156.005 110.715 156.635 ;
        RECT 110.885 156.035 114.395 156.805 ;
        RECT 114.565 156.080 114.855 156.805 ;
        RECT 115.025 156.055 116.235 156.805 ;
        RECT 108.080 155.615 108.410 155.815 ;
        RECT 108.580 155.615 108.910 155.815 ;
        RECT 109.080 155.615 109.500 155.815 ;
        RECT 109.675 155.645 110.370 155.815 ;
        RECT 109.675 155.395 109.845 155.645 ;
        RECT 110.540 155.395 110.715 156.005 ;
        RECT 101.685 154.255 103.355 155.345 ;
        RECT 103.525 154.425 103.865 155.395 ;
        RECT 104.035 154.255 104.205 155.395 ;
        RECT 104.395 155.225 106.830 155.395 ;
        RECT 104.475 154.255 104.725 155.055 ;
        RECT 105.370 154.425 105.700 155.225 ;
        RECT 106.000 154.255 106.330 155.055 ;
        RECT 106.500 154.425 106.830 155.225 ;
        RECT 107.410 155.225 109.845 155.395 ;
        RECT 107.410 154.425 107.740 155.225 ;
        RECT 107.910 154.255 108.240 155.055 ;
        RECT 108.540 154.425 108.870 155.225 ;
        RECT 109.515 154.255 109.765 155.055 ;
        RECT 110.035 154.255 110.205 155.395 ;
        RECT 110.375 154.425 110.715 155.395 ;
        RECT 110.885 155.345 112.575 155.865 ;
        RECT 112.745 155.515 114.395 156.035 ;
        RECT 110.885 154.255 114.395 155.345 ;
        RECT 114.565 154.255 114.855 155.420 ;
        RECT 115.025 155.345 115.545 155.885 ;
        RECT 115.715 155.515 116.235 156.055 ;
        RECT 116.495 156.155 116.665 156.635 ;
        RECT 116.845 156.325 117.085 156.805 ;
        RECT 117.335 156.155 117.505 156.635 ;
        RECT 117.675 156.325 118.005 156.805 ;
        RECT 118.175 156.155 118.345 156.635 ;
        RECT 116.495 155.985 117.130 156.155 ;
        RECT 117.335 155.985 118.345 156.155 ;
        RECT 118.515 156.005 118.845 156.805 ;
        RECT 119.165 156.035 120.835 156.805 ;
        RECT 121.010 156.260 126.355 156.805 ;
        RECT 116.960 155.815 117.130 155.985 ;
        RECT 116.410 155.575 116.790 155.815 ;
        RECT 116.960 155.645 117.460 155.815 ;
        RECT 116.960 155.405 117.130 155.645 ;
        RECT 117.850 155.445 118.345 155.985 ;
        RECT 115.025 154.255 116.235 155.345 ;
        RECT 116.415 155.235 117.130 155.405 ;
        RECT 117.335 155.275 118.345 155.445 ;
        RECT 116.415 154.425 116.745 155.235 ;
        RECT 116.915 154.255 117.155 155.055 ;
        RECT 117.335 154.425 117.505 155.275 ;
        RECT 117.675 154.255 118.005 155.055 ;
        RECT 118.175 154.425 118.345 155.275 ;
        RECT 118.515 154.255 118.845 155.405 ;
        RECT 119.165 155.345 119.915 155.865 ;
        RECT 120.085 155.515 120.835 156.035 ;
        RECT 119.165 154.255 120.835 155.345 ;
        RECT 122.600 154.690 122.950 155.940 ;
        RECT 124.430 155.430 124.770 156.260 ;
        RECT 126.525 156.055 127.735 156.805 ;
        RECT 126.525 155.345 127.045 155.885 ;
        RECT 127.215 155.515 127.735 156.055 ;
        RECT 121.010 154.255 126.355 154.690 ;
        RECT 126.525 154.255 127.735 155.345 ;
        RECT 14.660 154.085 127.820 154.255 ;
        RECT 14.745 152.995 15.955 154.085 ;
        RECT 14.745 152.285 15.265 152.825 ;
        RECT 15.435 152.455 15.955 152.995 ;
        RECT 16.585 152.995 20.095 154.085 ;
        RECT 20.265 153.325 20.780 153.735 ;
        RECT 21.015 153.325 21.185 154.085 ;
        RECT 21.355 153.745 23.385 153.915 ;
        RECT 16.585 152.475 18.275 152.995 ;
        RECT 18.445 152.305 20.095 152.825 ;
        RECT 20.265 152.515 20.605 153.325 ;
        RECT 21.355 153.080 21.525 153.745 ;
        RECT 21.920 153.405 23.045 153.575 ;
        RECT 20.775 152.890 21.525 153.080 ;
        RECT 21.695 153.065 22.705 153.235 ;
        RECT 20.265 152.345 21.495 152.515 ;
        RECT 14.745 151.535 15.955 152.285 ;
        RECT 16.585 151.535 20.095 152.305 ;
        RECT 20.540 151.740 20.785 152.345 ;
        RECT 21.005 151.535 21.515 152.070 ;
        RECT 21.695 151.705 21.885 153.065 ;
        RECT 22.055 152.045 22.330 152.865 ;
        RECT 22.535 152.265 22.705 153.065 ;
        RECT 22.875 152.275 23.045 153.405 ;
        RECT 23.215 152.775 23.385 153.745 ;
        RECT 23.555 152.945 23.725 154.085 ;
        RECT 23.895 152.945 24.230 153.915 ;
        RECT 23.215 152.445 23.410 152.775 ;
        RECT 23.635 152.445 23.890 152.775 ;
        RECT 23.635 152.275 23.805 152.445 ;
        RECT 24.060 152.275 24.230 152.945 ;
        RECT 24.405 152.920 24.695 154.085 ;
        RECT 24.865 152.995 26.075 154.085 ;
        RECT 26.245 152.995 29.755 154.085 ;
        RECT 30.300 153.105 30.555 153.775 ;
        RECT 30.735 153.285 31.020 154.085 ;
        RECT 31.200 153.365 31.530 153.875 ;
        RECT 24.865 152.455 25.385 152.995 ;
        RECT 25.555 152.285 26.075 152.825 ;
        RECT 26.245 152.475 27.935 152.995 ;
        RECT 28.105 152.305 29.755 152.825 ;
        RECT 22.875 152.105 23.805 152.275 ;
        RECT 22.875 152.070 23.050 152.105 ;
        RECT 22.055 151.875 22.335 152.045 ;
        RECT 22.055 151.705 22.330 151.875 ;
        RECT 22.520 151.705 23.050 152.070 ;
        RECT 23.475 151.535 23.805 151.935 ;
        RECT 23.975 151.705 24.230 152.275 ;
        RECT 24.405 151.535 24.695 152.260 ;
        RECT 24.865 151.535 26.075 152.285 ;
        RECT 26.245 151.535 29.755 152.305 ;
        RECT 30.300 152.245 30.480 153.105 ;
        RECT 31.200 152.775 31.450 153.365 ;
        RECT 31.800 153.215 31.970 153.825 ;
        RECT 32.140 153.395 32.470 154.085 ;
        RECT 32.700 153.535 32.940 153.825 ;
        RECT 33.140 153.705 33.560 154.085 ;
        RECT 33.740 153.615 34.370 153.865 ;
        RECT 34.840 153.705 35.170 154.085 ;
        RECT 33.740 153.535 33.910 153.615 ;
        RECT 35.340 153.535 35.510 153.825 ;
        RECT 35.690 153.705 36.070 154.085 ;
        RECT 36.310 153.700 37.140 153.870 ;
        RECT 32.700 153.365 33.910 153.535 ;
        RECT 30.650 152.445 31.450 152.775 ;
        RECT 30.300 152.045 30.555 152.245 ;
        RECT 30.215 151.875 30.555 152.045 ;
        RECT 30.300 151.715 30.555 151.875 ;
        RECT 30.735 151.535 31.020 151.995 ;
        RECT 31.200 151.795 31.450 152.445 ;
        RECT 31.650 153.195 31.970 153.215 ;
        RECT 31.650 153.025 33.570 153.195 ;
        RECT 31.650 152.130 31.840 153.025 ;
        RECT 33.740 152.855 33.910 153.365 ;
        RECT 34.080 153.105 34.600 153.415 ;
        RECT 32.010 152.685 33.910 152.855 ;
        RECT 32.010 152.625 32.340 152.685 ;
        RECT 32.490 152.455 32.820 152.515 ;
        RECT 32.160 152.185 32.820 152.455 ;
        RECT 31.650 151.800 31.970 152.130 ;
        RECT 32.150 151.535 32.810 152.015 ;
        RECT 33.010 151.925 33.180 152.685 ;
        RECT 34.080 152.515 34.260 152.925 ;
        RECT 33.350 152.345 33.680 152.465 ;
        RECT 34.430 152.345 34.600 153.105 ;
        RECT 33.350 152.175 34.600 152.345 ;
        RECT 34.770 153.285 36.140 153.535 ;
        RECT 34.770 152.515 34.960 153.285 ;
        RECT 35.890 153.025 36.140 153.285 ;
        RECT 35.130 152.855 35.380 153.015 ;
        RECT 36.310 152.855 36.480 153.700 ;
        RECT 37.375 153.415 37.545 153.915 ;
        RECT 37.715 153.585 38.045 154.085 ;
        RECT 36.650 153.025 37.150 153.405 ;
        RECT 37.375 153.245 38.070 153.415 ;
        RECT 35.130 152.685 36.480 152.855 ;
        RECT 36.060 152.645 36.480 152.685 ;
        RECT 34.770 152.175 35.190 152.515 ;
        RECT 35.480 152.185 35.890 152.515 ;
        RECT 33.010 151.755 33.860 151.925 ;
        RECT 34.420 151.535 34.740 151.995 ;
        RECT 34.940 151.745 35.190 152.175 ;
        RECT 35.480 151.535 35.890 151.975 ;
        RECT 36.060 151.915 36.230 152.645 ;
        RECT 36.400 152.095 36.750 152.465 ;
        RECT 36.930 152.155 37.150 153.025 ;
        RECT 37.320 152.455 37.730 153.075 ;
        RECT 37.900 152.275 38.070 153.245 ;
        RECT 37.375 152.085 38.070 152.275 ;
        RECT 36.060 151.715 37.075 151.915 ;
        RECT 37.375 151.755 37.545 152.085 ;
        RECT 37.715 151.535 38.045 151.915 ;
        RECT 38.260 151.795 38.485 153.915 ;
        RECT 38.655 153.585 38.985 154.085 ;
        RECT 39.155 153.415 39.325 153.915 ;
        RECT 38.660 153.245 39.325 153.415 ;
        RECT 38.660 152.255 38.890 153.245 ;
        RECT 39.060 152.425 39.410 153.075 ;
        RECT 39.585 152.945 39.925 153.915 ;
        RECT 40.095 152.945 40.265 154.085 ;
        RECT 40.535 153.285 40.785 154.085 ;
        RECT 41.430 153.115 41.760 153.915 ;
        RECT 42.060 153.285 42.390 154.085 ;
        RECT 42.560 153.115 42.890 153.915 ;
        RECT 40.455 152.945 42.890 153.115 ;
        RECT 43.265 152.995 44.475 154.085 ;
        RECT 44.650 153.650 49.995 154.085 ;
        RECT 39.585 152.335 39.760 152.945 ;
        RECT 40.455 152.695 40.625 152.945 ;
        RECT 39.930 152.525 40.625 152.695 ;
        RECT 40.800 152.525 41.220 152.725 ;
        RECT 41.390 152.525 41.720 152.725 ;
        RECT 41.890 152.525 42.220 152.725 ;
        RECT 38.660 152.085 39.325 152.255 ;
        RECT 38.655 151.535 38.985 151.915 ;
        RECT 39.155 151.795 39.325 152.085 ;
        RECT 39.585 151.705 39.925 152.335 ;
        RECT 40.095 151.535 40.345 152.335 ;
        RECT 40.535 152.185 41.760 152.355 ;
        RECT 40.535 151.705 40.865 152.185 ;
        RECT 41.035 151.535 41.260 151.995 ;
        RECT 41.430 151.705 41.760 152.185 ;
        RECT 42.390 152.315 42.560 152.945 ;
        RECT 42.745 152.525 43.095 152.775 ;
        RECT 43.265 152.455 43.785 152.995 ;
        RECT 42.390 151.705 42.890 152.315 ;
        RECT 43.955 152.285 44.475 152.825 ;
        RECT 46.240 152.400 46.590 153.650 ;
        RECT 50.165 152.920 50.455 154.085 ;
        RECT 51.550 153.650 56.895 154.085 ;
        RECT 43.265 151.535 44.475 152.285 ;
        RECT 48.070 152.080 48.410 152.910 ;
        RECT 53.140 152.400 53.490 153.650 ;
        RECT 57.105 152.945 57.335 154.085 ;
        RECT 57.505 152.935 57.835 153.915 ;
        RECT 58.005 152.945 58.215 154.085 ;
        RECT 58.820 153.105 59.075 153.775 ;
        RECT 59.255 153.285 59.540 154.085 ;
        RECT 59.720 153.365 60.050 153.875 ;
        RECT 44.650 151.535 49.995 152.080 ;
        RECT 50.165 151.535 50.455 152.260 ;
        RECT 54.970 152.080 55.310 152.910 ;
        RECT 57.085 152.525 57.415 152.775 ;
        RECT 51.550 151.535 56.895 152.080 ;
        RECT 57.105 151.535 57.335 152.355 ;
        RECT 57.585 152.335 57.835 152.935 ;
        RECT 57.505 151.705 57.835 152.335 ;
        RECT 58.005 151.535 58.215 152.355 ;
        RECT 58.820 152.245 59.000 153.105 ;
        RECT 59.720 152.775 59.970 153.365 ;
        RECT 60.320 153.215 60.490 153.825 ;
        RECT 60.660 153.395 60.990 154.085 ;
        RECT 61.220 153.535 61.460 153.825 ;
        RECT 61.660 153.705 62.080 154.085 ;
        RECT 62.260 153.615 62.890 153.865 ;
        RECT 63.360 153.705 63.690 154.085 ;
        RECT 62.260 153.535 62.430 153.615 ;
        RECT 63.860 153.535 64.030 153.825 ;
        RECT 64.210 153.705 64.590 154.085 ;
        RECT 64.830 153.700 65.660 153.870 ;
        RECT 61.220 153.365 62.430 153.535 ;
        RECT 59.170 152.445 59.970 152.775 ;
        RECT 58.820 152.045 59.075 152.245 ;
        RECT 58.735 151.875 59.075 152.045 ;
        RECT 58.820 151.715 59.075 151.875 ;
        RECT 59.255 151.535 59.540 151.995 ;
        RECT 59.720 151.795 59.970 152.445 ;
        RECT 60.170 153.195 60.490 153.215 ;
        RECT 60.170 153.025 62.090 153.195 ;
        RECT 60.170 152.130 60.360 153.025 ;
        RECT 62.260 152.855 62.430 153.365 ;
        RECT 62.600 153.105 63.120 153.415 ;
        RECT 60.530 152.685 62.430 152.855 ;
        RECT 60.530 152.625 60.860 152.685 ;
        RECT 61.010 152.455 61.340 152.515 ;
        RECT 60.680 152.185 61.340 152.455 ;
        RECT 60.170 151.800 60.490 152.130 ;
        RECT 60.670 151.535 61.330 152.015 ;
        RECT 61.530 151.925 61.700 152.685 ;
        RECT 62.600 152.515 62.780 152.925 ;
        RECT 61.870 152.345 62.200 152.465 ;
        RECT 62.950 152.345 63.120 153.105 ;
        RECT 61.870 152.175 63.120 152.345 ;
        RECT 63.290 153.285 64.660 153.535 ;
        RECT 63.290 152.515 63.480 153.285 ;
        RECT 64.410 153.025 64.660 153.285 ;
        RECT 63.650 152.855 63.900 153.015 ;
        RECT 64.830 152.855 65.000 153.700 ;
        RECT 65.895 153.415 66.065 153.915 ;
        RECT 66.235 153.585 66.565 154.085 ;
        RECT 65.170 153.025 65.670 153.405 ;
        RECT 65.895 153.245 66.590 153.415 ;
        RECT 63.650 152.685 65.000 152.855 ;
        RECT 64.580 152.645 65.000 152.685 ;
        RECT 63.290 152.175 63.710 152.515 ;
        RECT 64.000 152.185 64.410 152.515 ;
        RECT 61.530 151.755 62.380 151.925 ;
        RECT 62.940 151.535 63.260 151.995 ;
        RECT 63.460 151.745 63.710 152.175 ;
        RECT 64.000 151.535 64.410 151.975 ;
        RECT 64.580 151.915 64.750 152.645 ;
        RECT 64.920 152.095 65.270 152.465 ;
        RECT 65.450 152.155 65.670 153.025 ;
        RECT 65.840 152.455 66.250 153.075 ;
        RECT 66.420 152.275 66.590 153.245 ;
        RECT 65.895 152.085 66.590 152.275 ;
        RECT 64.580 151.715 65.595 151.915 ;
        RECT 65.895 151.755 66.065 152.085 ;
        RECT 66.235 151.535 66.565 151.915 ;
        RECT 66.780 151.795 67.005 153.915 ;
        RECT 67.175 153.585 67.505 154.085 ;
        RECT 67.675 153.415 67.845 153.915 ;
        RECT 67.180 153.245 67.845 153.415 ;
        RECT 67.180 152.255 67.410 153.245 ;
        RECT 67.580 152.425 67.930 153.075 ;
        RECT 68.565 152.995 71.155 154.085 ;
        RECT 71.415 153.155 71.585 153.915 ;
        RECT 71.800 153.325 72.130 154.085 ;
        RECT 68.565 152.475 69.775 152.995 ;
        RECT 71.415 152.985 72.130 153.155 ;
        RECT 72.300 153.010 72.555 153.915 ;
        RECT 69.945 152.305 71.155 152.825 ;
        RECT 71.325 152.435 71.680 152.805 ;
        RECT 71.960 152.775 72.130 152.985 ;
        RECT 71.960 152.445 72.215 152.775 ;
        RECT 67.180 152.085 67.845 152.255 ;
        RECT 67.175 151.535 67.505 151.915 ;
        RECT 67.675 151.795 67.845 152.085 ;
        RECT 68.565 151.535 71.155 152.305 ;
        RECT 71.960 152.255 72.130 152.445 ;
        RECT 72.385 152.280 72.555 153.010 ;
        RECT 72.730 152.935 72.990 154.085 ;
        RECT 73.175 153.025 73.505 154.085 ;
        RECT 73.685 152.775 73.855 153.745 ;
        RECT 74.025 153.495 74.355 153.895 ;
        RECT 74.525 153.725 74.855 154.085 ;
        RECT 75.055 153.495 75.755 153.915 ;
        RECT 74.025 153.265 75.755 153.495 ;
        RECT 74.025 153.045 74.355 153.265 ;
        RECT 74.550 152.775 74.875 153.065 ;
        RECT 73.165 152.445 73.475 152.775 ;
        RECT 73.685 152.445 74.060 152.775 ;
        RECT 74.380 152.445 74.875 152.775 ;
        RECT 75.050 152.525 75.380 153.065 ;
        RECT 71.415 152.085 72.130 152.255 ;
        RECT 71.415 151.705 71.585 152.085 ;
        RECT 71.800 151.535 72.130 151.915 ;
        RECT 72.300 151.705 72.555 152.280 ;
        RECT 72.730 151.535 72.990 152.375 ;
        RECT 75.550 152.295 75.755 153.265 ;
        RECT 75.925 152.920 76.215 154.085 ;
        RECT 77.305 152.995 80.815 154.085 ;
        RECT 80.990 153.650 86.335 154.085 ;
        RECT 77.305 152.475 78.995 152.995 ;
        RECT 79.165 152.305 80.815 152.825 ;
        RECT 82.580 152.400 82.930 153.650 ;
        RECT 86.880 153.105 87.135 153.775 ;
        RECT 87.315 153.285 87.600 154.085 ;
        RECT 87.780 153.365 88.110 153.875 ;
        RECT 73.175 152.065 74.535 152.275 ;
        RECT 73.175 151.705 73.505 152.065 ;
        RECT 73.675 151.535 74.005 151.895 ;
        RECT 74.205 151.705 74.535 152.065 ;
        RECT 75.045 151.705 75.755 152.295 ;
        RECT 75.925 151.535 76.215 152.260 ;
        RECT 77.305 151.535 80.815 152.305 ;
        RECT 84.410 152.080 84.750 152.910 ;
        RECT 86.880 152.245 87.060 153.105 ;
        RECT 87.780 152.775 88.030 153.365 ;
        RECT 88.380 153.215 88.550 153.825 ;
        RECT 88.720 153.395 89.050 154.085 ;
        RECT 89.280 153.535 89.520 153.825 ;
        RECT 89.720 153.705 90.140 154.085 ;
        RECT 90.320 153.615 90.950 153.865 ;
        RECT 91.420 153.705 91.750 154.085 ;
        RECT 90.320 153.535 90.490 153.615 ;
        RECT 91.920 153.535 92.090 153.825 ;
        RECT 92.270 153.705 92.650 154.085 ;
        RECT 92.890 153.700 93.720 153.870 ;
        RECT 89.280 153.365 90.490 153.535 ;
        RECT 87.230 152.445 88.030 152.775 ;
        RECT 80.990 151.535 86.335 152.080 ;
        RECT 86.880 152.045 87.135 152.245 ;
        RECT 86.795 151.875 87.135 152.045 ;
        RECT 86.880 151.715 87.135 151.875 ;
        RECT 87.315 151.535 87.600 151.995 ;
        RECT 87.780 151.795 88.030 152.445 ;
        RECT 88.230 153.195 88.550 153.215 ;
        RECT 88.230 153.025 90.150 153.195 ;
        RECT 88.230 152.130 88.420 153.025 ;
        RECT 90.320 152.855 90.490 153.365 ;
        RECT 90.660 153.105 91.180 153.415 ;
        RECT 88.590 152.685 90.490 152.855 ;
        RECT 88.590 152.625 88.920 152.685 ;
        RECT 89.070 152.455 89.400 152.515 ;
        RECT 88.740 152.185 89.400 152.455 ;
        RECT 88.230 151.800 88.550 152.130 ;
        RECT 88.730 151.535 89.390 152.015 ;
        RECT 89.590 151.925 89.760 152.685 ;
        RECT 90.660 152.515 90.840 152.925 ;
        RECT 89.930 152.345 90.260 152.465 ;
        RECT 91.010 152.345 91.180 153.105 ;
        RECT 89.930 152.175 91.180 152.345 ;
        RECT 91.350 153.285 92.720 153.535 ;
        RECT 91.350 152.515 91.540 153.285 ;
        RECT 92.470 153.025 92.720 153.285 ;
        RECT 91.710 152.855 91.960 153.015 ;
        RECT 92.890 152.855 93.060 153.700 ;
        RECT 93.955 153.415 94.125 153.915 ;
        RECT 94.295 153.585 94.625 154.085 ;
        RECT 93.230 153.025 93.730 153.405 ;
        RECT 93.955 153.245 94.650 153.415 ;
        RECT 91.710 152.685 93.060 152.855 ;
        RECT 92.640 152.645 93.060 152.685 ;
        RECT 91.350 152.175 91.770 152.515 ;
        RECT 92.060 152.185 92.470 152.515 ;
        RECT 89.590 151.755 90.440 151.925 ;
        RECT 91.000 151.535 91.320 151.995 ;
        RECT 91.520 151.745 91.770 152.175 ;
        RECT 92.060 151.535 92.470 151.975 ;
        RECT 92.640 151.915 92.810 152.645 ;
        RECT 92.980 152.095 93.330 152.465 ;
        RECT 93.510 152.155 93.730 153.025 ;
        RECT 93.900 152.455 94.310 153.075 ;
        RECT 94.480 152.275 94.650 153.245 ;
        RECT 93.955 152.085 94.650 152.275 ;
        RECT 92.640 151.715 93.655 151.915 ;
        RECT 93.955 151.755 94.125 152.085 ;
        RECT 94.295 151.535 94.625 151.915 ;
        RECT 94.840 151.795 95.065 153.915 ;
        RECT 95.235 153.585 95.565 154.085 ;
        RECT 95.735 153.415 95.905 153.915 ;
        RECT 96.170 153.650 101.515 154.085 ;
        RECT 95.240 153.245 95.905 153.415 ;
        RECT 95.240 152.255 95.470 153.245 ;
        RECT 95.640 152.425 95.990 153.075 ;
        RECT 97.760 152.400 98.110 153.650 ;
        RECT 101.685 152.920 101.975 154.085 ;
        RECT 102.605 152.945 102.875 153.915 ;
        RECT 103.085 153.285 103.365 154.085 ;
        RECT 103.535 153.575 105.190 153.865 ;
        RECT 103.600 153.235 105.190 153.405 ;
        RECT 103.600 153.115 103.770 153.235 ;
        RECT 103.045 152.945 103.770 153.115 ;
        RECT 95.240 152.085 95.905 152.255 ;
        RECT 95.235 151.535 95.565 151.915 ;
        RECT 95.735 151.795 95.905 152.085 ;
        RECT 99.590 152.080 99.930 152.910 ;
        RECT 96.170 151.535 101.515 152.080 ;
        RECT 101.685 151.535 101.975 152.260 ;
        RECT 102.605 152.210 102.775 152.945 ;
        RECT 103.045 152.775 103.215 152.945 ;
        RECT 103.960 152.895 104.675 153.065 ;
        RECT 104.870 152.945 105.190 153.235 ;
        RECT 105.365 152.945 105.705 153.915 ;
        RECT 105.875 152.945 106.045 154.085 ;
        RECT 106.315 153.285 106.565 154.085 ;
        RECT 107.210 153.115 107.540 153.915 ;
        RECT 107.840 153.285 108.170 154.085 ;
        RECT 108.340 153.115 108.670 153.915 ;
        RECT 106.235 152.945 108.670 153.115 ;
        RECT 109.045 152.945 109.385 153.915 ;
        RECT 109.555 152.945 109.725 154.085 ;
        RECT 109.995 153.285 110.245 154.085 ;
        RECT 110.890 153.115 111.220 153.915 ;
        RECT 111.520 153.285 111.850 154.085 ;
        RECT 112.020 153.115 112.350 153.915 ;
        RECT 113.190 153.650 118.535 154.085 ;
        RECT 109.915 152.945 112.350 153.115 ;
        RECT 102.945 152.445 103.215 152.775 ;
        RECT 103.385 152.445 103.790 152.775 ;
        RECT 103.960 152.445 104.670 152.895 ;
        RECT 103.045 152.275 103.215 152.445 ;
        RECT 102.605 151.865 102.875 152.210 ;
        RECT 103.045 152.105 104.655 152.275 ;
        RECT 104.840 152.205 105.190 152.775 ;
        RECT 105.365 152.335 105.540 152.945 ;
        RECT 106.235 152.695 106.405 152.945 ;
        RECT 105.710 152.525 106.405 152.695 ;
        RECT 106.580 152.525 107.000 152.725 ;
        RECT 107.170 152.525 107.500 152.725 ;
        RECT 107.670 152.525 108.000 152.725 ;
        RECT 103.065 151.535 103.445 151.935 ;
        RECT 103.615 151.755 103.785 152.105 ;
        RECT 103.955 151.535 104.285 151.935 ;
        RECT 104.485 151.755 104.655 152.105 ;
        RECT 104.855 151.535 105.185 152.035 ;
        RECT 105.365 151.705 105.705 152.335 ;
        RECT 105.875 151.535 106.125 152.335 ;
        RECT 106.315 152.185 107.540 152.355 ;
        RECT 106.315 151.705 106.645 152.185 ;
        RECT 106.815 151.535 107.040 151.995 ;
        RECT 107.210 151.705 107.540 152.185 ;
        RECT 108.170 152.315 108.340 152.945 ;
        RECT 108.525 152.525 108.875 152.775 ;
        RECT 109.045 152.385 109.220 152.945 ;
        RECT 109.915 152.695 110.085 152.945 ;
        RECT 109.390 152.525 110.085 152.695 ;
        RECT 110.260 152.525 110.680 152.725 ;
        RECT 110.850 152.525 111.180 152.725 ;
        RECT 111.350 152.525 111.680 152.725 ;
        RECT 109.045 152.335 109.275 152.385 ;
        RECT 108.170 151.705 108.670 152.315 ;
        RECT 109.045 151.705 109.385 152.335 ;
        RECT 109.555 151.535 109.805 152.335 ;
        RECT 109.995 152.185 111.220 152.355 ;
        RECT 109.995 151.705 110.325 152.185 ;
        RECT 110.495 151.535 110.720 151.995 ;
        RECT 110.890 151.705 111.220 152.185 ;
        RECT 111.850 152.315 112.020 152.945 ;
        RECT 112.205 152.525 112.555 152.775 ;
        RECT 114.780 152.400 115.130 153.650 ;
        RECT 118.765 152.945 118.975 154.085 ;
        RECT 119.145 152.935 119.475 153.915 ;
        RECT 119.645 152.945 119.875 154.085 ;
        RECT 120.635 153.155 120.805 153.915 ;
        RECT 120.985 153.325 121.315 154.085 ;
        RECT 120.635 152.985 121.300 153.155 ;
        RECT 121.485 153.010 121.755 153.915 ;
        RECT 111.850 151.705 112.350 152.315 ;
        RECT 116.610 152.080 116.950 152.910 ;
        RECT 113.190 151.535 118.535 152.080 ;
        RECT 118.765 151.535 118.975 152.355 ;
        RECT 119.145 152.335 119.395 152.935 ;
        RECT 121.130 152.840 121.300 152.985 ;
        RECT 119.565 152.525 119.895 152.775 ;
        RECT 120.565 152.435 120.895 152.805 ;
        RECT 121.130 152.510 121.415 152.840 ;
        RECT 119.145 151.705 119.475 152.335 ;
        RECT 119.645 151.535 119.875 152.355 ;
        RECT 121.130 152.255 121.300 152.510 ;
        RECT 120.635 152.085 121.300 152.255 ;
        RECT 121.585 152.210 121.755 153.010 ;
        RECT 122.845 152.995 126.355 154.085 ;
        RECT 126.525 152.995 127.735 154.085 ;
        RECT 122.845 152.475 124.535 152.995 ;
        RECT 124.705 152.305 126.355 152.825 ;
        RECT 126.525 152.455 127.045 152.995 ;
        RECT 120.635 151.705 120.805 152.085 ;
        RECT 120.985 151.535 121.315 151.915 ;
        RECT 121.495 151.705 121.755 152.210 ;
        RECT 122.845 151.535 126.355 152.305 ;
        RECT 127.215 152.285 127.735 152.825 ;
        RECT 126.525 151.535 127.735 152.285 ;
        RECT 14.660 151.365 127.820 151.535 ;
        RECT 14.745 150.615 15.955 151.365 ;
        RECT 16.960 150.655 17.215 151.185 ;
        RECT 17.395 150.905 17.680 151.365 ;
        RECT 14.745 150.075 15.265 150.615 ;
        RECT 15.435 149.905 15.955 150.445 ;
        RECT 16.960 150.005 17.140 150.655 ;
        RECT 17.860 150.455 18.110 151.105 ;
        RECT 17.310 150.125 18.110 150.455 ;
        RECT 14.745 148.815 15.955 149.905 ;
        RECT 16.875 149.835 17.140 150.005 ;
        RECT 16.960 149.795 17.140 149.835 ;
        RECT 16.960 149.125 17.215 149.795 ;
        RECT 17.395 148.815 17.680 149.615 ;
        RECT 17.860 149.535 18.110 150.125 ;
        RECT 18.310 150.770 18.630 151.100 ;
        RECT 18.810 150.885 19.470 151.365 ;
        RECT 19.670 150.975 20.520 151.145 ;
        RECT 18.310 149.875 18.500 150.770 ;
        RECT 18.820 150.445 19.480 150.715 ;
        RECT 19.150 150.385 19.480 150.445 ;
        RECT 18.670 150.215 19.000 150.275 ;
        RECT 19.670 150.215 19.840 150.975 ;
        RECT 21.080 150.905 21.400 151.365 ;
        RECT 21.600 150.725 21.850 151.155 ;
        RECT 22.140 150.925 22.550 151.365 ;
        RECT 22.720 150.985 23.735 151.185 ;
        RECT 20.010 150.555 21.260 150.725 ;
        RECT 20.010 150.435 20.340 150.555 ;
        RECT 18.670 150.045 20.570 150.215 ;
        RECT 18.310 149.705 20.230 149.875 ;
        RECT 18.310 149.685 18.630 149.705 ;
        RECT 17.860 149.025 18.190 149.535 ;
        RECT 18.460 149.075 18.630 149.685 ;
        RECT 20.400 149.535 20.570 150.045 ;
        RECT 20.740 149.975 20.920 150.385 ;
        RECT 21.090 149.795 21.260 150.555 ;
        RECT 18.800 148.815 19.130 149.505 ;
        RECT 19.360 149.365 20.570 149.535 ;
        RECT 20.740 149.485 21.260 149.795 ;
        RECT 21.430 150.385 21.850 150.725 ;
        RECT 22.140 150.385 22.550 150.715 ;
        RECT 21.430 149.615 21.620 150.385 ;
        RECT 22.720 150.255 22.890 150.985 ;
        RECT 24.035 150.815 24.205 151.145 ;
        RECT 24.375 150.985 24.705 151.365 ;
        RECT 23.060 150.435 23.410 150.805 ;
        RECT 22.720 150.215 23.140 150.255 ;
        RECT 21.790 150.045 23.140 150.215 ;
        RECT 21.790 149.885 22.040 150.045 ;
        RECT 22.550 149.615 22.800 149.875 ;
        RECT 21.430 149.365 22.800 149.615 ;
        RECT 19.360 149.075 19.600 149.365 ;
        RECT 20.400 149.285 20.570 149.365 ;
        RECT 19.800 148.815 20.220 149.195 ;
        RECT 20.400 149.035 21.030 149.285 ;
        RECT 21.500 148.815 21.830 149.195 ;
        RECT 22.000 149.075 22.170 149.365 ;
        RECT 22.970 149.200 23.140 150.045 ;
        RECT 23.590 149.875 23.810 150.745 ;
        RECT 24.035 150.625 24.730 150.815 ;
        RECT 23.310 149.495 23.810 149.875 ;
        RECT 23.980 149.825 24.390 150.445 ;
        RECT 24.560 149.655 24.730 150.625 ;
        RECT 24.035 149.485 24.730 149.655 ;
        RECT 22.350 148.815 22.730 149.195 ;
        RECT 22.970 149.030 23.800 149.200 ;
        RECT 24.035 148.985 24.205 149.485 ;
        RECT 24.375 148.815 24.705 149.315 ;
        RECT 24.920 148.985 25.145 151.105 ;
        RECT 25.315 150.985 25.645 151.365 ;
        RECT 25.815 150.815 25.985 151.105 ;
        RECT 25.320 150.645 25.985 150.815 ;
        RECT 25.320 149.655 25.550 150.645 ;
        RECT 26.245 150.615 27.455 151.365 ;
        RECT 27.630 150.820 32.975 151.365 ;
        RECT 25.720 149.825 26.070 150.475 ;
        RECT 26.245 149.905 26.765 150.445 ;
        RECT 26.935 150.075 27.455 150.615 ;
        RECT 25.320 149.485 25.985 149.655 ;
        RECT 25.315 148.815 25.645 149.315 ;
        RECT 25.815 148.985 25.985 149.485 ;
        RECT 26.245 148.815 27.455 149.905 ;
        RECT 29.220 149.250 29.570 150.500 ;
        RECT 31.050 149.990 31.390 150.820 ;
        RECT 33.185 150.545 33.415 151.365 ;
        RECT 33.585 150.565 33.915 151.195 ;
        RECT 33.165 150.125 33.495 150.375 ;
        RECT 33.665 149.965 33.915 150.565 ;
        RECT 34.085 150.545 34.295 151.365 ;
        RECT 34.525 150.615 35.735 151.365 ;
        RECT 35.995 150.815 36.165 151.195 ;
        RECT 36.345 150.985 36.675 151.365 ;
        RECT 35.995 150.645 36.660 150.815 ;
        RECT 36.855 150.690 37.115 151.195 ;
        RECT 27.630 148.815 32.975 149.250 ;
        RECT 33.185 148.815 33.415 149.955 ;
        RECT 33.585 148.985 33.915 149.965 ;
        RECT 34.085 148.815 34.295 149.955 ;
        RECT 34.525 149.905 35.045 150.445 ;
        RECT 35.215 150.075 35.735 150.615 ;
        RECT 35.925 150.095 36.255 150.465 ;
        RECT 36.490 150.390 36.660 150.645 ;
        RECT 36.490 150.060 36.775 150.390 ;
        RECT 36.490 149.915 36.660 150.060 ;
        RECT 34.525 148.815 35.735 149.905 ;
        RECT 35.995 149.745 36.660 149.915 ;
        RECT 36.945 149.890 37.115 150.690 ;
        RECT 37.285 150.640 37.575 151.365 ;
        RECT 37.745 150.595 41.255 151.365 ;
        RECT 35.995 148.985 36.165 149.745 ;
        RECT 36.345 148.815 36.675 149.575 ;
        RECT 36.845 148.985 37.115 149.890 ;
        RECT 37.285 148.815 37.575 149.980 ;
        RECT 37.745 149.905 39.435 150.425 ;
        RECT 39.605 150.075 41.255 150.595 ;
        RECT 41.425 150.565 41.765 151.195 ;
        RECT 41.935 150.565 42.185 151.365 ;
        RECT 42.375 150.715 42.705 151.195 ;
        RECT 42.875 150.905 43.100 151.365 ;
        RECT 43.270 150.715 43.600 151.195 ;
        RECT 41.425 149.955 41.600 150.565 ;
        RECT 42.375 150.545 43.600 150.715 ;
        RECT 44.230 150.585 44.730 151.195 ;
        RECT 45.105 150.595 48.615 151.365 ;
        RECT 48.795 150.865 49.125 151.365 ;
        RECT 49.325 150.795 49.495 151.145 ;
        RECT 49.695 150.965 50.025 151.365 ;
        RECT 50.195 150.795 50.365 151.145 ;
        RECT 50.535 150.965 50.915 151.365 ;
        RECT 41.770 150.205 42.465 150.375 ;
        RECT 42.295 149.955 42.465 150.205 ;
        RECT 42.640 150.175 43.060 150.375 ;
        RECT 43.230 150.175 43.560 150.375 ;
        RECT 43.730 150.175 44.060 150.375 ;
        RECT 44.230 149.955 44.400 150.585 ;
        RECT 44.585 150.125 44.935 150.375 ;
        RECT 37.745 148.815 41.255 149.905 ;
        RECT 41.425 148.985 41.765 149.955 ;
        RECT 41.935 148.815 42.105 149.955 ;
        RECT 42.295 149.785 44.730 149.955 ;
        RECT 42.375 148.815 42.625 149.615 ;
        RECT 43.270 148.985 43.600 149.785 ;
        RECT 43.900 148.815 44.230 149.615 ;
        RECT 44.400 148.985 44.730 149.785 ;
        RECT 45.105 149.905 46.795 150.425 ;
        RECT 46.965 150.075 48.615 150.595 ;
        RECT 48.790 150.125 49.140 150.695 ;
        RECT 49.325 150.625 50.935 150.795 ;
        RECT 51.105 150.690 51.375 151.035 ;
        RECT 50.765 150.455 50.935 150.625 ;
        RECT 45.105 148.815 48.615 149.905 ;
        RECT 48.790 149.665 49.110 149.955 ;
        RECT 49.310 149.835 50.020 150.455 ;
        RECT 50.190 150.125 50.595 150.455 ;
        RECT 50.765 150.125 51.035 150.455 ;
        RECT 50.765 149.955 50.935 150.125 ;
        RECT 51.205 149.955 51.375 150.690 ;
        RECT 50.210 149.785 50.935 149.955 ;
        RECT 50.210 149.665 50.380 149.785 ;
        RECT 48.790 149.495 50.380 149.665 ;
        RECT 48.790 149.035 50.445 149.325 ;
        RECT 50.615 148.815 50.895 149.615 ;
        RECT 51.105 148.985 51.375 149.955 ;
        RECT 51.545 150.565 51.885 151.195 ;
        RECT 52.055 150.565 52.305 151.365 ;
        RECT 52.495 150.715 52.825 151.195 ;
        RECT 52.995 150.905 53.220 151.365 ;
        RECT 53.390 150.715 53.720 151.195 ;
        RECT 51.545 149.955 51.720 150.565 ;
        RECT 52.495 150.545 53.720 150.715 ;
        RECT 54.350 150.585 54.850 151.195 ;
        RECT 55.225 150.595 56.895 151.365 ;
        RECT 51.890 150.205 52.585 150.375 ;
        RECT 52.415 149.955 52.585 150.205 ;
        RECT 52.760 150.175 53.180 150.375 ;
        RECT 53.350 150.175 53.680 150.375 ;
        RECT 53.850 150.175 54.180 150.375 ;
        RECT 54.350 149.955 54.520 150.585 ;
        RECT 54.705 150.125 55.055 150.375 ;
        RECT 51.545 148.985 51.885 149.955 ;
        RECT 52.055 148.815 52.225 149.955 ;
        RECT 52.415 149.785 54.850 149.955 ;
        RECT 52.495 148.815 52.745 149.615 ;
        RECT 53.390 148.985 53.720 149.785 ;
        RECT 54.020 148.815 54.350 149.615 ;
        RECT 54.520 148.985 54.850 149.785 ;
        RECT 55.225 149.905 55.975 150.425 ;
        RECT 56.145 150.075 56.895 150.595 ;
        RECT 57.340 150.555 57.585 151.160 ;
        RECT 57.805 150.830 58.315 151.365 ;
        RECT 57.065 150.385 58.295 150.555 ;
        RECT 55.225 148.815 56.895 149.905 ;
        RECT 57.065 149.575 57.405 150.385 ;
        RECT 57.575 149.820 58.325 150.010 ;
        RECT 57.065 149.165 57.580 149.575 ;
        RECT 57.815 148.815 57.985 149.575 ;
        RECT 58.155 149.155 58.325 149.820 ;
        RECT 58.495 149.835 58.685 151.195 ;
        RECT 58.855 150.345 59.130 151.195 ;
        RECT 59.320 150.830 59.850 151.195 ;
        RECT 60.275 150.965 60.605 151.365 ;
        RECT 59.675 150.795 59.850 150.830 ;
        RECT 58.855 150.175 59.135 150.345 ;
        RECT 58.855 150.035 59.130 150.175 ;
        RECT 59.335 149.835 59.505 150.635 ;
        RECT 58.495 149.665 59.505 149.835 ;
        RECT 59.675 150.625 60.605 150.795 ;
        RECT 60.775 150.625 61.030 151.195 ;
        RECT 59.675 149.495 59.845 150.625 ;
        RECT 60.435 150.455 60.605 150.625 ;
        RECT 58.720 149.325 59.845 149.495 ;
        RECT 60.015 150.125 60.210 150.455 ;
        RECT 60.435 150.125 60.690 150.455 ;
        RECT 60.015 149.155 60.185 150.125 ;
        RECT 60.860 149.955 61.030 150.625 ;
        RECT 58.155 148.985 60.185 149.155 ;
        RECT 60.355 148.815 60.525 149.955 ;
        RECT 60.695 148.985 61.030 149.955 ;
        RECT 61.665 150.690 61.925 151.195 ;
        RECT 62.105 150.985 62.435 151.365 ;
        RECT 62.615 150.815 62.785 151.195 ;
        RECT 61.665 149.890 61.835 150.690 ;
        RECT 62.120 150.645 62.785 150.815 ;
        RECT 62.120 150.390 62.290 150.645 ;
        RECT 63.045 150.640 63.335 151.365 ;
        RECT 64.055 150.815 64.225 151.195 ;
        RECT 64.405 150.985 64.735 151.365 ;
        RECT 64.055 150.645 64.720 150.815 ;
        RECT 64.915 150.690 65.175 151.195 ;
        RECT 62.005 150.060 62.290 150.390 ;
        RECT 62.525 150.095 62.855 150.465 ;
        RECT 63.985 150.095 64.315 150.465 ;
        RECT 64.550 150.390 64.720 150.645 ;
        RECT 62.120 149.915 62.290 150.060 ;
        RECT 64.550 150.060 64.835 150.390 ;
        RECT 61.665 148.985 61.935 149.890 ;
        RECT 62.120 149.745 62.785 149.915 ;
        RECT 62.105 148.815 62.435 149.575 ;
        RECT 62.615 148.985 62.785 149.745 ;
        RECT 63.045 148.815 63.335 149.980 ;
        RECT 64.550 149.915 64.720 150.060 ;
        RECT 64.055 149.745 64.720 149.915 ;
        RECT 65.005 149.890 65.175 150.690 ;
        RECT 65.805 150.595 67.475 151.365 ;
        RECT 67.735 150.815 67.905 151.195 ;
        RECT 68.120 150.985 68.450 151.365 ;
        RECT 67.735 150.645 68.450 150.815 ;
        RECT 64.055 148.985 64.225 149.745 ;
        RECT 64.405 148.815 64.735 149.575 ;
        RECT 64.905 148.985 65.175 149.890 ;
        RECT 65.805 149.905 66.555 150.425 ;
        RECT 66.725 150.075 67.475 150.595 ;
        RECT 67.645 150.095 68.000 150.465 ;
        RECT 68.280 150.455 68.450 150.645 ;
        RECT 68.620 150.620 68.875 151.195 ;
        RECT 68.280 150.125 68.535 150.455 ;
        RECT 68.280 149.915 68.450 150.125 ;
        RECT 65.805 148.815 67.475 149.905 ;
        RECT 67.735 149.745 68.450 149.915 ;
        RECT 68.705 149.890 68.875 150.620 ;
        RECT 69.050 150.525 69.310 151.365 ;
        RECT 69.490 150.525 69.750 151.365 ;
        RECT 69.925 150.620 70.180 151.195 ;
        RECT 70.350 150.985 70.680 151.365 ;
        RECT 70.895 150.815 71.065 151.195 ;
        RECT 71.385 150.885 71.665 151.365 ;
        RECT 70.350 150.645 71.065 150.815 ;
        RECT 71.835 150.715 72.095 151.105 ;
        RECT 72.270 150.885 72.525 151.365 ;
        RECT 72.695 150.715 72.990 151.105 ;
        RECT 73.170 150.885 73.445 151.365 ;
        RECT 73.615 150.865 73.915 151.195 ;
        RECT 67.735 148.985 67.905 149.745 ;
        RECT 68.120 148.815 68.450 149.575 ;
        RECT 68.620 148.985 68.875 149.890 ;
        RECT 69.050 148.815 69.310 149.965 ;
        RECT 69.490 148.815 69.750 149.965 ;
        RECT 69.925 149.890 70.095 150.620 ;
        RECT 70.350 150.455 70.520 150.645 ;
        RECT 71.340 150.545 72.990 150.715 ;
        RECT 70.265 150.125 70.520 150.455 ;
        RECT 70.350 149.915 70.520 150.125 ;
        RECT 70.800 150.095 71.155 150.465 ;
        RECT 71.340 150.035 71.745 150.545 ;
        RECT 71.915 150.205 73.055 150.375 ;
        RECT 69.925 148.985 70.180 149.890 ;
        RECT 70.350 149.745 71.065 149.915 ;
        RECT 71.340 149.865 72.095 150.035 ;
        RECT 70.350 148.815 70.680 149.575 ;
        RECT 70.895 148.985 71.065 149.745 ;
        RECT 71.380 148.815 71.665 149.685 ;
        RECT 71.835 149.615 72.095 149.865 ;
        RECT 72.885 149.955 73.055 150.205 ;
        RECT 73.225 150.125 73.575 150.695 ;
        RECT 73.745 149.955 73.915 150.865 ;
        RECT 72.885 149.785 73.915 149.955 ;
        RECT 71.835 149.445 72.955 149.615 ;
        RECT 71.835 148.985 72.095 149.445 ;
        RECT 72.270 148.815 72.525 149.275 ;
        RECT 72.695 148.985 72.955 149.445 ;
        RECT 73.125 148.815 73.435 149.615 ;
        RECT 73.605 148.985 73.915 149.785 ;
        RECT 75.005 150.865 75.305 151.195 ;
        RECT 75.475 150.885 75.750 151.365 ;
        RECT 75.005 149.955 75.175 150.865 ;
        RECT 75.930 150.715 76.225 151.105 ;
        RECT 76.395 150.885 76.650 151.365 ;
        RECT 76.825 150.715 77.085 151.105 ;
        RECT 77.255 150.885 77.535 151.365 ;
        RECT 75.345 150.125 75.695 150.695 ;
        RECT 75.930 150.545 77.580 150.715 ;
        RECT 75.865 150.205 77.005 150.375 ;
        RECT 75.865 149.955 76.035 150.205 ;
        RECT 77.175 150.035 77.580 150.545 ;
        RECT 75.005 149.785 76.035 149.955 ;
        RECT 76.825 149.865 77.580 150.035 ;
        RECT 77.765 150.690 78.035 151.035 ;
        RECT 78.225 150.965 78.605 151.365 ;
        RECT 78.775 150.795 78.945 151.145 ;
        RECT 79.115 150.965 79.445 151.365 ;
        RECT 79.645 150.795 79.815 151.145 ;
        RECT 80.015 150.865 80.345 151.365 ;
        RECT 77.765 149.955 77.935 150.690 ;
        RECT 78.205 150.625 79.815 150.795 ;
        RECT 78.205 150.455 78.375 150.625 ;
        RECT 78.105 150.125 78.375 150.455 ;
        RECT 78.545 150.125 78.950 150.455 ;
        RECT 78.205 149.955 78.375 150.125 ;
        RECT 79.120 150.005 79.830 150.455 ;
        RECT 80.000 150.125 80.350 150.695 ;
        RECT 80.985 150.595 84.495 151.365 ;
        RECT 75.005 148.985 75.315 149.785 ;
        RECT 76.825 149.615 77.085 149.865 ;
        RECT 75.485 148.815 75.795 149.615 ;
        RECT 75.965 149.445 77.085 149.615 ;
        RECT 75.965 148.985 76.225 149.445 ;
        RECT 76.395 148.815 76.650 149.275 ;
        RECT 76.825 148.985 77.085 149.445 ;
        RECT 77.255 148.815 77.540 149.685 ;
        RECT 77.765 148.985 78.035 149.955 ;
        RECT 78.205 149.785 78.930 149.955 ;
        RECT 79.120 149.835 79.835 150.005 ;
        RECT 78.760 149.665 78.930 149.785 ;
        RECT 80.030 149.665 80.350 149.955 ;
        RECT 78.245 148.815 78.525 149.615 ;
        RECT 78.760 149.495 80.350 149.665 ;
        RECT 80.985 149.905 82.675 150.425 ;
        RECT 82.845 150.075 84.495 150.595 ;
        RECT 84.940 150.555 85.185 151.160 ;
        RECT 85.405 150.830 85.915 151.365 ;
        RECT 84.665 150.385 85.895 150.555 ;
        RECT 78.695 149.035 80.350 149.325 ;
        RECT 80.985 148.815 84.495 149.905 ;
        RECT 84.665 149.575 85.005 150.385 ;
        RECT 85.175 149.820 85.925 150.010 ;
        RECT 84.665 149.165 85.180 149.575 ;
        RECT 85.415 148.815 85.585 149.575 ;
        RECT 85.755 149.155 85.925 149.820 ;
        RECT 86.095 149.835 86.285 151.195 ;
        RECT 86.455 150.345 86.730 151.195 ;
        RECT 86.920 150.830 87.450 151.195 ;
        RECT 87.875 150.965 88.205 151.365 ;
        RECT 87.275 150.795 87.450 150.830 ;
        RECT 86.455 150.175 86.735 150.345 ;
        RECT 86.455 150.035 86.730 150.175 ;
        RECT 86.935 149.835 87.105 150.635 ;
        RECT 86.095 149.665 87.105 149.835 ;
        RECT 87.275 150.625 88.205 150.795 ;
        RECT 88.375 150.625 88.630 151.195 ;
        RECT 88.805 150.640 89.095 151.365 ;
        RECT 87.275 149.495 87.445 150.625 ;
        RECT 88.035 150.455 88.205 150.625 ;
        RECT 86.320 149.325 87.445 149.495 ;
        RECT 87.615 150.125 87.810 150.455 ;
        RECT 88.035 150.125 88.290 150.455 ;
        RECT 87.615 149.155 87.785 150.125 ;
        RECT 88.460 149.955 88.630 150.625 ;
        RECT 89.785 150.545 89.995 151.365 ;
        RECT 90.165 150.565 90.495 151.195 ;
        RECT 85.755 148.985 87.785 149.155 ;
        RECT 87.955 148.815 88.125 149.955 ;
        RECT 88.295 148.985 88.630 149.955 ;
        RECT 88.805 148.815 89.095 149.980 ;
        RECT 90.165 149.965 90.415 150.565 ;
        RECT 90.665 150.545 90.895 151.365 ;
        RECT 92.115 150.815 92.285 151.195 ;
        RECT 92.465 150.985 92.795 151.365 ;
        RECT 92.115 150.645 92.780 150.815 ;
        RECT 92.975 150.690 93.235 151.195 ;
        RECT 90.585 150.125 90.915 150.375 ;
        RECT 92.045 150.095 92.375 150.465 ;
        RECT 92.610 150.390 92.780 150.645 ;
        RECT 92.610 150.060 92.895 150.390 ;
        RECT 89.785 148.815 89.995 149.955 ;
        RECT 90.165 148.985 90.495 149.965 ;
        RECT 90.665 148.815 90.895 149.955 ;
        RECT 92.610 149.915 92.780 150.060 ;
        RECT 92.115 149.745 92.780 149.915 ;
        RECT 93.065 149.890 93.235 150.690 ;
        RECT 93.465 150.545 93.675 151.365 ;
        RECT 93.845 150.565 94.175 151.195 ;
        RECT 93.845 149.965 94.095 150.565 ;
        RECT 94.345 150.545 94.575 151.365 ;
        RECT 94.785 150.595 96.455 151.365 ;
        RECT 94.265 150.125 94.595 150.375 ;
        RECT 92.115 148.985 92.285 149.745 ;
        RECT 92.465 148.815 92.795 149.575 ;
        RECT 92.965 148.985 93.235 149.890 ;
        RECT 93.465 148.815 93.675 149.955 ;
        RECT 93.845 148.985 94.175 149.965 ;
        RECT 94.345 148.815 94.575 149.955 ;
        RECT 94.785 149.905 95.535 150.425 ;
        RECT 95.705 150.075 96.455 150.595 ;
        RECT 96.630 150.655 96.885 151.185 ;
        RECT 97.055 150.905 97.360 151.365 ;
        RECT 97.605 150.985 98.675 151.155 ;
        RECT 96.630 150.005 96.840 150.655 ;
        RECT 97.605 150.630 97.925 150.985 ;
        RECT 97.600 150.455 97.925 150.630 ;
        RECT 97.010 150.155 97.925 150.455 ;
        RECT 98.095 150.415 98.335 150.815 ;
        RECT 98.505 150.755 98.675 150.985 ;
        RECT 98.845 150.925 99.035 151.365 ;
        RECT 99.205 150.915 100.155 151.195 ;
        RECT 100.375 151.005 100.725 151.175 ;
        RECT 98.505 150.585 99.035 150.755 ;
        RECT 97.010 150.125 97.750 150.155 ;
        RECT 94.785 148.815 96.455 149.905 ;
        RECT 96.630 149.125 96.885 150.005 ;
        RECT 97.055 148.815 97.360 149.955 ;
        RECT 97.580 149.535 97.750 150.125 ;
        RECT 98.095 150.045 98.635 150.415 ;
        RECT 98.815 150.305 99.035 150.585 ;
        RECT 99.205 150.135 99.375 150.915 ;
        RECT 98.970 149.965 99.375 150.135 ;
        RECT 99.545 150.125 99.895 150.745 ;
        RECT 98.970 149.875 99.140 149.965 ;
        RECT 100.065 149.955 100.275 150.745 ;
        RECT 97.920 149.705 99.140 149.875 ;
        RECT 99.600 149.795 100.275 149.955 ;
        RECT 97.580 149.365 98.380 149.535 ;
        RECT 97.700 148.815 98.030 149.195 ;
        RECT 98.210 149.075 98.380 149.365 ;
        RECT 98.970 149.325 99.140 149.705 ;
        RECT 99.310 149.785 100.275 149.795 ;
        RECT 100.465 150.615 100.725 151.005 ;
        RECT 100.935 150.905 101.265 151.365 ;
        RECT 102.140 150.975 102.995 151.145 ;
        RECT 103.200 150.975 103.695 151.145 ;
        RECT 103.865 151.005 104.195 151.365 ;
        RECT 100.465 149.925 100.635 150.615 ;
        RECT 100.805 150.265 100.975 150.445 ;
        RECT 101.145 150.435 101.935 150.685 ;
        RECT 102.140 150.265 102.310 150.975 ;
        RECT 102.480 150.465 102.835 150.685 ;
        RECT 100.805 150.095 102.495 150.265 ;
        RECT 99.310 149.495 99.770 149.785 ;
        RECT 100.465 149.755 101.965 149.925 ;
        RECT 100.465 149.615 100.635 149.755 ;
        RECT 100.075 149.445 100.635 149.615 ;
        RECT 98.550 148.815 98.800 149.275 ;
        RECT 98.970 148.985 99.840 149.325 ;
        RECT 100.075 148.985 100.245 149.445 ;
        RECT 101.080 149.415 102.155 149.585 ;
        RECT 100.415 148.815 100.785 149.275 ;
        RECT 101.080 149.075 101.250 149.415 ;
        RECT 101.420 148.815 101.750 149.245 ;
        RECT 101.985 149.075 102.155 149.415 ;
        RECT 102.325 149.315 102.495 150.095 ;
        RECT 102.665 149.875 102.835 150.465 ;
        RECT 103.005 150.065 103.355 150.685 ;
        RECT 102.665 149.485 103.130 149.875 ;
        RECT 103.525 149.615 103.695 150.975 ;
        RECT 103.865 149.785 104.325 150.835 ;
        RECT 103.300 149.445 103.695 149.615 ;
        RECT 103.300 149.315 103.470 149.445 ;
        RECT 102.325 148.985 103.005 149.315 ;
        RECT 103.220 148.985 103.470 149.315 ;
        RECT 103.640 148.815 103.890 149.275 ;
        RECT 104.060 149.000 104.385 149.785 ;
        RECT 104.555 148.985 104.725 151.105 ;
        RECT 104.895 150.985 105.225 151.365 ;
        RECT 105.395 150.815 105.650 151.105 ;
        RECT 104.900 150.645 105.650 150.815 ;
        RECT 104.900 149.655 105.130 150.645 ;
        RECT 105.825 150.615 107.035 151.365 ;
        RECT 105.300 149.825 105.650 150.475 ;
        RECT 105.825 149.905 106.345 150.445 ;
        RECT 106.515 150.075 107.035 150.615 ;
        RECT 107.205 150.565 107.545 151.195 ;
        RECT 107.715 150.565 107.965 151.365 ;
        RECT 108.155 150.715 108.485 151.195 ;
        RECT 108.655 150.905 108.880 151.365 ;
        RECT 109.050 150.715 109.380 151.195 ;
        RECT 107.205 149.955 107.380 150.565 ;
        RECT 108.155 150.545 109.380 150.715 ;
        RECT 110.010 150.585 110.510 151.195 ;
        RECT 111.000 150.735 111.285 151.195 ;
        RECT 111.455 150.905 111.725 151.365 ;
        RECT 107.550 150.205 108.245 150.375 ;
        RECT 108.075 149.955 108.245 150.205 ;
        RECT 108.420 150.175 108.840 150.375 ;
        RECT 109.010 150.175 109.340 150.375 ;
        RECT 109.510 150.175 109.840 150.375 ;
        RECT 110.010 149.955 110.180 150.585 ;
        RECT 111.000 150.565 111.955 150.735 ;
        RECT 110.365 150.125 110.715 150.375 ;
        RECT 104.900 149.485 105.650 149.655 ;
        RECT 104.895 148.815 105.225 149.315 ;
        RECT 105.395 148.985 105.650 149.485 ;
        RECT 105.825 148.815 107.035 149.905 ;
        RECT 107.205 148.985 107.545 149.955 ;
        RECT 107.715 148.815 107.885 149.955 ;
        RECT 108.075 149.785 110.510 149.955 ;
        RECT 110.885 149.835 111.575 150.395 ;
        RECT 108.155 148.815 108.405 149.615 ;
        RECT 109.050 148.985 109.380 149.785 ;
        RECT 109.680 148.815 110.010 149.615 ;
        RECT 110.180 148.985 110.510 149.785 ;
        RECT 111.745 149.665 111.955 150.565 ;
        RECT 111.000 149.445 111.955 149.665 ;
        RECT 112.125 150.395 112.525 151.195 ;
        RECT 112.715 150.735 112.995 151.195 ;
        RECT 113.515 150.905 113.840 151.365 ;
        RECT 112.715 150.565 113.840 150.735 ;
        RECT 114.010 150.625 114.395 151.195 ;
        RECT 114.565 150.640 114.855 151.365 ;
        RECT 115.950 150.655 116.205 151.185 ;
        RECT 116.375 150.905 116.680 151.365 ;
        RECT 116.925 150.985 117.995 151.155 ;
        RECT 113.390 150.455 113.840 150.565 ;
        RECT 112.125 149.835 113.220 150.395 ;
        RECT 113.390 150.125 113.945 150.455 ;
        RECT 111.000 148.985 111.285 149.445 ;
        RECT 111.455 148.815 111.725 149.275 ;
        RECT 112.125 148.985 112.525 149.835 ;
        RECT 113.390 149.665 113.840 150.125 ;
        RECT 114.115 149.955 114.395 150.625 ;
        RECT 115.950 150.005 116.160 150.655 ;
        RECT 116.925 150.630 117.245 150.985 ;
        RECT 116.920 150.455 117.245 150.630 ;
        RECT 116.330 150.155 117.245 150.455 ;
        RECT 117.415 150.415 117.655 150.815 ;
        RECT 117.825 150.755 117.995 150.985 ;
        RECT 118.165 150.925 118.355 151.365 ;
        RECT 118.525 150.915 119.475 151.195 ;
        RECT 119.695 151.005 120.045 151.175 ;
        RECT 117.825 150.585 118.355 150.755 ;
        RECT 116.330 150.125 117.070 150.155 ;
        RECT 112.715 149.445 113.840 149.665 ;
        RECT 112.715 148.985 112.995 149.445 ;
        RECT 113.515 148.815 113.840 149.275 ;
        RECT 114.010 148.985 114.395 149.955 ;
        RECT 114.565 148.815 114.855 149.980 ;
        RECT 115.950 149.125 116.205 150.005 ;
        RECT 116.375 148.815 116.680 149.955 ;
        RECT 116.900 149.535 117.070 150.125 ;
        RECT 117.415 150.045 117.955 150.415 ;
        RECT 118.135 150.305 118.355 150.585 ;
        RECT 118.525 150.135 118.695 150.915 ;
        RECT 118.290 149.965 118.695 150.135 ;
        RECT 118.865 150.125 119.215 150.745 ;
        RECT 118.290 149.875 118.460 149.965 ;
        RECT 119.385 149.955 119.595 150.745 ;
        RECT 117.240 149.705 118.460 149.875 ;
        RECT 118.920 149.795 119.595 149.955 ;
        RECT 116.900 149.365 117.700 149.535 ;
        RECT 117.020 148.815 117.350 149.195 ;
        RECT 117.530 149.075 117.700 149.365 ;
        RECT 118.290 149.325 118.460 149.705 ;
        RECT 118.630 149.785 119.595 149.795 ;
        RECT 119.785 150.615 120.045 151.005 ;
        RECT 120.255 150.905 120.585 151.365 ;
        RECT 121.460 150.975 122.315 151.145 ;
        RECT 122.520 150.975 123.015 151.145 ;
        RECT 123.185 151.005 123.515 151.365 ;
        RECT 119.785 149.925 119.955 150.615 ;
        RECT 120.125 150.265 120.295 150.445 ;
        RECT 120.465 150.435 121.255 150.685 ;
        RECT 121.460 150.265 121.630 150.975 ;
        RECT 121.800 150.465 122.155 150.685 ;
        RECT 120.125 150.095 121.815 150.265 ;
        RECT 118.630 149.495 119.090 149.785 ;
        RECT 119.785 149.755 121.285 149.925 ;
        RECT 119.785 149.615 119.955 149.755 ;
        RECT 119.395 149.445 119.955 149.615 ;
        RECT 117.870 148.815 118.120 149.275 ;
        RECT 118.290 148.985 119.160 149.325 ;
        RECT 119.395 148.985 119.565 149.445 ;
        RECT 120.400 149.415 121.475 149.585 ;
        RECT 119.735 148.815 120.105 149.275 ;
        RECT 120.400 149.075 120.570 149.415 ;
        RECT 120.740 148.815 121.070 149.245 ;
        RECT 121.305 149.075 121.475 149.415 ;
        RECT 121.645 149.315 121.815 150.095 ;
        RECT 121.985 149.875 122.155 150.465 ;
        RECT 122.325 150.065 122.675 150.685 ;
        RECT 121.985 149.485 122.450 149.875 ;
        RECT 122.845 149.615 123.015 150.975 ;
        RECT 123.185 149.785 123.645 150.835 ;
        RECT 122.620 149.445 123.015 149.615 ;
        RECT 122.620 149.315 122.790 149.445 ;
        RECT 121.645 148.985 122.325 149.315 ;
        RECT 122.540 148.985 122.790 149.315 ;
        RECT 122.960 148.815 123.210 149.275 ;
        RECT 123.380 149.000 123.705 149.785 ;
        RECT 123.875 148.985 124.045 151.105 ;
        RECT 124.215 150.985 124.545 151.365 ;
        RECT 124.715 150.815 124.970 151.105 ;
        RECT 124.220 150.645 124.970 150.815 ;
        RECT 124.220 149.655 124.450 150.645 ;
        RECT 125.145 150.615 126.355 151.365 ;
        RECT 126.525 150.615 127.735 151.365 ;
        RECT 124.620 149.825 124.970 150.475 ;
        RECT 125.145 149.905 125.665 150.445 ;
        RECT 125.835 150.075 126.355 150.615 ;
        RECT 126.525 149.905 127.045 150.445 ;
        RECT 127.215 150.075 127.735 150.615 ;
        RECT 124.220 149.485 124.970 149.655 ;
        RECT 124.215 148.815 124.545 149.315 ;
        RECT 124.715 148.985 124.970 149.485 ;
        RECT 125.145 148.815 126.355 149.905 ;
        RECT 126.525 148.815 127.735 149.905 ;
        RECT 14.660 148.645 127.820 148.815 ;
        RECT 14.745 147.555 15.955 148.645 ;
        RECT 14.745 146.845 15.265 147.385 ;
        RECT 15.435 147.015 15.955 147.555 ;
        RECT 16.585 147.555 20.095 148.645 ;
        RECT 20.265 147.885 20.780 148.295 ;
        RECT 21.015 147.885 21.185 148.645 ;
        RECT 21.355 148.305 23.385 148.475 ;
        RECT 16.585 147.035 18.275 147.555 ;
        RECT 18.445 146.865 20.095 147.385 ;
        RECT 20.265 147.075 20.605 147.885 ;
        RECT 21.355 147.640 21.525 148.305 ;
        RECT 21.920 147.965 23.045 148.135 ;
        RECT 20.775 147.450 21.525 147.640 ;
        RECT 21.695 147.625 22.705 147.795 ;
        RECT 20.265 146.905 21.495 147.075 ;
        RECT 14.745 146.095 15.955 146.845 ;
        RECT 16.585 146.095 20.095 146.865 ;
        RECT 20.540 146.300 20.785 146.905 ;
        RECT 21.005 146.095 21.515 146.630 ;
        RECT 21.695 146.265 21.885 147.625 ;
        RECT 22.055 146.945 22.330 147.425 ;
        RECT 22.055 146.775 22.335 146.945 ;
        RECT 22.535 146.825 22.705 147.625 ;
        RECT 22.875 146.835 23.045 147.965 ;
        RECT 23.215 147.335 23.385 148.305 ;
        RECT 23.555 147.505 23.725 148.645 ;
        RECT 23.895 147.505 24.230 148.475 ;
        RECT 23.215 147.005 23.410 147.335 ;
        RECT 23.635 147.005 23.890 147.335 ;
        RECT 23.635 146.835 23.805 147.005 ;
        RECT 24.060 146.835 24.230 147.505 ;
        RECT 24.405 147.480 24.695 148.645 ;
        RECT 24.865 147.570 25.135 148.475 ;
        RECT 25.305 147.885 25.635 148.645 ;
        RECT 25.815 147.715 25.985 148.475 ;
        RECT 22.055 146.265 22.330 146.775 ;
        RECT 22.875 146.665 23.805 146.835 ;
        RECT 22.875 146.630 23.050 146.665 ;
        RECT 22.520 146.265 23.050 146.630 ;
        RECT 23.475 146.095 23.805 146.495 ;
        RECT 23.975 146.265 24.230 146.835 ;
        RECT 24.405 146.095 24.695 146.820 ;
        RECT 24.865 146.770 25.035 147.570 ;
        RECT 25.320 147.545 25.985 147.715 ;
        RECT 26.245 147.555 27.915 148.645 ;
        RECT 28.175 147.715 28.345 148.475 ;
        RECT 28.525 147.885 28.855 148.645 ;
        RECT 25.320 147.400 25.490 147.545 ;
        RECT 25.205 147.070 25.490 147.400 ;
        RECT 25.320 146.815 25.490 147.070 ;
        RECT 25.725 146.995 26.055 147.365 ;
        RECT 26.245 147.035 26.995 147.555 ;
        RECT 28.175 147.545 28.840 147.715 ;
        RECT 29.025 147.570 29.295 148.475 ;
        RECT 28.670 147.400 28.840 147.545 ;
        RECT 27.165 146.865 27.915 147.385 ;
        RECT 28.105 146.995 28.435 147.365 ;
        RECT 28.670 147.070 28.955 147.400 ;
        RECT 24.865 146.265 25.125 146.770 ;
        RECT 25.320 146.645 25.985 146.815 ;
        RECT 25.305 146.095 25.635 146.475 ;
        RECT 25.815 146.265 25.985 146.645 ;
        RECT 26.245 146.095 27.915 146.865 ;
        RECT 28.670 146.815 28.840 147.070 ;
        RECT 28.175 146.645 28.840 146.815 ;
        RECT 29.125 146.770 29.295 147.570 ;
        RECT 28.175 146.265 28.345 146.645 ;
        RECT 28.525 146.095 28.855 146.475 ;
        RECT 29.035 146.265 29.295 146.770 ;
        RECT 29.470 147.505 29.805 148.475 ;
        RECT 29.975 147.505 30.145 148.645 ;
        RECT 30.315 148.305 32.345 148.475 ;
        RECT 29.470 146.835 29.640 147.505 ;
        RECT 30.315 147.335 30.485 148.305 ;
        RECT 29.810 147.005 30.065 147.335 ;
        RECT 30.290 147.005 30.485 147.335 ;
        RECT 30.655 147.965 31.780 148.135 ;
        RECT 29.895 146.835 30.065 147.005 ;
        RECT 30.655 146.835 30.825 147.965 ;
        RECT 29.470 146.265 29.725 146.835 ;
        RECT 29.895 146.665 30.825 146.835 ;
        RECT 30.995 147.625 32.005 147.795 ;
        RECT 30.995 146.825 31.165 147.625 ;
        RECT 31.370 147.285 31.645 147.425 ;
        RECT 31.365 147.115 31.645 147.285 ;
        RECT 30.650 146.630 30.825 146.665 ;
        RECT 29.895 146.095 30.225 146.495 ;
        RECT 30.650 146.265 31.180 146.630 ;
        RECT 31.370 146.265 31.645 147.115 ;
        RECT 31.815 146.265 32.005 147.625 ;
        RECT 32.175 147.640 32.345 148.305 ;
        RECT 32.515 147.885 32.685 148.645 ;
        RECT 32.920 147.885 33.435 148.295 ;
        RECT 32.175 147.450 32.925 147.640 ;
        RECT 33.095 147.075 33.435 147.885 ;
        RECT 32.205 146.905 33.435 147.075 ;
        RECT 34.065 147.555 35.735 148.645 ;
        RECT 36.110 147.675 36.440 148.475 ;
        RECT 36.610 147.845 36.940 148.645 ;
        RECT 37.240 147.675 37.570 148.475 ;
        RECT 38.215 147.845 38.465 148.645 ;
        RECT 34.065 147.035 34.815 147.555 ;
        RECT 36.110 147.505 38.545 147.675 ;
        RECT 38.735 147.505 38.905 148.645 ;
        RECT 39.075 147.505 39.415 148.475 ;
        RECT 32.185 146.095 32.695 146.630 ;
        RECT 32.915 146.300 33.160 146.905 ;
        RECT 34.985 146.865 35.735 147.385 ;
        RECT 35.905 147.085 36.255 147.335 ;
        RECT 36.440 146.875 36.610 147.505 ;
        RECT 36.780 147.085 37.110 147.285 ;
        RECT 37.280 147.085 37.610 147.285 ;
        RECT 37.780 147.085 38.200 147.285 ;
        RECT 38.375 147.255 38.545 147.505 ;
        RECT 38.375 147.085 39.070 147.255 ;
        RECT 34.065 146.095 35.735 146.865 ;
        RECT 36.110 146.265 36.610 146.875 ;
        RECT 37.240 146.745 38.465 146.915 ;
        RECT 39.240 146.895 39.415 147.505 ;
        RECT 37.240 146.265 37.570 146.745 ;
        RECT 37.740 146.095 37.965 146.555 ;
        RECT 38.135 146.265 38.465 146.745 ;
        RECT 38.655 146.095 38.905 146.895 ;
        RECT 39.075 146.265 39.415 146.895 ;
        RECT 39.585 147.505 39.925 148.475 ;
        RECT 40.095 147.505 40.265 148.645 ;
        RECT 40.535 147.845 40.785 148.645 ;
        RECT 41.430 147.675 41.760 148.475 ;
        RECT 42.060 147.845 42.390 148.645 ;
        RECT 42.560 147.675 42.890 148.475 ;
        RECT 40.455 147.505 42.890 147.675 ;
        RECT 43.725 147.555 47.235 148.645 ;
        RECT 47.410 148.135 49.065 148.425 ;
        RECT 47.410 147.795 49.000 147.965 ;
        RECT 49.235 147.845 49.515 148.645 ;
        RECT 39.585 146.945 39.760 147.505 ;
        RECT 40.455 147.255 40.625 147.505 ;
        RECT 39.930 147.085 40.625 147.255 ;
        RECT 40.800 147.085 41.220 147.285 ;
        RECT 41.390 147.085 41.720 147.285 ;
        RECT 41.890 147.085 42.220 147.285 ;
        RECT 39.585 146.895 39.815 146.945 ;
        RECT 39.585 146.265 39.925 146.895 ;
        RECT 40.095 146.095 40.345 146.895 ;
        RECT 40.535 146.745 41.760 146.915 ;
        RECT 40.535 146.265 40.865 146.745 ;
        RECT 41.035 146.095 41.260 146.555 ;
        RECT 41.430 146.265 41.760 146.745 ;
        RECT 42.390 146.875 42.560 147.505 ;
        RECT 42.745 147.085 43.095 147.335 ;
        RECT 43.725 147.035 45.415 147.555 ;
        RECT 47.410 147.505 47.730 147.795 ;
        RECT 48.830 147.675 49.000 147.795 ;
        RECT 42.390 146.265 42.890 146.875 ;
        RECT 45.585 146.865 47.235 147.385 ;
        RECT 43.725 146.095 47.235 146.865 ;
        RECT 47.410 146.765 47.760 147.335 ;
        RECT 47.930 147.005 48.640 147.625 ;
        RECT 48.830 147.505 49.555 147.675 ;
        RECT 49.725 147.505 49.995 148.475 ;
        RECT 49.385 147.335 49.555 147.505 ;
        RECT 48.810 147.005 49.215 147.335 ;
        RECT 49.385 147.005 49.655 147.335 ;
        RECT 49.385 146.835 49.555 147.005 ;
        RECT 47.945 146.665 49.555 146.835 ;
        RECT 49.825 146.770 49.995 147.505 ;
        RECT 50.165 147.480 50.455 148.645 ;
        RECT 51.085 147.570 51.355 148.475 ;
        RECT 51.525 147.885 51.855 148.645 ;
        RECT 52.035 147.715 52.205 148.475 ;
        RECT 47.415 146.095 47.745 146.595 ;
        RECT 47.945 146.315 48.115 146.665 ;
        RECT 48.315 146.095 48.645 146.495 ;
        RECT 48.815 146.315 48.985 146.665 ;
        RECT 49.155 146.095 49.535 146.495 ;
        RECT 49.725 146.425 49.995 146.770 ;
        RECT 50.165 146.095 50.455 146.820 ;
        RECT 51.085 146.770 51.255 147.570 ;
        RECT 51.540 147.545 52.205 147.715 ;
        RECT 51.540 147.400 51.710 147.545 ;
        RECT 51.425 147.070 51.710 147.400 ;
        RECT 53.385 147.505 53.725 148.475 ;
        RECT 53.895 147.505 54.065 148.645 ;
        RECT 54.335 147.845 54.585 148.645 ;
        RECT 55.230 147.675 55.560 148.475 ;
        RECT 55.860 147.845 56.190 148.645 ;
        RECT 56.360 147.675 56.690 148.475 ;
        RECT 54.255 147.505 56.690 147.675 ;
        RECT 57.065 147.555 59.655 148.645 ;
        RECT 59.825 147.885 60.340 148.295 ;
        RECT 60.575 147.885 60.745 148.645 ;
        RECT 60.915 148.305 62.945 148.475 ;
        RECT 51.540 146.815 51.710 147.070 ;
        RECT 51.945 146.995 52.275 147.365 ;
        RECT 53.385 146.895 53.560 147.505 ;
        RECT 54.255 147.255 54.425 147.505 ;
        RECT 53.730 147.085 54.425 147.255 ;
        RECT 54.600 147.085 55.020 147.285 ;
        RECT 55.190 147.085 55.520 147.285 ;
        RECT 55.690 147.085 56.020 147.285 ;
        RECT 51.085 146.265 51.345 146.770 ;
        RECT 51.540 146.645 52.205 146.815 ;
        RECT 51.525 146.095 51.855 146.475 ;
        RECT 52.035 146.265 52.205 146.645 ;
        RECT 53.385 146.265 53.725 146.895 ;
        RECT 53.895 146.095 54.145 146.895 ;
        RECT 54.335 146.745 55.560 146.915 ;
        RECT 54.335 146.265 54.665 146.745 ;
        RECT 54.835 146.095 55.060 146.555 ;
        RECT 55.230 146.265 55.560 146.745 ;
        RECT 56.190 146.875 56.360 147.505 ;
        RECT 56.545 147.085 56.895 147.335 ;
        RECT 57.065 147.035 58.275 147.555 ;
        RECT 56.190 146.265 56.690 146.875 ;
        RECT 58.445 146.865 59.655 147.385 ;
        RECT 59.825 147.075 60.165 147.885 ;
        RECT 60.915 147.640 61.085 148.305 ;
        RECT 61.480 147.965 62.605 148.135 ;
        RECT 60.335 147.450 61.085 147.640 ;
        RECT 61.255 147.625 62.265 147.795 ;
        RECT 59.825 146.905 61.055 147.075 ;
        RECT 57.065 146.095 59.655 146.865 ;
        RECT 60.100 146.300 60.345 146.905 ;
        RECT 60.565 146.095 61.075 146.630 ;
        RECT 61.255 146.265 61.445 147.625 ;
        RECT 61.615 146.605 61.890 147.425 ;
        RECT 62.095 146.825 62.265 147.625 ;
        RECT 62.435 146.835 62.605 147.965 ;
        RECT 62.775 147.335 62.945 148.305 ;
        RECT 63.115 147.505 63.285 148.645 ;
        RECT 63.455 147.505 63.790 148.475 ;
        RECT 62.775 147.005 62.970 147.335 ;
        RECT 63.195 147.005 63.450 147.335 ;
        RECT 63.195 146.835 63.365 147.005 ;
        RECT 63.620 146.835 63.790 147.505 ;
        RECT 63.965 147.555 65.175 148.645 ;
        RECT 65.350 148.210 70.695 148.645 ;
        RECT 63.965 147.015 64.485 147.555 ;
        RECT 64.655 146.845 65.175 147.385 ;
        RECT 66.940 146.960 67.290 148.210 ;
        RECT 70.870 147.495 71.130 148.645 ;
        RECT 71.305 147.570 71.560 148.475 ;
        RECT 71.730 147.885 72.060 148.645 ;
        RECT 72.275 147.715 72.445 148.475 ;
        RECT 62.435 146.665 63.365 146.835 ;
        RECT 62.435 146.630 62.610 146.665 ;
        RECT 61.615 146.435 61.895 146.605 ;
        RECT 61.615 146.265 61.890 146.435 ;
        RECT 62.080 146.265 62.610 146.630 ;
        RECT 63.035 146.095 63.365 146.495 ;
        RECT 63.535 146.265 63.790 146.835 ;
        RECT 63.965 146.095 65.175 146.845 ;
        RECT 68.770 146.640 69.110 147.470 ;
        RECT 65.350 146.095 70.695 146.640 ;
        RECT 70.870 146.095 71.130 146.935 ;
        RECT 71.305 146.840 71.475 147.570 ;
        RECT 71.730 147.545 72.445 147.715 ;
        RECT 72.795 147.715 72.965 148.475 ;
        RECT 73.180 147.885 73.510 148.645 ;
        RECT 72.795 147.545 73.510 147.715 ;
        RECT 73.680 147.570 73.935 148.475 ;
        RECT 71.730 147.335 71.900 147.545 ;
        RECT 71.645 147.005 71.900 147.335 ;
        RECT 71.305 146.265 71.560 146.840 ;
        RECT 71.730 146.815 71.900 147.005 ;
        RECT 72.180 146.995 72.535 147.365 ;
        RECT 72.705 146.995 73.060 147.365 ;
        RECT 73.340 147.335 73.510 147.545 ;
        RECT 73.340 147.005 73.595 147.335 ;
        RECT 73.340 146.815 73.510 147.005 ;
        RECT 73.765 146.840 73.935 147.570 ;
        RECT 74.110 147.495 74.370 148.645 ;
        RECT 74.545 147.555 75.755 148.645 ;
        RECT 74.545 147.015 75.065 147.555 ;
        RECT 75.925 147.480 76.215 148.645 ;
        RECT 76.590 147.675 76.920 148.475 ;
        RECT 77.090 147.845 77.420 148.645 ;
        RECT 77.720 147.675 78.050 148.475 ;
        RECT 78.695 147.845 78.945 148.645 ;
        RECT 76.590 147.505 79.025 147.675 ;
        RECT 79.215 147.505 79.385 148.645 ;
        RECT 79.555 147.505 79.895 148.475 ;
        RECT 71.730 146.645 72.445 146.815 ;
        RECT 71.730 146.095 72.060 146.475 ;
        RECT 72.275 146.265 72.445 146.645 ;
        RECT 72.795 146.645 73.510 146.815 ;
        RECT 72.795 146.265 72.965 146.645 ;
        RECT 73.180 146.095 73.510 146.475 ;
        RECT 73.680 146.265 73.935 146.840 ;
        RECT 74.110 146.095 74.370 146.935 ;
        RECT 75.235 146.845 75.755 147.385 ;
        RECT 76.385 147.085 76.735 147.335 ;
        RECT 76.920 146.875 77.090 147.505 ;
        RECT 77.260 147.085 77.590 147.285 ;
        RECT 77.760 147.085 78.090 147.285 ;
        RECT 78.260 147.085 78.680 147.285 ;
        RECT 78.855 147.255 79.025 147.505 ;
        RECT 78.855 147.085 79.550 147.255 ;
        RECT 74.545 146.095 75.755 146.845 ;
        RECT 75.925 146.095 76.215 146.820 ;
        RECT 76.590 146.265 77.090 146.875 ;
        RECT 77.720 146.745 78.945 146.915 ;
        RECT 79.720 146.895 79.895 147.505 ;
        RECT 77.720 146.265 78.050 146.745 ;
        RECT 78.220 146.095 78.445 146.555 ;
        RECT 78.615 146.265 78.945 146.745 ;
        RECT 79.135 146.095 79.385 146.895 ;
        RECT 79.555 146.265 79.895 146.895 ;
        RECT 80.065 147.505 80.405 148.475 ;
        RECT 80.575 147.505 80.745 148.645 ;
        RECT 81.015 147.845 81.265 148.645 ;
        RECT 81.910 147.675 82.240 148.475 ;
        RECT 82.540 147.845 82.870 148.645 ;
        RECT 83.040 147.675 83.370 148.475 ;
        RECT 80.935 147.505 83.370 147.675 ;
        RECT 83.745 147.555 84.955 148.645 ;
        RECT 85.500 147.665 85.755 148.335 ;
        RECT 85.935 147.845 86.220 148.645 ;
        RECT 86.400 147.925 86.730 148.435 ;
        RECT 80.065 146.895 80.240 147.505 ;
        RECT 80.935 147.255 81.105 147.505 ;
        RECT 80.410 147.085 81.105 147.255 ;
        RECT 81.280 147.085 81.700 147.285 ;
        RECT 81.870 147.085 82.200 147.285 ;
        RECT 82.370 147.085 82.700 147.285 ;
        RECT 80.065 146.265 80.405 146.895 ;
        RECT 80.575 146.095 80.825 146.895 ;
        RECT 81.015 146.745 82.240 146.915 ;
        RECT 81.015 146.265 81.345 146.745 ;
        RECT 81.515 146.095 81.740 146.555 ;
        RECT 81.910 146.265 82.240 146.745 ;
        RECT 82.870 146.875 83.040 147.505 ;
        RECT 83.225 147.085 83.575 147.335 ;
        RECT 83.745 147.015 84.265 147.555 ;
        RECT 82.870 146.265 83.370 146.875 ;
        RECT 84.435 146.845 84.955 147.385 ;
        RECT 83.745 146.095 84.955 146.845 ;
        RECT 85.500 146.805 85.680 147.665 ;
        RECT 86.400 147.335 86.650 147.925 ;
        RECT 87.000 147.775 87.170 148.385 ;
        RECT 87.340 147.955 87.670 148.645 ;
        RECT 87.900 148.095 88.140 148.385 ;
        RECT 88.340 148.265 88.760 148.645 ;
        RECT 88.940 148.175 89.570 148.425 ;
        RECT 90.040 148.265 90.370 148.645 ;
        RECT 88.940 148.095 89.110 148.175 ;
        RECT 90.540 148.095 90.710 148.385 ;
        RECT 90.890 148.265 91.270 148.645 ;
        RECT 91.510 148.260 92.340 148.430 ;
        RECT 87.900 147.925 89.110 148.095 ;
        RECT 85.850 147.005 86.650 147.335 ;
        RECT 85.500 146.605 85.755 146.805 ;
        RECT 85.415 146.435 85.755 146.605 ;
        RECT 85.500 146.275 85.755 146.435 ;
        RECT 85.935 146.095 86.220 146.555 ;
        RECT 86.400 146.355 86.650 147.005 ;
        RECT 86.850 147.755 87.170 147.775 ;
        RECT 86.850 147.585 88.770 147.755 ;
        RECT 86.850 146.690 87.040 147.585 ;
        RECT 88.940 147.415 89.110 147.925 ;
        RECT 89.280 147.665 89.800 147.975 ;
        RECT 87.210 147.245 89.110 147.415 ;
        RECT 87.210 147.185 87.540 147.245 ;
        RECT 87.690 147.015 88.020 147.075 ;
        RECT 87.360 146.745 88.020 147.015 ;
        RECT 86.850 146.360 87.170 146.690 ;
        RECT 87.350 146.095 88.010 146.575 ;
        RECT 88.210 146.485 88.380 147.245 ;
        RECT 89.280 147.075 89.460 147.485 ;
        RECT 88.550 146.905 88.880 147.025 ;
        RECT 89.630 146.905 89.800 147.665 ;
        RECT 88.550 146.735 89.800 146.905 ;
        RECT 89.970 147.845 91.340 148.095 ;
        RECT 89.970 147.075 90.160 147.845 ;
        RECT 91.090 147.585 91.340 147.845 ;
        RECT 90.330 147.415 90.580 147.575 ;
        RECT 91.510 147.415 91.680 148.260 ;
        RECT 92.575 147.975 92.745 148.475 ;
        RECT 92.915 148.145 93.245 148.645 ;
        RECT 91.850 147.585 92.350 147.965 ;
        RECT 92.575 147.805 93.270 147.975 ;
        RECT 90.330 147.245 91.680 147.415 ;
        RECT 91.260 147.205 91.680 147.245 ;
        RECT 89.970 146.735 90.390 147.075 ;
        RECT 90.680 146.745 91.090 147.075 ;
        RECT 88.210 146.315 89.060 146.485 ;
        RECT 89.620 146.095 89.940 146.555 ;
        RECT 90.140 146.305 90.390 146.735 ;
        RECT 90.680 146.095 91.090 146.535 ;
        RECT 91.260 146.475 91.430 147.205 ;
        RECT 91.600 146.655 91.950 147.025 ;
        RECT 92.130 146.715 92.350 147.585 ;
        RECT 92.520 147.015 92.930 147.635 ;
        RECT 93.100 146.835 93.270 147.805 ;
        RECT 92.575 146.645 93.270 146.835 ;
        RECT 91.260 146.275 92.275 146.475 ;
        RECT 92.575 146.315 92.745 146.645 ;
        RECT 92.915 146.095 93.245 146.475 ;
        RECT 93.460 146.355 93.685 148.475 ;
        RECT 93.855 148.145 94.185 148.645 ;
        RECT 94.355 147.975 94.525 148.475 ;
        RECT 93.860 147.805 94.525 147.975 ;
        RECT 93.860 146.815 94.090 147.805 ;
        RECT 94.260 146.985 94.610 147.635 ;
        RECT 95.285 147.505 95.515 148.645 ;
        RECT 95.685 147.495 96.015 148.475 ;
        RECT 96.185 147.505 96.395 148.645 ;
        RECT 96.625 147.885 97.140 148.295 ;
        RECT 97.375 147.885 97.545 148.645 ;
        RECT 97.715 148.305 99.745 148.475 ;
        RECT 95.265 147.085 95.595 147.335 ;
        RECT 93.860 146.645 94.525 146.815 ;
        RECT 93.855 146.095 94.185 146.475 ;
        RECT 94.355 146.355 94.525 146.645 ;
        RECT 95.285 146.095 95.515 146.915 ;
        RECT 95.765 146.895 96.015 147.495 ;
        RECT 96.625 147.075 96.965 147.885 ;
        RECT 97.715 147.640 97.885 148.305 ;
        RECT 98.280 147.965 99.405 148.135 ;
        RECT 97.135 147.450 97.885 147.640 ;
        RECT 98.055 147.625 99.065 147.795 ;
        RECT 95.685 146.265 96.015 146.895 ;
        RECT 96.185 146.095 96.395 146.915 ;
        RECT 96.625 146.905 97.855 147.075 ;
        RECT 96.900 146.300 97.145 146.905 ;
        RECT 97.365 146.095 97.875 146.630 ;
        RECT 98.055 146.265 98.245 147.625 ;
        RECT 98.415 147.285 98.690 147.425 ;
        RECT 98.415 147.115 98.695 147.285 ;
        RECT 98.415 146.265 98.690 147.115 ;
        RECT 98.895 146.825 99.065 147.625 ;
        RECT 99.235 146.835 99.405 147.965 ;
        RECT 99.575 147.335 99.745 148.305 ;
        RECT 99.915 147.505 100.085 148.645 ;
        RECT 100.255 147.505 100.590 148.475 ;
        RECT 99.575 147.005 99.770 147.335 ;
        RECT 99.995 147.005 100.250 147.335 ;
        RECT 99.995 146.835 100.165 147.005 ;
        RECT 100.420 146.835 100.590 147.505 ;
        RECT 101.685 147.480 101.975 148.645 ;
        RECT 102.235 147.715 102.405 148.475 ;
        RECT 102.585 147.885 102.915 148.645 ;
        RECT 102.235 147.545 102.900 147.715 ;
        RECT 103.085 147.570 103.355 148.475 ;
        RECT 102.730 147.400 102.900 147.545 ;
        RECT 102.165 146.995 102.495 147.365 ;
        RECT 102.730 147.070 103.015 147.400 ;
        RECT 99.235 146.665 100.165 146.835 ;
        RECT 99.235 146.630 99.410 146.665 ;
        RECT 98.880 146.265 99.410 146.630 ;
        RECT 99.835 146.095 100.165 146.495 ;
        RECT 100.335 146.265 100.590 146.835 ;
        RECT 101.685 146.095 101.975 146.820 ;
        RECT 102.730 146.815 102.900 147.070 ;
        RECT 102.235 146.645 102.900 146.815 ;
        RECT 103.185 146.770 103.355 147.570 ;
        RECT 102.235 146.265 102.405 146.645 ;
        RECT 102.585 146.095 102.915 146.475 ;
        RECT 103.095 146.265 103.355 146.770 ;
        RECT 103.985 147.505 104.255 148.475 ;
        RECT 104.465 147.845 104.745 148.645 ;
        RECT 104.915 148.135 106.570 148.425 ;
        RECT 104.980 147.795 106.570 147.965 ;
        RECT 104.980 147.675 105.150 147.795 ;
        RECT 104.425 147.505 105.150 147.675 ;
        RECT 103.985 146.770 104.155 147.505 ;
        RECT 104.425 147.335 104.595 147.505 ;
        RECT 105.340 147.455 106.055 147.625 ;
        RECT 106.250 147.505 106.570 147.795 ;
        RECT 106.745 147.505 107.085 148.475 ;
        RECT 107.255 147.505 107.425 148.645 ;
        RECT 107.695 147.845 107.945 148.645 ;
        RECT 108.590 147.675 108.920 148.475 ;
        RECT 109.220 147.845 109.550 148.645 ;
        RECT 109.720 147.675 110.050 148.475 ;
        RECT 107.615 147.505 110.050 147.675 ;
        RECT 110.425 147.555 112.095 148.645 ;
        RECT 112.265 147.885 112.780 148.295 ;
        RECT 113.015 147.885 113.185 148.645 ;
        RECT 113.355 148.305 115.385 148.475 ;
        RECT 104.325 147.005 104.595 147.335 ;
        RECT 104.765 147.005 105.170 147.335 ;
        RECT 105.340 147.005 106.050 147.455 ;
        RECT 104.425 146.835 104.595 147.005 ;
        RECT 103.985 146.425 104.255 146.770 ;
        RECT 104.425 146.665 106.035 146.835 ;
        RECT 106.220 146.765 106.570 147.335 ;
        RECT 106.745 146.945 106.920 147.505 ;
        RECT 107.615 147.255 107.785 147.505 ;
        RECT 107.090 147.085 107.785 147.255 ;
        RECT 107.960 147.085 108.380 147.285 ;
        RECT 108.550 147.085 108.880 147.285 ;
        RECT 109.050 147.085 109.380 147.285 ;
        RECT 106.745 146.895 106.975 146.945 ;
        RECT 104.445 146.095 104.825 146.495 ;
        RECT 104.995 146.315 105.165 146.665 ;
        RECT 105.335 146.095 105.665 146.495 ;
        RECT 105.865 146.315 106.035 146.665 ;
        RECT 106.235 146.095 106.565 146.595 ;
        RECT 106.745 146.265 107.085 146.895 ;
        RECT 107.255 146.095 107.505 146.895 ;
        RECT 107.695 146.745 108.920 146.915 ;
        RECT 107.695 146.265 108.025 146.745 ;
        RECT 108.195 146.095 108.420 146.555 ;
        RECT 108.590 146.265 108.920 146.745 ;
        RECT 109.550 146.875 109.720 147.505 ;
        RECT 109.905 147.085 110.255 147.335 ;
        RECT 110.425 147.035 111.175 147.555 ;
        RECT 109.550 146.265 110.050 146.875 ;
        RECT 111.345 146.865 112.095 147.385 ;
        RECT 112.265 147.075 112.605 147.885 ;
        RECT 113.355 147.640 113.525 148.305 ;
        RECT 113.920 147.965 115.045 148.135 ;
        RECT 112.775 147.450 113.525 147.640 ;
        RECT 113.695 147.625 114.705 147.795 ;
        RECT 112.265 146.905 113.495 147.075 ;
        RECT 110.425 146.095 112.095 146.865 ;
        RECT 112.540 146.300 112.785 146.905 ;
        RECT 113.005 146.095 113.515 146.630 ;
        RECT 113.695 146.265 113.885 147.625 ;
        RECT 114.055 147.285 114.330 147.425 ;
        RECT 114.055 147.115 114.335 147.285 ;
        RECT 114.055 146.265 114.330 147.115 ;
        RECT 114.535 146.825 114.705 147.625 ;
        RECT 114.875 146.835 115.045 147.965 ;
        RECT 115.215 147.335 115.385 148.305 ;
        RECT 115.555 147.505 115.725 148.645 ;
        RECT 115.895 147.505 116.230 148.475 ;
        RECT 115.215 147.005 115.410 147.335 ;
        RECT 115.635 147.005 115.890 147.335 ;
        RECT 115.635 146.835 115.805 147.005 ;
        RECT 116.060 146.835 116.230 147.505 ;
        RECT 116.780 147.665 117.035 148.335 ;
        RECT 117.215 147.845 117.500 148.645 ;
        RECT 117.680 147.925 118.010 148.435 ;
        RECT 116.780 146.945 116.960 147.665 ;
        RECT 117.680 147.335 117.930 147.925 ;
        RECT 118.280 147.775 118.450 148.385 ;
        RECT 118.620 147.955 118.950 148.645 ;
        RECT 119.180 148.095 119.420 148.385 ;
        RECT 119.620 148.265 120.040 148.645 ;
        RECT 120.220 148.175 120.850 148.425 ;
        RECT 121.320 148.265 121.650 148.645 ;
        RECT 120.220 148.095 120.390 148.175 ;
        RECT 121.820 148.095 121.990 148.385 ;
        RECT 122.170 148.265 122.550 148.645 ;
        RECT 122.790 148.260 123.620 148.430 ;
        RECT 119.180 147.925 120.390 148.095 ;
        RECT 117.130 147.005 117.930 147.335 ;
        RECT 114.875 146.665 115.805 146.835 ;
        RECT 114.875 146.630 115.050 146.665 ;
        RECT 114.520 146.265 115.050 146.630 ;
        RECT 115.475 146.095 115.805 146.495 ;
        RECT 115.975 146.265 116.230 146.835 ;
        RECT 116.695 146.805 116.960 146.945 ;
        RECT 116.695 146.775 117.035 146.805 ;
        RECT 116.780 146.275 117.035 146.775 ;
        RECT 117.215 146.095 117.500 146.555 ;
        RECT 117.680 146.355 117.930 147.005 ;
        RECT 118.130 147.755 118.450 147.775 ;
        RECT 118.130 147.585 120.050 147.755 ;
        RECT 118.130 146.690 118.320 147.585 ;
        RECT 120.220 147.415 120.390 147.925 ;
        RECT 120.560 147.665 121.080 147.975 ;
        RECT 118.490 147.245 120.390 147.415 ;
        RECT 118.490 147.185 118.820 147.245 ;
        RECT 118.970 147.015 119.300 147.075 ;
        RECT 118.640 146.745 119.300 147.015 ;
        RECT 118.130 146.360 118.450 146.690 ;
        RECT 118.630 146.095 119.290 146.575 ;
        RECT 119.490 146.485 119.660 147.245 ;
        RECT 120.560 147.075 120.740 147.485 ;
        RECT 119.830 146.905 120.160 147.025 ;
        RECT 120.910 146.905 121.080 147.665 ;
        RECT 119.830 146.735 121.080 146.905 ;
        RECT 121.250 147.845 122.620 148.095 ;
        RECT 121.250 147.075 121.440 147.845 ;
        RECT 122.370 147.585 122.620 147.845 ;
        RECT 121.610 147.415 121.860 147.575 ;
        RECT 122.790 147.415 122.960 148.260 ;
        RECT 123.855 147.975 124.025 148.475 ;
        RECT 124.195 148.145 124.525 148.645 ;
        RECT 123.130 147.585 123.630 147.965 ;
        RECT 123.855 147.805 124.550 147.975 ;
        RECT 121.610 147.245 122.960 147.415 ;
        RECT 122.540 147.205 122.960 147.245 ;
        RECT 121.250 146.735 121.670 147.075 ;
        RECT 121.960 146.745 122.370 147.075 ;
        RECT 119.490 146.315 120.340 146.485 ;
        RECT 120.900 146.095 121.220 146.555 ;
        RECT 121.420 146.305 121.670 146.735 ;
        RECT 121.960 146.095 122.370 146.535 ;
        RECT 122.540 146.475 122.710 147.205 ;
        RECT 122.880 146.655 123.230 147.025 ;
        RECT 123.410 146.715 123.630 147.585 ;
        RECT 123.800 147.015 124.210 147.635 ;
        RECT 124.380 146.835 124.550 147.805 ;
        RECT 123.855 146.645 124.550 146.835 ;
        RECT 122.540 146.275 123.555 146.475 ;
        RECT 123.855 146.315 124.025 146.645 ;
        RECT 124.195 146.095 124.525 146.475 ;
        RECT 124.740 146.355 124.965 148.475 ;
        RECT 125.135 148.145 125.465 148.645 ;
        RECT 125.635 147.975 125.805 148.475 ;
        RECT 125.140 147.805 125.805 147.975 ;
        RECT 125.140 146.815 125.370 147.805 ;
        RECT 125.540 146.985 125.890 147.635 ;
        RECT 126.525 147.555 127.735 148.645 ;
        RECT 126.525 147.015 127.045 147.555 ;
        RECT 127.215 146.845 127.735 147.385 ;
        RECT 125.140 146.645 125.805 146.815 ;
        RECT 125.135 146.095 125.465 146.475 ;
        RECT 125.635 146.355 125.805 146.645 ;
        RECT 126.525 146.095 127.735 146.845 ;
        RECT 14.660 145.925 127.820 146.095 ;
        RECT 14.745 145.175 15.955 145.925 ;
        RECT 14.745 144.635 15.265 145.175 ;
        RECT 16.125 145.155 19.635 145.925 ;
        RECT 15.435 144.465 15.955 145.005 ;
        RECT 14.745 143.375 15.955 144.465 ;
        RECT 16.125 144.465 17.815 144.985 ;
        RECT 17.985 144.635 19.635 145.155 ;
        RECT 19.845 145.105 20.075 145.925 ;
        RECT 20.245 145.125 20.575 145.755 ;
        RECT 19.825 144.685 20.155 144.935 ;
        RECT 20.325 144.525 20.575 145.125 ;
        RECT 20.745 145.105 20.955 145.925 ;
        RECT 21.225 145.105 21.455 145.925 ;
        RECT 21.625 145.125 21.955 145.755 ;
        RECT 21.205 144.685 21.535 144.935 ;
        RECT 21.705 144.525 21.955 145.125 ;
        RECT 22.125 145.105 22.335 145.925 ;
        RECT 22.940 145.585 23.195 145.745 ;
        RECT 22.855 145.415 23.195 145.585 ;
        RECT 23.375 145.465 23.660 145.925 ;
        RECT 22.940 145.215 23.195 145.415 ;
        RECT 16.125 143.375 19.635 144.465 ;
        RECT 19.845 143.375 20.075 144.515 ;
        RECT 20.245 143.545 20.575 144.525 ;
        RECT 20.745 143.375 20.955 144.515 ;
        RECT 21.225 143.375 21.455 144.515 ;
        RECT 21.625 143.545 21.955 144.525 ;
        RECT 22.125 143.375 22.335 144.515 ;
        RECT 22.940 144.355 23.120 145.215 ;
        RECT 23.840 145.015 24.090 145.665 ;
        RECT 23.290 144.685 24.090 145.015 ;
        RECT 22.940 143.685 23.195 144.355 ;
        RECT 23.375 143.375 23.660 144.175 ;
        RECT 23.840 144.095 24.090 144.685 ;
        RECT 24.290 145.330 24.610 145.660 ;
        RECT 24.790 145.445 25.450 145.925 ;
        RECT 25.650 145.535 26.500 145.705 ;
        RECT 24.290 144.435 24.480 145.330 ;
        RECT 24.800 145.005 25.460 145.275 ;
        RECT 25.130 144.945 25.460 145.005 ;
        RECT 24.650 144.775 24.980 144.835 ;
        RECT 25.650 144.775 25.820 145.535 ;
        RECT 27.060 145.465 27.380 145.925 ;
        RECT 27.580 145.285 27.830 145.715 ;
        RECT 28.120 145.485 28.530 145.925 ;
        RECT 28.700 145.545 29.715 145.745 ;
        RECT 25.990 145.115 27.240 145.285 ;
        RECT 25.990 144.995 26.320 145.115 ;
        RECT 24.650 144.605 26.550 144.775 ;
        RECT 24.290 144.265 26.210 144.435 ;
        RECT 24.290 144.245 24.610 144.265 ;
        RECT 23.840 143.585 24.170 144.095 ;
        RECT 24.440 143.635 24.610 144.245 ;
        RECT 26.380 144.095 26.550 144.605 ;
        RECT 26.720 144.535 26.900 144.945 ;
        RECT 27.070 144.355 27.240 145.115 ;
        RECT 24.780 143.375 25.110 144.065 ;
        RECT 25.340 143.925 26.550 144.095 ;
        RECT 26.720 144.045 27.240 144.355 ;
        RECT 27.410 144.945 27.830 145.285 ;
        RECT 28.120 144.945 28.530 145.275 ;
        RECT 27.410 144.175 27.600 144.945 ;
        RECT 28.700 144.815 28.870 145.545 ;
        RECT 30.015 145.375 30.185 145.705 ;
        RECT 30.355 145.545 30.685 145.925 ;
        RECT 29.040 144.995 29.390 145.365 ;
        RECT 28.700 144.775 29.120 144.815 ;
        RECT 27.770 144.605 29.120 144.775 ;
        RECT 27.770 144.445 28.020 144.605 ;
        RECT 28.530 144.175 28.780 144.435 ;
        RECT 27.410 143.925 28.780 144.175 ;
        RECT 25.340 143.635 25.580 143.925 ;
        RECT 26.380 143.845 26.550 143.925 ;
        RECT 25.780 143.375 26.200 143.755 ;
        RECT 26.380 143.595 27.010 143.845 ;
        RECT 27.480 143.375 27.810 143.755 ;
        RECT 27.980 143.635 28.150 143.925 ;
        RECT 28.950 143.760 29.120 144.605 ;
        RECT 29.570 144.435 29.790 145.305 ;
        RECT 30.015 145.185 30.710 145.375 ;
        RECT 29.290 144.055 29.790 144.435 ;
        RECT 29.960 144.385 30.370 145.005 ;
        RECT 30.540 144.215 30.710 145.185 ;
        RECT 30.015 144.045 30.710 144.215 ;
        RECT 28.330 143.375 28.710 143.755 ;
        RECT 28.950 143.590 29.780 143.760 ;
        RECT 30.015 143.545 30.185 144.045 ;
        RECT 30.355 143.375 30.685 143.875 ;
        RECT 30.900 143.545 31.125 145.665 ;
        RECT 31.295 145.545 31.625 145.925 ;
        RECT 31.795 145.375 31.965 145.665 ;
        RECT 31.300 145.205 31.965 145.375 ;
        RECT 31.300 144.215 31.530 145.205 ;
        RECT 32.225 145.175 33.435 145.925 ;
        RECT 31.700 144.385 32.050 145.035 ;
        RECT 32.225 144.465 32.745 145.005 ;
        RECT 32.915 144.635 33.435 145.175 ;
        RECT 33.605 145.155 37.115 145.925 ;
        RECT 37.285 145.200 37.575 145.925 ;
        RECT 38.205 145.155 40.795 145.925 ;
        RECT 33.605 144.465 35.295 144.985 ;
        RECT 35.465 144.635 37.115 145.155 ;
        RECT 31.300 144.045 31.965 144.215 ;
        RECT 31.295 143.375 31.625 143.875 ;
        RECT 31.795 143.545 31.965 144.045 ;
        RECT 32.225 143.375 33.435 144.465 ;
        RECT 33.605 143.375 37.115 144.465 ;
        RECT 37.285 143.375 37.575 144.540 ;
        RECT 38.205 144.465 39.415 144.985 ;
        RECT 39.585 144.635 40.795 145.155 ;
        RECT 41.005 145.105 41.235 145.925 ;
        RECT 41.405 145.125 41.735 145.755 ;
        RECT 40.985 144.685 41.315 144.935 ;
        RECT 41.485 144.525 41.735 145.125 ;
        RECT 41.905 145.105 42.115 145.925 ;
        RECT 42.720 145.215 42.975 145.745 ;
        RECT 43.155 145.465 43.440 145.925 ;
        RECT 42.720 144.565 42.900 145.215 ;
        RECT 43.620 145.015 43.870 145.665 ;
        RECT 43.070 144.685 43.870 145.015 ;
        RECT 38.205 143.375 40.795 144.465 ;
        RECT 41.005 143.375 41.235 144.515 ;
        RECT 41.405 143.545 41.735 144.525 ;
        RECT 41.905 143.375 42.115 144.515 ;
        RECT 42.635 144.395 42.900 144.565 ;
        RECT 42.720 144.355 42.900 144.395 ;
        RECT 42.720 143.685 42.975 144.355 ;
        RECT 43.155 143.375 43.440 144.175 ;
        RECT 43.620 144.095 43.870 144.685 ;
        RECT 44.070 145.330 44.390 145.660 ;
        RECT 44.570 145.445 45.230 145.925 ;
        RECT 45.430 145.535 46.280 145.705 ;
        RECT 44.070 144.435 44.260 145.330 ;
        RECT 44.580 145.005 45.240 145.275 ;
        RECT 44.910 144.945 45.240 145.005 ;
        RECT 44.430 144.775 44.760 144.835 ;
        RECT 45.430 144.775 45.600 145.535 ;
        RECT 46.840 145.465 47.160 145.925 ;
        RECT 47.360 145.285 47.610 145.715 ;
        RECT 47.900 145.485 48.310 145.925 ;
        RECT 48.480 145.545 49.495 145.745 ;
        RECT 45.770 145.115 47.020 145.285 ;
        RECT 45.770 144.995 46.100 145.115 ;
        RECT 44.430 144.605 46.330 144.775 ;
        RECT 44.070 144.265 45.990 144.435 ;
        RECT 44.070 144.245 44.390 144.265 ;
        RECT 43.620 143.585 43.950 144.095 ;
        RECT 44.220 143.635 44.390 144.245 ;
        RECT 46.160 144.095 46.330 144.605 ;
        RECT 46.500 144.535 46.680 144.945 ;
        RECT 46.850 144.355 47.020 145.115 ;
        RECT 44.560 143.375 44.890 144.065 ;
        RECT 45.120 143.925 46.330 144.095 ;
        RECT 46.500 144.045 47.020 144.355 ;
        RECT 47.190 144.945 47.610 145.285 ;
        RECT 47.900 144.945 48.310 145.275 ;
        RECT 47.190 144.175 47.380 144.945 ;
        RECT 48.480 144.815 48.650 145.545 ;
        RECT 49.795 145.375 49.965 145.705 ;
        RECT 50.135 145.545 50.465 145.925 ;
        RECT 48.820 144.995 49.170 145.365 ;
        RECT 48.480 144.775 48.900 144.815 ;
        RECT 47.550 144.605 48.900 144.775 ;
        RECT 47.550 144.445 47.800 144.605 ;
        RECT 48.310 144.175 48.560 144.435 ;
        RECT 47.190 143.925 48.560 144.175 ;
        RECT 45.120 143.635 45.360 143.925 ;
        RECT 46.160 143.845 46.330 143.925 ;
        RECT 45.560 143.375 45.980 143.755 ;
        RECT 46.160 143.595 46.790 143.845 ;
        RECT 47.260 143.375 47.590 143.755 ;
        RECT 47.760 143.635 47.930 143.925 ;
        RECT 48.730 143.760 48.900 144.605 ;
        RECT 49.350 144.435 49.570 145.305 ;
        RECT 49.795 145.185 50.490 145.375 ;
        RECT 49.070 144.055 49.570 144.435 ;
        RECT 49.740 144.385 50.150 145.005 ;
        RECT 50.320 144.215 50.490 145.185 ;
        RECT 49.795 144.045 50.490 144.215 ;
        RECT 48.110 143.375 48.490 143.755 ;
        RECT 48.730 143.590 49.560 143.760 ;
        RECT 49.795 143.545 49.965 144.045 ;
        RECT 50.135 143.375 50.465 143.875 ;
        RECT 50.680 143.545 50.905 145.665 ;
        RECT 51.075 145.545 51.405 145.925 ;
        RECT 51.575 145.375 51.745 145.665 ;
        RECT 51.080 145.205 51.745 145.375 ;
        RECT 51.080 144.215 51.310 145.205 ;
        RECT 52.010 145.185 52.265 145.755 ;
        RECT 52.435 145.525 52.765 145.925 ;
        RECT 53.190 145.390 53.720 145.755 ;
        RECT 53.910 145.585 54.185 145.755 ;
        RECT 53.905 145.415 54.185 145.585 ;
        RECT 53.190 145.355 53.365 145.390 ;
        RECT 52.435 145.185 53.365 145.355 ;
        RECT 51.480 144.385 51.830 145.035 ;
        RECT 52.010 144.515 52.180 145.185 ;
        RECT 52.435 145.015 52.605 145.185 ;
        RECT 52.350 144.685 52.605 145.015 ;
        RECT 52.830 144.685 53.025 145.015 ;
        RECT 51.080 144.045 51.745 144.215 ;
        RECT 51.075 143.375 51.405 143.875 ;
        RECT 51.575 143.545 51.745 144.045 ;
        RECT 52.010 143.545 52.345 144.515 ;
        RECT 52.515 143.375 52.685 144.515 ;
        RECT 52.855 143.715 53.025 144.685 ;
        RECT 53.195 144.055 53.365 145.185 ;
        RECT 53.535 144.395 53.705 145.195 ;
        RECT 53.910 144.595 54.185 145.415 ;
        RECT 54.355 144.395 54.545 145.755 ;
        RECT 54.725 145.390 55.235 145.925 ;
        RECT 55.455 145.115 55.700 145.720 ;
        RECT 56.605 145.155 58.275 145.925 ;
        RECT 54.745 144.945 55.975 145.115 ;
        RECT 53.535 144.225 54.545 144.395 ;
        RECT 54.715 144.380 55.465 144.570 ;
        RECT 53.195 143.885 54.320 144.055 ;
        RECT 54.715 143.715 54.885 144.380 ;
        RECT 55.635 144.135 55.975 144.945 ;
        RECT 52.855 143.545 54.885 143.715 ;
        RECT 55.055 143.375 55.225 144.135 ;
        RECT 55.460 143.725 55.975 144.135 ;
        RECT 56.605 144.465 57.355 144.985 ;
        RECT 57.525 144.635 58.275 145.155 ;
        RECT 58.485 145.105 58.715 145.925 ;
        RECT 58.885 145.125 59.215 145.755 ;
        RECT 58.465 144.685 58.795 144.935 ;
        RECT 58.965 144.525 59.215 145.125 ;
        RECT 59.385 145.105 59.595 145.925 ;
        RECT 60.285 145.155 62.875 145.925 ;
        RECT 63.045 145.200 63.335 145.925 ;
        RECT 56.605 143.375 58.275 144.465 ;
        RECT 58.485 143.375 58.715 144.515 ;
        RECT 58.885 143.545 59.215 144.525 ;
        RECT 59.385 143.375 59.595 144.515 ;
        RECT 60.285 144.465 61.495 144.985 ;
        RECT 61.665 144.635 62.875 145.155 ;
        RECT 64.240 145.115 64.485 145.720 ;
        RECT 64.705 145.390 65.215 145.925 ;
        RECT 63.965 144.945 65.195 145.115 ;
        RECT 60.285 143.375 62.875 144.465 ;
        RECT 63.045 143.375 63.335 144.540 ;
        RECT 63.965 144.135 64.305 144.945 ;
        RECT 64.475 144.380 65.225 144.570 ;
        RECT 63.965 143.725 64.480 144.135 ;
        RECT 64.715 143.375 64.885 144.135 ;
        RECT 65.055 143.715 65.225 144.380 ;
        RECT 65.395 144.395 65.585 145.755 ;
        RECT 65.755 144.905 66.030 145.755 ;
        RECT 66.220 145.390 66.750 145.755 ;
        RECT 67.175 145.525 67.505 145.925 ;
        RECT 66.575 145.355 66.750 145.390 ;
        RECT 65.755 144.735 66.035 144.905 ;
        RECT 65.755 144.595 66.030 144.735 ;
        RECT 66.235 144.395 66.405 145.195 ;
        RECT 65.395 144.225 66.405 144.395 ;
        RECT 66.575 145.185 67.505 145.355 ;
        RECT 67.675 145.185 67.930 145.755 ;
        RECT 68.570 145.380 73.915 145.925 ;
        RECT 74.090 145.380 79.435 145.925 ;
        RECT 79.615 145.425 79.945 145.925 ;
        RECT 66.575 144.055 66.745 145.185 ;
        RECT 67.335 145.015 67.505 145.185 ;
        RECT 65.620 143.885 66.745 144.055 ;
        RECT 66.915 144.685 67.110 145.015 ;
        RECT 67.335 144.685 67.590 145.015 ;
        RECT 66.915 143.715 67.085 144.685 ;
        RECT 67.760 144.515 67.930 145.185 ;
        RECT 65.055 143.545 67.085 143.715 ;
        RECT 67.255 143.375 67.425 144.515 ;
        RECT 67.595 143.545 67.930 144.515 ;
        RECT 70.160 143.810 70.510 145.060 ;
        RECT 71.990 144.550 72.330 145.380 ;
        RECT 75.680 143.810 76.030 145.060 ;
        RECT 77.510 144.550 77.850 145.380 ;
        RECT 80.145 145.355 80.315 145.705 ;
        RECT 80.515 145.525 80.845 145.925 ;
        RECT 81.015 145.355 81.185 145.705 ;
        RECT 81.355 145.525 81.735 145.925 ;
        RECT 79.610 144.685 79.960 145.255 ;
        RECT 80.145 145.185 81.755 145.355 ;
        RECT 81.925 145.250 82.195 145.595 ;
        RECT 81.585 145.015 81.755 145.185 ;
        RECT 79.610 144.225 79.930 144.515 ;
        RECT 80.130 144.395 80.840 145.015 ;
        RECT 81.010 144.685 81.415 145.015 ;
        RECT 81.585 144.685 81.855 145.015 ;
        RECT 81.585 144.515 81.755 144.685 ;
        RECT 82.025 144.515 82.195 145.250 ;
        RECT 82.825 145.155 84.495 145.925 ;
        RECT 81.030 144.345 81.755 144.515 ;
        RECT 81.030 144.225 81.200 144.345 ;
        RECT 79.610 144.055 81.200 144.225 ;
        RECT 68.570 143.375 73.915 143.810 ;
        RECT 74.090 143.375 79.435 143.810 ;
        RECT 79.610 143.595 81.265 143.885 ;
        RECT 81.435 143.375 81.715 144.175 ;
        RECT 81.925 143.545 82.195 144.515 ;
        RECT 82.825 144.465 83.575 144.985 ;
        RECT 83.745 144.635 84.495 145.155 ;
        RECT 84.940 145.115 85.185 145.720 ;
        RECT 85.405 145.390 85.915 145.925 ;
        RECT 84.665 144.945 85.895 145.115 ;
        RECT 82.825 143.375 84.495 144.465 ;
        RECT 84.665 144.135 85.005 144.945 ;
        RECT 85.175 144.380 85.925 144.570 ;
        RECT 84.665 143.725 85.180 144.135 ;
        RECT 85.415 143.375 85.585 144.135 ;
        RECT 85.755 143.715 85.925 144.380 ;
        RECT 86.095 144.395 86.285 145.755 ;
        RECT 86.455 144.905 86.730 145.755 ;
        RECT 86.920 145.390 87.450 145.755 ;
        RECT 87.875 145.525 88.205 145.925 ;
        RECT 87.275 145.355 87.450 145.390 ;
        RECT 86.455 144.735 86.735 144.905 ;
        RECT 86.455 144.595 86.730 144.735 ;
        RECT 86.935 144.395 87.105 145.195 ;
        RECT 86.095 144.225 87.105 144.395 ;
        RECT 87.275 145.185 88.205 145.355 ;
        RECT 88.375 145.185 88.630 145.755 ;
        RECT 88.805 145.200 89.095 145.925 ;
        RECT 90.275 145.375 90.445 145.755 ;
        RECT 90.625 145.545 90.955 145.925 ;
        RECT 90.275 145.205 90.940 145.375 ;
        RECT 91.135 145.250 91.395 145.755 ;
        RECT 87.275 144.055 87.445 145.185 ;
        RECT 88.035 145.015 88.205 145.185 ;
        RECT 86.320 143.885 87.445 144.055 ;
        RECT 87.615 144.685 87.810 145.015 ;
        RECT 88.035 144.685 88.290 145.015 ;
        RECT 87.615 143.715 87.785 144.685 ;
        RECT 88.460 144.515 88.630 145.185 ;
        RECT 90.205 144.655 90.535 145.025 ;
        RECT 90.770 144.950 90.940 145.205 ;
        RECT 90.770 144.620 91.055 144.950 ;
        RECT 85.755 143.545 87.785 143.715 ;
        RECT 87.955 143.375 88.125 144.515 ;
        RECT 88.295 143.545 88.630 144.515 ;
        RECT 88.805 143.375 89.095 144.540 ;
        RECT 90.770 144.475 90.940 144.620 ;
        RECT 90.275 144.305 90.940 144.475 ;
        RECT 91.225 144.450 91.395 145.250 ;
        RECT 92.025 145.155 93.695 145.925 ;
        RECT 90.275 143.545 90.445 144.305 ;
        RECT 90.625 143.375 90.955 144.135 ;
        RECT 91.125 143.545 91.395 144.450 ;
        RECT 92.025 144.465 92.775 144.985 ;
        RECT 92.945 144.635 93.695 145.155 ;
        RECT 93.980 145.295 94.265 145.755 ;
        RECT 94.435 145.465 94.705 145.925 ;
        RECT 93.980 145.125 94.935 145.295 ;
        RECT 92.025 143.375 93.695 144.465 ;
        RECT 93.865 144.395 94.555 144.955 ;
        RECT 94.725 144.225 94.935 145.125 ;
        RECT 93.980 144.005 94.935 144.225 ;
        RECT 95.105 144.955 95.505 145.755 ;
        RECT 95.695 145.295 95.975 145.755 ;
        RECT 96.495 145.465 96.820 145.925 ;
        RECT 95.695 145.125 96.820 145.295 ;
        RECT 96.990 145.185 97.375 145.755 ;
        RECT 96.370 145.015 96.820 145.125 ;
        RECT 95.105 144.395 96.200 144.955 ;
        RECT 96.370 144.685 96.925 145.015 ;
        RECT 93.980 143.545 94.265 144.005 ;
        RECT 94.435 143.375 94.705 143.835 ;
        RECT 95.105 143.545 95.505 144.395 ;
        RECT 96.370 144.225 96.820 144.685 ;
        RECT 97.095 144.515 97.375 145.185 ;
        RECT 98.005 145.155 101.515 145.925 ;
        RECT 101.690 145.380 107.035 145.925 ;
        RECT 107.215 145.425 107.545 145.925 ;
        RECT 95.695 144.005 96.820 144.225 ;
        RECT 95.695 143.545 95.975 144.005 ;
        RECT 96.495 143.375 96.820 143.835 ;
        RECT 96.990 143.545 97.375 144.515 ;
        RECT 98.005 144.465 99.695 144.985 ;
        RECT 99.865 144.635 101.515 145.155 ;
        RECT 98.005 143.375 101.515 144.465 ;
        RECT 103.280 143.810 103.630 145.060 ;
        RECT 105.110 144.550 105.450 145.380 ;
        RECT 107.745 145.355 107.915 145.705 ;
        RECT 108.115 145.525 108.445 145.925 ;
        RECT 108.615 145.355 108.785 145.705 ;
        RECT 108.955 145.525 109.335 145.925 ;
        RECT 107.210 144.685 107.560 145.255 ;
        RECT 107.745 145.185 109.355 145.355 ;
        RECT 109.525 145.250 109.795 145.595 ;
        RECT 109.185 145.015 109.355 145.185 ;
        RECT 107.210 144.225 107.530 144.515 ;
        RECT 107.730 144.395 108.440 145.015 ;
        RECT 108.610 144.685 109.015 145.015 ;
        RECT 109.185 144.685 109.455 145.015 ;
        RECT 109.185 144.515 109.355 144.685 ;
        RECT 109.625 144.515 109.795 145.250 ;
        RECT 108.630 144.345 109.355 144.515 ;
        RECT 108.630 144.225 108.800 144.345 ;
        RECT 107.210 144.055 108.800 144.225 ;
        RECT 101.690 143.375 107.035 143.810 ;
        RECT 107.210 143.595 108.865 143.885 ;
        RECT 109.035 143.375 109.315 144.175 ;
        RECT 109.525 143.545 109.795 144.515 ;
        RECT 109.965 145.125 110.305 145.755 ;
        RECT 110.475 145.125 110.725 145.925 ;
        RECT 110.915 145.275 111.245 145.755 ;
        RECT 111.415 145.465 111.640 145.925 ;
        RECT 111.810 145.275 112.140 145.755 ;
        RECT 109.965 145.075 110.195 145.125 ;
        RECT 110.915 145.105 112.140 145.275 ;
        RECT 112.770 145.145 113.270 145.755 ;
        RECT 114.565 145.200 114.855 145.925 ;
        RECT 109.965 144.515 110.140 145.075 ;
        RECT 110.310 144.765 111.005 144.935 ;
        RECT 110.835 144.515 111.005 144.765 ;
        RECT 111.180 144.735 111.600 144.935 ;
        RECT 111.770 144.735 112.100 144.935 ;
        RECT 112.270 144.735 112.600 144.935 ;
        RECT 112.770 144.515 112.940 145.145 ;
        RECT 115.760 145.115 116.005 145.720 ;
        RECT 116.225 145.390 116.735 145.925 ;
        RECT 115.485 144.945 116.715 145.115 ;
        RECT 113.125 144.685 113.475 144.935 ;
        RECT 109.965 143.545 110.305 144.515 ;
        RECT 110.475 143.375 110.645 144.515 ;
        RECT 110.835 144.345 113.270 144.515 ;
        RECT 110.915 143.375 111.165 144.175 ;
        RECT 111.810 143.545 112.140 144.345 ;
        RECT 112.440 143.375 112.770 144.175 ;
        RECT 112.940 143.545 113.270 144.345 ;
        RECT 114.565 143.375 114.855 144.540 ;
        RECT 115.485 144.135 115.825 144.945 ;
        RECT 115.995 144.380 116.745 144.570 ;
        RECT 115.485 143.725 116.000 144.135 ;
        RECT 116.235 143.375 116.405 144.135 ;
        RECT 116.575 143.715 116.745 144.380 ;
        RECT 116.915 144.395 117.105 145.755 ;
        RECT 117.275 145.585 117.550 145.755 ;
        RECT 117.275 145.415 117.555 145.585 ;
        RECT 117.275 144.595 117.550 145.415 ;
        RECT 117.740 145.390 118.270 145.755 ;
        RECT 118.695 145.525 119.025 145.925 ;
        RECT 118.095 145.355 118.270 145.390 ;
        RECT 117.755 144.395 117.925 145.195 ;
        RECT 116.915 144.225 117.925 144.395 ;
        RECT 118.095 145.185 119.025 145.355 ;
        RECT 119.195 145.185 119.450 145.755 ;
        RECT 118.095 144.055 118.265 145.185 ;
        RECT 118.855 145.015 119.025 145.185 ;
        RECT 117.140 143.885 118.265 144.055 ;
        RECT 118.435 144.685 118.630 145.015 ;
        RECT 118.855 144.685 119.110 145.015 ;
        RECT 118.435 143.715 118.605 144.685 ;
        RECT 119.280 144.515 119.450 145.185 ;
        RECT 119.665 145.105 119.895 145.925 ;
        RECT 120.065 145.125 120.395 145.755 ;
        RECT 119.645 144.685 119.975 144.935 ;
        RECT 120.145 144.525 120.395 145.125 ;
        RECT 120.565 145.105 120.775 145.925 ;
        RECT 121.555 145.375 121.725 145.755 ;
        RECT 121.905 145.545 122.235 145.925 ;
        RECT 121.555 145.205 122.220 145.375 ;
        RECT 122.415 145.250 122.675 145.755 ;
        RECT 121.485 144.655 121.815 145.025 ;
        RECT 122.050 144.950 122.220 145.205 ;
        RECT 116.575 143.545 118.605 143.715 ;
        RECT 118.775 143.375 118.945 144.515 ;
        RECT 119.115 143.545 119.450 144.515 ;
        RECT 119.665 143.375 119.895 144.515 ;
        RECT 120.065 143.545 120.395 144.525 ;
        RECT 122.050 144.620 122.335 144.950 ;
        RECT 120.565 143.375 120.775 144.515 ;
        RECT 122.050 144.475 122.220 144.620 ;
        RECT 121.555 144.305 122.220 144.475 ;
        RECT 122.505 144.450 122.675 145.250 ;
        RECT 122.845 145.155 126.355 145.925 ;
        RECT 126.525 145.175 127.735 145.925 ;
        RECT 121.555 143.545 121.725 144.305 ;
        RECT 121.905 143.375 122.235 144.135 ;
        RECT 122.405 143.545 122.675 144.450 ;
        RECT 122.845 144.465 124.535 144.985 ;
        RECT 124.705 144.635 126.355 145.155 ;
        RECT 126.525 144.465 127.045 145.005 ;
        RECT 127.215 144.635 127.735 145.175 ;
        RECT 122.845 143.375 126.355 144.465 ;
        RECT 126.525 143.375 127.735 144.465 ;
        RECT 14.660 143.205 127.820 143.375 ;
        RECT 14.745 142.115 15.955 143.205 ;
        RECT 14.745 141.405 15.265 141.945 ;
        RECT 15.435 141.575 15.955 142.115 ;
        RECT 16.125 142.115 18.715 143.205 ;
        RECT 18.890 142.770 24.235 143.205 ;
        RECT 16.125 141.595 17.335 142.115 ;
        RECT 17.505 141.425 18.715 141.945 ;
        RECT 20.480 141.520 20.830 142.770 ;
        RECT 24.405 142.040 24.695 143.205 ;
        RECT 25.325 142.115 28.835 143.205 ;
        RECT 29.010 142.770 34.355 143.205 ;
        RECT 14.745 140.655 15.955 141.405 ;
        RECT 16.125 140.655 18.715 141.425 ;
        RECT 22.310 141.200 22.650 142.030 ;
        RECT 25.325 141.595 27.015 142.115 ;
        RECT 27.185 141.425 28.835 141.945 ;
        RECT 30.600 141.520 30.950 142.770 ;
        RECT 34.525 142.065 34.795 143.035 ;
        RECT 35.005 142.405 35.285 143.205 ;
        RECT 35.455 142.695 37.110 142.985 ;
        RECT 35.520 142.355 37.110 142.525 ;
        RECT 35.520 142.235 35.690 142.355 ;
        RECT 34.965 142.065 35.690 142.235 ;
        RECT 18.890 140.655 24.235 141.200 ;
        RECT 24.405 140.655 24.695 141.380 ;
        RECT 25.325 140.655 28.835 141.425 ;
        RECT 32.430 141.200 32.770 142.030 ;
        RECT 34.525 141.330 34.695 142.065 ;
        RECT 34.965 141.895 35.135 142.065 ;
        RECT 34.865 141.565 35.135 141.895 ;
        RECT 35.305 141.565 35.710 141.895 ;
        RECT 35.880 141.565 36.590 142.185 ;
        RECT 36.790 142.065 37.110 142.355 ;
        RECT 38.205 142.115 41.715 143.205 ;
        RECT 41.890 142.770 47.235 143.205 ;
        RECT 34.965 141.395 35.135 141.565 ;
        RECT 29.010 140.655 34.355 141.200 ;
        RECT 34.525 140.985 34.795 141.330 ;
        RECT 34.965 141.225 36.575 141.395 ;
        RECT 36.760 141.325 37.110 141.895 ;
        RECT 38.205 141.595 39.895 142.115 ;
        RECT 40.065 141.425 41.715 141.945 ;
        RECT 43.480 141.520 43.830 142.770 ;
        RECT 47.405 142.065 47.675 143.035 ;
        RECT 47.885 142.405 48.165 143.205 ;
        RECT 48.335 142.695 49.990 142.985 ;
        RECT 48.400 142.355 49.990 142.525 ;
        RECT 48.400 142.235 48.570 142.355 ;
        RECT 47.845 142.065 48.570 142.235 ;
        RECT 34.985 140.655 35.365 141.055 ;
        RECT 35.535 140.875 35.705 141.225 ;
        RECT 35.875 140.655 36.205 141.055 ;
        RECT 36.405 140.875 36.575 141.225 ;
        RECT 36.775 140.655 37.105 141.155 ;
        RECT 38.205 140.655 41.715 141.425 ;
        RECT 45.310 141.200 45.650 142.030 ;
        RECT 47.405 141.330 47.575 142.065 ;
        RECT 47.845 141.895 48.015 142.065 ;
        RECT 47.745 141.565 48.015 141.895 ;
        RECT 48.185 141.565 48.590 141.895 ;
        RECT 48.760 141.565 49.470 142.185 ;
        RECT 49.670 142.065 49.990 142.355 ;
        RECT 50.165 142.040 50.455 143.205 ;
        RECT 50.625 142.115 52.295 143.205 ;
        RECT 47.845 141.395 48.015 141.565 ;
        RECT 41.890 140.655 47.235 141.200 ;
        RECT 47.405 140.985 47.675 141.330 ;
        RECT 47.845 141.225 49.455 141.395 ;
        RECT 49.640 141.325 49.990 141.895 ;
        RECT 50.625 141.595 51.375 142.115 ;
        RECT 52.465 142.065 52.805 143.035 ;
        RECT 52.975 142.065 53.145 143.205 ;
        RECT 53.415 142.405 53.665 143.205 ;
        RECT 54.310 142.235 54.640 143.035 ;
        RECT 54.940 142.405 55.270 143.205 ;
        RECT 55.440 142.235 55.770 143.035 ;
        RECT 56.260 142.575 56.545 143.035 ;
        RECT 56.715 142.745 56.985 143.205 ;
        RECT 56.260 142.355 57.215 142.575 ;
        RECT 53.335 142.065 55.770 142.235 ;
        RECT 51.545 141.425 52.295 141.945 ;
        RECT 47.865 140.655 48.245 141.055 ;
        RECT 48.415 140.875 48.585 141.225 ;
        RECT 48.755 140.655 49.085 141.055 ;
        RECT 49.285 140.875 49.455 141.225 ;
        RECT 49.655 140.655 49.985 141.155 ;
        RECT 50.165 140.655 50.455 141.380 ;
        RECT 50.625 140.655 52.295 141.425 ;
        RECT 52.465 141.505 52.640 142.065 ;
        RECT 53.335 141.815 53.505 142.065 ;
        RECT 52.810 141.645 53.505 141.815 ;
        RECT 53.680 141.645 54.100 141.845 ;
        RECT 54.270 141.645 54.600 141.845 ;
        RECT 54.770 141.645 55.100 141.845 ;
        RECT 52.465 141.455 52.695 141.505 ;
        RECT 52.465 140.825 52.805 141.455 ;
        RECT 52.975 140.655 53.225 141.455 ;
        RECT 53.415 141.305 54.640 141.475 ;
        RECT 53.415 140.825 53.745 141.305 ;
        RECT 53.915 140.655 54.140 141.115 ;
        RECT 54.310 140.825 54.640 141.305 ;
        RECT 55.270 141.435 55.440 142.065 ;
        RECT 55.625 141.645 55.975 141.895 ;
        RECT 56.145 141.625 56.835 142.185 ;
        RECT 57.005 141.455 57.215 142.355 ;
        RECT 55.270 140.825 55.770 141.435 ;
        RECT 56.260 141.285 57.215 141.455 ;
        RECT 57.385 142.185 57.785 143.035 ;
        RECT 57.975 142.575 58.255 143.035 ;
        RECT 58.775 142.745 59.100 143.205 ;
        RECT 57.975 142.355 59.100 142.575 ;
        RECT 57.385 141.625 58.480 142.185 ;
        RECT 58.650 141.895 59.100 142.355 ;
        RECT 59.270 142.065 59.655 143.035 ;
        RECT 56.260 140.825 56.545 141.285 ;
        RECT 56.715 140.655 56.985 141.115 ;
        RECT 57.385 140.825 57.785 141.625 ;
        RECT 58.650 141.565 59.205 141.895 ;
        RECT 58.650 141.455 59.100 141.565 ;
        RECT 57.975 141.285 59.100 141.455 ;
        RECT 59.375 141.395 59.655 142.065 ;
        RECT 57.975 140.825 58.255 141.285 ;
        RECT 58.775 140.655 59.100 141.115 ;
        RECT 59.270 140.825 59.655 141.395 ;
        RECT 59.830 142.015 60.085 142.895 ;
        RECT 60.255 142.065 60.560 143.205 ;
        RECT 60.900 142.825 61.230 143.205 ;
        RECT 61.410 142.655 61.580 142.945 ;
        RECT 61.750 142.745 62.000 143.205 ;
        RECT 60.780 142.485 61.580 142.655 ;
        RECT 62.170 142.695 63.040 143.035 ;
        RECT 59.830 141.365 60.040 142.015 ;
        RECT 60.780 141.895 60.950 142.485 ;
        RECT 62.170 142.315 62.340 142.695 ;
        RECT 63.275 142.575 63.445 143.035 ;
        RECT 63.615 142.745 63.985 143.205 ;
        RECT 64.280 142.605 64.450 142.945 ;
        RECT 64.620 142.775 64.950 143.205 ;
        RECT 65.185 142.605 65.355 142.945 ;
        RECT 61.120 142.145 62.340 142.315 ;
        RECT 62.510 142.235 62.970 142.525 ;
        RECT 63.275 142.405 63.835 142.575 ;
        RECT 64.280 142.435 65.355 142.605 ;
        RECT 65.525 142.705 66.205 143.035 ;
        RECT 66.420 142.705 66.670 143.035 ;
        RECT 66.840 142.745 67.090 143.205 ;
        RECT 63.665 142.265 63.835 142.405 ;
        RECT 62.510 142.225 63.475 142.235 ;
        RECT 62.170 142.055 62.340 142.145 ;
        RECT 62.800 142.065 63.475 142.225 ;
        RECT 60.210 141.865 60.950 141.895 ;
        RECT 60.210 141.565 61.125 141.865 ;
        RECT 60.800 141.390 61.125 141.565 ;
        RECT 59.830 140.835 60.085 141.365 ;
        RECT 60.255 140.655 60.560 141.115 ;
        RECT 60.805 141.035 61.125 141.390 ;
        RECT 61.295 141.605 61.835 141.975 ;
        RECT 62.170 141.885 62.575 142.055 ;
        RECT 61.295 141.205 61.535 141.605 ;
        RECT 62.015 141.435 62.235 141.715 ;
        RECT 61.705 141.265 62.235 141.435 ;
        RECT 61.705 141.035 61.875 141.265 ;
        RECT 62.405 141.105 62.575 141.885 ;
        RECT 62.745 141.275 63.095 141.895 ;
        RECT 63.265 141.275 63.475 142.065 ;
        RECT 63.665 142.095 65.165 142.265 ;
        RECT 63.665 141.405 63.835 142.095 ;
        RECT 65.525 141.925 65.695 142.705 ;
        RECT 66.500 142.575 66.670 142.705 ;
        RECT 64.005 141.755 65.695 141.925 ;
        RECT 65.865 142.145 66.330 142.535 ;
        RECT 66.500 142.405 66.895 142.575 ;
        RECT 64.005 141.575 64.175 141.755 ;
        RECT 60.805 140.865 61.875 141.035 ;
        RECT 62.045 140.655 62.235 141.095 ;
        RECT 62.405 140.825 63.355 141.105 ;
        RECT 63.665 141.015 63.925 141.405 ;
        RECT 64.345 141.335 65.135 141.585 ;
        RECT 63.575 140.845 63.925 141.015 ;
        RECT 64.135 140.655 64.465 141.115 ;
        RECT 65.340 141.045 65.510 141.755 ;
        RECT 65.865 141.555 66.035 142.145 ;
        RECT 65.680 141.335 66.035 141.555 ;
        RECT 66.205 141.335 66.555 141.955 ;
        RECT 66.725 141.045 66.895 142.405 ;
        RECT 67.260 142.235 67.585 143.020 ;
        RECT 67.065 141.185 67.525 142.235 ;
        RECT 65.340 140.875 66.195 141.045 ;
        RECT 66.400 140.875 66.895 141.045 ;
        RECT 67.065 140.655 67.395 141.015 ;
        RECT 67.755 140.915 67.925 143.035 ;
        RECT 68.095 142.705 68.425 143.205 ;
        RECT 68.595 142.535 68.850 143.035 ;
        RECT 68.100 142.365 68.850 142.535 ;
        RECT 68.100 141.375 68.330 142.365 ;
        RECT 68.500 141.545 68.850 142.195 ;
        RECT 69.025 142.130 69.295 143.035 ;
        RECT 69.465 142.445 69.795 143.205 ;
        RECT 69.975 142.275 70.145 143.035 ;
        RECT 68.100 141.205 68.850 141.375 ;
        RECT 68.095 140.655 68.425 141.035 ;
        RECT 68.595 140.915 68.850 141.205 ;
        RECT 69.025 141.330 69.195 142.130 ;
        RECT 69.480 142.105 70.145 142.275 ;
        RECT 70.405 142.115 71.615 143.205 ;
        RECT 69.480 141.960 69.650 142.105 ;
        RECT 69.365 141.630 69.650 141.960 ;
        RECT 69.480 141.375 69.650 141.630 ;
        RECT 69.885 141.555 70.215 141.925 ;
        RECT 70.405 141.575 70.925 142.115 ;
        RECT 71.845 142.065 72.055 143.205 ;
        RECT 72.225 142.055 72.555 143.035 ;
        RECT 72.725 142.065 72.955 143.205 ;
        RECT 73.165 142.115 75.755 143.205 ;
        RECT 71.095 141.405 71.615 141.945 ;
        RECT 69.025 140.825 69.285 141.330 ;
        RECT 69.480 141.205 70.145 141.375 ;
        RECT 69.465 140.655 69.795 141.035 ;
        RECT 69.975 140.825 70.145 141.205 ;
        RECT 70.405 140.655 71.615 141.405 ;
        RECT 71.845 140.655 72.055 141.475 ;
        RECT 72.225 141.455 72.475 142.055 ;
        RECT 72.645 141.645 72.975 141.895 ;
        RECT 73.165 141.595 74.375 142.115 ;
        RECT 75.925 142.040 76.215 143.205 ;
        RECT 76.845 142.115 79.435 143.205 ;
        RECT 79.610 142.770 84.955 143.205 ;
        RECT 85.130 142.770 90.475 143.205 ;
        RECT 90.650 142.770 95.995 143.205 ;
        RECT 96.170 142.770 101.515 143.205 ;
        RECT 72.225 140.825 72.555 141.455 ;
        RECT 72.725 140.655 72.955 141.475 ;
        RECT 74.545 141.425 75.755 141.945 ;
        RECT 76.845 141.595 78.055 142.115 ;
        RECT 78.225 141.425 79.435 141.945 ;
        RECT 81.200 141.520 81.550 142.770 ;
        RECT 73.165 140.655 75.755 141.425 ;
        RECT 75.925 140.655 76.215 141.380 ;
        RECT 76.845 140.655 79.435 141.425 ;
        RECT 83.030 141.200 83.370 142.030 ;
        RECT 86.720 141.520 87.070 142.770 ;
        RECT 88.550 141.200 88.890 142.030 ;
        RECT 92.240 141.520 92.590 142.770 ;
        RECT 94.070 141.200 94.410 142.030 ;
        RECT 97.760 141.520 98.110 142.770 ;
        RECT 101.685 142.040 101.975 143.205 ;
        RECT 102.145 142.115 104.735 143.205 ;
        RECT 104.910 142.770 110.255 143.205 ;
        RECT 110.430 142.770 115.775 143.205 ;
        RECT 99.590 141.200 99.930 142.030 ;
        RECT 102.145 141.595 103.355 142.115 ;
        RECT 103.525 141.425 104.735 141.945 ;
        RECT 106.500 141.520 106.850 142.770 ;
        RECT 79.610 140.655 84.955 141.200 ;
        RECT 85.130 140.655 90.475 141.200 ;
        RECT 90.650 140.655 95.995 141.200 ;
        RECT 96.170 140.655 101.515 141.200 ;
        RECT 101.685 140.655 101.975 141.380 ;
        RECT 102.145 140.655 104.735 141.425 ;
        RECT 108.330 141.200 108.670 142.030 ;
        RECT 112.020 141.520 112.370 142.770 ;
        RECT 115.945 142.445 116.460 142.855 ;
        RECT 116.695 142.445 116.865 143.205 ;
        RECT 117.035 142.865 119.065 143.035 ;
        RECT 113.850 141.200 114.190 142.030 ;
        RECT 115.945 141.635 116.285 142.445 ;
        RECT 117.035 142.200 117.205 142.865 ;
        RECT 117.600 142.525 118.725 142.695 ;
        RECT 116.455 142.010 117.205 142.200 ;
        RECT 117.375 142.185 118.385 142.355 ;
        RECT 115.945 141.465 117.175 141.635 ;
        RECT 104.910 140.655 110.255 141.200 ;
        RECT 110.430 140.655 115.775 141.200 ;
        RECT 116.220 140.860 116.465 141.465 ;
        RECT 116.685 140.655 117.195 141.190 ;
        RECT 117.375 140.825 117.565 142.185 ;
        RECT 117.735 141.845 118.010 141.985 ;
        RECT 117.735 141.675 118.015 141.845 ;
        RECT 117.735 140.825 118.010 141.675 ;
        RECT 118.215 141.385 118.385 142.185 ;
        RECT 118.555 141.395 118.725 142.525 ;
        RECT 118.895 141.895 119.065 142.865 ;
        RECT 119.235 142.065 119.405 143.205 ;
        RECT 119.575 142.065 119.910 143.035 ;
        RECT 120.125 142.065 120.355 143.205 ;
        RECT 118.895 141.565 119.090 141.895 ;
        RECT 119.315 141.565 119.570 141.895 ;
        RECT 119.315 141.395 119.485 141.565 ;
        RECT 119.740 141.395 119.910 142.065 ;
        RECT 120.525 142.055 120.855 143.035 ;
        RECT 121.025 142.065 121.235 143.205 ;
        RECT 121.465 142.115 122.675 143.205 ;
        RECT 122.845 142.115 126.355 143.205 ;
        RECT 126.525 142.115 127.735 143.205 ;
        RECT 120.105 141.645 120.435 141.895 ;
        RECT 118.555 141.225 119.485 141.395 ;
        RECT 118.555 141.190 118.730 141.225 ;
        RECT 118.200 140.825 118.730 141.190 ;
        RECT 119.155 140.655 119.485 141.055 ;
        RECT 119.655 140.825 119.910 141.395 ;
        RECT 120.125 140.655 120.355 141.475 ;
        RECT 120.605 141.455 120.855 142.055 ;
        RECT 121.465 141.575 121.985 142.115 ;
        RECT 120.525 140.825 120.855 141.455 ;
        RECT 121.025 140.655 121.235 141.475 ;
        RECT 122.155 141.405 122.675 141.945 ;
        RECT 122.845 141.595 124.535 142.115 ;
        RECT 124.705 141.425 126.355 141.945 ;
        RECT 126.525 141.575 127.045 142.115 ;
        RECT 121.465 140.655 122.675 141.405 ;
        RECT 122.845 140.655 126.355 141.425 ;
        RECT 127.215 141.405 127.735 141.945 ;
        RECT 126.525 140.655 127.735 141.405 ;
        RECT 14.660 140.485 127.820 140.655 ;
        RECT 14.745 139.735 15.955 140.485 ;
        RECT 16.500 139.775 16.755 140.305 ;
        RECT 16.935 140.025 17.220 140.485 ;
        RECT 14.745 139.195 15.265 139.735 ;
        RECT 15.435 139.025 15.955 139.565 ;
        RECT 14.745 137.935 15.955 139.025 ;
        RECT 16.500 138.915 16.680 139.775 ;
        RECT 17.400 139.575 17.650 140.225 ;
        RECT 16.850 139.245 17.650 139.575 ;
        RECT 16.500 138.445 16.755 138.915 ;
        RECT 16.415 138.275 16.755 138.445 ;
        RECT 16.500 138.245 16.755 138.275 ;
        RECT 16.935 137.935 17.220 138.735 ;
        RECT 17.400 138.655 17.650 139.245 ;
        RECT 17.850 139.890 18.170 140.220 ;
        RECT 18.350 140.005 19.010 140.485 ;
        RECT 19.210 140.095 20.060 140.265 ;
        RECT 17.850 138.995 18.040 139.890 ;
        RECT 18.360 139.565 19.020 139.835 ;
        RECT 18.690 139.505 19.020 139.565 ;
        RECT 18.210 139.335 18.540 139.395 ;
        RECT 19.210 139.335 19.380 140.095 ;
        RECT 20.620 140.025 20.940 140.485 ;
        RECT 21.140 139.845 21.390 140.275 ;
        RECT 21.680 140.045 22.090 140.485 ;
        RECT 22.260 140.105 23.275 140.305 ;
        RECT 19.550 139.675 20.800 139.845 ;
        RECT 19.550 139.555 19.880 139.675 ;
        RECT 18.210 139.165 20.110 139.335 ;
        RECT 17.850 138.825 19.770 138.995 ;
        RECT 17.850 138.805 18.170 138.825 ;
        RECT 17.400 138.145 17.730 138.655 ;
        RECT 18.000 138.195 18.170 138.805 ;
        RECT 19.940 138.655 20.110 139.165 ;
        RECT 20.280 139.095 20.460 139.505 ;
        RECT 20.630 138.915 20.800 139.675 ;
        RECT 18.340 137.935 18.670 138.625 ;
        RECT 18.900 138.485 20.110 138.655 ;
        RECT 20.280 138.605 20.800 138.915 ;
        RECT 20.970 139.505 21.390 139.845 ;
        RECT 21.680 139.505 22.090 139.835 ;
        RECT 20.970 138.735 21.160 139.505 ;
        RECT 22.260 139.375 22.430 140.105 ;
        RECT 23.575 139.935 23.745 140.265 ;
        RECT 23.915 140.105 24.245 140.485 ;
        RECT 22.600 139.555 22.950 139.925 ;
        RECT 22.260 139.335 22.680 139.375 ;
        RECT 21.330 139.165 22.680 139.335 ;
        RECT 21.330 139.005 21.580 139.165 ;
        RECT 22.090 138.735 22.340 138.995 ;
        RECT 20.970 138.485 22.340 138.735 ;
        RECT 18.900 138.195 19.140 138.485 ;
        RECT 19.940 138.405 20.110 138.485 ;
        RECT 19.340 137.935 19.760 138.315 ;
        RECT 19.940 138.155 20.570 138.405 ;
        RECT 21.040 137.935 21.370 138.315 ;
        RECT 21.540 138.195 21.710 138.485 ;
        RECT 22.510 138.320 22.680 139.165 ;
        RECT 23.130 138.995 23.350 139.865 ;
        RECT 23.575 139.745 24.270 139.935 ;
        RECT 22.850 138.615 23.350 138.995 ;
        RECT 23.520 138.945 23.930 139.565 ;
        RECT 24.100 138.775 24.270 139.745 ;
        RECT 23.575 138.605 24.270 138.775 ;
        RECT 21.890 137.935 22.270 138.315 ;
        RECT 22.510 138.150 23.340 138.320 ;
        RECT 23.575 138.105 23.745 138.605 ;
        RECT 23.915 137.935 24.245 138.435 ;
        RECT 24.460 138.105 24.685 140.225 ;
        RECT 24.855 140.105 25.185 140.485 ;
        RECT 25.355 139.935 25.525 140.225 ;
        RECT 24.860 139.765 25.525 139.935 ;
        RECT 24.860 138.775 25.090 139.765 ;
        RECT 25.785 139.715 28.375 140.485 ;
        RECT 28.550 139.940 33.895 140.485 ;
        RECT 25.260 138.945 25.610 139.595 ;
        RECT 25.785 139.025 26.995 139.545 ;
        RECT 27.165 139.195 28.375 139.715 ;
        RECT 24.860 138.605 25.525 138.775 ;
        RECT 24.855 137.935 25.185 138.435 ;
        RECT 25.355 138.105 25.525 138.605 ;
        RECT 25.785 137.935 28.375 139.025 ;
        RECT 30.140 138.370 30.490 139.620 ;
        RECT 31.970 139.110 32.310 139.940 ;
        RECT 34.265 139.855 34.595 140.215 ;
        RECT 35.215 140.025 35.465 140.485 ;
        RECT 35.635 140.025 36.195 140.315 ;
        RECT 34.265 139.665 35.655 139.855 ;
        RECT 35.485 139.575 35.655 139.665 ;
        RECT 34.080 139.245 34.755 139.495 ;
        RECT 34.975 139.245 35.315 139.495 ;
        RECT 35.485 139.245 35.775 139.575 ;
        RECT 34.080 138.885 34.345 139.245 ;
        RECT 35.485 138.995 35.655 139.245 ;
        RECT 34.715 138.825 35.655 138.995 ;
        RECT 28.550 137.935 33.895 138.370 ;
        RECT 34.265 137.935 34.545 138.605 ;
        RECT 34.715 138.275 35.015 138.825 ;
        RECT 35.945 138.655 36.195 140.025 ;
        RECT 37.285 139.760 37.575 140.485 ;
        RECT 38.665 139.810 38.935 140.155 ;
        RECT 39.125 140.085 39.505 140.485 ;
        RECT 39.675 139.915 39.845 140.265 ;
        RECT 40.015 140.085 40.345 140.485 ;
        RECT 40.545 139.915 40.715 140.265 ;
        RECT 40.915 139.985 41.245 140.485 ;
        RECT 35.215 137.935 35.545 138.655 ;
        RECT 35.735 138.105 36.195 138.655 ;
        RECT 37.285 137.935 37.575 139.100 ;
        RECT 38.665 139.075 38.835 139.810 ;
        RECT 39.105 139.745 40.715 139.915 ;
        RECT 39.105 139.575 39.275 139.745 ;
        RECT 39.005 139.245 39.275 139.575 ;
        RECT 39.445 139.245 39.850 139.575 ;
        RECT 39.105 139.075 39.275 139.245 ;
        RECT 38.665 138.105 38.935 139.075 ;
        RECT 39.105 138.905 39.830 139.075 ;
        RECT 40.020 138.955 40.730 139.575 ;
        RECT 40.900 139.245 41.250 139.815 ;
        RECT 41.885 139.715 44.475 140.485 ;
        RECT 44.650 139.940 49.995 140.485 ;
        RECT 50.170 139.940 55.515 140.485 ;
        RECT 39.660 138.785 39.830 138.905 ;
        RECT 40.930 138.785 41.250 139.075 ;
        RECT 39.145 137.935 39.425 138.735 ;
        RECT 39.660 138.615 41.250 138.785 ;
        RECT 41.885 139.025 43.095 139.545 ;
        RECT 43.265 139.195 44.475 139.715 ;
        RECT 39.595 138.155 41.250 138.445 ;
        RECT 41.885 137.935 44.475 139.025 ;
        RECT 46.240 138.370 46.590 139.620 ;
        RECT 48.070 139.110 48.410 139.940 ;
        RECT 51.760 138.370 52.110 139.620 ;
        RECT 53.590 139.110 53.930 139.940 ;
        RECT 55.725 139.665 55.955 140.485 ;
        RECT 56.125 139.685 56.455 140.315 ;
        RECT 55.705 139.245 56.035 139.495 ;
        RECT 56.205 139.085 56.455 139.685 ;
        RECT 56.625 139.665 56.835 140.485 ;
        RECT 57.525 139.715 59.195 140.485 ;
        RECT 44.650 137.935 49.995 138.370 ;
        RECT 50.170 137.935 55.515 138.370 ;
        RECT 55.725 137.935 55.955 139.075 ;
        RECT 56.125 138.105 56.455 139.085 ;
        RECT 56.625 137.935 56.835 139.075 ;
        RECT 57.525 139.025 58.275 139.545 ;
        RECT 58.445 139.195 59.195 139.715 ;
        RECT 59.365 139.685 59.705 140.315 ;
        RECT 59.875 139.685 60.125 140.485 ;
        RECT 60.315 139.835 60.645 140.315 ;
        RECT 60.815 140.025 61.040 140.485 ;
        RECT 61.210 139.835 61.540 140.315 ;
        RECT 59.365 139.075 59.540 139.685 ;
        RECT 60.315 139.665 61.540 139.835 ;
        RECT 62.170 139.705 62.670 140.315 ;
        RECT 63.045 139.760 63.335 140.485 ;
        RECT 59.710 139.325 60.405 139.495 ;
        RECT 60.235 139.075 60.405 139.325 ;
        RECT 60.580 139.295 61.000 139.495 ;
        RECT 61.170 139.295 61.500 139.495 ;
        RECT 61.670 139.295 62.000 139.495 ;
        RECT 62.170 139.075 62.340 139.705 ;
        RECT 63.965 139.685 64.305 140.315 ;
        RECT 64.475 139.685 64.725 140.485 ;
        RECT 64.915 139.835 65.245 140.315 ;
        RECT 65.415 140.025 65.640 140.485 ;
        RECT 65.810 139.835 66.140 140.315 ;
        RECT 62.525 139.245 62.875 139.495 ;
        RECT 57.525 137.935 59.195 139.025 ;
        RECT 59.365 138.105 59.705 139.075 ;
        RECT 59.875 137.935 60.045 139.075 ;
        RECT 60.235 138.905 62.670 139.075 ;
        RECT 60.315 137.935 60.565 138.735 ;
        RECT 61.210 138.105 61.540 138.905 ;
        RECT 61.840 137.935 62.170 138.735 ;
        RECT 62.340 138.105 62.670 138.905 ;
        RECT 63.045 137.935 63.335 139.100 ;
        RECT 63.965 139.075 64.140 139.685 ;
        RECT 64.915 139.665 66.140 139.835 ;
        RECT 66.770 139.705 67.270 140.315 ;
        RECT 68.020 140.145 68.275 140.305 ;
        RECT 67.935 139.975 68.275 140.145 ;
        RECT 68.455 140.025 68.740 140.485 ;
        RECT 68.020 139.775 68.275 139.975 ;
        RECT 64.310 139.325 65.005 139.495 ;
        RECT 64.835 139.075 65.005 139.325 ;
        RECT 65.180 139.295 65.600 139.495 ;
        RECT 65.770 139.295 66.100 139.495 ;
        RECT 66.270 139.295 66.600 139.495 ;
        RECT 66.770 139.075 66.940 139.705 ;
        RECT 67.125 139.245 67.475 139.495 ;
        RECT 63.965 138.105 64.305 139.075 ;
        RECT 64.475 137.935 64.645 139.075 ;
        RECT 64.835 138.905 67.270 139.075 ;
        RECT 64.915 137.935 65.165 138.735 ;
        RECT 65.810 138.105 66.140 138.905 ;
        RECT 66.440 137.935 66.770 138.735 ;
        RECT 66.940 138.105 67.270 138.905 ;
        RECT 68.020 138.915 68.200 139.775 ;
        RECT 68.920 139.575 69.170 140.225 ;
        RECT 68.370 139.245 69.170 139.575 ;
        RECT 68.020 138.245 68.275 138.915 ;
        RECT 68.455 137.935 68.740 138.735 ;
        RECT 68.920 138.655 69.170 139.245 ;
        RECT 69.370 139.890 69.690 140.220 ;
        RECT 69.870 140.005 70.530 140.485 ;
        RECT 70.730 140.095 71.580 140.265 ;
        RECT 69.370 138.995 69.560 139.890 ;
        RECT 69.880 139.565 70.540 139.835 ;
        RECT 70.210 139.505 70.540 139.565 ;
        RECT 69.730 139.335 70.060 139.395 ;
        RECT 70.730 139.335 70.900 140.095 ;
        RECT 72.140 140.025 72.460 140.485 ;
        RECT 72.660 139.845 72.910 140.275 ;
        RECT 73.200 140.045 73.610 140.485 ;
        RECT 73.780 140.105 74.795 140.305 ;
        RECT 71.070 139.675 72.320 139.845 ;
        RECT 71.070 139.555 71.400 139.675 ;
        RECT 69.730 139.165 71.630 139.335 ;
        RECT 69.370 138.825 71.290 138.995 ;
        RECT 69.370 138.805 69.690 138.825 ;
        RECT 68.920 138.145 69.250 138.655 ;
        RECT 69.520 138.195 69.690 138.805 ;
        RECT 71.460 138.655 71.630 139.165 ;
        RECT 71.800 139.095 71.980 139.505 ;
        RECT 72.150 138.915 72.320 139.675 ;
        RECT 69.860 137.935 70.190 138.625 ;
        RECT 70.420 138.485 71.630 138.655 ;
        RECT 71.800 138.605 72.320 138.915 ;
        RECT 72.490 139.505 72.910 139.845 ;
        RECT 73.200 139.505 73.610 139.835 ;
        RECT 72.490 138.735 72.680 139.505 ;
        RECT 73.780 139.375 73.950 140.105 ;
        RECT 75.095 139.935 75.265 140.265 ;
        RECT 75.435 140.105 75.765 140.485 ;
        RECT 74.120 139.555 74.470 139.925 ;
        RECT 73.780 139.335 74.200 139.375 ;
        RECT 72.850 139.165 74.200 139.335 ;
        RECT 72.850 139.005 73.100 139.165 ;
        RECT 73.610 138.735 73.860 138.995 ;
        RECT 72.490 138.485 73.860 138.735 ;
        RECT 70.420 138.195 70.660 138.485 ;
        RECT 71.460 138.405 71.630 138.485 ;
        RECT 70.860 137.935 71.280 138.315 ;
        RECT 71.460 138.155 72.090 138.405 ;
        RECT 72.560 137.935 72.890 138.315 ;
        RECT 73.060 138.195 73.230 138.485 ;
        RECT 74.030 138.320 74.200 139.165 ;
        RECT 74.650 138.995 74.870 139.865 ;
        RECT 75.095 139.745 75.790 139.935 ;
        RECT 74.370 138.615 74.870 138.995 ;
        RECT 75.040 138.945 75.450 139.565 ;
        RECT 75.620 138.775 75.790 139.745 ;
        RECT 75.095 138.605 75.790 138.775 ;
        RECT 73.410 137.935 73.790 138.315 ;
        RECT 74.030 138.150 74.860 138.320 ;
        RECT 75.095 138.105 75.265 138.605 ;
        RECT 75.435 137.935 75.765 138.435 ;
        RECT 75.980 138.105 76.205 140.225 ;
        RECT 76.375 140.105 76.705 140.485 ;
        RECT 76.875 139.935 77.045 140.225 ;
        RECT 76.380 139.765 77.045 139.935 ;
        RECT 76.380 138.775 76.610 139.765 ;
        RECT 77.765 139.715 79.435 140.485 ;
        RECT 76.780 138.945 77.130 139.595 ;
        RECT 77.765 139.025 78.515 139.545 ;
        RECT 78.685 139.195 79.435 139.715 ;
        RECT 79.605 139.685 79.945 140.315 ;
        RECT 80.115 139.685 80.365 140.485 ;
        RECT 80.555 139.835 80.885 140.315 ;
        RECT 81.055 140.025 81.280 140.485 ;
        RECT 81.450 139.835 81.780 140.315 ;
        RECT 79.605 139.075 79.780 139.685 ;
        RECT 80.555 139.665 81.780 139.835 ;
        RECT 82.410 139.705 82.910 140.315 ;
        RECT 83.285 139.735 84.495 140.485 ;
        RECT 79.950 139.325 80.645 139.495 ;
        RECT 80.475 139.075 80.645 139.325 ;
        RECT 80.820 139.295 81.240 139.495 ;
        RECT 81.410 139.295 81.740 139.495 ;
        RECT 81.910 139.295 82.240 139.495 ;
        RECT 82.410 139.075 82.580 139.705 ;
        RECT 82.765 139.245 83.115 139.495 ;
        RECT 76.380 138.605 77.045 138.775 ;
        RECT 76.375 137.935 76.705 138.435 ;
        RECT 76.875 138.105 77.045 138.605 ;
        RECT 77.765 137.935 79.435 139.025 ;
        RECT 79.605 138.105 79.945 139.075 ;
        RECT 80.115 137.935 80.285 139.075 ;
        RECT 80.475 138.905 82.910 139.075 ;
        RECT 80.555 137.935 80.805 138.735 ;
        RECT 81.450 138.105 81.780 138.905 ;
        RECT 82.080 137.935 82.410 138.735 ;
        RECT 82.580 138.105 82.910 138.905 ;
        RECT 83.285 139.025 83.805 139.565 ;
        RECT 83.975 139.195 84.495 139.735 ;
        RECT 84.940 139.675 85.185 140.280 ;
        RECT 85.405 139.950 85.915 140.485 ;
        RECT 84.665 139.505 85.895 139.675 ;
        RECT 83.285 137.935 84.495 139.025 ;
        RECT 84.665 138.695 85.005 139.505 ;
        RECT 85.175 138.940 85.925 139.130 ;
        RECT 84.665 138.285 85.180 138.695 ;
        RECT 85.415 137.935 85.585 138.695 ;
        RECT 85.755 138.275 85.925 138.940 ;
        RECT 86.095 138.955 86.285 140.315 ;
        RECT 86.455 139.465 86.730 140.315 ;
        RECT 86.920 139.950 87.450 140.315 ;
        RECT 87.875 140.085 88.205 140.485 ;
        RECT 87.275 139.915 87.450 139.950 ;
        RECT 86.455 139.295 86.735 139.465 ;
        RECT 86.455 139.155 86.730 139.295 ;
        RECT 86.935 138.955 87.105 139.755 ;
        RECT 86.095 138.785 87.105 138.955 ;
        RECT 87.275 139.745 88.205 139.915 ;
        RECT 88.375 139.745 88.630 140.315 ;
        RECT 88.805 139.760 89.095 140.485 ;
        RECT 89.355 139.935 89.525 140.315 ;
        RECT 89.705 140.105 90.035 140.485 ;
        RECT 89.355 139.765 90.020 139.935 ;
        RECT 90.215 139.810 90.475 140.315 ;
        RECT 87.275 138.615 87.445 139.745 ;
        RECT 88.035 139.575 88.205 139.745 ;
        RECT 86.320 138.445 87.445 138.615 ;
        RECT 87.615 139.245 87.810 139.575 ;
        RECT 88.035 139.245 88.290 139.575 ;
        RECT 87.615 138.275 87.785 139.245 ;
        RECT 88.460 139.075 88.630 139.745 ;
        RECT 89.285 139.215 89.615 139.585 ;
        RECT 89.850 139.510 90.020 139.765 ;
        RECT 89.850 139.180 90.135 139.510 ;
        RECT 85.755 138.105 87.785 138.275 ;
        RECT 87.955 137.935 88.125 139.075 ;
        RECT 88.295 138.105 88.630 139.075 ;
        RECT 88.805 137.935 89.095 139.100 ;
        RECT 89.850 139.035 90.020 139.180 ;
        RECT 89.355 138.865 90.020 139.035 ;
        RECT 90.305 139.010 90.475 139.810 ;
        RECT 90.645 139.715 92.315 140.485 ;
        RECT 92.490 139.940 97.835 140.485 ;
        RECT 89.355 138.105 89.525 138.865 ;
        RECT 89.705 137.935 90.035 138.695 ;
        RECT 90.205 138.105 90.475 139.010 ;
        RECT 90.645 139.025 91.395 139.545 ;
        RECT 91.565 139.195 92.315 139.715 ;
        RECT 90.645 137.935 92.315 139.025 ;
        RECT 94.080 138.370 94.430 139.620 ;
        RECT 95.910 139.110 96.250 139.940 ;
        RECT 98.380 139.775 98.635 140.305 ;
        RECT 98.815 140.025 99.100 140.485 ;
        RECT 98.380 139.125 98.560 139.775 ;
        RECT 99.280 139.575 99.530 140.225 ;
        RECT 98.730 139.245 99.530 139.575 ;
        RECT 98.295 138.955 98.560 139.125 ;
        RECT 98.380 138.915 98.560 138.955 ;
        RECT 92.490 137.935 97.835 138.370 ;
        RECT 98.380 138.245 98.635 138.915 ;
        RECT 98.815 137.935 99.100 138.735 ;
        RECT 99.280 138.655 99.530 139.245 ;
        RECT 99.730 139.890 100.050 140.220 ;
        RECT 100.230 140.005 100.890 140.485 ;
        RECT 101.090 140.095 101.940 140.265 ;
        RECT 99.730 138.995 99.920 139.890 ;
        RECT 100.240 139.565 100.900 139.835 ;
        RECT 100.570 139.505 100.900 139.565 ;
        RECT 100.090 139.335 100.420 139.395 ;
        RECT 101.090 139.335 101.260 140.095 ;
        RECT 102.500 140.025 102.820 140.485 ;
        RECT 103.020 139.845 103.270 140.275 ;
        RECT 103.560 140.045 103.970 140.485 ;
        RECT 104.140 140.105 105.155 140.305 ;
        RECT 101.430 139.675 102.680 139.845 ;
        RECT 101.430 139.555 101.760 139.675 ;
        RECT 100.090 139.165 101.990 139.335 ;
        RECT 99.730 138.825 101.650 138.995 ;
        RECT 99.730 138.805 100.050 138.825 ;
        RECT 99.280 138.145 99.610 138.655 ;
        RECT 99.880 138.195 100.050 138.805 ;
        RECT 101.820 138.655 101.990 139.165 ;
        RECT 102.160 139.095 102.340 139.505 ;
        RECT 102.510 138.915 102.680 139.675 ;
        RECT 100.220 137.935 100.550 138.625 ;
        RECT 100.780 138.485 101.990 138.655 ;
        RECT 102.160 138.605 102.680 138.915 ;
        RECT 102.850 139.505 103.270 139.845 ;
        RECT 103.560 139.505 103.970 139.835 ;
        RECT 102.850 138.735 103.040 139.505 ;
        RECT 104.140 139.375 104.310 140.105 ;
        RECT 105.455 139.935 105.625 140.265 ;
        RECT 105.795 140.105 106.125 140.485 ;
        RECT 104.480 139.555 104.830 139.925 ;
        RECT 104.140 139.335 104.560 139.375 ;
        RECT 103.210 139.165 104.560 139.335 ;
        RECT 103.210 139.005 103.460 139.165 ;
        RECT 103.970 138.735 104.220 138.995 ;
        RECT 102.850 138.485 104.220 138.735 ;
        RECT 100.780 138.195 101.020 138.485 ;
        RECT 101.820 138.405 101.990 138.485 ;
        RECT 101.220 137.935 101.640 138.315 ;
        RECT 101.820 138.155 102.450 138.405 ;
        RECT 102.920 137.935 103.250 138.315 ;
        RECT 103.420 138.195 103.590 138.485 ;
        RECT 104.390 138.320 104.560 139.165 ;
        RECT 105.010 138.995 105.230 139.865 ;
        RECT 105.455 139.745 106.150 139.935 ;
        RECT 104.730 138.615 105.230 138.995 ;
        RECT 105.400 138.945 105.810 139.565 ;
        RECT 105.980 138.775 106.150 139.745 ;
        RECT 105.455 138.605 106.150 138.775 ;
        RECT 103.770 137.935 104.150 138.315 ;
        RECT 104.390 138.150 105.220 138.320 ;
        RECT 105.455 138.105 105.625 138.605 ;
        RECT 105.795 137.935 106.125 138.435 ;
        RECT 106.340 138.105 106.565 140.225 ;
        RECT 106.735 140.105 107.065 140.485 ;
        RECT 107.235 139.935 107.405 140.225 ;
        RECT 106.740 139.765 107.405 139.935 ;
        RECT 106.740 138.775 106.970 139.765 ;
        RECT 108.125 139.715 109.795 140.485 ;
        RECT 107.140 138.945 107.490 139.595 ;
        RECT 108.125 139.025 108.875 139.545 ;
        RECT 109.045 139.195 109.795 139.715 ;
        RECT 110.170 139.705 110.670 140.315 ;
        RECT 109.965 139.245 110.315 139.495 ;
        RECT 110.500 139.075 110.670 139.705 ;
        RECT 111.300 139.835 111.630 140.315 ;
        RECT 111.800 140.025 112.025 140.485 ;
        RECT 112.195 139.835 112.525 140.315 ;
        RECT 111.300 139.665 112.525 139.835 ;
        RECT 112.715 139.685 112.965 140.485 ;
        RECT 113.135 139.685 113.475 140.315 ;
        RECT 114.565 139.760 114.855 140.485 ;
        RECT 113.245 139.635 113.475 139.685 ;
        RECT 115.525 139.665 115.755 140.485 ;
        RECT 115.925 139.685 116.255 140.315 ;
        RECT 110.840 139.295 111.170 139.495 ;
        RECT 111.340 139.295 111.670 139.495 ;
        RECT 111.840 139.295 112.260 139.495 ;
        RECT 112.435 139.325 113.130 139.495 ;
        RECT 112.435 139.075 112.605 139.325 ;
        RECT 113.300 139.075 113.475 139.635 ;
        RECT 115.505 139.245 115.835 139.495 ;
        RECT 106.740 138.605 107.405 138.775 ;
        RECT 106.735 137.935 107.065 138.435 ;
        RECT 107.235 138.105 107.405 138.605 ;
        RECT 108.125 137.935 109.795 139.025 ;
        RECT 110.170 138.905 112.605 139.075 ;
        RECT 110.170 138.105 110.500 138.905 ;
        RECT 110.670 137.935 111.000 138.735 ;
        RECT 111.300 138.105 111.630 138.905 ;
        RECT 112.275 137.935 112.525 138.735 ;
        RECT 112.795 137.935 112.965 139.075 ;
        RECT 113.135 138.105 113.475 139.075 ;
        RECT 114.565 137.935 114.855 139.100 ;
        RECT 116.005 139.085 116.255 139.685 ;
        RECT 116.425 139.665 116.635 140.485 ;
        RECT 117.240 139.805 117.495 140.305 ;
        RECT 117.675 140.025 117.960 140.485 ;
        RECT 117.155 139.775 117.495 139.805 ;
        RECT 117.155 139.635 117.420 139.775 ;
        RECT 115.525 137.935 115.755 139.075 ;
        RECT 115.925 138.105 116.255 139.085 ;
        RECT 116.425 137.935 116.635 139.075 ;
        RECT 117.240 138.915 117.420 139.635 ;
        RECT 118.140 139.575 118.390 140.225 ;
        RECT 117.590 139.245 118.390 139.575 ;
        RECT 117.240 138.245 117.495 138.915 ;
        RECT 117.675 137.935 117.960 138.735 ;
        RECT 118.140 138.655 118.390 139.245 ;
        RECT 118.590 139.890 118.910 140.220 ;
        RECT 119.090 140.005 119.750 140.485 ;
        RECT 119.950 140.095 120.800 140.265 ;
        RECT 118.590 138.995 118.780 139.890 ;
        RECT 119.100 139.565 119.760 139.835 ;
        RECT 119.430 139.505 119.760 139.565 ;
        RECT 118.950 139.335 119.280 139.395 ;
        RECT 119.950 139.335 120.120 140.095 ;
        RECT 121.360 140.025 121.680 140.485 ;
        RECT 121.880 139.845 122.130 140.275 ;
        RECT 122.420 140.045 122.830 140.485 ;
        RECT 123.000 140.105 124.015 140.305 ;
        RECT 120.290 139.675 121.540 139.845 ;
        RECT 120.290 139.555 120.620 139.675 ;
        RECT 118.950 139.165 120.850 139.335 ;
        RECT 118.590 138.825 120.510 138.995 ;
        RECT 118.590 138.805 118.910 138.825 ;
        RECT 118.140 138.145 118.470 138.655 ;
        RECT 118.740 138.195 118.910 138.805 ;
        RECT 120.680 138.655 120.850 139.165 ;
        RECT 121.020 139.095 121.200 139.505 ;
        RECT 121.370 138.915 121.540 139.675 ;
        RECT 119.080 137.935 119.410 138.625 ;
        RECT 119.640 138.485 120.850 138.655 ;
        RECT 121.020 138.605 121.540 138.915 ;
        RECT 121.710 139.505 122.130 139.845 ;
        RECT 122.420 139.505 122.830 139.835 ;
        RECT 121.710 138.735 121.900 139.505 ;
        RECT 123.000 139.375 123.170 140.105 ;
        RECT 124.315 139.935 124.485 140.265 ;
        RECT 124.655 140.105 124.985 140.485 ;
        RECT 123.340 139.555 123.690 139.925 ;
        RECT 123.000 139.335 123.420 139.375 ;
        RECT 122.070 139.165 123.420 139.335 ;
        RECT 122.070 139.005 122.320 139.165 ;
        RECT 122.830 138.735 123.080 138.995 ;
        RECT 121.710 138.485 123.080 138.735 ;
        RECT 119.640 138.195 119.880 138.485 ;
        RECT 120.680 138.405 120.850 138.485 ;
        RECT 120.080 137.935 120.500 138.315 ;
        RECT 120.680 138.155 121.310 138.405 ;
        RECT 121.780 137.935 122.110 138.315 ;
        RECT 122.280 138.195 122.450 138.485 ;
        RECT 123.250 138.320 123.420 139.165 ;
        RECT 123.870 138.995 124.090 139.865 ;
        RECT 124.315 139.745 125.010 139.935 ;
        RECT 123.590 138.615 124.090 138.995 ;
        RECT 124.260 138.945 124.670 139.565 ;
        RECT 124.840 138.775 125.010 139.745 ;
        RECT 124.315 138.605 125.010 138.775 ;
        RECT 122.630 137.935 123.010 138.315 ;
        RECT 123.250 138.150 124.080 138.320 ;
        RECT 124.315 138.105 124.485 138.605 ;
        RECT 124.655 137.935 124.985 138.435 ;
        RECT 125.200 138.105 125.425 140.225 ;
        RECT 125.595 140.105 125.925 140.485 ;
        RECT 126.095 139.935 126.265 140.225 ;
        RECT 125.600 139.765 126.265 139.935 ;
        RECT 125.600 138.775 125.830 139.765 ;
        RECT 126.525 139.735 127.735 140.485 ;
        RECT 126.000 138.945 126.350 139.595 ;
        RECT 126.525 139.025 127.045 139.565 ;
        RECT 127.215 139.195 127.735 139.735 ;
        RECT 125.600 138.605 126.265 138.775 ;
        RECT 125.595 137.935 125.925 138.435 ;
        RECT 126.095 138.105 126.265 138.605 ;
        RECT 126.525 137.935 127.735 139.025 ;
        RECT 14.660 137.765 127.820 137.935 ;
        RECT 14.745 136.675 15.955 137.765 ;
        RECT 14.745 135.965 15.265 136.505 ;
        RECT 15.435 136.135 15.955 136.675 ;
        RECT 16.585 136.675 20.095 137.765 ;
        RECT 16.585 136.155 18.275 136.675 ;
        RECT 20.270 136.625 20.605 137.595 ;
        RECT 20.775 136.625 20.945 137.765 ;
        RECT 21.115 137.425 23.145 137.595 ;
        RECT 18.445 135.985 20.095 136.505 ;
        RECT 14.745 135.215 15.955 135.965 ;
        RECT 16.585 135.215 20.095 135.985 ;
        RECT 20.270 135.955 20.440 136.625 ;
        RECT 21.115 136.455 21.285 137.425 ;
        RECT 20.610 136.125 20.865 136.455 ;
        RECT 21.090 136.125 21.285 136.455 ;
        RECT 21.455 137.085 22.580 137.255 ;
        RECT 20.695 135.955 20.865 136.125 ;
        RECT 21.455 135.955 21.625 137.085 ;
        RECT 20.270 135.385 20.525 135.955 ;
        RECT 20.695 135.785 21.625 135.955 ;
        RECT 21.795 136.745 22.805 136.915 ;
        RECT 21.795 135.945 21.965 136.745 ;
        RECT 22.170 136.405 22.445 136.545 ;
        RECT 22.165 136.235 22.445 136.405 ;
        RECT 21.450 135.750 21.625 135.785 ;
        RECT 20.695 135.215 21.025 135.615 ;
        RECT 21.450 135.385 21.980 135.750 ;
        RECT 22.170 135.385 22.445 136.235 ;
        RECT 22.615 135.385 22.805 136.745 ;
        RECT 22.975 136.760 23.145 137.425 ;
        RECT 23.315 137.005 23.485 137.765 ;
        RECT 23.720 137.005 24.235 137.415 ;
        RECT 22.975 136.570 23.725 136.760 ;
        RECT 23.895 136.195 24.235 137.005 ;
        RECT 24.405 136.600 24.695 137.765 ;
        RECT 24.865 136.675 28.375 137.765 ;
        RECT 23.005 136.025 24.235 136.195 ;
        RECT 24.865 136.155 26.555 136.675 ;
        RECT 28.550 136.625 28.885 137.595 ;
        RECT 29.055 136.625 29.225 137.765 ;
        RECT 29.395 137.425 31.425 137.595 ;
        RECT 22.985 135.215 23.495 135.750 ;
        RECT 23.715 135.420 23.960 136.025 ;
        RECT 26.725 135.985 28.375 136.505 ;
        RECT 24.405 135.215 24.695 135.940 ;
        RECT 24.865 135.215 28.375 135.985 ;
        RECT 28.550 135.955 28.720 136.625 ;
        RECT 29.395 136.455 29.565 137.425 ;
        RECT 28.890 136.125 29.145 136.455 ;
        RECT 29.370 136.125 29.565 136.455 ;
        RECT 29.735 137.085 30.860 137.255 ;
        RECT 28.975 135.955 29.145 136.125 ;
        RECT 29.735 135.955 29.905 137.085 ;
        RECT 28.550 135.385 28.805 135.955 ;
        RECT 28.975 135.785 29.905 135.955 ;
        RECT 30.075 136.745 31.085 136.915 ;
        RECT 30.075 135.945 30.245 136.745 ;
        RECT 30.450 136.065 30.725 136.545 ;
        RECT 30.445 135.895 30.725 136.065 ;
        RECT 29.730 135.750 29.905 135.785 ;
        RECT 28.975 135.215 29.305 135.615 ;
        RECT 29.730 135.385 30.260 135.750 ;
        RECT 30.450 135.385 30.725 135.895 ;
        RECT 30.895 135.385 31.085 136.745 ;
        RECT 31.255 136.760 31.425 137.425 ;
        RECT 31.595 137.005 31.765 137.765 ;
        RECT 32.000 137.005 32.515 137.415 ;
        RECT 32.885 137.095 33.165 137.765 ;
        RECT 31.255 136.570 32.005 136.760 ;
        RECT 32.175 136.195 32.515 137.005 ;
        RECT 33.335 136.875 33.635 137.425 ;
        RECT 33.835 137.045 34.165 137.765 ;
        RECT 34.355 137.045 34.815 137.595 ;
        RECT 32.700 136.455 32.965 136.815 ;
        RECT 33.335 136.705 34.275 136.875 ;
        RECT 34.105 136.455 34.275 136.705 ;
        RECT 32.700 136.205 33.375 136.455 ;
        RECT 33.595 136.205 33.935 136.455 ;
        RECT 31.285 136.025 32.515 136.195 ;
        RECT 34.105 136.125 34.395 136.455 ;
        RECT 34.105 136.035 34.275 136.125 ;
        RECT 31.265 135.215 31.775 135.750 ;
        RECT 31.995 135.420 32.240 136.025 ;
        RECT 32.885 135.845 34.275 136.035 ;
        RECT 32.885 135.485 33.215 135.845 ;
        RECT 34.565 135.675 34.815 137.045 ;
        RECT 33.835 135.215 34.085 135.675 ;
        RECT 34.255 135.385 34.815 135.675 ;
        RECT 34.985 136.625 35.255 137.595 ;
        RECT 35.465 136.965 35.745 137.765 ;
        RECT 35.915 137.255 37.570 137.545 ;
        RECT 35.980 136.915 37.570 137.085 ;
        RECT 35.980 136.795 36.150 136.915 ;
        RECT 35.425 136.625 36.150 136.795 ;
        RECT 34.985 135.890 35.155 136.625 ;
        RECT 35.425 136.455 35.595 136.625 ;
        RECT 35.325 136.125 35.595 136.455 ;
        RECT 35.765 136.125 36.170 136.455 ;
        RECT 36.340 136.125 37.050 136.745 ;
        RECT 37.250 136.625 37.570 136.915 ;
        RECT 37.745 136.625 38.015 137.595 ;
        RECT 38.225 136.965 38.505 137.765 ;
        RECT 38.675 137.255 40.330 137.545 ;
        RECT 38.740 136.915 40.330 137.085 ;
        RECT 38.740 136.795 38.910 136.915 ;
        RECT 38.185 136.625 38.910 136.795 ;
        RECT 35.425 135.955 35.595 136.125 ;
        RECT 34.985 135.545 35.255 135.890 ;
        RECT 35.425 135.785 37.035 135.955 ;
        RECT 37.220 135.885 37.570 136.455 ;
        RECT 37.745 135.890 37.915 136.625 ;
        RECT 38.185 136.455 38.355 136.625 ;
        RECT 38.085 136.125 38.355 136.455 ;
        RECT 38.525 136.125 38.930 136.455 ;
        RECT 39.100 136.125 39.810 136.745 ;
        RECT 40.010 136.625 40.330 136.915 ;
        RECT 40.965 136.675 43.555 137.765 ;
        RECT 38.185 135.955 38.355 136.125 ;
        RECT 35.445 135.215 35.825 135.615 ;
        RECT 35.995 135.435 36.165 135.785 ;
        RECT 36.335 135.215 36.665 135.615 ;
        RECT 36.865 135.435 37.035 135.785 ;
        RECT 37.235 135.215 37.565 135.715 ;
        RECT 37.745 135.545 38.015 135.890 ;
        RECT 38.185 135.785 39.795 135.955 ;
        RECT 39.980 135.885 40.330 136.455 ;
        RECT 40.965 136.155 42.175 136.675 ;
        RECT 43.725 136.625 43.995 137.595 ;
        RECT 44.205 136.965 44.485 137.765 ;
        RECT 44.655 137.255 46.310 137.545 ;
        RECT 44.720 136.915 46.310 137.085 ;
        RECT 44.720 136.795 44.890 136.915 ;
        RECT 44.165 136.625 44.890 136.795 ;
        RECT 42.345 135.985 43.555 136.505 ;
        RECT 38.205 135.215 38.585 135.615 ;
        RECT 38.755 135.435 38.925 135.785 ;
        RECT 39.095 135.215 39.425 135.615 ;
        RECT 39.625 135.435 39.795 135.785 ;
        RECT 39.995 135.215 40.325 135.715 ;
        RECT 40.965 135.215 43.555 135.985 ;
        RECT 43.725 135.890 43.895 136.625 ;
        RECT 44.165 136.455 44.335 136.625 ;
        RECT 45.080 136.575 45.795 136.745 ;
        RECT 45.990 136.625 46.310 136.915 ;
        RECT 46.485 136.625 46.825 137.595 ;
        RECT 46.995 136.625 47.165 137.765 ;
        RECT 47.435 136.965 47.685 137.765 ;
        RECT 48.330 136.795 48.660 137.595 ;
        RECT 48.960 136.965 49.290 137.765 ;
        RECT 49.460 136.795 49.790 137.595 ;
        RECT 47.355 136.625 49.790 136.795 ;
        RECT 44.065 136.125 44.335 136.455 ;
        RECT 44.505 136.125 44.910 136.455 ;
        RECT 45.080 136.125 45.790 136.575 ;
        RECT 44.165 135.955 44.335 136.125 ;
        RECT 43.725 135.545 43.995 135.890 ;
        RECT 44.165 135.785 45.775 135.955 ;
        RECT 45.960 135.885 46.310 136.455 ;
        RECT 46.485 136.065 46.660 136.625 ;
        RECT 47.355 136.375 47.525 136.625 ;
        RECT 46.830 136.205 47.525 136.375 ;
        RECT 47.700 136.205 48.120 136.405 ;
        RECT 48.290 136.205 48.620 136.405 ;
        RECT 48.790 136.205 49.120 136.405 ;
        RECT 46.485 136.015 46.715 136.065 ;
        RECT 44.185 135.215 44.565 135.615 ;
        RECT 44.735 135.435 44.905 135.785 ;
        RECT 45.075 135.215 45.405 135.615 ;
        RECT 45.605 135.435 45.775 135.785 ;
        RECT 45.975 135.215 46.305 135.715 ;
        RECT 46.485 135.385 46.825 136.015 ;
        RECT 46.995 135.215 47.245 136.015 ;
        RECT 47.435 135.865 48.660 136.035 ;
        RECT 47.435 135.385 47.765 135.865 ;
        RECT 47.935 135.215 48.160 135.675 ;
        RECT 48.330 135.385 48.660 135.865 ;
        RECT 49.290 135.995 49.460 136.625 ;
        RECT 50.165 136.600 50.455 137.765 ;
        RECT 50.625 136.675 53.215 137.765 ;
        RECT 53.385 137.005 53.900 137.415 ;
        RECT 54.135 137.005 54.305 137.765 ;
        RECT 54.475 137.425 56.505 137.595 ;
        RECT 49.645 136.205 49.995 136.455 ;
        RECT 50.625 136.155 51.835 136.675 ;
        RECT 49.290 135.385 49.790 135.995 ;
        RECT 52.005 135.985 53.215 136.505 ;
        RECT 53.385 136.195 53.725 137.005 ;
        RECT 54.475 136.760 54.645 137.425 ;
        RECT 55.040 137.085 56.165 137.255 ;
        RECT 53.895 136.570 54.645 136.760 ;
        RECT 54.815 136.745 55.825 136.915 ;
        RECT 53.385 136.025 54.615 136.195 ;
        RECT 50.165 135.215 50.455 135.940 ;
        RECT 50.625 135.215 53.215 135.985 ;
        RECT 53.660 135.420 53.905 136.025 ;
        RECT 54.125 135.215 54.635 135.750 ;
        RECT 54.815 135.385 55.005 136.745 ;
        RECT 55.175 136.405 55.450 136.545 ;
        RECT 55.175 136.235 55.455 136.405 ;
        RECT 55.175 135.385 55.450 136.235 ;
        RECT 55.655 135.945 55.825 136.745 ;
        RECT 55.995 135.955 56.165 137.085 ;
        RECT 56.335 136.455 56.505 137.425 ;
        RECT 56.675 136.625 56.845 137.765 ;
        RECT 57.015 136.625 57.350 137.595 ;
        RECT 58.075 136.835 58.245 137.595 ;
        RECT 58.425 137.005 58.755 137.765 ;
        RECT 58.075 136.665 58.740 136.835 ;
        RECT 58.925 136.690 59.195 137.595 ;
        RECT 56.335 136.125 56.530 136.455 ;
        RECT 56.755 136.125 57.010 136.455 ;
        RECT 56.755 135.955 56.925 136.125 ;
        RECT 57.180 135.955 57.350 136.625 ;
        RECT 58.570 136.520 58.740 136.665 ;
        RECT 58.005 136.115 58.335 136.485 ;
        RECT 58.570 136.190 58.855 136.520 ;
        RECT 55.995 135.785 56.925 135.955 ;
        RECT 55.995 135.750 56.170 135.785 ;
        RECT 55.640 135.385 56.170 135.750 ;
        RECT 56.595 135.215 56.925 135.615 ;
        RECT 57.095 135.385 57.350 135.955 ;
        RECT 58.570 135.935 58.740 136.190 ;
        RECT 58.075 135.765 58.740 135.935 ;
        RECT 59.025 135.890 59.195 136.690 ;
        RECT 59.365 136.675 61.035 137.765 ;
        RECT 59.365 136.155 60.115 136.675 ;
        RECT 61.205 136.625 61.545 137.595 ;
        RECT 61.715 136.625 61.885 137.765 ;
        RECT 62.155 136.965 62.405 137.765 ;
        RECT 63.050 136.795 63.380 137.595 ;
        RECT 63.680 136.965 64.010 137.765 ;
        RECT 64.180 136.795 64.510 137.595 ;
        RECT 65.000 137.135 65.285 137.595 ;
        RECT 65.455 137.305 65.725 137.765 ;
        RECT 65.000 136.915 65.955 137.135 ;
        RECT 62.075 136.625 64.510 136.795 ;
        RECT 60.285 135.985 61.035 136.505 ;
        RECT 58.075 135.385 58.245 135.765 ;
        RECT 58.425 135.215 58.755 135.595 ;
        RECT 58.935 135.385 59.195 135.890 ;
        RECT 59.365 135.215 61.035 135.985 ;
        RECT 61.205 136.015 61.380 136.625 ;
        RECT 62.075 136.375 62.245 136.625 ;
        RECT 61.550 136.205 62.245 136.375 ;
        RECT 62.420 136.205 62.840 136.405 ;
        RECT 63.010 136.205 63.340 136.405 ;
        RECT 63.510 136.205 63.840 136.405 ;
        RECT 61.205 135.385 61.545 136.015 ;
        RECT 61.715 135.215 61.965 136.015 ;
        RECT 62.155 135.865 63.380 136.035 ;
        RECT 62.155 135.385 62.485 135.865 ;
        RECT 62.655 135.215 62.880 135.675 ;
        RECT 63.050 135.385 63.380 135.865 ;
        RECT 64.010 135.995 64.180 136.625 ;
        RECT 64.365 136.205 64.715 136.455 ;
        RECT 64.885 136.185 65.575 136.745 ;
        RECT 65.745 136.015 65.955 136.915 ;
        RECT 64.010 135.385 64.510 135.995 ;
        RECT 65.000 135.845 65.955 136.015 ;
        RECT 66.125 136.745 66.525 137.595 ;
        RECT 66.715 137.135 66.995 137.595 ;
        RECT 67.515 137.305 67.840 137.765 ;
        RECT 66.715 136.915 67.840 137.135 ;
        RECT 66.125 136.185 67.220 136.745 ;
        RECT 67.390 136.455 67.840 136.915 ;
        RECT 68.010 136.625 68.395 137.595 ;
        RECT 65.000 135.385 65.285 135.845 ;
        RECT 65.455 135.215 65.725 135.675 ;
        RECT 66.125 135.385 66.525 136.185 ;
        RECT 67.390 136.125 67.945 136.455 ;
        RECT 67.390 136.015 67.840 136.125 ;
        RECT 66.715 135.845 67.840 136.015 ;
        RECT 68.115 135.955 68.395 136.625 ;
        RECT 68.570 137.375 68.905 137.595 ;
        RECT 69.910 137.385 70.265 137.765 ;
        RECT 68.570 136.755 68.825 137.375 ;
        RECT 69.075 137.215 69.305 137.255 ;
        RECT 70.435 137.215 70.685 137.595 ;
        RECT 69.075 137.015 70.685 137.215 ;
        RECT 69.075 136.925 69.260 137.015 ;
        RECT 69.850 137.005 70.685 137.015 ;
        RECT 70.935 136.985 71.185 137.765 ;
        RECT 71.355 136.915 71.615 137.595 ;
        RECT 69.415 136.815 69.745 136.845 ;
        RECT 69.415 136.755 71.215 136.815 ;
        RECT 68.570 136.645 71.275 136.755 ;
        RECT 68.570 136.585 69.745 136.645 ;
        RECT 71.075 136.610 71.275 136.645 ;
        RECT 68.565 136.205 69.055 136.405 ;
        RECT 69.245 136.205 69.720 136.415 ;
        RECT 66.715 135.385 66.995 135.845 ;
        RECT 67.515 135.215 67.840 135.675 ;
        RECT 68.010 135.385 68.395 135.955 ;
        RECT 68.570 135.215 69.025 135.980 ;
        RECT 69.500 135.805 69.720 136.205 ;
        RECT 69.965 136.205 70.295 136.415 ;
        RECT 69.965 135.805 70.175 136.205 ;
        RECT 70.465 136.170 70.875 136.475 ;
        RECT 71.105 136.035 71.275 136.610 ;
        RECT 71.005 135.915 71.275 136.035 ;
        RECT 70.430 135.870 71.275 135.915 ;
        RECT 70.430 135.745 71.185 135.870 ;
        RECT 70.430 135.595 70.600 135.745 ;
        RECT 71.445 135.715 71.615 136.915 ;
        RECT 72.245 136.675 75.755 137.765 ;
        RECT 72.245 136.155 73.935 136.675 ;
        RECT 75.925 136.600 76.215 137.765 ;
        RECT 77.305 136.625 77.575 137.595 ;
        RECT 77.785 136.965 78.065 137.765 ;
        RECT 78.235 137.255 79.890 137.545 ;
        RECT 78.300 136.915 79.890 137.085 ;
        RECT 78.300 136.795 78.470 136.915 ;
        RECT 77.745 136.625 78.470 136.795 ;
        RECT 74.105 135.985 75.755 136.505 ;
        RECT 69.300 135.385 70.600 135.595 ;
        RECT 70.855 135.215 71.185 135.575 ;
        RECT 71.355 135.385 71.615 135.715 ;
        RECT 72.245 135.215 75.755 135.985 ;
        RECT 75.925 135.215 76.215 135.940 ;
        RECT 77.305 135.890 77.475 136.625 ;
        RECT 77.745 136.455 77.915 136.625 ;
        RECT 77.645 136.125 77.915 136.455 ;
        RECT 78.085 136.125 78.490 136.455 ;
        RECT 78.660 136.125 79.370 136.745 ;
        RECT 79.570 136.625 79.890 136.915 ;
        RECT 80.065 136.625 80.405 137.595 ;
        RECT 80.575 136.625 80.745 137.765 ;
        RECT 81.015 136.965 81.265 137.765 ;
        RECT 81.910 136.795 82.240 137.595 ;
        RECT 82.540 136.965 82.870 137.765 ;
        RECT 83.040 136.795 83.370 137.595 ;
        RECT 84.120 137.425 84.375 137.455 ;
        RECT 84.035 137.255 84.375 137.425 ;
        RECT 80.935 136.625 83.370 136.795 ;
        RECT 84.120 136.785 84.375 137.255 ;
        RECT 84.555 136.965 84.840 137.765 ;
        RECT 85.020 137.045 85.350 137.555 ;
        RECT 77.745 135.955 77.915 136.125 ;
        RECT 77.305 135.545 77.575 135.890 ;
        RECT 77.745 135.785 79.355 135.955 ;
        RECT 79.540 135.885 79.890 136.455 ;
        RECT 80.065 136.015 80.240 136.625 ;
        RECT 80.935 136.375 81.105 136.625 ;
        RECT 80.410 136.205 81.105 136.375 ;
        RECT 81.280 136.205 81.700 136.405 ;
        RECT 81.870 136.205 82.200 136.405 ;
        RECT 82.370 136.205 82.700 136.405 ;
        RECT 77.765 135.215 78.145 135.615 ;
        RECT 78.315 135.435 78.485 135.785 ;
        RECT 78.655 135.215 78.985 135.615 ;
        RECT 79.185 135.435 79.355 135.785 ;
        RECT 79.555 135.215 79.885 135.715 ;
        RECT 80.065 135.385 80.405 136.015 ;
        RECT 80.575 135.215 80.825 136.015 ;
        RECT 81.015 135.865 82.240 136.035 ;
        RECT 81.015 135.385 81.345 135.865 ;
        RECT 81.515 135.215 81.740 135.675 ;
        RECT 81.910 135.385 82.240 135.865 ;
        RECT 82.870 135.995 83.040 136.625 ;
        RECT 83.225 136.205 83.575 136.455 ;
        RECT 82.870 135.385 83.370 135.995 ;
        RECT 84.120 135.925 84.300 136.785 ;
        RECT 85.020 136.455 85.270 137.045 ;
        RECT 85.620 136.895 85.790 137.505 ;
        RECT 85.960 137.075 86.290 137.765 ;
        RECT 86.520 137.215 86.760 137.505 ;
        RECT 86.960 137.385 87.380 137.765 ;
        RECT 87.560 137.295 88.190 137.545 ;
        RECT 88.660 137.385 88.990 137.765 ;
        RECT 87.560 137.215 87.730 137.295 ;
        RECT 89.160 137.215 89.330 137.505 ;
        RECT 89.510 137.385 89.890 137.765 ;
        RECT 90.130 137.380 90.960 137.550 ;
        RECT 86.520 137.045 87.730 137.215 ;
        RECT 84.470 136.125 85.270 136.455 ;
        RECT 84.120 135.395 84.375 135.925 ;
        RECT 84.555 135.215 84.840 135.675 ;
        RECT 85.020 135.475 85.270 136.125 ;
        RECT 85.470 136.875 85.790 136.895 ;
        RECT 85.470 136.705 87.390 136.875 ;
        RECT 85.470 135.810 85.660 136.705 ;
        RECT 87.560 136.535 87.730 137.045 ;
        RECT 87.900 136.785 88.420 137.095 ;
        RECT 85.830 136.365 87.730 136.535 ;
        RECT 85.830 136.305 86.160 136.365 ;
        RECT 86.310 136.135 86.640 136.195 ;
        RECT 85.980 135.865 86.640 136.135 ;
        RECT 85.470 135.480 85.790 135.810 ;
        RECT 85.970 135.215 86.630 135.695 ;
        RECT 86.830 135.605 87.000 136.365 ;
        RECT 87.900 136.195 88.080 136.605 ;
        RECT 87.170 136.025 87.500 136.145 ;
        RECT 88.250 136.025 88.420 136.785 ;
        RECT 87.170 135.855 88.420 136.025 ;
        RECT 88.590 136.965 89.960 137.215 ;
        RECT 88.590 136.195 88.780 136.965 ;
        RECT 89.710 136.705 89.960 136.965 ;
        RECT 88.950 136.535 89.200 136.695 ;
        RECT 90.130 136.535 90.300 137.380 ;
        RECT 91.195 137.095 91.365 137.595 ;
        RECT 91.535 137.265 91.865 137.765 ;
        RECT 90.470 136.705 90.970 137.085 ;
        RECT 91.195 136.925 91.890 137.095 ;
        RECT 88.950 136.365 90.300 136.535 ;
        RECT 89.880 136.325 90.300 136.365 ;
        RECT 88.590 135.855 89.010 136.195 ;
        RECT 89.300 135.865 89.710 136.195 ;
        RECT 86.830 135.435 87.680 135.605 ;
        RECT 88.240 135.215 88.560 135.675 ;
        RECT 88.760 135.425 89.010 135.855 ;
        RECT 89.300 135.215 89.710 135.655 ;
        RECT 89.880 135.595 90.050 136.325 ;
        RECT 90.220 135.775 90.570 136.145 ;
        RECT 90.750 135.835 90.970 136.705 ;
        RECT 91.140 136.135 91.550 136.755 ;
        RECT 91.720 135.955 91.890 136.925 ;
        RECT 91.195 135.765 91.890 135.955 ;
        RECT 89.880 135.395 90.895 135.595 ;
        RECT 91.195 135.435 91.365 135.765 ;
        RECT 91.535 135.215 91.865 135.595 ;
        RECT 92.080 135.475 92.305 137.595 ;
        RECT 92.475 137.265 92.805 137.765 ;
        RECT 92.975 137.095 93.145 137.595 ;
        RECT 92.480 136.925 93.145 137.095 ;
        RECT 92.480 135.935 92.710 136.925 ;
        RECT 92.880 136.105 93.230 136.755 ;
        RECT 93.410 136.625 93.745 137.595 ;
        RECT 93.915 136.625 94.085 137.765 ;
        RECT 94.255 137.425 96.285 137.595 ;
        RECT 93.410 135.955 93.580 136.625 ;
        RECT 94.255 136.455 94.425 137.425 ;
        RECT 93.750 136.125 94.005 136.455 ;
        RECT 94.230 136.125 94.425 136.455 ;
        RECT 94.595 137.085 95.720 137.255 ;
        RECT 93.835 135.955 94.005 136.125 ;
        RECT 94.595 135.955 94.765 137.085 ;
        RECT 92.480 135.765 93.145 135.935 ;
        RECT 92.475 135.215 92.805 135.595 ;
        RECT 92.975 135.475 93.145 135.765 ;
        RECT 93.410 135.385 93.665 135.955 ;
        RECT 93.835 135.785 94.765 135.955 ;
        RECT 94.935 136.745 95.945 136.915 ;
        RECT 94.935 135.945 95.105 136.745 ;
        RECT 94.590 135.750 94.765 135.785 ;
        RECT 93.835 135.215 94.165 135.615 ;
        RECT 94.590 135.385 95.120 135.750 ;
        RECT 95.310 135.725 95.585 136.545 ;
        RECT 95.305 135.555 95.585 135.725 ;
        RECT 95.310 135.385 95.585 135.555 ;
        RECT 95.755 135.385 95.945 136.745 ;
        RECT 96.115 136.760 96.285 137.425 ;
        RECT 96.455 137.005 96.625 137.765 ;
        RECT 96.860 137.005 97.375 137.415 ;
        RECT 96.115 136.570 96.865 136.760 ;
        RECT 97.035 136.195 97.375 137.005 ;
        RECT 98.210 136.795 98.540 137.595 ;
        RECT 98.710 136.965 99.040 137.765 ;
        RECT 99.340 136.795 99.670 137.595 ;
        RECT 100.315 136.965 100.565 137.765 ;
        RECT 98.210 136.625 100.645 136.795 ;
        RECT 100.835 136.625 101.005 137.765 ;
        RECT 101.175 136.625 101.515 137.595 ;
        RECT 98.005 136.205 98.355 136.455 ;
        RECT 96.145 136.025 97.375 136.195 ;
        RECT 96.125 135.215 96.635 135.750 ;
        RECT 96.855 135.420 97.100 136.025 ;
        RECT 98.540 135.995 98.710 136.625 ;
        RECT 98.880 136.205 99.210 136.405 ;
        RECT 99.380 136.205 99.710 136.405 ;
        RECT 99.880 136.205 100.300 136.405 ;
        RECT 100.475 136.375 100.645 136.625 ;
        RECT 100.475 136.205 101.170 136.375 ;
        RECT 98.210 135.385 98.710 135.995 ;
        RECT 99.340 135.865 100.565 136.035 ;
        RECT 101.340 136.015 101.515 136.625 ;
        RECT 101.685 136.600 101.975 137.765 ;
        RECT 103.065 137.005 103.580 137.415 ;
        RECT 103.815 137.005 103.985 137.765 ;
        RECT 104.155 137.425 106.185 137.595 ;
        RECT 103.065 136.195 103.405 137.005 ;
        RECT 104.155 136.760 104.325 137.425 ;
        RECT 104.720 137.085 105.845 137.255 ;
        RECT 103.575 136.570 104.325 136.760 ;
        RECT 104.495 136.745 105.505 136.915 ;
        RECT 103.065 136.025 104.295 136.195 ;
        RECT 99.340 135.385 99.670 135.865 ;
        RECT 99.840 135.215 100.065 135.675 ;
        RECT 100.235 135.385 100.565 135.865 ;
        RECT 100.755 135.215 101.005 136.015 ;
        RECT 101.175 135.385 101.515 136.015 ;
        RECT 101.685 135.215 101.975 135.940 ;
        RECT 103.340 135.420 103.585 136.025 ;
        RECT 103.805 135.215 104.315 135.750 ;
        RECT 104.495 135.385 104.685 136.745 ;
        RECT 104.855 136.405 105.130 136.545 ;
        RECT 104.855 136.235 105.135 136.405 ;
        RECT 104.855 135.385 105.130 136.235 ;
        RECT 105.335 135.945 105.505 136.745 ;
        RECT 105.675 135.955 105.845 137.085 ;
        RECT 106.015 136.455 106.185 137.425 ;
        RECT 106.355 136.625 106.525 137.765 ;
        RECT 106.695 136.625 107.030 137.595 ;
        RECT 106.015 136.125 106.210 136.455 ;
        RECT 106.435 136.125 106.690 136.455 ;
        RECT 106.435 135.955 106.605 136.125 ;
        RECT 106.860 135.955 107.030 136.625 ;
        RECT 105.675 135.785 106.605 135.955 ;
        RECT 105.675 135.750 105.850 135.785 ;
        RECT 105.320 135.385 105.850 135.750 ;
        RECT 106.275 135.215 106.605 135.615 ;
        RECT 106.775 135.385 107.030 135.955 ;
        RECT 107.205 136.690 107.475 137.595 ;
        RECT 107.645 137.005 107.975 137.765 ;
        RECT 108.155 136.835 108.325 137.595 ;
        RECT 107.205 135.890 107.375 136.690 ;
        RECT 107.660 136.665 108.325 136.835 ;
        RECT 109.505 137.005 110.020 137.415 ;
        RECT 110.255 137.005 110.425 137.765 ;
        RECT 110.595 137.425 112.625 137.595 ;
        RECT 107.660 136.520 107.830 136.665 ;
        RECT 107.545 136.190 107.830 136.520 ;
        RECT 107.660 135.935 107.830 136.190 ;
        RECT 108.065 136.115 108.395 136.485 ;
        RECT 109.505 136.195 109.845 137.005 ;
        RECT 110.595 136.760 110.765 137.425 ;
        RECT 111.160 137.085 112.285 137.255 ;
        RECT 110.015 136.570 110.765 136.760 ;
        RECT 110.935 136.745 111.945 136.915 ;
        RECT 109.505 136.025 110.735 136.195 ;
        RECT 107.205 135.385 107.465 135.890 ;
        RECT 107.660 135.765 108.325 135.935 ;
        RECT 107.645 135.215 107.975 135.595 ;
        RECT 108.155 135.385 108.325 135.765 ;
        RECT 109.780 135.420 110.025 136.025 ;
        RECT 110.245 135.215 110.755 135.750 ;
        RECT 110.935 135.385 111.125 136.745 ;
        RECT 111.295 136.405 111.570 136.545 ;
        RECT 111.295 136.235 111.575 136.405 ;
        RECT 111.295 135.385 111.570 136.235 ;
        RECT 111.775 135.945 111.945 136.745 ;
        RECT 112.115 135.955 112.285 137.085 ;
        RECT 112.455 136.455 112.625 137.425 ;
        RECT 112.795 136.625 112.965 137.765 ;
        RECT 113.135 136.625 113.470 137.595 ;
        RECT 112.455 136.125 112.650 136.455 ;
        RECT 112.875 136.125 113.130 136.455 ;
        RECT 112.875 135.955 113.045 136.125 ;
        RECT 113.300 135.955 113.470 136.625 ;
        RECT 114.020 136.785 114.275 137.455 ;
        RECT 114.455 136.965 114.740 137.765 ;
        RECT 114.920 137.045 115.250 137.555 ;
        RECT 114.020 136.065 114.200 136.785 ;
        RECT 114.920 136.455 115.170 137.045 ;
        RECT 115.520 136.895 115.690 137.505 ;
        RECT 115.860 137.075 116.190 137.765 ;
        RECT 116.420 137.215 116.660 137.505 ;
        RECT 116.860 137.385 117.280 137.765 ;
        RECT 117.460 137.295 118.090 137.545 ;
        RECT 118.560 137.385 118.890 137.765 ;
        RECT 117.460 137.215 117.630 137.295 ;
        RECT 119.060 137.215 119.230 137.505 ;
        RECT 119.410 137.385 119.790 137.765 ;
        RECT 120.030 137.380 120.860 137.550 ;
        RECT 116.420 137.045 117.630 137.215 ;
        RECT 114.370 136.125 115.170 136.455 ;
        RECT 112.115 135.785 113.045 135.955 ;
        RECT 112.115 135.750 112.290 135.785 ;
        RECT 111.760 135.385 112.290 135.750 ;
        RECT 112.715 135.215 113.045 135.615 ;
        RECT 113.215 135.385 113.470 135.955 ;
        RECT 113.935 135.925 114.200 136.065 ;
        RECT 113.935 135.895 114.275 135.925 ;
        RECT 114.020 135.395 114.275 135.895 ;
        RECT 114.455 135.215 114.740 135.675 ;
        RECT 114.920 135.475 115.170 136.125 ;
        RECT 115.370 136.875 115.690 136.895 ;
        RECT 115.370 136.705 117.290 136.875 ;
        RECT 115.370 135.810 115.560 136.705 ;
        RECT 117.460 136.535 117.630 137.045 ;
        RECT 117.800 136.785 118.320 137.095 ;
        RECT 115.730 136.365 117.630 136.535 ;
        RECT 115.730 136.305 116.060 136.365 ;
        RECT 116.210 136.135 116.540 136.195 ;
        RECT 115.880 135.865 116.540 136.135 ;
        RECT 115.370 135.480 115.690 135.810 ;
        RECT 115.870 135.215 116.530 135.695 ;
        RECT 116.730 135.605 116.900 136.365 ;
        RECT 117.800 136.195 117.980 136.605 ;
        RECT 117.070 136.025 117.400 136.145 ;
        RECT 118.150 136.025 118.320 136.785 ;
        RECT 117.070 135.855 118.320 136.025 ;
        RECT 118.490 136.965 119.860 137.215 ;
        RECT 118.490 136.195 118.680 136.965 ;
        RECT 119.610 136.705 119.860 136.965 ;
        RECT 118.850 136.535 119.100 136.695 ;
        RECT 120.030 136.535 120.200 137.380 ;
        RECT 121.095 137.095 121.265 137.595 ;
        RECT 121.435 137.265 121.765 137.765 ;
        RECT 120.370 136.705 120.870 137.085 ;
        RECT 121.095 136.925 121.790 137.095 ;
        RECT 118.850 136.365 120.200 136.535 ;
        RECT 119.780 136.325 120.200 136.365 ;
        RECT 118.490 135.855 118.910 136.195 ;
        RECT 119.200 135.865 119.610 136.195 ;
        RECT 116.730 135.435 117.580 135.605 ;
        RECT 118.140 135.215 118.460 135.675 ;
        RECT 118.660 135.425 118.910 135.855 ;
        RECT 119.200 135.215 119.610 135.655 ;
        RECT 119.780 135.595 119.950 136.325 ;
        RECT 120.120 135.775 120.470 136.145 ;
        RECT 120.650 135.835 120.870 136.705 ;
        RECT 121.040 136.135 121.450 136.755 ;
        RECT 121.620 135.955 121.790 136.925 ;
        RECT 121.095 135.765 121.790 135.955 ;
        RECT 119.780 135.395 120.795 135.595 ;
        RECT 121.095 135.435 121.265 135.765 ;
        RECT 121.435 135.215 121.765 135.595 ;
        RECT 121.980 135.475 122.205 137.595 ;
        RECT 122.375 137.265 122.705 137.765 ;
        RECT 122.875 137.095 123.045 137.595 ;
        RECT 122.380 136.925 123.045 137.095 ;
        RECT 122.380 135.935 122.610 136.925 ;
        RECT 123.395 136.835 123.565 137.595 ;
        RECT 123.745 137.005 124.075 137.765 ;
        RECT 122.780 136.105 123.130 136.755 ;
        RECT 123.395 136.665 124.060 136.835 ;
        RECT 124.245 136.690 124.515 137.595 ;
        RECT 123.890 136.520 124.060 136.665 ;
        RECT 123.325 136.115 123.655 136.485 ;
        RECT 123.890 136.190 124.175 136.520 ;
        RECT 123.890 135.935 124.060 136.190 ;
        RECT 122.380 135.765 123.045 135.935 ;
        RECT 122.375 135.215 122.705 135.595 ;
        RECT 122.875 135.475 123.045 135.765 ;
        RECT 123.395 135.765 124.060 135.935 ;
        RECT 124.345 135.890 124.515 136.690 ;
        RECT 124.685 136.675 126.355 137.765 ;
        RECT 126.525 136.675 127.735 137.765 ;
        RECT 124.685 136.155 125.435 136.675 ;
        RECT 125.605 135.985 126.355 136.505 ;
        RECT 126.525 136.135 127.045 136.675 ;
        RECT 123.395 135.385 123.565 135.765 ;
        RECT 123.745 135.215 124.075 135.595 ;
        RECT 124.255 135.385 124.515 135.890 ;
        RECT 124.685 135.215 126.355 135.985 ;
        RECT 127.215 135.965 127.735 136.505 ;
        RECT 126.525 135.215 127.735 135.965 ;
        RECT 14.660 135.045 127.820 135.215 ;
        RECT 14.745 134.295 15.955 135.045 ;
        RECT 14.745 133.755 15.265 134.295 ;
        RECT 16.645 134.225 16.855 135.045 ;
        RECT 17.025 134.245 17.355 134.875 ;
        RECT 15.435 133.585 15.955 134.125 ;
        RECT 17.025 133.645 17.275 134.245 ;
        RECT 17.525 134.225 17.755 135.045 ;
        RECT 18.055 134.495 18.225 134.875 ;
        RECT 18.405 134.665 18.735 135.045 ;
        RECT 18.055 134.325 18.720 134.495 ;
        RECT 18.915 134.370 19.175 134.875 ;
        RECT 17.445 133.805 17.775 134.055 ;
        RECT 17.985 133.775 18.315 134.145 ;
        RECT 18.550 134.070 18.720 134.325 ;
        RECT 18.550 133.740 18.835 134.070 ;
        RECT 14.745 132.495 15.955 133.585 ;
        RECT 16.645 132.495 16.855 133.635 ;
        RECT 17.025 132.665 17.355 133.645 ;
        RECT 17.525 132.495 17.755 133.635 ;
        RECT 18.550 133.595 18.720 133.740 ;
        RECT 18.055 133.425 18.720 133.595 ;
        RECT 19.005 133.570 19.175 134.370 ;
        RECT 19.385 134.225 19.615 135.045 ;
        RECT 19.785 134.245 20.115 134.875 ;
        RECT 19.365 133.805 19.695 134.055 ;
        RECT 19.865 133.645 20.115 134.245 ;
        RECT 20.285 134.225 20.495 135.045 ;
        RECT 21.100 134.705 21.355 134.865 ;
        RECT 21.015 134.535 21.355 134.705 ;
        RECT 21.535 134.585 21.820 135.045 ;
        RECT 21.100 134.335 21.355 134.535 ;
        RECT 18.055 132.665 18.225 133.425 ;
        RECT 18.405 132.495 18.735 133.255 ;
        RECT 18.905 132.665 19.175 133.570 ;
        RECT 19.385 132.495 19.615 133.635 ;
        RECT 19.785 132.665 20.115 133.645 ;
        RECT 20.285 132.495 20.495 133.635 ;
        RECT 21.100 133.475 21.280 134.335 ;
        RECT 22.000 134.135 22.250 134.785 ;
        RECT 21.450 133.805 22.250 134.135 ;
        RECT 21.100 132.805 21.355 133.475 ;
        RECT 21.535 132.495 21.820 133.295 ;
        RECT 22.000 133.215 22.250 133.805 ;
        RECT 22.450 134.450 22.770 134.780 ;
        RECT 22.950 134.565 23.610 135.045 ;
        RECT 23.810 134.655 24.660 134.825 ;
        RECT 22.450 133.555 22.640 134.450 ;
        RECT 22.960 134.125 23.620 134.395 ;
        RECT 23.290 134.065 23.620 134.125 ;
        RECT 22.810 133.895 23.140 133.955 ;
        RECT 23.810 133.895 23.980 134.655 ;
        RECT 25.220 134.585 25.540 135.045 ;
        RECT 25.740 134.405 25.990 134.835 ;
        RECT 26.280 134.605 26.690 135.045 ;
        RECT 26.860 134.665 27.875 134.865 ;
        RECT 24.150 134.235 25.400 134.405 ;
        RECT 24.150 134.115 24.480 134.235 ;
        RECT 22.810 133.725 24.710 133.895 ;
        RECT 22.450 133.385 24.370 133.555 ;
        RECT 22.450 133.365 22.770 133.385 ;
        RECT 22.000 132.705 22.330 133.215 ;
        RECT 22.600 132.755 22.770 133.365 ;
        RECT 24.540 133.215 24.710 133.725 ;
        RECT 24.880 133.655 25.060 134.065 ;
        RECT 25.230 133.475 25.400 134.235 ;
        RECT 22.940 132.495 23.270 133.185 ;
        RECT 23.500 133.045 24.710 133.215 ;
        RECT 24.880 133.165 25.400 133.475 ;
        RECT 25.570 134.065 25.990 134.405 ;
        RECT 26.280 134.065 26.690 134.395 ;
        RECT 25.570 133.295 25.760 134.065 ;
        RECT 26.860 133.935 27.030 134.665 ;
        RECT 28.175 134.495 28.345 134.825 ;
        RECT 28.515 134.665 28.845 135.045 ;
        RECT 27.200 134.115 27.550 134.485 ;
        RECT 26.860 133.895 27.280 133.935 ;
        RECT 25.930 133.725 27.280 133.895 ;
        RECT 25.930 133.565 26.180 133.725 ;
        RECT 26.690 133.295 26.940 133.555 ;
        RECT 25.570 133.045 26.940 133.295 ;
        RECT 23.500 132.755 23.740 133.045 ;
        RECT 24.540 132.965 24.710 133.045 ;
        RECT 23.940 132.495 24.360 132.875 ;
        RECT 24.540 132.715 25.170 132.965 ;
        RECT 25.640 132.495 25.970 132.875 ;
        RECT 26.140 132.755 26.310 133.045 ;
        RECT 27.110 132.880 27.280 133.725 ;
        RECT 27.730 133.555 27.950 134.425 ;
        RECT 28.175 134.305 28.870 134.495 ;
        RECT 27.450 133.175 27.950 133.555 ;
        RECT 28.120 133.505 28.530 134.125 ;
        RECT 28.700 133.335 28.870 134.305 ;
        RECT 28.175 133.165 28.870 133.335 ;
        RECT 26.490 132.495 26.870 132.875 ;
        RECT 27.110 132.710 27.940 132.880 ;
        RECT 28.175 132.665 28.345 133.165 ;
        RECT 28.515 132.495 28.845 132.995 ;
        RECT 29.060 132.665 29.285 134.785 ;
        RECT 29.455 134.665 29.785 135.045 ;
        RECT 29.955 134.495 30.125 134.785 ;
        RECT 29.460 134.325 30.125 134.495 ;
        RECT 31.045 134.415 31.375 134.775 ;
        RECT 31.995 134.585 32.245 135.045 ;
        RECT 32.415 134.585 32.975 134.875 ;
        RECT 29.460 133.335 29.690 134.325 ;
        RECT 31.045 134.225 32.435 134.415 ;
        RECT 29.860 133.505 30.210 134.155 ;
        RECT 32.265 134.135 32.435 134.225 ;
        RECT 30.860 133.805 31.535 134.055 ;
        RECT 31.755 133.805 32.095 134.055 ;
        RECT 32.265 133.805 32.555 134.135 ;
        RECT 30.860 133.445 31.125 133.805 ;
        RECT 32.265 133.555 32.435 133.805 ;
        RECT 31.495 133.385 32.435 133.555 ;
        RECT 29.460 133.165 30.125 133.335 ;
        RECT 29.455 132.495 29.785 132.995 ;
        RECT 29.955 132.665 30.125 133.165 ;
        RECT 31.045 132.495 31.325 133.165 ;
        RECT 31.495 132.835 31.795 133.385 ;
        RECT 32.725 133.215 32.975 134.585 ;
        RECT 33.420 134.235 33.665 134.840 ;
        RECT 33.885 134.510 34.395 135.045 ;
        RECT 31.995 132.495 32.325 133.215 ;
        RECT 32.515 132.665 32.975 133.215 ;
        RECT 33.145 134.065 34.375 134.235 ;
        RECT 33.145 133.255 33.485 134.065 ;
        RECT 33.655 133.500 34.405 133.690 ;
        RECT 33.145 132.845 33.660 133.255 ;
        RECT 33.895 132.495 34.065 133.255 ;
        RECT 34.235 132.835 34.405 133.500 ;
        RECT 34.575 133.515 34.765 134.875 ;
        RECT 34.935 134.025 35.210 134.875 ;
        RECT 35.400 134.510 35.930 134.875 ;
        RECT 36.355 134.645 36.685 135.045 ;
        RECT 35.755 134.475 35.930 134.510 ;
        RECT 34.935 133.855 35.215 134.025 ;
        RECT 34.935 133.715 35.210 133.855 ;
        RECT 35.415 133.515 35.585 134.315 ;
        RECT 34.575 133.345 35.585 133.515 ;
        RECT 35.755 134.305 36.685 134.475 ;
        RECT 36.855 134.305 37.110 134.875 ;
        RECT 37.285 134.320 37.575 135.045 ;
        RECT 35.755 133.175 35.925 134.305 ;
        RECT 36.515 134.135 36.685 134.305 ;
        RECT 34.800 133.005 35.925 133.175 ;
        RECT 36.095 133.805 36.290 134.135 ;
        RECT 36.515 133.805 36.770 134.135 ;
        RECT 36.095 132.835 36.265 133.805 ;
        RECT 36.940 133.635 37.110 134.305 ;
        RECT 37.745 134.275 39.415 135.045 ;
        RECT 39.595 134.545 39.925 135.045 ;
        RECT 40.125 134.475 40.295 134.825 ;
        RECT 40.495 134.645 40.825 135.045 ;
        RECT 40.995 134.475 41.165 134.825 ;
        RECT 41.335 134.645 41.715 135.045 ;
        RECT 34.235 132.665 36.265 132.835 ;
        RECT 36.435 132.495 36.605 133.635 ;
        RECT 36.775 132.665 37.110 133.635 ;
        RECT 37.285 132.495 37.575 133.660 ;
        RECT 37.745 133.585 38.495 134.105 ;
        RECT 38.665 133.755 39.415 134.275 ;
        RECT 39.590 133.805 39.940 134.375 ;
        RECT 40.125 134.305 41.735 134.475 ;
        RECT 41.905 134.370 42.175 134.715 ;
        RECT 42.355 134.545 42.685 135.045 ;
        RECT 42.885 134.475 43.055 134.825 ;
        RECT 43.255 134.645 43.585 135.045 ;
        RECT 43.755 134.475 43.925 134.825 ;
        RECT 44.095 134.645 44.475 135.045 ;
        RECT 41.565 134.135 41.735 134.305 ;
        RECT 37.745 132.495 39.415 133.585 ;
        RECT 39.590 133.345 39.910 133.635 ;
        RECT 40.110 133.515 40.820 134.135 ;
        RECT 40.990 133.805 41.395 134.135 ;
        RECT 41.565 133.805 41.835 134.135 ;
        RECT 41.565 133.635 41.735 133.805 ;
        RECT 42.005 133.635 42.175 134.370 ;
        RECT 42.350 133.805 42.700 134.375 ;
        RECT 42.885 134.305 44.495 134.475 ;
        RECT 44.665 134.370 44.935 134.715 ;
        RECT 44.325 134.135 44.495 134.305 ;
        RECT 41.010 133.465 41.735 133.635 ;
        RECT 41.010 133.345 41.180 133.465 ;
        RECT 39.590 133.175 41.180 133.345 ;
        RECT 39.590 132.715 41.245 133.005 ;
        RECT 41.415 132.495 41.695 133.295 ;
        RECT 41.905 132.665 42.175 133.635 ;
        RECT 42.350 133.345 42.670 133.635 ;
        RECT 42.870 133.515 43.580 134.135 ;
        RECT 43.750 133.805 44.155 134.135 ;
        RECT 44.325 133.805 44.595 134.135 ;
        RECT 44.325 133.635 44.495 133.805 ;
        RECT 44.765 133.635 44.935 134.370 ;
        RECT 43.770 133.465 44.495 133.635 ;
        RECT 43.770 133.345 43.940 133.465 ;
        RECT 42.350 133.175 43.940 133.345 ;
        RECT 42.350 132.715 44.005 133.005 ;
        RECT 44.175 132.495 44.455 133.295 ;
        RECT 44.665 132.665 44.935 133.635 ;
        RECT 45.105 134.245 45.445 134.875 ;
        RECT 45.615 134.245 45.865 135.045 ;
        RECT 46.055 134.395 46.385 134.875 ;
        RECT 46.555 134.585 46.780 135.045 ;
        RECT 46.950 134.395 47.280 134.875 ;
        RECT 45.105 133.685 45.280 134.245 ;
        RECT 46.055 134.225 47.280 134.395 ;
        RECT 47.910 134.265 48.410 134.875 ;
        RECT 45.450 133.885 46.145 134.055 ;
        RECT 45.105 133.635 45.335 133.685 ;
        RECT 45.975 133.635 46.145 133.885 ;
        RECT 46.320 133.855 46.740 134.055 ;
        RECT 46.910 133.855 47.240 134.055 ;
        RECT 47.410 133.855 47.740 134.055 ;
        RECT 47.910 133.635 48.080 134.265 ;
        RECT 48.785 134.245 49.125 134.875 ;
        RECT 49.295 134.245 49.545 135.045 ;
        RECT 49.735 134.395 50.065 134.875 ;
        RECT 50.235 134.585 50.460 135.045 ;
        RECT 50.630 134.395 50.960 134.875 ;
        RECT 48.785 134.195 49.015 134.245 ;
        RECT 49.735 134.225 50.960 134.395 ;
        RECT 51.590 134.265 52.090 134.875 ;
        RECT 52.840 134.705 53.095 134.865 ;
        RECT 52.755 134.535 53.095 134.705 ;
        RECT 53.275 134.585 53.560 135.045 ;
        RECT 52.840 134.335 53.095 134.535 ;
        RECT 48.265 133.805 48.615 134.055 ;
        RECT 48.785 133.635 48.960 134.195 ;
        RECT 49.130 133.885 49.825 134.055 ;
        RECT 49.655 133.635 49.825 133.885 ;
        RECT 50.000 133.855 50.420 134.055 ;
        RECT 50.590 133.855 50.920 134.055 ;
        RECT 51.090 133.855 51.420 134.055 ;
        RECT 51.590 133.635 51.760 134.265 ;
        RECT 51.945 133.805 52.295 134.055 ;
        RECT 45.105 132.665 45.445 133.635 ;
        RECT 45.615 132.495 45.785 133.635 ;
        RECT 45.975 133.465 48.410 133.635 ;
        RECT 46.055 132.495 46.305 133.295 ;
        RECT 46.950 132.665 47.280 133.465 ;
        RECT 47.580 132.495 47.910 133.295 ;
        RECT 48.080 132.665 48.410 133.465 ;
        RECT 48.785 132.665 49.125 133.635 ;
        RECT 49.295 132.495 49.465 133.635 ;
        RECT 49.655 133.465 52.090 133.635 ;
        RECT 49.735 132.495 49.985 133.295 ;
        RECT 50.630 132.665 50.960 133.465 ;
        RECT 51.260 132.495 51.590 133.295 ;
        RECT 51.760 132.665 52.090 133.465 ;
        RECT 52.840 133.475 53.020 134.335 ;
        RECT 53.740 134.135 53.990 134.785 ;
        RECT 53.190 133.805 53.990 134.135 ;
        RECT 52.840 132.805 53.095 133.475 ;
        RECT 53.275 132.495 53.560 133.295 ;
        RECT 53.740 133.215 53.990 133.805 ;
        RECT 54.190 134.450 54.510 134.780 ;
        RECT 54.690 134.565 55.350 135.045 ;
        RECT 55.550 134.655 56.400 134.825 ;
        RECT 54.190 133.555 54.380 134.450 ;
        RECT 54.700 134.125 55.360 134.395 ;
        RECT 55.030 134.065 55.360 134.125 ;
        RECT 54.550 133.895 54.880 133.955 ;
        RECT 55.550 133.895 55.720 134.655 ;
        RECT 56.960 134.585 57.280 135.045 ;
        RECT 57.480 134.405 57.730 134.835 ;
        RECT 58.020 134.605 58.430 135.045 ;
        RECT 58.600 134.665 59.615 134.865 ;
        RECT 55.890 134.235 57.140 134.405 ;
        RECT 55.890 134.115 56.220 134.235 ;
        RECT 54.550 133.725 56.450 133.895 ;
        RECT 54.190 133.385 56.110 133.555 ;
        RECT 54.190 133.365 54.510 133.385 ;
        RECT 53.740 132.705 54.070 133.215 ;
        RECT 54.340 132.755 54.510 133.365 ;
        RECT 56.280 133.215 56.450 133.725 ;
        RECT 56.620 133.655 56.800 134.065 ;
        RECT 56.970 133.475 57.140 134.235 ;
        RECT 54.680 132.495 55.010 133.185 ;
        RECT 55.240 133.045 56.450 133.215 ;
        RECT 56.620 133.165 57.140 133.475 ;
        RECT 57.310 134.065 57.730 134.405 ;
        RECT 58.020 134.065 58.430 134.395 ;
        RECT 57.310 133.295 57.500 134.065 ;
        RECT 58.600 133.935 58.770 134.665 ;
        RECT 59.915 134.495 60.085 134.825 ;
        RECT 60.255 134.665 60.585 135.045 ;
        RECT 58.940 134.115 59.290 134.485 ;
        RECT 58.600 133.895 59.020 133.935 ;
        RECT 57.670 133.725 59.020 133.895 ;
        RECT 57.670 133.565 57.920 133.725 ;
        RECT 58.430 133.295 58.680 133.555 ;
        RECT 57.310 133.045 58.680 133.295 ;
        RECT 55.240 132.755 55.480 133.045 ;
        RECT 56.280 132.965 56.450 133.045 ;
        RECT 55.680 132.495 56.100 132.875 ;
        RECT 56.280 132.715 56.910 132.965 ;
        RECT 57.380 132.495 57.710 132.875 ;
        RECT 57.880 132.755 58.050 133.045 ;
        RECT 58.850 132.880 59.020 133.725 ;
        RECT 59.470 133.555 59.690 134.425 ;
        RECT 59.915 134.305 60.610 134.495 ;
        RECT 59.190 133.175 59.690 133.555 ;
        RECT 59.860 133.505 60.270 134.125 ;
        RECT 60.440 133.335 60.610 134.305 ;
        RECT 59.915 133.165 60.610 133.335 ;
        RECT 58.230 132.495 58.610 132.875 ;
        RECT 58.850 132.710 59.680 132.880 ;
        RECT 59.915 132.665 60.085 133.165 ;
        RECT 60.255 132.495 60.585 132.995 ;
        RECT 60.800 132.665 61.025 134.785 ;
        RECT 61.195 134.665 61.525 135.045 ;
        RECT 61.695 134.495 61.865 134.785 ;
        RECT 61.200 134.325 61.865 134.495 ;
        RECT 61.200 133.335 61.430 134.325 ;
        RECT 63.045 134.320 63.335 135.045 ;
        RECT 63.505 134.245 63.845 134.875 ;
        RECT 64.015 134.245 64.265 135.045 ;
        RECT 64.455 134.395 64.785 134.875 ;
        RECT 64.955 134.585 65.180 135.045 ;
        RECT 65.350 134.395 65.680 134.875 ;
        RECT 61.600 133.505 61.950 134.155 ;
        RECT 63.505 133.685 63.680 134.245 ;
        RECT 64.455 134.225 65.680 134.395 ;
        RECT 66.310 134.265 66.810 134.875 ;
        RECT 68.110 134.500 73.455 135.045 ;
        RECT 73.630 134.500 78.975 135.045 ;
        RECT 79.155 134.545 79.485 135.045 ;
        RECT 63.850 133.885 64.545 134.055 ;
        RECT 61.200 133.165 61.865 133.335 ;
        RECT 61.195 132.495 61.525 132.995 ;
        RECT 61.695 132.665 61.865 133.165 ;
        RECT 63.045 132.495 63.335 133.660 ;
        RECT 63.505 133.635 63.735 133.685 ;
        RECT 64.375 133.635 64.545 133.885 ;
        RECT 64.720 133.855 65.140 134.055 ;
        RECT 65.310 133.855 65.640 134.055 ;
        RECT 65.810 133.855 66.140 134.055 ;
        RECT 66.310 133.635 66.480 134.265 ;
        RECT 66.665 133.805 67.015 134.055 ;
        RECT 63.505 132.665 63.845 133.635 ;
        RECT 64.015 132.495 64.185 133.635 ;
        RECT 64.375 133.465 66.810 133.635 ;
        RECT 64.455 132.495 64.705 133.295 ;
        RECT 65.350 132.665 65.680 133.465 ;
        RECT 65.980 132.495 66.310 133.295 ;
        RECT 66.480 132.665 66.810 133.465 ;
        RECT 69.700 132.930 70.050 134.180 ;
        RECT 71.530 133.670 71.870 134.500 ;
        RECT 75.220 132.930 75.570 134.180 ;
        RECT 77.050 133.670 77.390 134.500 ;
        RECT 79.685 134.475 79.855 134.825 ;
        RECT 80.055 134.645 80.385 135.045 ;
        RECT 80.555 134.475 80.725 134.825 ;
        RECT 80.895 134.645 81.275 135.045 ;
        RECT 79.150 133.805 79.500 134.375 ;
        RECT 79.685 134.305 81.295 134.475 ;
        RECT 81.465 134.370 81.735 134.715 ;
        RECT 81.910 134.500 87.255 135.045 ;
        RECT 81.125 134.135 81.295 134.305 ;
        RECT 79.150 133.345 79.470 133.635 ;
        RECT 79.670 133.515 80.380 134.135 ;
        RECT 80.550 133.805 80.955 134.135 ;
        RECT 81.125 133.805 81.395 134.135 ;
        RECT 81.125 133.635 81.295 133.805 ;
        RECT 81.565 133.635 81.735 134.370 ;
        RECT 80.570 133.465 81.295 133.635 ;
        RECT 80.570 133.345 80.740 133.465 ;
        RECT 79.150 133.175 80.740 133.345 ;
        RECT 68.110 132.495 73.455 132.930 ;
        RECT 73.630 132.495 78.975 132.930 ;
        RECT 79.150 132.715 80.805 133.005 ;
        RECT 80.975 132.495 81.255 133.295 ;
        RECT 81.465 132.665 81.735 133.635 ;
        RECT 83.500 132.930 83.850 134.180 ;
        RECT 85.330 133.670 85.670 134.500 ;
        RECT 87.485 134.225 87.695 135.045 ;
        RECT 87.865 134.245 88.195 134.875 ;
        RECT 87.865 133.645 88.115 134.245 ;
        RECT 88.365 134.225 88.595 135.045 ;
        RECT 88.805 134.320 89.095 135.045 ;
        RECT 89.640 134.335 89.895 134.865 ;
        RECT 90.075 134.585 90.360 135.045 ;
        RECT 88.285 133.805 88.615 134.055 ;
        RECT 89.640 133.685 89.820 134.335 ;
        RECT 90.540 134.135 90.790 134.785 ;
        RECT 89.990 133.805 90.790 134.135 ;
        RECT 81.910 132.495 87.255 132.930 ;
        RECT 87.485 132.495 87.695 133.635 ;
        RECT 87.865 132.665 88.195 133.645 ;
        RECT 88.365 132.495 88.595 133.635 ;
        RECT 88.805 132.495 89.095 133.660 ;
        RECT 89.555 133.515 89.820 133.685 ;
        RECT 89.640 133.475 89.820 133.515 ;
        RECT 89.640 132.805 89.895 133.475 ;
        RECT 90.075 132.495 90.360 133.295 ;
        RECT 90.540 133.215 90.790 133.805 ;
        RECT 90.990 134.450 91.310 134.780 ;
        RECT 91.490 134.565 92.150 135.045 ;
        RECT 92.350 134.655 93.200 134.825 ;
        RECT 90.990 133.555 91.180 134.450 ;
        RECT 91.500 134.125 92.160 134.395 ;
        RECT 91.830 134.065 92.160 134.125 ;
        RECT 91.350 133.895 91.680 133.955 ;
        RECT 92.350 133.895 92.520 134.655 ;
        RECT 93.760 134.585 94.080 135.045 ;
        RECT 94.280 134.405 94.530 134.835 ;
        RECT 94.820 134.605 95.230 135.045 ;
        RECT 95.400 134.665 96.415 134.865 ;
        RECT 92.690 134.235 93.940 134.405 ;
        RECT 92.690 134.115 93.020 134.235 ;
        RECT 91.350 133.725 93.250 133.895 ;
        RECT 90.990 133.385 92.910 133.555 ;
        RECT 90.990 133.365 91.310 133.385 ;
        RECT 90.540 132.705 90.870 133.215 ;
        RECT 91.140 132.755 91.310 133.365 ;
        RECT 93.080 133.215 93.250 133.725 ;
        RECT 93.420 133.655 93.600 134.065 ;
        RECT 93.770 133.475 93.940 134.235 ;
        RECT 91.480 132.495 91.810 133.185 ;
        RECT 92.040 133.045 93.250 133.215 ;
        RECT 93.420 133.165 93.940 133.475 ;
        RECT 94.110 134.065 94.530 134.405 ;
        RECT 94.820 134.065 95.230 134.395 ;
        RECT 94.110 133.295 94.300 134.065 ;
        RECT 95.400 133.935 95.570 134.665 ;
        RECT 96.715 134.495 96.885 134.825 ;
        RECT 97.055 134.665 97.385 135.045 ;
        RECT 95.740 134.115 96.090 134.485 ;
        RECT 95.400 133.895 95.820 133.935 ;
        RECT 94.470 133.725 95.820 133.895 ;
        RECT 94.470 133.565 94.720 133.725 ;
        RECT 95.230 133.295 95.480 133.555 ;
        RECT 94.110 133.045 95.480 133.295 ;
        RECT 92.040 132.755 92.280 133.045 ;
        RECT 93.080 132.965 93.250 133.045 ;
        RECT 92.480 132.495 92.900 132.875 ;
        RECT 93.080 132.715 93.710 132.965 ;
        RECT 94.180 132.495 94.510 132.875 ;
        RECT 94.680 132.755 94.850 133.045 ;
        RECT 95.650 132.880 95.820 133.725 ;
        RECT 96.270 133.555 96.490 134.425 ;
        RECT 96.715 134.305 97.410 134.495 ;
        RECT 95.990 133.175 96.490 133.555 ;
        RECT 96.660 133.505 97.070 134.125 ;
        RECT 97.240 133.335 97.410 134.305 ;
        RECT 96.715 133.165 97.410 133.335 ;
        RECT 95.030 132.495 95.410 132.875 ;
        RECT 95.650 132.710 96.480 132.880 ;
        RECT 96.715 132.665 96.885 133.165 ;
        RECT 97.055 132.495 97.385 132.995 ;
        RECT 97.600 132.665 97.825 134.785 ;
        RECT 97.995 134.665 98.325 135.045 ;
        RECT 98.495 134.495 98.665 134.785 ;
        RECT 98.000 134.325 98.665 134.495 ;
        RECT 98.925 134.370 99.195 134.715 ;
        RECT 99.385 134.645 99.765 135.045 ;
        RECT 99.935 134.475 100.105 134.825 ;
        RECT 100.275 134.645 100.605 135.045 ;
        RECT 100.805 134.475 100.975 134.825 ;
        RECT 101.175 134.545 101.505 135.045 ;
        RECT 98.000 133.335 98.230 134.325 ;
        RECT 98.400 133.505 98.750 134.155 ;
        RECT 98.925 133.635 99.095 134.370 ;
        RECT 99.365 134.305 100.975 134.475 ;
        RECT 99.365 134.135 99.535 134.305 ;
        RECT 99.265 133.805 99.535 134.135 ;
        RECT 99.705 133.805 100.110 134.135 ;
        RECT 99.365 133.635 99.535 133.805 ;
        RECT 100.280 133.685 100.990 134.135 ;
        RECT 101.160 133.805 101.510 134.375 ;
        RECT 101.745 134.225 101.955 135.045 ;
        RECT 102.125 134.245 102.455 134.875 ;
        RECT 98.000 133.165 98.665 133.335 ;
        RECT 97.995 132.495 98.325 132.995 ;
        RECT 98.495 132.665 98.665 133.165 ;
        RECT 98.925 132.665 99.195 133.635 ;
        RECT 99.365 133.465 100.090 133.635 ;
        RECT 100.280 133.515 100.995 133.685 ;
        RECT 102.125 133.645 102.375 134.245 ;
        RECT 102.625 134.225 102.855 135.045 ;
        RECT 103.525 134.370 103.795 134.715 ;
        RECT 103.985 134.645 104.365 135.045 ;
        RECT 104.535 134.475 104.705 134.825 ;
        RECT 104.875 134.645 105.205 135.045 ;
        RECT 105.405 134.475 105.575 134.825 ;
        RECT 105.775 134.545 106.105 135.045 ;
        RECT 102.545 133.805 102.875 134.055 ;
        RECT 99.920 133.345 100.090 133.465 ;
        RECT 101.190 133.345 101.510 133.635 ;
        RECT 99.405 132.495 99.685 133.295 ;
        RECT 99.920 133.175 101.510 133.345 ;
        RECT 99.855 132.715 101.510 133.005 ;
        RECT 101.745 132.495 101.955 133.635 ;
        RECT 102.125 132.665 102.455 133.645 ;
        RECT 103.525 133.635 103.695 134.370 ;
        RECT 103.965 134.305 105.575 134.475 ;
        RECT 103.965 134.135 104.135 134.305 ;
        RECT 103.865 133.805 104.135 134.135 ;
        RECT 104.305 133.805 104.710 134.135 ;
        RECT 103.965 133.635 104.135 133.805 ;
        RECT 102.625 132.495 102.855 133.635 ;
        RECT 103.525 132.665 103.795 133.635 ;
        RECT 103.965 133.465 104.690 133.635 ;
        RECT 104.880 133.515 105.590 134.135 ;
        RECT 105.760 133.805 106.110 134.375 ;
        RECT 106.285 134.245 106.625 134.875 ;
        RECT 106.795 134.245 107.045 135.045 ;
        RECT 107.235 134.395 107.565 134.875 ;
        RECT 107.735 134.585 107.960 135.045 ;
        RECT 108.130 134.395 108.460 134.875 ;
        RECT 106.285 134.195 106.515 134.245 ;
        RECT 107.235 134.225 108.460 134.395 ;
        RECT 109.090 134.265 109.590 134.875 ;
        RECT 109.965 134.370 110.235 134.715 ;
        RECT 110.425 134.645 110.805 135.045 ;
        RECT 110.975 134.475 111.145 134.825 ;
        RECT 111.315 134.645 111.645 135.045 ;
        RECT 111.845 134.475 112.015 134.825 ;
        RECT 112.215 134.545 112.545 135.045 ;
        RECT 106.285 133.635 106.460 134.195 ;
        RECT 106.630 133.885 107.325 134.055 ;
        RECT 107.155 133.635 107.325 133.885 ;
        RECT 107.500 133.855 107.920 134.055 ;
        RECT 108.090 133.855 108.420 134.055 ;
        RECT 108.590 133.855 108.920 134.055 ;
        RECT 109.090 133.635 109.260 134.265 ;
        RECT 109.445 133.805 109.795 134.055 ;
        RECT 109.965 133.635 110.135 134.370 ;
        RECT 110.405 134.305 112.015 134.475 ;
        RECT 110.405 134.135 110.575 134.305 ;
        RECT 110.305 133.805 110.575 134.135 ;
        RECT 110.745 133.805 111.150 134.135 ;
        RECT 110.405 133.635 110.575 133.805 ;
        RECT 104.520 133.345 104.690 133.465 ;
        RECT 105.790 133.345 106.110 133.635 ;
        RECT 104.005 132.495 104.285 133.295 ;
        RECT 104.520 133.175 106.110 133.345 ;
        RECT 104.455 132.715 106.110 133.005 ;
        RECT 106.285 132.665 106.625 133.635 ;
        RECT 106.795 132.495 106.965 133.635 ;
        RECT 107.155 133.465 109.590 133.635 ;
        RECT 107.235 132.495 107.485 133.295 ;
        RECT 108.130 132.665 108.460 133.465 ;
        RECT 108.760 132.495 109.090 133.295 ;
        RECT 109.260 132.665 109.590 133.465 ;
        RECT 109.965 132.665 110.235 133.635 ;
        RECT 110.405 133.465 111.130 133.635 ;
        RECT 111.320 133.515 112.030 134.135 ;
        RECT 112.200 133.805 112.550 134.375 ;
        RECT 112.725 134.275 114.395 135.045 ;
        RECT 114.565 134.320 114.855 135.045 ;
        RECT 115.485 134.275 118.995 135.045 ;
        RECT 119.255 134.495 119.425 134.875 ;
        RECT 119.605 134.665 119.935 135.045 ;
        RECT 119.255 134.325 119.920 134.495 ;
        RECT 120.115 134.370 120.375 134.875 ;
        RECT 121.010 134.500 126.355 135.045 ;
        RECT 110.960 133.345 111.130 133.465 ;
        RECT 112.230 133.345 112.550 133.635 ;
        RECT 110.445 132.495 110.725 133.295 ;
        RECT 110.960 133.175 112.550 133.345 ;
        RECT 112.725 133.585 113.475 134.105 ;
        RECT 113.645 133.755 114.395 134.275 ;
        RECT 110.895 132.715 112.550 133.005 ;
        RECT 112.725 132.495 114.395 133.585 ;
        RECT 114.565 132.495 114.855 133.660 ;
        RECT 115.485 133.585 117.175 134.105 ;
        RECT 117.345 133.755 118.995 134.275 ;
        RECT 119.185 133.775 119.515 134.145 ;
        RECT 119.750 134.070 119.920 134.325 ;
        RECT 119.750 133.740 120.035 134.070 ;
        RECT 119.750 133.595 119.920 133.740 ;
        RECT 115.485 132.495 118.995 133.585 ;
        RECT 119.255 133.425 119.920 133.595 ;
        RECT 120.205 133.570 120.375 134.370 ;
        RECT 119.255 132.665 119.425 133.425 ;
        RECT 119.605 132.495 119.935 133.255 ;
        RECT 120.105 132.665 120.375 133.570 ;
        RECT 122.600 132.930 122.950 134.180 ;
        RECT 124.430 133.670 124.770 134.500 ;
        RECT 126.525 134.295 127.735 135.045 ;
        RECT 126.525 133.585 127.045 134.125 ;
        RECT 127.215 133.755 127.735 134.295 ;
        RECT 121.010 132.495 126.355 132.930 ;
        RECT 126.525 132.495 127.735 133.585 ;
        RECT 14.660 132.325 127.820 132.495 ;
        RECT 14.745 131.235 15.955 132.325 ;
        RECT 14.745 130.525 15.265 131.065 ;
        RECT 15.435 130.695 15.955 131.235 ;
        RECT 16.585 131.235 20.095 132.325 ;
        RECT 20.265 131.565 20.780 131.975 ;
        RECT 21.015 131.565 21.185 132.325 ;
        RECT 21.355 131.985 23.385 132.155 ;
        RECT 16.585 130.715 18.275 131.235 ;
        RECT 18.445 130.545 20.095 131.065 ;
        RECT 20.265 130.755 20.605 131.565 ;
        RECT 21.355 131.320 21.525 131.985 ;
        RECT 21.920 131.645 23.045 131.815 ;
        RECT 20.775 131.130 21.525 131.320 ;
        RECT 21.695 131.305 22.705 131.475 ;
        RECT 20.265 130.585 21.495 130.755 ;
        RECT 14.745 129.775 15.955 130.525 ;
        RECT 16.585 129.775 20.095 130.545 ;
        RECT 20.540 129.980 20.785 130.585 ;
        RECT 21.005 129.775 21.515 130.310 ;
        RECT 21.695 129.945 21.885 131.305 ;
        RECT 22.055 130.625 22.330 131.105 ;
        RECT 22.055 130.455 22.335 130.625 ;
        RECT 22.535 130.505 22.705 131.305 ;
        RECT 22.875 130.515 23.045 131.645 ;
        RECT 23.215 131.015 23.385 131.985 ;
        RECT 23.555 131.185 23.725 132.325 ;
        RECT 23.895 131.185 24.230 132.155 ;
        RECT 23.215 130.685 23.410 131.015 ;
        RECT 23.635 130.685 23.890 131.015 ;
        RECT 23.635 130.515 23.805 130.685 ;
        RECT 24.060 130.515 24.230 131.185 ;
        RECT 24.405 131.160 24.695 132.325 ;
        RECT 25.325 131.235 28.835 132.325 ;
        RECT 29.005 131.250 29.275 132.155 ;
        RECT 29.445 131.565 29.775 132.325 ;
        RECT 29.955 131.395 30.125 132.155 ;
        RECT 30.760 131.985 31.015 132.015 ;
        RECT 30.675 131.815 31.015 131.985 ;
        RECT 25.325 130.715 27.015 131.235 ;
        RECT 27.185 130.545 28.835 131.065 ;
        RECT 22.055 129.945 22.330 130.455 ;
        RECT 22.875 130.345 23.805 130.515 ;
        RECT 22.875 130.310 23.050 130.345 ;
        RECT 22.520 129.945 23.050 130.310 ;
        RECT 23.475 129.775 23.805 130.175 ;
        RECT 23.975 129.945 24.230 130.515 ;
        RECT 24.405 129.775 24.695 130.500 ;
        RECT 25.325 129.775 28.835 130.545 ;
        RECT 29.005 130.450 29.175 131.250 ;
        RECT 29.460 131.225 30.125 131.395 ;
        RECT 30.760 131.345 31.015 131.815 ;
        RECT 31.195 131.525 31.480 132.325 ;
        RECT 31.660 131.605 31.990 132.115 ;
        RECT 29.460 131.080 29.630 131.225 ;
        RECT 29.345 130.750 29.630 131.080 ;
        RECT 29.460 130.495 29.630 130.750 ;
        RECT 29.865 130.675 30.195 131.045 ;
        RECT 29.005 129.945 29.265 130.450 ;
        RECT 29.460 130.325 30.125 130.495 ;
        RECT 29.445 129.775 29.775 130.155 ;
        RECT 29.955 129.945 30.125 130.325 ;
        RECT 30.760 130.485 30.940 131.345 ;
        RECT 31.660 131.015 31.910 131.605 ;
        RECT 32.260 131.455 32.430 132.065 ;
        RECT 32.600 131.635 32.930 132.325 ;
        RECT 33.160 131.775 33.400 132.065 ;
        RECT 33.600 131.945 34.020 132.325 ;
        RECT 34.200 131.855 34.830 132.105 ;
        RECT 35.300 131.945 35.630 132.325 ;
        RECT 34.200 131.775 34.370 131.855 ;
        RECT 35.800 131.775 35.970 132.065 ;
        RECT 36.150 131.945 36.530 132.325 ;
        RECT 36.770 131.940 37.600 132.110 ;
        RECT 33.160 131.605 34.370 131.775 ;
        RECT 31.110 130.685 31.910 131.015 ;
        RECT 30.760 129.955 31.015 130.485 ;
        RECT 31.195 129.775 31.480 130.235 ;
        RECT 31.660 130.035 31.910 130.685 ;
        RECT 32.110 131.435 32.430 131.455 ;
        RECT 32.110 131.265 34.030 131.435 ;
        RECT 32.110 130.370 32.300 131.265 ;
        RECT 34.200 131.095 34.370 131.605 ;
        RECT 34.540 131.345 35.060 131.655 ;
        RECT 32.470 130.925 34.370 131.095 ;
        RECT 32.470 130.865 32.800 130.925 ;
        RECT 32.950 130.695 33.280 130.755 ;
        RECT 32.620 130.425 33.280 130.695 ;
        RECT 32.110 130.040 32.430 130.370 ;
        RECT 32.610 129.775 33.270 130.255 ;
        RECT 33.470 130.165 33.640 130.925 ;
        RECT 34.540 130.755 34.720 131.165 ;
        RECT 33.810 130.585 34.140 130.705 ;
        RECT 34.890 130.585 35.060 131.345 ;
        RECT 33.810 130.415 35.060 130.585 ;
        RECT 35.230 131.525 36.600 131.775 ;
        RECT 35.230 130.755 35.420 131.525 ;
        RECT 36.350 131.265 36.600 131.525 ;
        RECT 35.590 131.095 35.840 131.255 ;
        RECT 36.770 131.095 36.940 131.940 ;
        RECT 37.835 131.655 38.005 132.155 ;
        RECT 38.175 131.825 38.505 132.325 ;
        RECT 37.110 131.265 37.610 131.645 ;
        RECT 37.835 131.485 38.530 131.655 ;
        RECT 35.590 130.925 36.940 131.095 ;
        RECT 36.520 130.885 36.940 130.925 ;
        RECT 35.230 130.415 35.650 130.755 ;
        RECT 35.940 130.425 36.350 130.755 ;
        RECT 33.470 129.995 34.320 130.165 ;
        RECT 34.880 129.775 35.200 130.235 ;
        RECT 35.400 129.985 35.650 130.415 ;
        RECT 35.940 129.775 36.350 130.215 ;
        RECT 36.520 130.155 36.690 130.885 ;
        RECT 36.860 130.335 37.210 130.705 ;
        RECT 37.390 130.395 37.610 131.265 ;
        RECT 37.780 130.695 38.190 131.315 ;
        RECT 38.360 130.515 38.530 131.485 ;
        RECT 37.835 130.325 38.530 130.515 ;
        RECT 36.520 129.955 37.535 130.155 ;
        RECT 37.835 129.995 38.005 130.325 ;
        RECT 38.175 129.775 38.505 130.155 ;
        RECT 38.720 130.035 38.945 132.155 ;
        RECT 39.115 131.825 39.445 132.325 ;
        RECT 39.615 131.655 39.785 132.155 ;
        RECT 39.120 131.485 39.785 131.655 ;
        RECT 40.135 131.580 40.405 132.325 ;
        RECT 41.035 132.320 47.310 132.325 ;
        RECT 39.120 130.495 39.350 131.485 ;
        RECT 40.575 131.410 40.865 132.150 ;
        RECT 41.035 131.595 41.290 132.320 ;
        RECT 41.475 131.425 41.735 132.150 ;
        RECT 41.905 131.595 42.150 132.320 ;
        RECT 42.335 131.425 42.595 132.150 ;
        RECT 42.765 131.595 43.010 132.320 ;
        RECT 43.195 131.425 43.455 132.150 ;
        RECT 43.625 131.595 43.870 132.320 ;
        RECT 44.040 131.425 44.300 132.150 ;
        RECT 44.470 131.595 44.730 132.320 ;
        RECT 44.900 131.425 45.160 132.150 ;
        RECT 45.330 131.595 45.590 132.320 ;
        RECT 45.760 131.425 46.020 132.150 ;
        RECT 46.190 131.595 46.450 132.320 ;
        RECT 46.620 131.425 46.880 132.150 ;
        RECT 47.050 131.525 47.310 132.320 ;
        RECT 41.475 131.410 46.880 131.425 ;
        RECT 39.520 130.665 39.870 131.315 ;
        RECT 40.135 131.185 46.880 131.410 ;
        RECT 40.135 130.595 41.300 131.185 ;
        RECT 47.480 131.015 47.730 132.150 ;
        RECT 47.910 131.515 48.170 132.325 ;
        RECT 48.345 131.015 48.590 132.155 ;
        RECT 48.770 131.515 49.065 132.325 ;
        RECT 50.165 131.160 50.455 132.325 ;
        RECT 51.085 131.235 54.595 132.325 ;
        RECT 54.770 131.890 60.115 132.325 ;
        RECT 60.290 131.890 65.635 132.325 ;
        RECT 41.470 130.765 48.590 131.015 ;
        RECT 39.120 130.325 39.785 130.495 ;
        RECT 40.135 130.425 46.880 130.595 ;
        RECT 39.115 129.775 39.445 130.155 ;
        RECT 39.615 130.035 39.785 130.325 ;
        RECT 40.135 129.775 40.435 130.255 ;
        RECT 40.605 129.970 40.865 130.425 ;
        RECT 41.035 129.775 41.295 130.255 ;
        RECT 41.475 129.970 41.735 130.425 ;
        RECT 41.905 129.775 42.155 130.255 ;
        RECT 42.335 129.970 42.595 130.425 ;
        RECT 42.765 129.775 43.015 130.255 ;
        RECT 43.195 129.970 43.455 130.425 ;
        RECT 43.625 129.775 43.870 130.255 ;
        RECT 44.040 129.970 44.315 130.425 ;
        RECT 44.485 129.775 44.730 130.255 ;
        RECT 44.900 129.970 45.160 130.425 ;
        RECT 45.330 129.775 45.590 130.255 ;
        RECT 45.760 129.970 46.020 130.425 ;
        RECT 46.190 129.775 46.450 130.255 ;
        RECT 46.620 129.970 46.880 130.425 ;
        RECT 47.050 129.775 47.310 130.335 ;
        RECT 47.480 129.955 47.730 130.765 ;
        RECT 47.910 129.775 48.170 130.300 ;
        RECT 48.340 129.955 48.590 130.765 ;
        RECT 48.760 130.455 49.075 131.015 ;
        RECT 51.085 130.715 52.775 131.235 ;
        RECT 52.945 130.545 54.595 131.065 ;
        RECT 56.360 130.640 56.710 131.890 ;
        RECT 48.770 129.775 49.075 130.285 ;
        RECT 50.165 129.775 50.455 130.500 ;
        RECT 51.085 129.775 54.595 130.545 ;
        RECT 58.190 130.320 58.530 131.150 ;
        RECT 61.880 130.640 62.230 131.890 ;
        RECT 65.805 131.565 66.320 131.975 ;
        RECT 66.555 131.565 66.725 132.325 ;
        RECT 66.895 131.985 68.925 132.155 ;
        RECT 63.710 130.320 64.050 131.150 ;
        RECT 65.805 130.755 66.145 131.565 ;
        RECT 66.895 131.320 67.065 131.985 ;
        RECT 67.460 131.645 68.585 131.815 ;
        RECT 66.315 131.130 67.065 131.320 ;
        RECT 67.235 131.305 68.245 131.475 ;
        RECT 65.805 130.585 67.035 130.755 ;
        RECT 54.770 129.775 60.115 130.320 ;
        RECT 60.290 129.775 65.635 130.320 ;
        RECT 66.080 129.980 66.325 130.585 ;
        RECT 66.545 129.775 67.055 130.310 ;
        RECT 67.235 129.945 67.425 131.305 ;
        RECT 67.595 130.625 67.870 131.105 ;
        RECT 67.595 130.455 67.875 130.625 ;
        RECT 68.075 130.505 68.245 131.305 ;
        RECT 68.415 130.515 68.585 131.645 ;
        RECT 68.755 131.015 68.925 131.985 ;
        RECT 69.095 131.185 69.265 132.325 ;
        RECT 69.435 131.185 69.770 132.155 ;
        RECT 69.950 131.900 70.285 132.325 ;
        RECT 70.455 131.720 70.640 132.125 ;
        RECT 68.755 130.685 68.950 131.015 ;
        RECT 69.175 130.685 69.430 131.015 ;
        RECT 69.175 130.515 69.345 130.685 ;
        RECT 69.600 130.515 69.770 131.185 ;
        RECT 67.595 129.945 67.870 130.455 ;
        RECT 68.415 130.345 69.345 130.515 ;
        RECT 68.415 130.310 68.590 130.345 ;
        RECT 68.060 129.945 68.590 130.310 ;
        RECT 69.015 129.775 69.345 130.175 ;
        RECT 69.515 129.945 69.770 130.515 ;
        RECT 69.975 131.545 70.640 131.720 ;
        RECT 70.845 131.545 71.175 132.325 ;
        RECT 69.975 130.515 70.315 131.545 ;
        RECT 71.345 131.355 71.615 132.125 ;
        RECT 70.485 131.185 71.615 131.355 ;
        RECT 70.485 130.685 70.735 131.185 ;
        RECT 69.975 130.345 70.660 130.515 ;
        RECT 70.915 130.435 71.275 131.015 ;
        RECT 69.950 129.775 70.285 130.175 ;
        RECT 70.455 129.945 70.660 130.345 ;
        RECT 71.445 130.275 71.615 131.185 ;
        RECT 70.870 129.775 71.145 130.255 ;
        RECT 71.355 129.945 71.615 130.275 ;
        RECT 71.785 131.605 72.245 132.155 ;
        RECT 72.435 131.605 72.765 132.325 ;
        RECT 71.785 130.235 72.035 131.605 ;
        RECT 72.965 131.435 73.265 131.985 ;
        RECT 73.435 131.655 73.715 132.325 ;
        RECT 72.325 131.265 73.265 131.435 ;
        RECT 72.325 131.015 72.495 131.265 ;
        RECT 73.635 131.015 73.900 131.375 ;
        RECT 72.205 130.685 72.495 131.015 ;
        RECT 72.665 130.765 73.005 131.015 ;
        RECT 73.225 130.765 73.900 131.015 ;
        RECT 74.085 131.355 74.355 132.125 ;
        RECT 74.525 131.545 74.855 132.325 ;
        RECT 75.060 131.720 75.245 132.125 ;
        RECT 75.415 131.900 75.750 132.325 ;
        RECT 75.060 131.545 75.725 131.720 ;
        RECT 74.085 131.185 75.215 131.355 ;
        RECT 72.325 130.595 72.495 130.685 ;
        RECT 72.325 130.405 73.715 130.595 ;
        RECT 71.785 129.945 72.345 130.235 ;
        RECT 72.515 129.775 72.765 130.235 ;
        RECT 73.385 130.045 73.715 130.405 ;
        RECT 74.085 130.275 74.255 131.185 ;
        RECT 74.425 130.435 74.785 131.015 ;
        RECT 74.965 130.685 75.215 131.185 ;
        RECT 75.385 130.515 75.725 131.545 ;
        RECT 75.925 131.160 76.215 132.325 ;
        RECT 76.845 131.235 78.515 132.325 ;
        RECT 78.685 131.605 79.145 132.155 ;
        RECT 79.335 131.605 79.665 132.325 ;
        RECT 76.845 130.715 77.595 131.235 ;
        RECT 77.765 130.545 78.515 131.065 ;
        RECT 75.040 130.345 75.725 130.515 ;
        RECT 74.085 129.945 74.345 130.275 ;
        RECT 74.555 129.775 74.830 130.255 ;
        RECT 75.040 129.945 75.245 130.345 ;
        RECT 75.415 129.775 75.750 130.175 ;
        RECT 75.925 129.775 76.215 130.500 ;
        RECT 76.845 129.775 78.515 130.545 ;
        RECT 78.685 130.235 78.935 131.605 ;
        RECT 79.865 131.435 80.165 131.985 ;
        RECT 80.335 131.655 80.615 132.325 ;
        RECT 79.225 131.265 80.165 131.435 ;
        RECT 79.225 131.015 79.395 131.265 ;
        RECT 80.535 131.015 80.800 131.375 ;
        RECT 79.105 130.685 79.395 131.015 ;
        RECT 79.565 130.765 79.905 131.015 ;
        RECT 80.125 130.765 80.800 131.015 ;
        RECT 80.985 131.235 83.575 132.325 ;
        RECT 83.750 131.890 89.095 132.325 ;
        RECT 80.985 130.715 82.195 131.235 ;
        RECT 79.225 130.595 79.395 130.685 ;
        RECT 79.225 130.405 80.615 130.595 ;
        RECT 82.365 130.545 83.575 131.065 ;
        RECT 85.340 130.640 85.690 131.890 ;
        RECT 89.305 131.185 89.535 132.325 ;
        RECT 89.705 131.175 90.035 132.155 ;
        RECT 90.205 131.185 90.415 132.325 ;
        RECT 90.755 131.525 90.925 132.325 ;
        RECT 91.095 131.305 91.425 132.155 ;
        RECT 91.595 131.525 91.765 132.325 ;
        RECT 91.935 131.305 92.265 132.155 ;
        RECT 92.435 131.525 92.605 132.325 ;
        RECT 92.775 131.305 93.105 132.155 ;
        RECT 93.275 131.525 93.445 132.325 ;
        RECT 93.615 131.305 93.945 132.155 ;
        RECT 94.115 131.525 94.285 132.325 ;
        RECT 94.455 131.305 94.785 132.155 ;
        RECT 94.955 131.525 95.125 132.325 ;
        RECT 95.295 131.305 95.625 132.155 ;
        RECT 95.795 131.525 95.965 132.325 ;
        RECT 96.135 131.305 96.465 132.155 ;
        RECT 96.635 131.525 96.805 132.325 ;
        RECT 96.975 131.305 97.305 132.155 ;
        RECT 97.475 131.525 97.645 132.325 ;
        RECT 97.815 131.305 98.145 132.155 ;
        RECT 98.315 131.525 98.485 132.325 ;
        RECT 98.655 131.305 98.985 132.155 ;
        RECT 99.155 131.525 99.325 132.325 ;
        RECT 99.495 131.305 99.825 132.155 ;
        RECT 99.995 131.475 100.165 132.325 ;
        RECT 100.335 131.305 100.665 132.155 ;
        RECT 100.835 131.475 101.005 132.325 ;
        RECT 101.175 131.305 101.505 132.155 ;
        RECT 78.685 129.945 79.245 130.235 ;
        RECT 79.415 129.775 79.665 130.235 ;
        RECT 80.285 130.045 80.615 130.405 ;
        RECT 80.985 129.775 83.575 130.545 ;
        RECT 87.170 130.320 87.510 131.150 ;
        RECT 89.285 130.765 89.615 131.015 ;
        RECT 83.750 129.775 89.095 130.320 ;
        RECT 89.305 129.775 89.535 130.595 ;
        RECT 89.785 130.575 90.035 131.175 ;
        RECT 90.645 131.135 97.305 131.305 ;
        RECT 97.475 131.135 99.825 131.305 ;
        RECT 99.995 131.135 101.505 131.305 ;
        RECT 101.685 131.160 101.975 132.325 ;
        RECT 102.605 131.235 104.275 132.325 ;
        RECT 104.450 131.890 109.795 132.325 ;
        RECT 90.645 130.595 90.920 131.135 ;
        RECT 97.475 130.965 97.650 131.135 ;
        RECT 99.995 130.965 100.165 131.135 ;
        RECT 91.090 130.765 97.650 130.965 ;
        RECT 97.855 130.765 100.165 130.965 ;
        RECT 100.335 130.765 101.510 130.965 ;
        RECT 97.475 130.595 97.650 130.765 ;
        RECT 99.995 130.595 100.165 130.765 ;
        RECT 102.605 130.715 103.355 131.235 ;
        RECT 89.705 129.945 90.035 130.575 ;
        RECT 90.205 129.775 90.415 130.595 ;
        RECT 90.645 130.425 97.305 130.595 ;
        RECT 97.475 130.425 99.825 130.595 ;
        RECT 99.995 130.425 101.505 130.595 ;
        RECT 103.525 130.545 104.275 131.065 ;
        RECT 106.040 130.640 106.390 131.890 ;
        RECT 109.965 131.605 110.425 132.155 ;
        RECT 110.615 131.605 110.945 132.325 ;
        RECT 90.755 129.775 90.925 130.255 ;
        RECT 91.095 129.950 91.425 130.425 ;
        RECT 91.595 129.775 91.765 130.255 ;
        RECT 91.935 129.950 92.265 130.425 ;
        RECT 92.435 129.775 92.605 130.255 ;
        RECT 92.775 129.950 93.105 130.425 ;
        RECT 93.275 129.775 93.445 130.255 ;
        RECT 93.615 129.950 93.945 130.425 ;
        RECT 94.115 129.775 94.285 130.255 ;
        RECT 94.455 129.950 94.785 130.425 ;
        RECT 94.955 129.775 95.125 130.255 ;
        RECT 95.295 129.950 95.625 130.425 ;
        RECT 95.375 129.945 95.545 129.950 ;
        RECT 95.795 129.775 95.965 130.255 ;
        RECT 96.135 129.950 96.465 130.425 ;
        RECT 96.215 129.945 96.385 129.950 ;
        RECT 96.635 129.775 96.805 130.255 ;
        RECT 96.975 129.950 97.305 130.425 ;
        RECT 97.055 129.945 97.305 129.950 ;
        RECT 97.475 129.775 97.645 130.255 ;
        RECT 97.815 129.950 98.145 130.425 ;
        RECT 98.315 129.775 98.485 130.255 ;
        RECT 98.655 129.950 98.985 130.425 ;
        RECT 99.155 129.775 99.325 130.255 ;
        RECT 99.495 129.950 99.825 130.425 ;
        RECT 99.995 129.775 100.165 130.255 ;
        RECT 100.335 129.950 100.665 130.425 ;
        RECT 100.835 129.775 101.005 130.255 ;
        RECT 101.175 129.950 101.505 130.425 ;
        RECT 101.685 129.775 101.975 130.500 ;
        RECT 102.605 129.775 104.275 130.545 ;
        RECT 107.870 130.320 108.210 131.150 ;
        RECT 104.450 129.775 109.795 130.320 ;
        RECT 109.965 130.235 110.215 131.605 ;
        RECT 111.145 131.435 111.445 131.985 ;
        RECT 111.615 131.655 111.895 132.325 ;
        RECT 110.505 131.265 111.445 131.435 ;
        RECT 110.505 131.015 110.675 131.265 ;
        RECT 111.815 131.015 112.080 131.375 ;
        RECT 110.385 130.685 110.675 131.015 ;
        RECT 110.845 130.765 111.185 131.015 ;
        RECT 111.405 130.765 112.080 131.015 ;
        RECT 112.725 131.235 115.315 132.325 ;
        RECT 115.490 131.890 120.835 132.325 ;
        RECT 121.010 131.890 126.355 132.325 ;
        RECT 112.725 130.715 113.935 131.235 ;
        RECT 110.505 130.595 110.675 130.685 ;
        RECT 110.505 130.405 111.895 130.595 ;
        RECT 114.105 130.545 115.315 131.065 ;
        RECT 117.080 130.640 117.430 131.890 ;
        RECT 109.965 129.945 110.525 130.235 ;
        RECT 110.695 129.775 110.945 130.235 ;
        RECT 111.565 130.045 111.895 130.405 ;
        RECT 112.725 129.775 115.315 130.545 ;
        RECT 118.910 130.320 119.250 131.150 ;
        RECT 122.600 130.640 122.950 131.890 ;
        RECT 126.525 131.235 127.735 132.325 ;
        RECT 124.430 130.320 124.770 131.150 ;
        RECT 126.525 130.695 127.045 131.235 ;
        RECT 127.215 130.525 127.735 131.065 ;
        RECT 115.490 129.775 120.835 130.320 ;
        RECT 121.010 129.775 126.355 130.320 ;
        RECT 126.525 129.775 127.735 130.525 ;
        RECT 14.660 129.605 127.820 129.775 ;
        RECT 14.745 128.855 15.955 129.605 ;
        RECT 16.125 128.855 17.335 129.605 ;
        RECT 17.880 129.265 18.135 129.425 ;
        RECT 17.795 129.095 18.135 129.265 ;
        RECT 18.315 129.145 18.600 129.605 ;
        RECT 14.745 128.315 15.265 128.855 ;
        RECT 15.435 128.145 15.955 128.685 ;
        RECT 14.745 127.055 15.955 128.145 ;
        RECT 16.125 128.145 16.645 128.685 ;
        RECT 16.815 128.315 17.335 128.855 ;
        RECT 17.880 128.895 18.135 129.095 ;
        RECT 16.125 127.055 17.335 128.145 ;
        RECT 17.880 128.035 18.060 128.895 ;
        RECT 18.780 128.695 19.030 129.345 ;
        RECT 18.230 128.365 19.030 128.695 ;
        RECT 17.880 127.365 18.135 128.035 ;
        RECT 18.315 127.055 18.600 127.855 ;
        RECT 18.780 127.775 19.030 128.365 ;
        RECT 19.230 129.010 19.550 129.340 ;
        RECT 19.730 129.125 20.390 129.605 ;
        RECT 20.590 129.215 21.440 129.385 ;
        RECT 19.230 128.115 19.420 129.010 ;
        RECT 19.740 128.685 20.400 128.955 ;
        RECT 20.070 128.625 20.400 128.685 ;
        RECT 19.590 128.455 19.920 128.515 ;
        RECT 20.590 128.455 20.760 129.215 ;
        RECT 22.000 129.145 22.320 129.605 ;
        RECT 22.520 128.965 22.770 129.395 ;
        RECT 23.060 129.165 23.470 129.605 ;
        RECT 23.640 129.225 24.655 129.425 ;
        RECT 20.930 128.795 22.180 128.965 ;
        RECT 20.930 128.675 21.260 128.795 ;
        RECT 19.590 128.285 21.490 128.455 ;
        RECT 19.230 127.945 21.150 128.115 ;
        RECT 19.230 127.925 19.550 127.945 ;
        RECT 18.780 127.265 19.110 127.775 ;
        RECT 19.380 127.315 19.550 127.925 ;
        RECT 21.320 127.775 21.490 128.285 ;
        RECT 21.660 128.215 21.840 128.625 ;
        RECT 22.010 128.035 22.180 128.795 ;
        RECT 19.720 127.055 20.050 127.745 ;
        RECT 20.280 127.605 21.490 127.775 ;
        RECT 21.660 127.725 22.180 128.035 ;
        RECT 22.350 128.625 22.770 128.965 ;
        RECT 23.060 128.625 23.470 128.955 ;
        RECT 22.350 127.855 22.540 128.625 ;
        RECT 23.640 128.495 23.810 129.225 ;
        RECT 24.955 129.055 25.125 129.385 ;
        RECT 25.295 129.225 25.625 129.605 ;
        RECT 23.980 128.675 24.330 129.045 ;
        RECT 23.640 128.455 24.060 128.495 ;
        RECT 22.710 128.285 24.060 128.455 ;
        RECT 22.710 128.125 22.960 128.285 ;
        RECT 23.470 127.855 23.720 128.115 ;
        RECT 22.350 127.605 23.720 127.855 ;
        RECT 20.280 127.315 20.520 127.605 ;
        RECT 21.320 127.525 21.490 127.605 ;
        RECT 20.720 127.055 21.140 127.435 ;
        RECT 21.320 127.275 21.950 127.525 ;
        RECT 22.420 127.055 22.750 127.435 ;
        RECT 22.920 127.315 23.090 127.605 ;
        RECT 23.890 127.440 24.060 128.285 ;
        RECT 24.510 128.115 24.730 128.985 ;
        RECT 24.955 128.865 25.650 129.055 ;
        RECT 24.230 127.735 24.730 128.115 ;
        RECT 24.900 128.065 25.310 128.685 ;
        RECT 25.480 127.895 25.650 128.865 ;
        RECT 24.955 127.725 25.650 127.895 ;
        RECT 23.270 127.055 23.650 127.435 ;
        RECT 23.890 127.270 24.720 127.440 ;
        RECT 24.955 127.225 25.125 127.725 ;
        RECT 25.295 127.055 25.625 127.555 ;
        RECT 25.840 127.225 26.065 129.345 ;
        RECT 26.235 129.225 26.565 129.605 ;
        RECT 26.735 129.055 26.905 129.345 ;
        RECT 28.090 129.060 33.435 129.605 ;
        RECT 26.240 128.885 26.905 129.055 ;
        RECT 26.240 127.895 26.470 128.885 ;
        RECT 26.640 128.065 26.990 128.715 ;
        RECT 26.240 127.725 26.905 127.895 ;
        RECT 26.235 127.055 26.565 127.555 ;
        RECT 26.735 127.225 26.905 127.725 ;
        RECT 29.680 127.490 30.030 128.740 ;
        RECT 31.510 128.230 31.850 129.060 ;
        RECT 33.645 128.785 33.875 129.605 ;
        RECT 34.045 128.805 34.375 129.435 ;
        RECT 33.625 128.365 33.955 128.615 ;
        RECT 34.125 128.205 34.375 128.805 ;
        RECT 34.545 128.785 34.755 129.605 ;
        RECT 35.445 128.835 37.115 129.605 ;
        RECT 37.285 128.880 37.575 129.605 ;
        RECT 38.665 128.930 38.925 129.435 ;
        RECT 39.105 129.225 39.435 129.605 ;
        RECT 39.615 129.055 39.785 129.435 ;
        RECT 28.090 127.055 33.435 127.490 ;
        RECT 33.645 127.055 33.875 128.195 ;
        RECT 34.045 127.225 34.375 128.205 ;
        RECT 34.545 127.055 34.755 128.195 ;
        RECT 35.445 128.145 36.195 128.665 ;
        RECT 36.365 128.315 37.115 128.835 ;
        RECT 35.445 127.055 37.115 128.145 ;
        RECT 37.285 127.055 37.575 128.220 ;
        RECT 38.665 128.130 38.835 128.930 ;
        RECT 39.120 128.885 39.785 129.055 ;
        RECT 40.245 128.975 40.575 129.335 ;
        RECT 41.195 129.145 41.445 129.605 ;
        RECT 41.615 129.145 42.175 129.435 ;
        RECT 39.120 128.630 39.290 128.885 ;
        RECT 40.245 128.785 41.635 128.975 ;
        RECT 39.005 128.300 39.290 128.630 ;
        RECT 39.525 128.335 39.855 128.705 ;
        RECT 41.465 128.695 41.635 128.785 ;
        RECT 40.060 128.365 40.735 128.615 ;
        RECT 40.955 128.365 41.295 128.615 ;
        RECT 41.465 128.365 41.755 128.695 ;
        RECT 39.120 128.155 39.290 128.300 ;
        RECT 38.665 127.225 38.935 128.130 ;
        RECT 39.120 127.985 39.785 128.155 ;
        RECT 40.060 128.005 40.325 128.365 ;
        RECT 41.465 128.115 41.635 128.365 ;
        RECT 39.105 127.055 39.435 127.815 ;
        RECT 39.615 127.225 39.785 127.985 ;
        RECT 40.695 127.945 41.635 128.115 ;
        RECT 40.245 127.055 40.525 127.725 ;
        RECT 40.695 127.395 40.995 127.945 ;
        RECT 41.925 127.775 42.175 129.145 ;
        RECT 42.545 128.975 42.875 129.335 ;
        RECT 43.495 129.145 43.745 129.605 ;
        RECT 43.915 129.145 44.475 129.435 ;
        RECT 42.545 128.785 43.935 128.975 ;
        RECT 43.765 128.695 43.935 128.785 ;
        RECT 42.360 128.365 43.035 128.615 ;
        RECT 43.255 128.365 43.595 128.615 ;
        RECT 43.765 128.365 44.055 128.695 ;
        RECT 42.360 128.005 42.625 128.365 ;
        RECT 43.765 128.115 43.935 128.365 ;
        RECT 41.195 127.055 41.525 127.775 ;
        RECT 41.715 127.225 42.175 127.775 ;
        RECT 42.995 127.945 43.935 128.115 ;
        RECT 42.545 127.055 42.825 127.725 ;
        RECT 42.995 127.395 43.295 127.945 ;
        RECT 44.225 127.775 44.475 129.145 ;
        RECT 45.315 128.915 45.645 129.605 ;
        RECT 46.105 129.010 46.725 129.435 ;
        RECT 46.895 129.115 47.225 129.605 ;
        RECT 46.365 128.675 46.725 129.010 ;
        RECT 47.605 128.975 47.935 129.335 ;
        RECT 48.555 129.145 48.805 129.605 ;
        RECT 48.975 129.145 49.535 129.435 ;
        RECT 45.305 128.395 46.725 128.675 ;
        RECT 43.495 127.055 43.825 127.775 ;
        RECT 44.015 127.225 44.475 127.775 ;
        RECT 44.775 127.055 45.105 128.225 ;
        RECT 45.305 127.225 45.635 128.395 ;
        RECT 45.835 127.055 46.165 128.225 ;
        RECT 46.365 127.225 46.725 128.395 ;
        RECT 46.895 128.365 47.235 128.945 ;
        RECT 47.605 128.785 48.995 128.975 ;
        RECT 48.825 128.695 48.995 128.785 ;
        RECT 47.420 128.365 48.095 128.615 ;
        RECT 48.315 128.365 48.655 128.615 ;
        RECT 48.825 128.365 49.115 128.695 ;
        RECT 46.895 127.055 47.225 128.195 ;
        RECT 47.420 128.005 47.685 128.365 ;
        RECT 48.825 128.115 48.995 128.365 ;
        RECT 48.055 127.945 48.995 128.115 ;
        RECT 47.605 127.055 47.885 127.725 ;
        RECT 48.055 127.395 48.355 127.945 ;
        RECT 49.285 127.775 49.535 129.145 ;
        RECT 49.705 128.855 50.915 129.605 ;
        RECT 48.555 127.055 48.885 127.775 ;
        RECT 49.075 127.225 49.535 127.775 ;
        RECT 49.705 128.145 50.225 128.685 ;
        RECT 50.395 128.315 50.915 128.855 ;
        RECT 51.085 128.835 54.595 129.605 ;
        RECT 51.085 128.145 52.775 128.665 ;
        RECT 52.945 128.315 54.595 128.835 ;
        RECT 55.040 128.795 55.285 129.400 ;
        RECT 55.505 129.070 56.015 129.605 ;
        RECT 54.765 128.625 55.995 128.795 ;
        RECT 49.705 127.055 50.915 128.145 ;
        RECT 51.085 127.055 54.595 128.145 ;
        RECT 54.765 127.815 55.105 128.625 ;
        RECT 55.275 128.060 56.025 128.250 ;
        RECT 54.765 127.405 55.280 127.815 ;
        RECT 55.515 127.055 55.685 127.815 ;
        RECT 55.855 127.395 56.025 128.060 ;
        RECT 56.195 128.075 56.385 129.435 ;
        RECT 56.555 129.265 56.830 129.435 ;
        RECT 56.555 129.095 56.835 129.265 ;
        RECT 56.555 128.275 56.830 129.095 ;
        RECT 57.020 129.070 57.550 129.435 ;
        RECT 57.975 129.205 58.305 129.605 ;
        RECT 57.375 129.035 57.550 129.070 ;
        RECT 57.035 128.075 57.205 128.875 ;
        RECT 56.195 127.905 57.205 128.075 ;
        RECT 57.375 128.865 58.305 129.035 ;
        RECT 58.475 128.865 58.730 129.435 ;
        RECT 57.375 127.735 57.545 128.865 ;
        RECT 58.135 128.695 58.305 128.865 ;
        RECT 56.420 127.565 57.545 127.735 ;
        RECT 57.715 128.365 57.910 128.695 ;
        RECT 58.135 128.365 58.390 128.695 ;
        RECT 57.715 127.395 57.885 128.365 ;
        RECT 58.560 128.195 58.730 128.865 ;
        RECT 59.365 128.835 62.875 129.605 ;
        RECT 63.045 128.880 63.335 129.605 ;
        RECT 63.505 128.855 64.715 129.605 ;
        RECT 65.260 129.265 65.515 129.425 ;
        RECT 65.175 129.095 65.515 129.265 ;
        RECT 65.695 129.145 65.980 129.605 ;
        RECT 55.855 127.225 57.885 127.395 ;
        RECT 58.055 127.055 58.225 128.195 ;
        RECT 58.395 127.225 58.730 128.195 ;
        RECT 59.365 128.145 61.055 128.665 ;
        RECT 61.225 128.315 62.875 128.835 ;
        RECT 59.365 127.055 62.875 128.145 ;
        RECT 63.045 127.055 63.335 128.220 ;
        RECT 63.505 128.145 64.025 128.685 ;
        RECT 64.195 128.315 64.715 128.855 ;
        RECT 65.260 128.895 65.515 129.095 ;
        RECT 63.505 127.055 64.715 128.145 ;
        RECT 65.260 128.035 65.440 128.895 ;
        RECT 66.160 128.695 66.410 129.345 ;
        RECT 65.610 128.365 66.410 128.695 ;
        RECT 65.260 127.365 65.515 128.035 ;
        RECT 65.695 127.055 65.980 127.855 ;
        RECT 66.160 127.775 66.410 128.365 ;
        RECT 66.610 129.010 66.930 129.340 ;
        RECT 67.110 129.125 67.770 129.605 ;
        RECT 67.970 129.215 68.820 129.385 ;
        RECT 66.610 128.115 66.800 129.010 ;
        RECT 67.120 128.685 67.780 128.955 ;
        RECT 67.450 128.625 67.780 128.685 ;
        RECT 66.970 128.455 67.300 128.515 ;
        RECT 67.970 128.455 68.140 129.215 ;
        RECT 69.380 129.145 69.700 129.605 ;
        RECT 69.900 128.965 70.150 129.395 ;
        RECT 70.440 129.165 70.850 129.605 ;
        RECT 71.020 129.225 72.035 129.425 ;
        RECT 68.310 128.795 69.560 128.965 ;
        RECT 68.310 128.675 68.640 128.795 ;
        RECT 66.970 128.285 68.870 128.455 ;
        RECT 66.610 127.945 68.530 128.115 ;
        RECT 66.610 127.925 66.930 127.945 ;
        RECT 66.160 127.265 66.490 127.775 ;
        RECT 66.760 127.315 66.930 127.925 ;
        RECT 68.700 127.775 68.870 128.285 ;
        RECT 69.040 128.215 69.220 128.625 ;
        RECT 69.390 128.035 69.560 128.795 ;
        RECT 67.100 127.055 67.430 127.745 ;
        RECT 67.660 127.605 68.870 127.775 ;
        RECT 69.040 127.725 69.560 128.035 ;
        RECT 69.730 128.625 70.150 128.965 ;
        RECT 70.440 128.625 70.850 128.955 ;
        RECT 69.730 127.855 69.920 128.625 ;
        RECT 71.020 128.495 71.190 129.225 ;
        RECT 72.335 129.055 72.505 129.385 ;
        RECT 72.675 129.225 73.005 129.605 ;
        RECT 71.360 128.675 71.710 129.045 ;
        RECT 71.020 128.455 71.440 128.495 ;
        RECT 70.090 128.285 71.440 128.455 ;
        RECT 70.090 128.125 70.340 128.285 ;
        RECT 70.850 127.855 71.100 128.115 ;
        RECT 69.730 127.605 71.100 127.855 ;
        RECT 67.660 127.315 67.900 127.605 ;
        RECT 68.700 127.525 68.870 127.605 ;
        RECT 68.100 127.055 68.520 127.435 ;
        RECT 68.700 127.275 69.330 127.525 ;
        RECT 69.800 127.055 70.130 127.435 ;
        RECT 70.300 127.315 70.470 127.605 ;
        RECT 71.270 127.440 71.440 128.285 ;
        RECT 71.890 128.115 72.110 128.985 ;
        RECT 72.335 128.865 73.030 129.055 ;
        RECT 71.610 127.735 72.110 128.115 ;
        RECT 72.280 128.065 72.690 128.685 ;
        RECT 72.860 127.895 73.030 128.865 ;
        RECT 72.335 127.725 73.030 127.895 ;
        RECT 70.650 127.055 71.030 127.435 ;
        RECT 71.270 127.270 72.100 127.440 ;
        RECT 72.335 127.225 72.505 127.725 ;
        RECT 72.675 127.055 73.005 127.555 ;
        RECT 73.220 127.225 73.445 129.345 ;
        RECT 73.615 129.225 73.945 129.605 ;
        RECT 74.115 129.055 74.285 129.345 ;
        RECT 73.620 128.885 74.285 129.055 ;
        RECT 74.745 128.975 75.075 129.335 ;
        RECT 75.695 129.145 75.945 129.605 ;
        RECT 76.115 129.145 76.675 129.435 ;
        RECT 73.620 127.895 73.850 128.885 ;
        RECT 74.745 128.785 76.135 128.975 ;
        RECT 74.020 128.065 74.370 128.715 ;
        RECT 75.965 128.695 76.135 128.785 ;
        RECT 74.560 128.365 75.235 128.615 ;
        RECT 75.455 128.365 75.795 128.615 ;
        RECT 75.965 128.365 76.255 128.695 ;
        RECT 74.560 128.005 74.825 128.365 ;
        RECT 75.965 128.115 76.135 128.365 ;
        RECT 75.195 127.945 76.135 128.115 ;
        RECT 73.620 127.725 74.285 127.895 ;
        RECT 73.615 127.055 73.945 127.555 ;
        RECT 74.115 127.225 74.285 127.725 ;
        RECT 74.745 127.055 75.025 127.725 ;
        RECT 75.195 127.395 75.495 127.945 ;
        RECT 76.425 127.775 76.675 129.145 ;
        RECT 77.045 128.975 77.375 129.335 ;
        RECT 77.995 129.145 78.245 129.605 ;
        RECT 78.415 129.145 78.975 129.435 ;
        RECT 77.045 128.785 78.435 128.975 ;
        RECT 78.265 128.695 78.435 128.785 ;
        RECT 76.860 128.365 77.535 128.615 ;
        RECT 77.755 128.365 78.095 128.615 ;
        RECT 78.265 128.365 78.555 128.695 ;
        RECT 76.860 128.005 77.125 128.365 ;
        RECT 78.265 128.115 78.435 128.365 ;
        RECT 75.695 127.055 76.025 127.775 ;
        RECT 76.215 127.225 76.675 127.775 ;
        RECT 77.495 127.945 78.435 128.115 ;
        RECT 77.045 127.055 77.325 127.725 ;
        RECT 77.495 127.395 77.795 127.945 ;
        RECT 78.725 127.775 78.975 129.145 ;
        RECT 79.420 128.795 79.665 129.400 ;
        RECT 79.885 129.070 80.395 129.605 ;
        RECT 77.995 127.055 78.325 127.775 ;
        RECT 78.515 127.225 78.975 127.775 ;
        RECT 79.145 128.625 80.375 128.795 ;
        RECT 79.145 127.815 79.485 128.625 ;
        RECT 79.655 128.060 80.405 128.250 ;
        RECT 79.145 127.405 79.660 127.815 ;
        RECT 79.895 127.055 80.065 127.815 ;
        RECT 80.235 127.395 80.405 128.060 ;
        RECT 80.575 128.075 80.765 129.435 ;
        RECT 80.935 128.585 81.210 129.435 ;
        RECT 81.400 129.070 81.930 129.435 ;
        RECT 82.355 129.205 82.685 129.605 ;
        RECT 81.755 129.035 81.930 129.070 ;
        RECT 80.935 128.415 81.215 128.585 ;
        RECT 80.935 128.275 81.210 128.415 ;
        RECT 81.415 128.075 81.585 128.875 ;
        RECT 80.575 127.905 81.585 128.075 ;
        RECT 81.755 128.865 82.685 129.035 ;
        RECT 82.855 128.865 83.110 129.435 ;
        RECT 81.755 127.735 81.925 128.865 ;
        RECT 82.515 128.695 82.685 128.865 ;
        RECT 80.800 127.565 81.925 127.735 ;
        RECT 82.095 128.365 82.290 128.695 ;
        RECT 82.515 128.365 82.770 128.695 ;
        RECT 82.095 127.395 82.265 128.365 ;
        RECT 82.940 128.195 83.110 128.865 ;
        RECT 80.235 127.225 82.265 127.395 ;
        RECT 82.435 127.055 82.605 128.195 ;
        RECT 82.775 127.225 83.110 128.195 ;
        RECT 83.285 129.145 83.845 129.435 ;
        RECT 84.015 129.145 84.265 129.605 ;
        RECT 83.285 127.775 83.535 129.145 ;
        RECT 84.885 128.975 85.215 129.335 ;
        RECT 83.825 128.785 85.215 128.975 ;
        RECT 85.585 128.835 87.255 129.605 ;
        RECT 87.515 129.055 87.685 129.435 ;
        RECT 87.865 129.225 88.195 129.605 ;
        RECT 87.515 128.885 88.180 129.055 ;
        RECT 88.375 128.930 88.635 129.435 ;
        RECT 83.825 128.695 83.995 128.785 ;
        RECT 83.705 128.365 83.995 128.695 ;
        RECT 84.165 128.365 84.505 128.615 ;
        RECT 84.725 128.365 85.400 128.615 ;
        RECT 83.825 128.115 83.995 128.365 ;
        RECT 83.825 127.945 84.765 128.115 ;
        RECT 85.135 128.005 85.400 128.365 ;
        RECT 85.585 128.145 86.335 128.665 ;
        RECT 86.505 128.315 87.255 128.835 ;
        RECT 87.445 128.335 87.775 128.705 ;
        RECT 88.010 128.630 88.180 128.885 ;
        RECT 88.010 128.300 88.295 128.630 ;
        RECT 88.010 128.155 88.180 128.300 ;
        RECT 83.285 127.225 83.745 127.775 ;
        RECT 83.935 127.055 84.265 127.775 ;
        RECT 84.465 127.395 84.765 127.945 ;
        RECT 84.935 127.055 85.215 127.725 ;
        RECT 85.585 127.055 87.255 128.145 ;
        RECT 87.515 127.985 88.180 128.155 ;
        RECT 88.465 128.130 88.635 128.930 ;
        RECT 88.805 128.880 89.095 129.605 ;
        RECT 89.730 128.865 89.985 129.435 ;
        RECT 90.155 129.205 90.485 129.605 ;
        RECT 90.910 129.070 91.440 129.435 ;
        RECT 90.910 129.035 91.085 129.070 ;
        RECT 90.155 128.865 91.085 129.035 ;
        RECT 87.515 127.225 87.685 127.985 ;
        RECT 87.865 127.055 88.195 127.815 ;
        RECT 88.365 127.225 88.635 128.130 ;
        RECT 88.805 127.055 89.095 128.220 ;
        RECT 89.730 128.195 89.900 128.865 ;
        RECT 90.155 128.695 90.325 128.865 ;
        RECT 90.070 128.365 90.325 128.695 ;
        RECT 90.550 128.365 90.745 128.695 ;
        RECT 89.730 127.225 90.065 128.195 ;
        RECT 90.235 127.055 90.405 128.195 ;
        RECT 90.575 127.395 90.745 128.365 ;
        RECT 90.915 127.735 91.085 128.865 ;
        RECT 91.255 128.075 91.425 128.875 ;
        RECT 91.630 128.585 91.905 129.435 ;
        RECT 91.625 128.415 91.905 128.585 ;
        RECT 91.630 128.275 91.905 128.415 ;
        RECT 92.075 128.075 92.265 129.435 ;
        RECT 92.445 129.070 92.955 129.605 ;
        RECT 93.175 128.795 93.420 129.400 ;
        RECT 94.415 129.055 94.585 129.435 ;
        RECT 94.765 129.225 95.095 129.605 ;
        RECT 94.415 128.885 95.080 129.055 ;
        RECT 95.275 128.930 95.535 129.435 ;
        RECT 95.705 129.095 96.010 129.605 ;
        RECT 92.465 128.625 93.695 128.795 ;
        RECT 91.255 127.905 92.265 128.075 ;
        RECT 92.435 128.060 93.185 128.250 ;
        RECT 90.915 127.565 92.040 127.735 ;
        RECT 92.435 127.395 92.605 128.060 ;
        RECT 93.355 127.815 93.695 128.625 ;
        RECT 94.345 128.335 94.675 128.705 ;
        RECT 94.910 128.630 95.080 128.885 ;
        RECT 94.910 128.300 95.195 128.630 ;
        RECT 94.910 128.155 95.080 128.300 ;
        RECT 90.575 127.225 92.605 127.395 ;
        RECT 92.775 127.055 92.945 127.815 ;
        RECT 93.180 127.405 93.695 127.815 ;
        RECT 94.415 127.985 95.080 128.155 ;
        RECT 95.365 128.130 95.535 128.930 ;
        RECT 95.705 128.365 96.020 128.925 ;
        RECT 96.190 128.615 96.440 129.425 ;
        RECT 96.610 129.080 96.870 129.605 ;
        RECT 97.050 128.615 97.300 129.425 ;
        RECT 97.470 129.045 97.730 129.605 ;
        RECT 97.900 128.955 98.160 129.410 ;
        RECT 98.330 129.125 98.590 129.605 ;
        RECT 98.760 128.955 99.020 129.410 ;
        RECT 99.190 129.125 99.450 129.605 ;
        RECT 99.620 128.955 99.880 129.410 ;
        RECT 100.050 129.125 100.295 129.605 ;
        RECT 100.465 128.955 100.740 129.410 ;
        RECT 100.910 129.125 101.155 129.605 ;
        RECT 101.325 128.955 101.585 129.410 ;
        RECT 101.765 129.125 102.015 129.605 ;
        RECT 102.185 128.955 102.445 129.410 ;
        RECT 102.625 129.125 102.875 129.605 ;
        RECT 103.045 128.955 103.305 129.410 ;
        RECT 103.485 129.125 103.745 129.605 ;
        RECT 103.915 128.955 104.175 129.410 ;
        RECT 104.345 129.125 104.645 129.605 ;
        RECT 104.905 129.145 105.465 129.435 ;
        RECT 105.635 129.145 105.885 129.605 ;
        RECT 97.900 128.785 104.645 128.955 ;
        RECT 96.190 128.365 103.310 128.615 ;
        RECT 94.415 127.225 94.585 127.985 ;
        RECT 94.765 127.055 95.095 127.815 ;
        RECT 95.265 127.225 95.535 128.130 ;
        RECT 95.715 127.055 96.010 127.865 ;
        RECT 96.190 127.225 96.435 128.365 ;
        RECT 96.610 127.055 96.870 127.865 ;
        RECT 97.050 127.230 97.300 128.365 ;
        RECT 103.480 128.195 104.645 128.785 ;
        RECT 97.900 127.970 104.645 128.195 ;
        RECT 97.900 127.955 103.305 127.970 ;
        RECT 97.470 127.060 97.730 127.855 ;
        RECT 97.900 127.230 98.160 127.955 ;
        RECT 98.330 127.060 98.590 127.785 ;
        RECT 98.760 127.230 99.020 127.955 ;
        RECT 99.190 127.060 99.450 127.785 ;
        RECT 99.620 127.230 99.880 127.955 ;
        RECT 100.050 127.060 100.310 127.785 ;
        RECT 100.480 127.230 100.740 127.955 ;
        RECT 100.910 127.060 101.155 127.785 ;
        RECT 101.325 127.230 101.585 127.955 ;
        RECT 101.770 127.060 102.015 127.785 ;
        RECT 102.185 127.230 102.445 127.955 ;
        RECT 102.630 127.060 102.875 127.785 ;
        RECT 103.045 127.230 103.305 127.955 ;
        RECT 103.490 127.060 103.745 127.785 ;
        RECT 103.915 127.230 104.205 127.970 ;
        RECT 97.470 127.055 103.745 127.060 ;
        RECT 104.375 127.055 104.645 127.800 ;
        RECT 104.905 127.775 105.155 129.145 ;
        RECT 106.505 128.975 106.835 129.335 ;
        RECT 105.445 128.785 106.835 128.975 ;
        RECT 107.205 129.145 107.765 129.435 ;
        RECT 107.935 129.145 108.185 129.605 ;
        RECT 105.445 128.695 105.615 128.785 ;
        RECT 105.325 128.365 105.615 128.695 ;
        RECT 105.785 128.365 106.125 128.615 ;
        RECT 106.345 128.365 107.020 128.615 ;
        RECT 105.445 128.115 105.615 128.365 ;
        RECT 105.445 127.945 106.385 128.115 ;
        RECT 106.755 128.005 107.020 128.365 ;
        RECT 104.905 127.225 105.365 127.775 ;
        RECT 105.555 127.055 105.885 127.775 ;
        RECT 106.085 127.395 106.385 127.945 ;
        RECT 107.205 127.775 107.455 129.145 ;
        RECT 108.805 128.975 109.135 129.335 ;
        RECT 107.745 128.785 109.135 128.975 ;
        RECT 109.705 128.975 110.035 129.335 ;
        RECT 110.655 129.145 110.905 129.605 ;
        RECT 111.075 129.145 111.635 129.435 ;
        RECT 109.705 128.785 111.095 128.975 ;
        RECT 107.745 128.695 107.915 128.785 ;
        RECT 107.625 128.365 107.915 128.695 ;
        RECT 110.925 128.695 111.095 128.785 ;
        RECT 108.085 128.365 108.425 128.615 ;
        RECT 108.645 128.365 109.320 128.615 ;
        RECT 107.745 128.115 107.915 128.365 ;
        RECT 107.745 127.945 108.685 128.115 ;
        RECT 109.055 128.005 109.320 128.365 ;
        RECT 109.520 128.365 110.195 128.615 ;
        RECT 110.415 128.365 110.755 128.615 ;
        RECT 110.925 128.365 111.215 128.695 ;
        RECT 109.520 128.005 109.785 128.365 ;
        RECT 110.925 128.115 111.095 128.365 ;
        RECT 106.555 127.055 106.835 127.725 ;
        RECT 107.205 127.225 107.665 127.775 ;
        RECT 107.855 127.055 108.185 127.775 ;
        RECT 108.385 127.395 108.685 127.945 ;
        RECT 110.155 127.945 111.095 128.115 ;
        RECT 108.855 127.055 109.135 127.725 ;
        RECT 109.705 127.055 109.985 127.725 ;
        RECT 110.155 127.395 110.455 127.945 ;
        RECT 111.385 127.775 111.635 129.145 ;
        RECT 110.655 127.055 110.985 127.775 ;
        RECT 111.175 127.225 111.635 127.775 ;
        RECT 111.805 129.145 112.365 129.435 ;
        RECT 112.535 129.145 112.785 129.605 ;
        RECT 111.805 127.775 112.055 129.145 ;
        RECT 113.405 128.975 113.735 129.335 ;
        RECT 112.345 128.785 113.735 128.975 ;
        RECT 114.565 128.880 114.855 129.605 ;
        RECT 115.485 128.835 118.075 129.605 ;
        RECT 112.345 128.695 112.515 128.785 ;
        RECT 112.225 128.365 112.515 128.695 ;
        RECT 112.685 128.365 113.025 128.615 ;
        RECT 113.245 128.365 113.920 128.615 ;
        RECT 112.345 128.115 112.515 128.365 ;
        RECT 112.345 127.945 113.285 128.115 ;
        RECT 113.655 128.005 113.920 128.365 ;
        RECT 111.805 127.225 112.265 127.775 ;
        RECT 112.455 127.055 112.785 127.775 ;
        RECT 112.985 127.395 113.285 127.945 ;
        RECT 113.455 127.055 113.735 127.725 ;
        RECT 114.565 127.055 114.855 128.220 ;
        RECT 115.485 128.145 116.695 128.665 ;
        RECT 116.865 128.315 118.075 128.835 ;
        RECT 118.285 128.785 118.515 129.605 ;
        RECT 118.685 128.805 119.015 129.435 ;
        RECT 118.265 128.365 118.595 128.615 ;
        RECT 118.765 128.205 119.015 128.805 ;
        RECT 119.185 128.785 119.395 129.605 ;
        RECT 119.715 129.055 119.885 129.435 ;
        RECT 120.065 129.225 120.395 129.605 ;
        RECT 119.715 128.885 120.380 129.055 ;
        RECT 120.575 128.930 120.835 129.435 ;
        RECT 121.010 129.060 126.355 129.605 ;
        RECT 119.645 128.335 119.975 128.705 ;
        RECT 120.210 128.630 120.380 128.885 ;
        RECT 115.485 127.055 118.075 128.145 ;
        RECT 118.285 127.055 118.515 128.195 ;
        RECT 118.685 127.225 119.015 128.205 ;
        RECT 120.210 128.300 120.495 128.630 ;
        RECT 119.185 127.055 119.395 128.195 ;
        RECT 120.210 128.155 120.380 128.300 ;
        RECT 119.715 127.985 120.380 128.155 ;
        RECT 120.665 128.130 120.835 128.930 ;
        RECT 119.715 127.225 119.885 127.985 ;
        RECT 120.065 127.055 120.395 127.815 ;
        RECT 120.565 127.225 120.835 128.130 ;
        RECT 122.600 127.490 122.950 128.740 ;
        RECT 124.430 128.230 124.770 129.060 ;
        RECT 126.525 128.855 127.735 129.605 ;
        RECT 126.525 128.145 127.045 128.685 ;
        RECT 127.215 128.315 127.735 128.855 ;
        RECT 121.010 127.055 126.355 127.490 ;
        RECT 126.525 127.055 127.735 128.145 ;
        RECT 14.660 126.885 127.820 127.055 ;
        RECT 14.745 125.795 15.955 126.885 ;
        RECT 14.745 125.085 15.265 125.625 ;
        RECT 15.435 125.255 15.955 125.795 ;
        RECT 16.125 125.795 17.335 126.885 ;
        RECT 17.505 125.795 21.015 126.885 ;
        RECT 16.125 125.255 16.645 125.795 ;
        RECT 16.815 125.085 17.335 125.625 ;
        RECT 17.505 125.275 19.195 125.795 ;
        RECT 21.245 125.745 21.455 126.885 ;
        RECT 21.625 125.735 21.955 126.715 ;
        RECT 22.125 125.745 22.355 126.885 ;
        RECT 23.115 125.955 23.285 126.715 ;
        RECT 23.465 126.125 23.795 126.885 ;
        RECT 23.115 125.785 23.780 125.955 ;
        RECT 23.965 125.810 24.235 126.715 ;
        RECT 19.365 125.105 21.015 125.625 ;
        RECT 14.745 124.335 15.955 125.085 ;
        RECT 16.125 124.335 17.335 125.085 ;
        RECT 17.505 124.335 21.015 125.105 ;
        RECT 21.245 124.335 21.455 125.155 ;
        RECT 21.625 125.135 21.875 125.735 ;
        RECT 23.610 125.640 23.780 125.785 ;
        RECT 22.045 125.325 22.375 125.575 ;
        RECT 23.045 125.235 23.375 125.605 ;
        RECT 23.610 125.310 23.895 125.640 ;
        RECT 21.625 124.505 21.955 125.135 ;
        RECT 22.125 124.335 22.355 125.155 ;
        RECT 23.610 125.055 23.780 125.310 ;
        RECT 23.115 124.885 23.780 125.055 ;
        RECT 24.065 125.010 24.235 125.810 ;
        RECT 24.405 125.720 24.695 126.885 ;
        RECT 25.790 126.450 31.135 126.885 ;
        RECT 31.310 126.450 36.655 126.885 ;
        RECT 27.380 125.200 27.730 126.450 ;
        RECT 23.115 124.505 23.285 124.885 ;
        RECT 23.465 124.335 23.795 124.715 ;
        RECT 23.975 124.505 24.235 125.010 ;
        RECT 24.405 124.335 24.695 125.060 ;
        RECT 29.210 124.880 29.550 125.710 ;
        RECT 32.900 125.200 33.250 126.450 ;
        RECT 37.025 126.215 37.305 126.885 ;
        RECT 37.475 125.995 37.775 126.545 ;
        RECT 37.975 126.165 38.305 126.885 ;
        RECT 38.495 126.165 38.955 126.715 ;
        RECT 34.730 124.880 35.070 125.710 ;
        RECT 36.840 125.575 37.105 125.935 ;
        RECT 37.475 125.825 38.415 125.995 ;
        RECT 38.245 125.575 38.415 125.825 ;
        RECT 36.840 125.325 37.515 125.575 ;
        RECT 37.735 125.325 38.075 125.575 ;
        RECT 38.245 125.245 38.535 125.575 ;
        RECT 38.245 125.155 38.415 125.245 ;
        RECT 37.025 124.965 38.415 125.155 ;
        RECT 25.790 124.335 31.135 124.880 ;
        RECT 31.310 124.335 36.655 124.880 ;
        RECT 37.025 124.605 37.355 124.965 ;
        RECT 38.705 124.795 38.955 126.165 ;
        RECT 39.125 125.795 40.335 126.885 ;
        RECT 40.505 126.165 40.965 126.715 ;
        RECT 41.155 126.165 41.485 126.885 ;
        RECT 39.125 125.255 39.645 125.795 ;
        RECT 39.815 125.085 40.335 125.625 ;
        RECT 37.975 124.335 38.225 124.795 ;
        RECT 38.395 124.505 38.955 124.795 ;
        RECT 39.125 124.335 40.335 125.085 ;
        RECT 40.505 124.795 40.755 126.165 ;
        RECT 41.685 125.995 41.985 126.545 ;
        RECT 42.155 126.215 42.435 126.885 ;
        RECT 43.005 126.215 43.285 126.885 ;
        RECT 41.045 125.825 41.985 125.995 ;
        RECT 43.455 125.995 43.755 126.545 ;
        RECT 43.955 126.165 44.285 126.885 ;
        RECT 44.475 126.165 44.935 126.715 ;
        RECT 41.045 125.575 41.215 125.825 ;
        RECT 42.355 125.575 42.620 125.935 ;
        RECT 40.925 125.245 41.215 125.575 ;
        RECT 41.385 125.325 41.725 125.575 ;
        RECT 41.945 125.325 42.620 125.575 ;
        RECT 42.820 125.575 43.085 125.935 ;
        RECT 43.455 125.825 44.395 125.995 ;
        RECT 44.225 125.575 44.395 125.825 ;
        RECT 42.820 125.325 43.495 125.575 ;
        RECT 43.715 125.325 44.055 125.575 ;
        RECT 41.045 125.155 41.215 125.245 ;
        RECT 44.225 125.245 44.515 125.575 ;
        RECT 44.225 125.155 44.395 125.245 ;
        RECT 41.045 124.965 42.435 125.155 ;
        RECT 40.505 124.505 41.065 124.795 ;
        RECT 41.235 124.335 41.485 124.795 ;
        RECT 42.105 124.605 42.435 124.965 ;
        RECT 43.005 124.965 44.395 125.155 ;
        RECT 43.005 124.605 43.335 124.965 ;
        RECT 44.685 124.795 44.935 126.165 ;
        RECT 43.955 124.335 44.205 124.795 ;
        RECT 44.375 124.505 44.935 124.795 ;
        RECT 45.105 126.165 45.565 126.715 ;
        RECT 45.755 126.165 46.085 126.885 ;
        RECT 45.105 124.795 45.355 126.165 ;
        RECT 46.285 125.995 46.585 126.545 ;
        RECT 46.755 126.215 47.035 126.885 ;
        RECT 47.460 126.015 47.745 126.885 ;
        RECT 47.915 126.255 48.175 126.715 ;
        RECT 48.350 126.425 48.605 126.885 ;
        RECT 48.775 126.255 49.035 126.715 ;
        RECT 47.915 126.085 49.035 126.255 ;
        RECT 49.205 126.085 49.515 126.885 ;
        RECT 45.645 125.825 46.585 125.995 ;
        RECT 45.645 125.575 45.815 125.825 ;
        RECT 46.955 125.575 47.220 125.935 ;
        RECT 47.915 125.835 48.175 126.085 ;
        RECT 49.685 125.915 49.995 126.715 ;
        RECT 45.525 125.245 45.815 125.575 ;
        RECT 45.985 125.325 46.325 125.575 ;
        RECT 46.545 125.325 47.220 125.575 ;
        RECT 47.420 125.665 48.175 125.835 ;
        RECT 48.965 125.745 49.995 125.915 ;
        RECT 45.645 125.155 45.815 125.245 ;
        RECT 47.420 125.155 47.825 125.665 ;
        RECT 48.965 125.495 49.135 125.745 ;
        RECT 47.995 125.325 49.135 125.495 ;
        RECT 45.645 124.965 47.035 125.155 ;
        RECT 47.420 124.985 49.070 125.155 ;
        RECT 49.305 125.005 49.655 125.575 ;
        RECT 45.105 124.505 45.665 124.795 ;
        RECT 45.835 124.335 46.085 124.795 ;
        RECT 46.705 124.605 47.035 124.965 ;
        RECT 47.465 124.335 47.745 124.815 ;
        RECT 47.915 124.595 48.175 124.985 ;
        RECT 48.350 124.335 48.605 124.815 ;
        RECT 48.775 124.595 49.070 124.985 ;
        RECT 49.825 124.835 49.995 125.745 ;
        RECT 50.165 125.720 50.455 126.885 ;
        RECT 50.625 125.795 52.295 126.885 ;
        RECT 52.470 126.450 57.815 126.885 ;
        RECT 50.625 125.275 51.375 125.795 ;
        RECT 51.545 125.105 52.295 125.625 ;
        RECT 54.060 125.200 54.410 126.450 ;
        RECT 58.075 125.955 58.245 126.715 ;
        RECT 58.425 126.125 58.755 126.885 ;
        RECT 58.075 125.785 58.740 125.955 ;
        RECT 58.925 125.810 59.195 126.715 ;
        RECT 49.250 124.335 49.525 124.815 ;
        RECT 49.695 124.505 49.995 124.835 ;
        RECT 50.165 124.335 50.455 125.060 ;
        RECT 50.625 124.335 52.295 125.105 ;
        RECT 55.890 124.880 56.230 125.710 ;
        RECT 58.570 125.640 58.740 125.785 ;
        RECT 58.005 125.235 58.335 125.605 ;
        RECT 58.570 125.310 58.855 125.640 ;
        RECT 58.570 125.055 58.740 125.310 ;
        RECT 58.075 124.885 58.740 125.055 ;
        RECT 59.025 125.010 59.195 125.810 ;
        RECT 59.365 126.125 59.880 126.535 ;
        RECT 60.115 126.125 60.285 126.885 ;
        RECT 60.455 126.545 62.485 126.715 ;
        RECT 59.365 125.315 59.705 126.125 ;
        RECT 60.455 125.880 60.625 126.545 ;
        RECT 61.020 126.205 62.145 126.375 ;
        RECT 59.875 125.690 60.625 125.880 ;
        RECT 60.795 125.865 61.805 126.035 ;
        RECT 59.365 125.145 60.595 125.315 ;
        RECT 52.470 124.335 57.815 124.880 ;
        RECT 58.075 124.505 58.245 124.885 ;
        RECT 58.425 124.335 58.755 124.715 ;
        RECT 58.935 124.505 59.195 125.010 ;
        RECT 59.640 124.540 59.885 125.145 ;
        RECT 60.105 124.335 60.615 124.870 ;
        RECT 60.795 124.505 60.985 125.865 ;
        RECT 61.155 125.525 61.430 125.665 ;
        RECT 61.155 125.355 61.435 125.525 ;
        RECT 61.155 124.505 61.430 125.355 ;
        RECT 61.635 125.065 61.805 125.865 ;
        RECT 61.975 125.075 62.145 126.205 ;
        RECT 62.315 125.575 62.485 126.545 ;
        RECT 62.655 125.745 62.825 126.885 ;
        RECT 62.995 125.745 63.330 126.715 ;
        RECT 62.315 125.245 62.510 125.575 ;
        RECT 62.735 125.245 62.990 125.575 ;
        RECT 62.735 125.075 62.905 125.245 ;
        RECT 63.160 125.075 63.330 125.745 ;
        RECT 63.505 125.795 64.715 126.885 ;
        RECT 64.885 125.795 68.395 126.885 ;
        RECT 63.505 125.255 64.025 125.795 ;
        RECT 64.195 125.085 64.715 125.625 ;
        RECT 64.885 125.275 66.575 125.795 ;
        RECT 68.625 125.745 68.835 126.885 ;
        RECT 69.005 125.735 69.335 126.715 ;
        RECT 69.505 125.745 69.735 126.885 ;
        RECT 70.495 125.955 70.665 126.715 ;
        RECT 70.845 126.125 71.175 126.885 ;
        RECT 70.495 125.785 71.160 125.955 ;
        RECT 71.345 125.810 71.615 126.715 ;
        RECT 66.745 125.105 68.395 125.625 ;
        RECT 61.975 124.905 62.905 125.075 ;
        RECT 61.975 124.870 62.150 124.905 ;
        RECT 61.620 124.505 62.150 124.870 ;
        RECT 62.575 124.335 62.905 124.735 ;
        RECT 63.075 124.505 63.330 125.075 ;
        RECT 63.505 124.335 64.715 125.085 ;
        RECT 64.885 124.335 68.395 125.105 ;
        RECT 68.625 124.335 68.835 125.155 ;
        RECT 69.005 125.135 69.255 125.735 ;
        RECT 70.990 125.640 71.160 125.785 ;
        RECT 69.425 125.325 69.755 125.575 ;
        RECT 70.425 125.235 70.755 125.605 ;
        RECT 70.990 125.310 71.275 125.640 ;
        RECT 69.005 124.505 69.335 125.135 ;
        RECT 69.505 124.335 69.735 125.155 ;
        RECT 70.990 125.055 71.160 125.310 ;
        RECT 70.495 124.885 71.160 125.055 ;
        RECT 71.445 125.010 71.615 125.810 ;
        RECT 70.495 124.505 70.665 124.885 ;
        RECT 70.845 124.335 71.175 124.715 ;
        RECT 71.355 124.505 71.615 125.010 ;
        RECT 72.705 125.915 73.015 126.715 ;
        RECT 73.185 126.085 73.495 126.885 ;
        RECT 73.665 126.255 73.925 126.715 ;
        RECT 74.095 126.425 74.350 126.885 ;
        RECT 74.525 126.255 74.785 126.715 ;
        RECT 73.665 126.085 74.785 126.255 ;
        RECT 72.705 125.745 73.735 125.915 ;
        RECT 72.705 124.835 72.875 125.745 ;
        RECT 73.045 125.005 73.395 125.575 ;
        RECT 73.565 125.495 73.735 125.745 ;
        RECT 74.525 125.835 74.785 126.085 ;
        RECT 74.955 126.015 75.240 126.885 ;
        RECT 74.525 125.665 75.280 125.835 ;
        RECT 75.925 125.720 76.215 126.885 ;
        RECT 76.385 125.795 78.055 126.885 ;
        RECT 78.600 126.545 78.855 126.575 ;
        RECT 78.515 126.375 78.855 126.545 ;
        RECT 78.600 125.905 78.855 126.375 ;
        RECT 79.035 126.085 79.320 126.885 ;
        RECT 79.500 126.165 79.830 126.675 ;
        RECT 73.565 125.325 74.705 125.495 ;
        RECT 74.875 125.155 75.280 125.665 ;
        RECT 76.385 125.275 77.135 125.795 ;
        RECT 73.630 124.985 75.280 125.155 ;
        RECT 77.305 125.105 78.055 125.625 ;
        RECT 72.705 124.505 73.005 124.835 ;
        RECT 73.175 124.335 73.450 124.815 ;
        RECT 73.630 124.595 73.925 124.985 ;
        RECT 74.095 124.335 74.350 124.815 ;
        RECT 74.525 124.595 74.785 124.985 ;
        RECT 74.955 124.335 75.235 124.815 ;
        RECT 75.925 124.335 76.215 125.060 ;
        RECT 76.385 124.335 78.055 125.105 ;
        RECT 78.600 125.045 78.780 125.905 ;
        RECT 79.500 125.575 79.750 126.165 ;
        RECT 80.100 126.015 80.270 126.625 ;
        RECT 80.440 126.195 80.770 126.885 ;
        RECT 81.000 126.335 81.240 126.625 ;
        RECT 81.440 126.505 81.860 126.885 ;
        RECT 82.040 126.415 82.670 126.665 ;
        RECT 83.140 126.505 83.470 126.885 ;
        RECT 82.040 126.335 82.210 126.415 ;
        RECT 83.640 126.335 83.810 126.625 ;
        RECT 83.990 126.505 84.370 126.885 ;
        RECT 84.610 126.500 85.440 126.670 ;
        RECT 81.000 126.165 82.210 126.335 ;
        RECT 78.950 125.245 79.750 125.575 ;
        RECT 78.600 124.515 78.855 125.045 ;
        RECT 79.035 124.335 79.320 124.795 ;
        RECT 79.500 124.595 79.750 125.245 ;
        RECT 79.950 125.995 80.270 126.015 ;
        RECT 79.950 125.825 81.870 125.995 ;
        RECT 79.950 124.930 80.140 125.825 ;
        RECT 82.040 125.655 82.210 126.165 ;
        RECT 82.380 125.905 82.900 126.215 ;
        RECT 80.310 125.485 82.210 125.655 ;
        RECT 80.310 125.425 80.640 125.485 ;
        RECT 80.790 125.255 81.120 125.315 ;
        RECT 80.460 124.985 81.120 125.255 ;
        RECT 79.950 124.600 80.270 124.930 ;
        RECT 80.450 124.335 81.110 124.815 ;
        RECT 81.310 124.725 81.480 125.485 ;
        RECT 82.380 125.315 82.560 125.725 ;
        RECT 81.650 125.145 81.980 125.265 ;
        RECT 82.730 125.145 82.900 125.905 ;
        RECT 81.650 124.975 82.900 125.145 ;
        RECT 83.070 126.085 84.440 126.335 ;
        RECT 83.070 125.315 83.260 126.085 ;
        RECT 84.190 125.825 84.440 126.085 ;
        RECT 83.430 125.655 83.680 125.815 ;
        RECT 84.610 125.655 84.780 126.500 ;
        RECT 85.675 126.215 85.845 126.715 ;
        RECT 86.015 126.385 86.345 126.885 ;
        RECT 84.950 125.825 85.450 126.205 ;
        RECT 85.675 126.045 86.370 126.215 ;
        RECT 83.430 125.485 84.780 125.655 ;
        RECT 84.360 125.445 84.780 125.485 ;
        RECT 83.070 124.975 83.490 125.315 ;
        RECT 83.780 124.985 84.190 125.315 ;
        RECT 81.310 124.555 82.160 124.725 ;
        RECT 82.720 124.335 83.040 124.795 ;
        RECT 83.240 124.545 83.490 124.975 ;
        RECT 83.780 124.335 84.190 124.775 ;
        RECT 84.360 124.715 84.530 125.445 ;
        RECT 84.700 124.895 85.050 125.265 ;
        RECT 85.230 124.955 85.450 125.825 ;
        RECT 85.620 125.255 86.030 125.875 ;
        RECT 86.200 125.075 86.370 126.045 ;
        RECT 85.675 124.885 86.370 125.075 ;
        RECT 84.360 124.515 85.375 124.715 ;
        RECT 85.675 124.555 85.845 124.885 ;
        RECT 86.015 124.335 86.345 124.715 ;
        RECT 86.560 124.595 86.785 126.715 ;
        RECT 86.955 126.385 87.285 126.885 ;
        RECT 87.455 126.215 87.625 126.715 ;
        RECT 86.960 126.045 87.625 126.215 ;
        RECT 86.960 125.055 87.190 126.045 ;
        RECT 87.360 125.225 87.710 125.875 ;
        RECT 87.885 125.795 89.555 126.885 ;
        RECT 89.815 126.215 89.985 126.715 ;
        RECT 90.155 126.385 90.485 126.885 ;
        RECT 89.815 126.045 90.480 126.215 ;
        RECT 87.885 125.275 88.635 125.795 ;
        RECT 88.805 125.105 89.555 125.625 ;
        RECT 89.730 125.225 90.080 125.875 ;
        RECT 86.960 124.885 87.625 125.055 ;
        RECT 86.955 124.335 87.285 124.715 ;
        RECT 87.455 124.595 87.625 124.885 ;
        RECT 87.885 124.335 89.555 125.105 ;
        RECT 90.250 125.055 90.480 126.045 ;
        RECT 89.815 124.885 90.480 125.055 ;
        RECT 89.815 124.595 89.985 124.885 ;
        RECT 90.155 124.335 90.485 124.715 ;
        RECT 90.655 124.595 90.880 126.715 ;
        RECT 91.095 126.385 91.425 126.885 ;
        RECT 91.595 126.215 91.765 126.715 ;
        RECT 92.000 126.500 92.830 126.670 ;
        RECT 93.070 126.505 93.450 126.885 ;
        RECT 91.070 126.045 91.765 126.215 ;
        RECT 91.070 125.075 91.240 126.045 ;
        RECT 91.410 125.255 91.820 125.875 ;
        RECT 91.990 125.825 92.490 126.205 ;
        RECT 91.070 124.885 91.765 125.075 ;
        RECT 91.990 124.955 92.210 125.825 ;
        RECT 92.660 125.655 92.830 126.500 ;
        RECT 93.630 126.335 93.800 126.625 ;
        RECT 93.970 126.505 94.300 126.885 ;
        RECT 94.770 126.415 95.400 126.665 ;
        RECT 95.580 126.505 96.000 126.885 ;
        RECT 95.230 126.335 95.400 126.415 ;
        RECT 96.200 126.335 96.440 126.625 ;
        RECT 93.000 126.085 94.370 126.335 ;
        RECT 93.000 125.825 93.250 126.085 ;
        RECT 93.760 125.655 94.010 125.815 ;
        RECT 92.660 125.485 94.010 125.655 ;
        RECT 92.660 125.445 93.080 125.485 ;
        RECT 92.390 124.895 92.740 125.265 ;
        RECT 91.095 124.335 91.425 124.715 ;
        RECT 91.595 124.555 91.765 124.885 ;
        RECT 92.910 124.715 93.080 125.445 ;
        RECT 94.180 125.315 94.370 126.085 ;
        RECT 93.250 124.985 93.660 125.315 ;
        RECT 93.950 124.975 94.370 125.315 ;
        RECT 94.540 125.905 95.060 126.215 ;
        RECT 95.230 126.165 96.440 126.335 ;
        RECT 96.670 126.195 97.000 126.885 ;
        RECT 94.540 125.145 94.710 125.905 ;
        RECT 94.880 125.315 95.060 125.725 ;
        RECT 95.230 125.655 95.400 126.165 ;
        RECT 97.170 126.015 97.340 126.625 ;
        RECT 97.610 126.165 97.940 126.675 ;
        RECT 97.170 125.995 97.490 126.015 ;
        RECT 95.570 125.825 97.490 125.995 ;
        RECT 95.230 125.485 97.130 125.655 ;
        RECT 95.460 125.145 95.790 125.265 ;
        RECT 94.540 124.975 95.790 125.145 ;
        RECT 92.065 124.515 93.080 124.715 ;
        RECT 93.250 124.335 93.660 124.775 ;
        RECT 93.950 124.545 94.200 124.975 ;
        RECT 94.400 124.335 94.720 124.795 ;
        RECT 95.960 124.725 96.130 125.485 ;
        RECT 96.800 125.425 97.130 125.485 ;
        RECT 96.320 125.255 96.650 125.315 ;
        RECT 96.320 124.985 96.980 125.255 ;
        RECT 97.300 124.930 97.490 125.825 ;
        RECT 95.280 124.555 96.130 124.725 ;
        RECT 96.330 124.335 96.990 124.815 ;
        RECT 97.170 124.600 97.490 124.930 ;
        RECT 97.690 125.575 97.940 126.165 ;
        RECT 98.120 126.085 98.405 126.885 ;
        RECT 98.585 126.545 98.840 126.575 ;
        RECT 98.585 126.375 98.925 126.545 ;
        RECT 98.585 125.905 98.840 126.375 ;
        RECT 99.585 126.215 99.865 126.885 ;
        RECT 100.035 125.995 100.335 126.545 ;
        RECT 100.535 126.165 100.865 126.885 ;
        RECT 101.055 126.165 101.515 126.715 ;
        RECT 97.690 125.245 98.490 125.575 ;
        RECT 97.690 124.595 97.940 125.245 ;
        RECT 98.660 125.045 98.840 125.905 ;
        RECT 99.400 125.575 99.665 125.935 ;
        RECT 100.035 125.825 100.975 125.995 ;
        RECT 100.805 125.575 100.975 125.825 ;
        RECT 99.400 125.325 100.075 125.575 ;
        RECT 100.295 125.325 100.635 125.575 ;
        RECT 100.805 125.245 101.095 125.575 ;
        RECT 100.805 125.155 100.975 125.245 ;
        RECT 98.120 124.335 98.405 124.795 ;
        RECT 98.585 124.515 98.840 125.045 ;
        RECT 99.585 124.965 100.975 125.155 ;
        RECT 99.585 124.605 99.915 124.965 ;
        RECT 101.265 124.795 101.515 126.165 ;
        RECT 101.685 125.720 101.975 126.885 ;
        RECT 102.145 125.795 105.655 126.885 ;
        RECT 105.830 126.450 111.175 126.885 ;
        RECT 102.145 125.275 103.835 125.795 ;
        RECT 104.005 125.105 105.655 125.625 ;
        RECT 107.420 125.200 107.770 126.450 ;
        RECT 111.345 126.125 111.860 126.535 ;
        RECT 112.095 126.125 112.265 126.885 ;
        RECT 112.435 126.545 114.465 126.715 ;
        RECT 100.535 124.335 100.785 124.795 ;
        RECT 100.955 124.505 101.515 124.795 ;
        RECT 101.685 124.335 101.975 125.060 ;
        RECT 102.145 124.335 105.655 125.105 ;
        RECT 109.250 124.880 109.590 125.710 ;
        RECT 111.345 125.315 111.685 126.125 ;
        RECT 112.435 125.880 112.605 126.545 ;
        RECT 113.000 126.205 114.125 126.375 ;
        RECT 111.855 125.690 112.605 125.880 ;
        RECT 112.775 125.865 113.785 126.035 ;
        RECT 111.345 125.145 112.575 125.315 ;
        RECT 105.830 124.335 111.175 124.880 ;
        RECT 111.620 124.540 111.865 125.145 ;
        RECT 112.085 124.335 112.595 124.870 ;
        RECT 112.775 124.505 112.965 125.865 ;
        RECT 113.135 124.845 113.410 125.665 ;
        RECT 113.615 125.065 113.785 125.865 ;
        RECT 113.955 125.075 114.125 126.205 ;
        RECT 114.295 125.575 114.465 126.545 ;
        RECT 114.635 125.745 114.805 126.885 ;
        RECT 114.975 125.745 115.310 126.715 ;
        RECT 114.295 125.245 114.490 125.575 ;
        RECT 114.715 125.245 114.970 125.575 ;
        RECT 114.715 125.075 114.885 125.245 ;
        RECT 115.140 125.075 115.310 125.745 ;
        RECT 113.955 124.905 114.885 125.075 ;
        RECT 113.955 124.870 114.130 124.905 ;
        RECT 113.135 124.675 113.415 124.845 ;
        RECT 113.135 124.505 113.410 124.675 ;
        RECT 113.600 124.505 114.130 124.870 ;
        RECT 114.555 124.335 114.885 124.735 ;
        RECT 115.055 124.505 115.310 125.075 ;
        RECT 115.860 125.905 116.115 126.575 ;
        RECT 116.295 126.085 116.580 126.885 ;
        RECT 116.760 126.165 117.090 126.675 ;
        RECT 115.860 125.045 116.040 125.905 ;
        RECT 116.760 125.575 117.010 126.165 ;
        RECT 117.360 126.015 117.530 126.625 ;
        RECT 117.700 126.195 118.030 126.885 ;
        RECT 118.260 126.335 118.500 126.625 ;
        RECT 118.700 126.505 119.120 126.885 ;
        RECT 119.300 126.415 119.930 126.665 ;
        RECT 120.400 126.505 120.730 126.885 ;
        RECT 119.300 126.335 119.470 126.415 ;
        RECT 120.900 126.335 121.070 126.625 ;
        RECT 121.250 126.505 121.630 126.885 ;
        RECT 121.870 126.500 122.700 126.670 ;
        RECT 118.260 126.165 119.470 126.335 ;
        RECT 116.210 125.245 117.010 125.575 ;
        RECT 115.860 124.845 116.115 125.045 ;
        RECT 115.775 124.675 116.115 124.845 ;
        RECT 115.860 124.515 116.115 124.675 ;
        RECT 116.295 124.335 116.580 124.795 ;
        RECT 116.760 124.595 117.010 125.245 ;
        RECT 117.210 125.995 117.530 126.015 ;
        RECT 117.210 125.825 119.130 125.995 ;
        RECT 117.210 124.930 117.400 125.825 ;
        RECT 119.300 125.655 119.470 126.165 ;
        RECT 119.640 125.905 120.160 126.215 ;
        RECT 117.570 125.485 119.470 125.655 ;
        RECT 117.570 125.425 117.900 125.485 ;
        RECT 118.050 125.255 118.380 125.315 ;
        RECT 117.720 124.985 118.380 125.255 ;
        RECT 117.210 124.600 117.530 124.930 ;
        RECT 117.710 124.335 118.370 124.815 ;
        RECT 118.570 124.725 118.740 125.485 ;
        RECT 119.640 125.315 119.820 125.725 ;
        RECT 118.910 125.145 119.240 125.265 ;
        RECT 119.990 125.145 120.160 125.905 ;
        RECT 118.910 124.975 120.160 125.145 ;
        RECT 120.330 126.085 121.700 126.335 ;
        RECT 120.330 125.315 120.520 126.085 ;
        RECT 121.450 125.825 121.700 126.085 ;
        RECT 120.690 125.655 120.940 125.815 ;
        RECT 121.870 125.655 122.040 126.500 ;
        RECT 122.935 126.215 123.105 126.715 ;
        RECT 123.275 126.385 123.605 126.885 ;
        RECT 122.210 125.825 122.710 126.205 ;
        RECT 122.935 126.045 123.630 126.215 ;
        RECT 120.690 125.485 122.040 125.655 ;
        RECT 121.620 125.445 122.040 125.485 ;
        RECT 120.330 124.975 120.750 125.315 ;
        RECT 121.040 124.985 121.450 125.315 ;
        RECT 118.570 124.555 119.420 124.725 ;
        RECT 119.980 124.335 120.300 124.795 ;
        RECT 120.500 124.545 120.750 124.975 ;
        RECT 121.040 124.335 121.450 124.775 ;
        RECT 121.620 124.715 121.790 125.445 ;
        RECT 121.960 124.895 122.310 125.265 ;
        RECT 122.490 124.955 122.710 125.825 ;
        RECT 122.880 125.255 123.290 125.875 ;
        RECT 123.460 125.075 123.630 126.045 ;
        RECT 122.935 124.885 123.630 125.075 ;
        RECT 121.620 124.515 122.635 124.715 ;
        RECT 122.935 124.555 123.105 124.885 ;
        RECT 123.275 124.335 123.605 124.715 ;
        RECT 123.820 124.595 124.045 126.715 ;
        RECT 124.215 126.385 124.545 126.885 ;
        RECT 124.715 126.215 124.885 126.715 ;
        RECT 124.220 126.045 124.885 126.215 ;
        RECT 124.220 125.055 124.450 126.045 ;
        RECT 124.620 125.225 124.970 125.875 ;
        RECT 125.145 125.795 126.355 126.885 ;
        RECT 126.525 125.795 127.735 126.885 ;
        RECT 125.145 125.255 125.665 125.795 ;
        RECT 125.835 125.085 126.355 125.625 ;
        RECT 126.525 125.255 127.045 125.795 ;
        RECT 127.215 125.085 127.735 125.625 ;
        RECT 124.220 124.885 124.885 125.055 ;
        RECT 124.215 124.335 124.545 124.715 ;
        RECT 124.715 124.595 124.885 124.885 ;
        RECT 125.145 124.335 126.355 125.085 ;
        RECT 126.525 124.335 127.735 125.085 ;
        RECT 14.660 124.165 127.820 124.335 ;
        RECT 14.745 123.415 15.955 124.165 ;
        RECT 16.125 123.415 17.335 124.165 ;
        RECT 17.510 123.620 22.855 124.165 ;
        RECT 14.745 122.875 15.265 123.415 ;
        RECT 15.435 122.705 15.955 123.245 ;
        RECT 14.745 121.615 15.955 122.705 ;
        RECT 16.125 122.705 16.645 123.245 ;
        RECT 16.815 122.875 17.335 123.415 ;
        RECT 16.125 121.615 17.335 122.705 ;
        RECT 19.100 122.050 19.450 123.300 ;
        RECT 20.930 122.790 21.270 123.620 ;
        RECT 23.300 123.355 23.545 123.960 ;
        RECT 23.765 123.630 24.275 124.165 ;
        RECT 23.025 123.185 24.255 123.355 ;
        RECT 23.025 122.375 23.365 123.185 ;
        RECT 23.535 122.620 24.285 122.810 ;
        RECT 17.510 121.615 22.855 122.050 ;
        RECT 23.025 121.965 23.540 122.375 ;
        RECT 23.775 121.615 23.945 122.375 ;
        RECT 24.115 121.955 24.285 122.620 ;
        RECT 24.455 122.635 24.645 123.995 ;
        RECT 24.815 123.825 25.090 123.995 ;
        RECT 24.815 123.655 25.095 123.825 ;
        RECT 24.815 122.835 25.090 123.655 ;
        RECT 25.280 123.630 25.810 123.995 ;
        RECT 26.235 123.765 26.565 124.165 ;
        RECT 25.635 123.595 25.810 123.630 ;
        RECT 25.295 122.635 25.465 123.435 ;
        RECT 24.455 122.465 25.465 122.635 ;
        RECT 25.635 123.425 26.565 123.595 ;
        RECT 26.735 123.425 26.990 123.995 ;
        RECT 27.630 123.620 32.975 124.165 ;
        RECT 25.635 122.295 25.805 123.425 ;
        RECT 26.395 123.255 26.565 123.425 ;
        RECT 24.680 122.125 25.805 122.295 ;
        RECT 25.975 122.925 26.170 123.255 ;
        RECT 26.395 122.925 26.650 123.255 ;
        RECT 25.975 121.955 26.145 122.925 ;
        RECT 26.820 122.755 26.990 123.425 ;
        RECT 24.115 121.785 26.145 121.955 ;
        RECT 26.315 121.615 26.485 122.755 ;
        RECT 26.655 121.785 26.990 122.755 ;
        RECT 29.220 122.050 29.570 123.300 ;
        RECT 31.050 122.790 31.390 123.620 ;
        RECT 33.420 123.355 33.665 123.960 ;
        RECT 33.885 123.630 34.395 124.165 ;
        RECT 33.145 123.185 34.375 123.355 ;
        RECT 33.145 122.375 33.485 123.185 ;
        RECT 33.655 122.620 34.405 122.810 ;
        RECT 27.630 121.615 32.975 122.050 ;
        RECT 33.145 121.965 33.660 122.375 ;
        RECT 33.895 121.615 34.065 122.375 ;
        RECT 34.235 121.955 34.405 122.620 ;
        RECT 34.575 122.635 34.765 123.995 ;
        RECT 34.935 123.145 35.210 123.995 ;
        RECT 35.400 123.630 35.930 123.995 ;
        RECT 36.355 123.765 36.685 124.165 ;
        RECT 35.755 123.595 35.930 123.630 ;
        RECT 34.935 122.975 35.215 123.145 ;
        RECT 34.935 122.835 35.210 122.975 ;
        RECT 35.415 122.635 35.585 123.435 ;
        RECT 34.575 122.465 35.585 122.635 ;
        RECT 35.755 123.425 36.685 123.595 ;
        RECT 36.855 123.425 37.110 123.995 ;
        RECT 37.285 123.440 37.575 124.165 ;
        RECT 35.755 122.295 35.925 123.425 ;
        RECT 36.515 123.255 36.685 123.425 ;
        RECT 34.800 122.125 35.925 122.295 ;
        RECT 36.095 122.925 36.290 123.255 ;
        RECT 36.515 122.925 36.770 123.255 ;
        RECT 36.095 121.955 36.265 122.925 ;
        RECT 36.940 122.755 37.110 123.425 ;
        RECT 38.205 123.395 41.715 124.165 ;
        RECT 41.890 123.620 47.235 124.165 ;
        RECT 47.410 123.620 52.755 124.165 ;
        RECT 53.300 123.825 53.555 123.985 ;
        RECT 53.215 123.655 53.555 123.825 ;
        RECT 53.735 123.705 54.020 124.165 ;
        RECT 34.235 121.785 36.265 121.955 ;
        RECT 36.435 121.615 36.605 122.755 ;
        RECT 36.775 121.785 37.110 122.755 ;
        RECT 37.285 121.615 37.575 122.780 ;
        RECT 38.205 122.705 39.895 123.225 ;
        RECT 40.065 122.875 41.715 123.395 ;
        RECT 38.205 121.615 41.715 122.705 ;
        RECT 43.480 122.050 43.830 123.300 ;
        RECT 45.310 122.790 45.650 123.620 ;
        RECT 49.000 122.050 49.350 123.300 ;
        RECT 50.830 122.790 51.170 123.620 ;
        RECT 53.300 123.455 53.555 123.655 ;
        RECT 53.300 122.595 53.480 123.455 ;
        RECT 54.200 123.255 54.450 123.905 ;
        RECT 53.650 122.925 54.450 123.255 ;
        RECT 41.890 121.615 47.235 122.050 ;
        RECT 47.410 121.615 52.755 122.050 ;
        RECT 53.300 121.925 53.555 122.595 ;
        RECT 53.735 121.615 54.020 122.415 ;
        RECT 54.200 122.335 54.450 122.925 ;
        RECT 54.650 123.570 54.970 123.900 ;
        RECT 55.150 123.685 55.810 124.165 ;
        RECT 56.010 123.775 56.860 123.945 ;
        RECT 54.650 122.675 54.840 123.570 ;
        RECT 55.160 123.245 55.820 123.515 ;
        RECT 55.490 123.185 55.820 123.245 ;
        RECT 55.010 123.015 55.340 123.075 ;
        RECT 56.010 123.015 56.180 123.775 ;
        RECT 57.420 123.705 57.740 124.165 ;
        RECT 57.940 123.525 58.190 123.955 ;
        RECT 58.480 123.725 58.890 124.165 ;
        RECT 59.060 123.785 60.075 123.985 ;
        RECT 56.350 123.355 57.600 123.525 ;
        RECT 56.350 123.235 56.680 123.355 ;
        RECT 55.010 122.845 56.910 123.015 ;
        RECT 54.650 122.505 56.570 122.675 ;
        RECT 54.650 122.485 54.970 122.505 ;
        RECT 54.200 121.825 54.530 122.335 ;
        RECT 54.800 121.875 54.970 122.485 ;
        RECT 56.740 122.335 56.910 122.845 ;
        RECT 57.080 122.775 57.260 123.185 ;
        RECT 57.430 122.595 57.600 123.355 ;
        RECT 55.140 121.615 55.470 122.305 ;
        RECT 55.700 122.165 56.910 122.335 ;
        RECT 57.080 122.285 57.600 122.595 ;
        RECT 57.770 123.185 58.190 123.525 ;
        RECT 58.480 123.185 58.890 123.515 ;
        RECT 57.770 122.415 57.960 123.185 ;
        RECT 59.060 123.055 59.230 123.785 ;
        RECT 60.375 123.615 60.545 123.945 ;
        RECT 60.715 123.785 61.045 124.165 ;
        RECT 59.400 123.235 59.750 123.605 ;
        RECT 59.060 123.015 59.480 123.055 ;
        RECT 58.130 122.845 59.480 123.015 ;
        RECT 58.130 122.685 58.380 122.845 ;
        RECT 58.890 122.415 59.140 122.675 ;
        RECT 57.770 122.165 59.140 122.415 ;
        RECT 55.700 121.875 55.940 122.165 ;
        RECT 56.740 122.085 56.910 122.165 ;
        RECT 56.140 121.615 56.560 121.995 ;
        RECT 56.740 121.835 57.370 122.085 ;
        RECT 57.840 121.615 58.170 121.995 ;
        RECT 58.340 121.875 58.510 122.165 ;
        RECT 59.310 122.000 59.480 122.845 ;
        RECT 59.930 122.675 60.150 123.545 ;
        RECT 60.375 123.425 61.070 123.615 ;
        RECT 59.650 122.295 60.150 122.675 ;
        RECT 60.320 122.625 60.730 123.245 ;
        RECT 60.900 122.455 61.070 123.425 ;
        RECT 60.375 122.285 61.070 122.455 ;
        RECT 58.690 121.615 59.070 121.995 ;
        RECT 59.310 121.830 60.140 122.000 ;
        RECT 60.375 121.785 60.545 122.285 ;
        RECT 60.715 121.615 61.045 122.115 ;
        RECT 61.260 121.785 61.485 123.905 ;
        RECT 61.655 123.785 61.985 124.165 ;
        RECT 62.155 123.615 62.325 123.905 ;
        RECT 61.660 123.445 62.325 123.615 ;
        RECT 61.660 122.455 61.890 123.445 ;
        RECT 63.045 123.440 63.335 124.165 ;
        RECT 64.240 123.355 64.485 123.960 ;
        RECT 64.705 123.630 65.215 124.165 ;
        RECT 62.060 122.625 62.410 123.275 ;
        RECT 63.965 123.185 65.195 123.355 ;
        RECT 61.660 122.285 62.325 122.455 ;
        RECT 61.655 121.615 61.985 122.115 ;
        RECT 62.155 121.785 62.325 122.285 ;
        RECT 63.045 121.615 63.335 122.780 ;
        RECT 63.965 122.375 64.305 123.185 ;
        RECT 64.475 122.620 65.225 122.810 ;
        RECT 63.965 121.965 64.480 122.375 ;
        RECT 64.715 121.615 64.885 122.375 ;
        RECT 65.055 121.955 65.225 122.620 ;
        RECT 65.395 122.635 65.585 123.995 ;
        RECT 65.755 123.825 66.030 123.995 ;
        RECT 65.755 123.655 66.035 123.825 ;
        RECT 65.755 122.835 66.030 123.655 ;
        RECT 66.220 123.630 66.750 123.995 ;
        RECT 67.175 123.765 67.505 124.165 ;
        RECT 66.575 123.595 66.750 123.630 ;
        RECT 66.235 122.635 66.405 123.435 ;
        RECT 65.395 122.465 66.405 122.635 ;
        RECT 66.575 123.425 67.505 123.595 ;
        RECT 67.675 123.425 67.930 123.995 ;
        RECT 66.575 122.295 66.745 123.425 ;
        RECT 67.335 123.255 67.505 123.425 ;
        RECT 65.620 122.125 66.745 122.295 ;
        RECT 66.915 122.925 67.110 123.255 ;
        RECT 67.335 122.925 67.590 123.255 ;
        RECT 66.915 121.955 67.085 122.925 ;
        RECT 67.760 122.755 67.930 123.425 ;
        RECT 68.105 123.395 70.695 124.165 ;
        RECT 70.870 123.620 76.215 124.165 ;
        RECT 76.390 123.620 81.735 124.165 ;
        RECT 65.055 121.785 67.085 121.955 ;
        RECT 67.255 121.615 67.425 122.755 ;
        RECT 67.595 121.785 67.930 122.755 ;
        RECT 68.105 122.705 69.315 123.225 ;
        RECT 69.485 122.875 70.695 123.395 ;
        RECT 68.105 121.615 70.695 122.705 ;
        RECT 72.460 122.050 72.810 123.300 ;
        RECT 74.290 122.790 74.630 123.620 ;
        RECT 77.980 122.050 78.330 123.300 ;
        RECT 79.810 122.790 80.150 123.620 ;
        RECT 81.965 123.345 82.175 124.165 ;
        RECT 82.345 123.365 82.675 123.995 ;
        RECT 82.345 122.765 82.595 123.365 ;
        RECT 82.845 123.345 83.075 124.165 ;
        RECT 83.835 123.615 84.005 123.995 ;
        RECT 84.185 123.785 84.515 124.165 ;
        RECT 83.835 123.445 84.500 123.615 ;
        RECT 84.695 123.490 84.955 123.995 ;
        RECT 82.765 122.925 83.095 123.175 ;
        RECT 83.765 122.895 84.095 123.265 ;
        RECT 84.330 123.190 84.500 123.445 ;
        RECT 84.330 122.860 84.615 123.190 ;
        RECT 70.870 121.615 76.215 122.050 ;
        RECT 76.390 121.615 81.735 122.050 ;
        RECT 81.965 121.615 82.175 122.755 ;
        RECT 82.345 121.785 82.675 122.765 ;
        RECT 82.845 121.615 83.075 122.755 ;
        RECT 84.330 122.715 84.500 122.860 ;
        RECT 83.835 122.545 84.500 122.715 ;
        RECT 84.785 122.690 84.955 123.490 ;
        RECT 85.125 123.395 88.635 124.165 ;
        RECT 88.805 123.440 89.095 124.165 ;
        RECT 89.265 123.395 92.775 124.165 ;
        RECT 83.835 121.785 84.005 122.545 ;
        RECT 84.185 121.615 84.515 122.375 ;
        RECT 84.685 121.785 84.955 122.690 ;
        RECT 85.125 122.705 86.815 123.225 ;
        RECT 86.985 122.875 88.635 123.395 ;
        RECT 85.125 121.615 88.635 122.705 ;
        RECT 88.805 121.615 89.095 122.780 ;
        RECT 89.265 122.705 90.955 123.225 ;
        RECT 91.125 122.875 92.775 123.395 ;
        RECT 92.985 123.345 93.215 124.165 ;
        RECT 93.385 123.365 93.715 123.995 ;
        RECT 92.965 122.925 93.295 123.175 ;
        RECT 93.465 122.765 93.715 123.365 ;
        RECT 93.885 123.345 94.095 124.165 ;
        RECT 94.325 123.415 95.535 124.165 ;
        RECT 89.265 121.615 92.775 122.705 ;
        RECT 92.985 121.615 93.215 122.755 ;
        RECT 93.385 121.785 93.715 122.765 ;
        RECT 93.885 121.615 94.095 122.755 ;
        RECT 94.325 122.705 94.845 123.245 ;
        RECT 95.015 122.875 95.535 123.415 ;
        RECT 95.705 123.395 99.215 124.165 ;
        RECT 99.390 123.620 104.735 124.165 ;
        RECT 104.910 123.620 110.255 124.165 ;
        RECT 95.705 122.705 97.395 123.225 ;
        RECT 97.565 122.875 99.215 123.395 ;
        RECT 94.325 121.615 95.535 122.705 ;
        RECT 95.705 121.615 99.215 122.705 ;
        RECT 100.980 122.050 101.330 123.300 ;
        RECT 102.810 122.790 103.150 123.620 ;
        RECT 106.500 122.050 106.850 123.300 ;
        RECT 108.330 122.790 108.670 123.620 ;
        RECT 110.700 123.355 110.945 123.960 ;
        RECT 111.165 123.630 111.675 124.165 ;
        RECT 110.425 123.185 111.655 123.355 ;
        RECT 110.425 122.375 110.765 123.185 ;
        RECT 110.935 122.620 111.685 122.810 ;
        RECT 99.390 121.615 104.735 122.050 ;
        RECT 104.910 121.615 110.255 122.050 ;
        RECT 110.425 121.965 110.940 122.375 ;
        RECT 111.175 121.615 111.345 122.375 ;
        RECT 111.515 121.955 111.685 122.620 ;
        RECT 111.855 122.635 112.045 123.995 ;
        RECT 112.215 123.145 112.490 123.995 ;
        RECT 112.680 123.630 113.210 123.995 ;
        RECT 113.635 123.765 113.965 124.165 ;
        RECT 113.035 123.595 113.210 123.630 ;
        RECT 112.215 122.975 112.495 123.145 ;
        RECT 112.215 122.835 112.490 122.975 ;
        RECT 112.695 122.635 112.865 123.435 ;
        RECT 111.855 122.465 112.865 122.635 ;
        RECT 113.035 123.425 113.965 123.595 ;
        RECT 114.135 123.425 114.390 123.995 ;
        RECT 114.565 123.440 114.855 124.165 ;
        RECT 115.860 123.455 116.115 123.985 ;
        RECT 116.295 123.705 116.580 124.165 ;
        RECT 113.035 122.295 113.205 123.425 ;
        RECT 113.795 123.255 113.965 123.425 ;
        RECT 112.080 122.125 113.205 122.295 ;
        RECT 113.375 122.925 113.570 123.255 ;
        RECT 113.795 122.925 114.050 123.255 ;
        RECT 113.375 121.955 113.545 122.925 ;
        RECT 114.220 122.755 114.390 123.425 ;
        RECT 115.860 123.145 116.040 123.455 ;
        RECT 116.760 123.255 117.010 123.905 ;
        RECT 115.775 122.975 116.040 123.145 ;
        RECT 111.515 121.785 113.545 121.955 ;
        RECT 113.715 121.615 113.885 122.755 ;
        RECT 114.055 121.785 114.390 122.755 ;
        RECT 114.565 121.615 114.855 122.780 ;
        RECT 115.860 122.595 116.040 122.975 ;
        RECT 116.210 122.925 117.010 123.255 ;
        RECT 115.860 121.925 116.115 122.595 ;
        RECT 116.295 121.615 116.580 122.415 ;
        RECT 116.760 122.335 117.010 122.925 ;
        RECT 117.210 123.570 117.530 123.900 ;
        RECT 117.710 123.685 118.370 124.165 ;
        RECT 118.570 123.775 119.420 123.945 ;
        RECT 117.210 122.675 117.400 123.570 ;
        RECT 117.720 123.245 118.380 123.515 ;
        RECT 118.050 123.185 118.380 123.245 ;
        RECT 117.570 123.015 117.900 123.075 ;
        RECT 118.570 123.015 118.740 123.775 ;
        RECT 119.980 123.705 120.300 124.165 ;
        RECT 120.500 123.525 120.750 123.955 ;
        RECT 121.040 123.725 121.450 124.165 ;
        RECT 121.620 123.785 122.635 123.985 ;
        RECT 118.910 123.355 120.160 123.525 ;
        RECT 118.910 123.235 119.240 123.355 ;
        RECT 117.570 122.845 119.470 123.015 ;
        RECT 117.210 122.505 119.130 122.675 ;
        RECT 117.210 122.485 117.530 122.505 ;
        RECT 116.760 121.825 117.090 122.335 ;
        RECT 117.360 121.875 117.530 122.485 ;
        RECT 119.300 122.335 119.470 122.845 ;
        RECT 119.640 122.775 119.820 123.185 ;
        RECT 119.990 122.595 120.160 123.355 ;
        RECT 117.700 121.615 118.030 122.305 ;
        RECT 118.260 122.165 119.470 122.335 ;
        RECT 119.640 122.285 120.160 122.595 ;
        RECT 120.330 123.185 120.750 123.525 ;
        RECT 121.040 123.185 121.450 123.515 ;
        RECT 120.330 122.415 120.520 123.185 ;
        RECT 121.620 123.055 121.790 123.785 ;
        RECT 122.935 123.615 123.105 123.945 ;
        RECT 123.275 123.785 123.605 124.165 ;
        RECT 121.960 123.235 122.310 123.605 ;
        RECT 121.620 123.015 122.040 123.055 ;
        RECT 120.690 122.845 122.040 123.015 ;
        RECT 120.690 122.685 120.940 122.845 ;
        RECT 121.450 122.415 121.700 122.675 ;
        RECT 120.330 122.165 121.700 122.415 ;
        RECT 118.260 121.875 118.500 122.165 ;
        RECT 119.300 122.085 119.470 122.165 ;
        RECT 118.700 121.615 119.120 121.995 ;
        RECT 119.300 121.835 119.930 122.085 ;
        RECT 120.400 121.615 120.730 121.995 ;
        RECT 120.900 121.875 121.070 122.165 ;
        RECT 121.870 122.000 122.040 122.845 ;
        RECT 122.490 122.675 122.710 123.545 ;
        RECT 122.935 123.425 123.630 123.615 ;
        RECT 122.210 122.295 122.710 122.675 ;
        RECT 122.880 122.625 123.290 123.245 ;
        RECT 123.460 122.455 123.630 123.425 ;
        RECT 122.935 122.285 123.630 122.455 ;
        RECT 121.250 121.615 121.630 121.995 ;
        RECT 121.870 121.830 122.700 122.000 ;
        RECT 122.935 121.785 123.105 122.285 ;
        RECT 123.275 121.615 123.605 122.115 ;
        RECT 123.820 121.785 124.045 123.905 ;
        RECT 124.215 123.785 124.545 124.165 ;
        RECT 124.715 123.615 124.885 123.905 ;
        RECT 124.220 123.445 124.885 123.615 ;
        RECT 124.220 122.455 124.450 123.445 ;
        RECT 125.145 123.415 126.355 124.165 ;
        RECT 126.525 123.415 127.735 124.165 ;
        RECT 124.620 122.625 124.970 123.275 ;
        RECT 125.145 122.705 125.665 123.245 ;
        RECT 125.835 122.875 126.355 123.415 ;
        RECT 126.525 122.705 127.045 123.245 ;
        RECT 127.215 122.875 127.735 123.415 ;
        RECT 124.220 122.285 124.885 122.455 ;
        RECT 124.215 121.615 124.545 122.115 ;
        RECT 124.715 121.785 124.885 122.285 ;
        RECT 125.145 121.615 126.355 122.705 ;
        RECT 126.525 121.615 127.735 122.705 ;
        RECT 14.660 121.445 127.820 121.615 ;
        RECT 14.745 120.355 15.955 121.445 ;
        RECT 14.745 119.645 15.265 120.185 ;
        RECT 15.435 119.815 15.955 120.355 ;
        RECT 16.585 120.355 20.095 121.445 ;
        RECT 16.585 119.835 18.275 120.355 ;
        RECT 20.270 120.305 20.605 121.275 ;
        RECT 20.775 120.305 20.945 121.445 ;
        RECT 21.115 121.105 23.145 121.275 ;
        RECT 18.445 119.665 20.095 120.185 ;
        RECT 14.745 118.895 15.955 119.645 ;
        RECT 16.585 118.895 20.095 119.665 ;
        RECT 20.270 119.635 20.440 120.305 ;
        RECT 21.115 120.135 21.285 121.105 ;
        RECT 20.610 119.805 20.865 120.135 ;
        RECT 21.090 119.805 21.285 120.135 ;
        RECT 21.455 120.765 22.580 120.935 ;
        RECT 20.695 119.635 20.865 119.805 ;
        RECT 21.455 119.635 21.625 120.765 ;
        RECT 20.270 119.065 20.525 119.635 ;
        RECT 20.695 119.465 21.625 119.635 ;
        RECT 21.795 120.425 22.805 120.595 ;
        RECT 21.795 119.625 21.965 120.425 ;
        RECT 22.170 119.745 22.445 120.225 ;
        RECT 22.165 119.575 22.445 119.745 ;
        RECT 21.450 119.430 21.625 119.465 ;
        RECT 20.695 118.895 21.025 119.295 ;
        RECT 21.450 119.065 21.980 119.430 ;
        RECT 22.170 119.065 22.445 119.575 ;
        RECT 22.615 119.065 22.805 120.425 ;
        RECT 22.975 120.440 23.145 121.105 ;
        RECT 23.315 120.685 23.485 121.445 ;
        RECT 23.720 120.685 24.235 121.095 ;
        RECT 22.975 120.250 23.725 120.440 ;
        RECT 23.895 119.875 24.235 120.685 ;
        RECT 24.405 120.280 24.695 121.445 ;
        RECT 24.865 120.355 26.075 121.445 ;
        RECT 26.245 120.370 26.515 121.275 ;
        RECT 26.685 120.685 27.015 121.445 ;
        RECT 27.195 120.515 27.365 121.275 ;
        RECT 23.005 119.705 24.235 119.875 ;
        RECT 24.865 119.815 25.385 120.355 ;
        RECT 22.985 118.895 23.495 119.430 ;
        RECT 23.715 119.100 23.960 119.705 ;
        RECT 25.555 119.645 26.075 120.185 ;
        RECT 24.405 118.895 24.695 119.620 ;
        RECT 24.865 118.895 26.075 119.645 ;
        RECT 26.245 119.570 26.415 120.370 ;
        RECT 26.700 120.345 27.365 120.515 ;
        RECT 27.625 120.355 30.215 121.445 ;
        RECT 30.760 121.105 31.015 121.135 ;
        RECT 30.675 120.935 31.015 121.105 ;
        RECT 30.760 120.465 31.015 120.935 ;
        RECT 31.195 120.645 31.480 121.445 ;
        RECT 31.660 120.725 31.990 121.235 ;
        RECT 26.700 120.200 26.870 120.345 ;
        RECT 26.585 119.870 26.870 120.200 ;
        RECT 26.700 119.615 26.870 119.870 ;
        RECT 27.105 119.795 27.435 120.165 ;
        RECT 27.625 119.835 28.835 120.355 ;
        RECT 29.005 119.665 30.215 120.185 ;
        RECT 26.245 119.065 26.505 119.570 ;
        RECT 26.700 119.445 27.365 119.615 ;
        RECT 26.685 118.895 27.015 119.275 ;
        RECT 27.195 119.065 27.365 119.445 ;
        RECT 27.625 118.895 30.215 119.665 ;
        RECT 30.760 119.605 30.940 120.465 ;
        RECT 31.660 120.135 31.910 120.725 ;
        RECT 32.260 120.575 32.430 121.185 ;
        RECT 32.600 120.755 32.930 121.445 ;
        RECT 33.160 120.895 33.400 121.185 ;
        RECT 33.600 121.065 34.020 121.445 ;
        RECT 34.200 120.975 34.830 121.225 ;
        RECT 35.300 121.065 35.630 121.445 ;
        RECT 34.200 120.895 34.370 120.975 ;
        RECT 35.800 120.895 35.970 121.185 ;
        RECT 36.150 121.065 36.530 121.445 ;
        RECT 36.770 121.060 37.600 121.230 ;
        RECT 33.160 120.725 34.370 120.895 ;
        RECT 31.110 119.805 31.910 120.135 ;
        RECT 30.760 119.075 31.015 119.605 ;
        RECT 31.195 118.895 31.480 119.355 ;
        RECT 31.660 119.155 31.910 119.805 ;
        RECT 32.110 120.555 32.430 120.575 ;
        RECT 32.110 120.385 34.030 120.555 ;
        RECT 32.110 119.490 32.300 120.385 ;
        RECT 34.200 120.215 34.370 120.725 ;
        RECT 34.540 120.465 35.060 120.775 ;
        RECT 32.470 120.045 34.370 120.215 ;
        RECT 32.470 119.985 32.800 120.045 ;
        RECT 32.950 119.815 33.280 119.875 ;
        RECT 32.620 119.545 33.280 119.815 ;
        RECT 32.110 119.160 32.430 119.490 ;
        RECT 32.610 118.895 33.270 119.375 ;
        RECT 33.470 119.285 33.640 120.045 ;
        RECT 34.540 119.875 34.720 120.285 ;
        RECT 33.810 119.705 34.140 119.825 ;
        RECT 34.890 119.705 35.060 120.465 ;
        RECT 33.810 119.535 35.060 119.705 ;
        RECT 35.230 120.645 36.600 120.895 ;
        RECT 35.230 119.875 35.420 120.645 ;
        RECT 36.350 120.385 36.600 120.645 ;
        RECT 35.590 120.215 35.840 120.375 ;
        RECT 36.770 120.215 36.940 121.060 ;
        RECT 37.835 120.775 38.005 121.275 ;
        RECT 38.175 120.945 38.505 121.445 ;
        RECT 37.110 120.385 37.610 120.765 ;
        RECT 37.835 120.605 38.530 120.775 ;
        RECT 35.590 120.045 36.940 120.215 ;
        RECT 36.520 120.005 36.940 120.045 ;
        RECT 35.230 119.535 35.650 119.875 ;
        RECT 35.940 119.545 36.350 119.875 ;
        RECT 33.470 119.115 34.320 119.285 ;
        RECT 34.880 118.895 35.200 119.355 ;
        RECT 35.400 119.105 35.650 119.535 ;
        RECT 35.940 118.895 36.350 119.335 ;
        RECT 36.520 119.275 36.690 120.005 ;
        RECT 36.860 119.455 37.210 119.825 ;
        RECT 37.390 119.515 37.610 120.385 ;
        RECT 37.780 119.815 38.190 120.435 ;
        RECT 38.360 119.635 38.530 120.605 ;
        RECT 37.835 119.445 38.530 119.635 ;
        RECT 36.520 119.075 37.535 119.275 ;
        RECT 37.835 119.115 38.005 119.445 ;
        RECT 38.175 118.895 38.505 119.275 ;
        RECT 38.720 119.155 38.945 121.275 ;
        RECT 39.115 120.945 39.445 121.445 ;
        RECT 39.615 120.775 39.785 121.275 ;
        RECT 39.120 120.605 39.785 120.775 ;
        RECT 39.120 119.615 39.350 120.605 ;
        RECT 39.520 119.785 39.870 120.435 ;
        RECT 40.050 120.305 40.385 121.275 ;
        RECT 40.555 120.305 40.725 121.445 ;
        RECT 40.895 121.105 42.925 121.275 ;
        RECT 40.050 119.635 40.220 120.305 ;
        RECT 40.895 120.135 41.065 121.105 ;
        RECT 40.390 119.805 40.645 120.135 ;
        RECT 40.870 119.805 41.065 120.135 ;
        RECT 41.235 120.765 42.360 120.935 ;
        RECT 40.475 119.635 40.645 119.805 ;
        RECT 41.235 119.635 41.405 120.765 ;
        RECT 39.120 119.445 39.785 119.615 ;
        RECT 39.115 118.895 39.445 119.275 ;
        RECT 39.615 119.155 39.785 119.445 ;
        RECT 40.050 119.065 40.305 119.635 ;
        RECT 40.475 119.465 41.405 119.635 ;
        RECT 41.575 120.425 42.585 120.595 ;
        RECT 41.575 119.625 41.745 120.425 ;
        RECT 41.950 120.085 42.225 120.225 ;
        RECT 41.945 119.915 42.225 120.085 ;
        RECT 41.230 119.430 41.405 119.465 ;
        RECT 40.475 118.895 40.805 119.295 ;
        RECT 41.230 119.065 41.760 119.430 ;
        RECT 41.950 119.065 42.225 119.915 ;
        RECT 42.395 119.065 42.585 120.425 ;
        RECT 42.755 120.440 42.925 121.105 ;
        RECT 43.095 120.685 43.265 121.445 ;
        RECT 43.500 120.685 44.015 121.095 ;
        RECT 42.755 120.250 43.505 120.440 ;
        RECT 43.675 119.875 44.015 120.685 ;
        RECT 42.785 119.705 44.015 119.875 ;
        RECT 44.645 120.370 44.915 121.275 ;
        RECT 45.085 120.685 45.415 121.445 ;
        RECT 45.595 120.515 45.765 121.275 ;
        RECT 42.765 118.895 43.275 119.430 ;
        RECT 43.495 119.100 43.740 119.705 ;
        RECT 44.645 119.570 44.815 120.370 ;
        RECT 45.100 120.345 45.765 120.515 ;
        RECT 46.025 120.685 46.540 121.095 ;
        RECT 46.775 120.685 46.945 121.445 ;
        RECT 47.115 121.105 49.145 121.275 ;
        RECT 45.100 120.200 45.270 120.345 ;
        RECT 44.985 119.870 45.270 120.200 ;
        RECT 45.100 119.615 45.270 119.870 ;
        RECT 45.505 119.795 45.835 120.165 ;
        RECT 46.025 119.875 46.365 120.685 ;
        RECT 47.115 120.440 47.285 121.105 ;
        RECT 47.680 120.765 48.805 120.935 ;
        RECT 46.535 120.250 47.285 120.440 ;
        RECT 47.455 120.425 48.465 120.595 ;
        RECT 46.025 119.705 47.255 119.875 ;
        RECT 44.645 119.065 44.905 119.570 ;
        RECT 45.100 119.445 45.765 119.615 ;
        RECT 45.085 118.895 45.415 119.275 ;
        RECT 45.595 119.065 45.765 119.445 ;
        RECT 46.300 119.100 46.545 119.705 ;
        RECT 46.765 118.895 47.275 119.430 ;
        RECT 47.455 119.065 47.645 120.425 ;
        RECT 47.815 120.085 48.090 120.225 ;
        RECT 47.815 119.915 48.095 120.085 ;
        RECT 47.815 119.065 48.090 119.915 ;
        RECT 48.295 119.625 48.465 120.425 ;
        RECT 48.635 119.635 48.805 120.765 ;
        RECT 48.975 120.135 49.145 121.105 ;
        RECT 49.315 120.305 49.485 121.445 ;
        RECT 49.655 120.305 49.990 121.275 ;
        RECT 48.975 119.805 49.170 120.135 ;
        RECT 49.395 119.805 49.650 120.135 ;
        RECT 49.395 119.635 49.565 119.805 ;
        RECT 49.820 119.635 49.990 120.305 ;
        RECT 50.165 120.280 50.455 121.445 ;
        RECT 50.665 120.305 50.895 121.445 ;
        RECT 51.065 120.295 51.395 121.275 ;
        RECT 51.565 120.305 51.775 121.445 ;
        RECT 52.005 120.355 53.215 121.445 ;
        RECT 50.645 119.885 50.975 120.135 ;
        RECT 48.635 119.465 49.565 119.635 ;
        RECT 48.635 119.430 48.810 119.465 ;
        RECT 48.280 119.065 48.810 119.430 ;
        RECT 49.235 118.895 49.565 119.295 ;
        RECT 49.735 119.065 49.990 119.635 ;
        RECT 50.165 118.895 50.455 119.620 ;
        RECT 50.665 118.895 50.895 119.715 ;
        RECT 51.145 119.695 51.395 120.295 ;
        RECT 52.005 119.815 52.525 120.355 ;
        RECT 53.535 120.295 53.865 121.445 ;
        RECT 54.035 120.425 54.205 121.275 ;
        RECT 54.375 120.645 54.705 121.445 ;
        RECT 54.875 120.425 55.045 121.275 ;
        RECT 55.225 120.645 55.465 121.445 ;
        RECT 55.635 120.465 55.965 121.275 ;
        RECT 54.035 120.255 55.045 120.425 ;
        RECT 55.250 120.295 55.965 120.465 ;
        RECT 57.125 120.305 57.335 121.445 ;
        RECT 57.505 120.295 57.835 121.275 ;
        RECT 58.005 120.305 58.235 121.445 ;
        RECT 59.740 121.105 59.995 121.135 ;
        RECT 59.655 120.935 59.995 121.105 ;
        RECT 59.740 120.465 59.995 120.935 ;
        RECT 60.175 120.645 60.460 121.445 ;
        RECT 60.640 120.725 60.970 121.235 ;
        RECT 51.065 119.065 51.395 119.695 ;
        RECT 51.565 118.895 51.775 119.715 ;
        RECT 52.695 119.645 53.215 120.185 ;
        RECT 54.035 120.085 54.530 120.255 ;
        RECT 54.035 119.915 54.535 120.085 ;
        RECT 55.250 120.055 55.420 120.295 ;
        RECT 54.035 119.715 54.530 119.915 ;
        RECT 54.920 119.885 55.420 120.055 ;
        RECT 55.590 119.885 55.970 120.125 ;
        RECT 55.250 119.715 55.420 119.885 ;
        RECT 52.005 118.895 53.215 119.645 ;
        RECT 53.535 118.895 53.865 119.695 ;
        RECT 54.035 119.545 55.045 119.715 ;
        RECT 55.250 119.545 55.885 119.715 ;
        RECT 54.035 119.065 54.205 119.545 ;
        RECT 54.375 118.895 54.705 119.375 ;
        RECT 54.875 119.065 55.045 119.545 ;
        RECT 55.295 118.895 55.535 119.375 ;
        RECT 55.715 119.065 55.885 119.545 ;
        RECT 57.125 118.895 57.335 119.715 ;
        RECT 57.505 119.695 57.755 120.295 ;
        RECT 57.925 119.885 58.255 120.135 ;
        RECT 57.505 119.065 57.835 119.695 ;
        RECT 58.005 118.895 58.235 119.715 ;
        RECT 59.740 119.605 59.920 120.465 ;
        RECT 60.640 120.135 60.890 120.725 ;
        RECT 61.240 120.575 61.410 121.185 ;
        RECT 61.580 120.755 61.910 121.445 ;
        RECT 62.140 120.895 62.380 121.185 ;
        RECT 62.580 121.065 63.000 121.445 ;
        RECT 63.180 120.975 63.810 121.225 ;
        RECT 64.280 121.065 64.610 121.445 ;
        RECT 63.180 120.895 63.350 120.975 ;
        RECT 64.780 120.895 64.950 121.185 ;
        RECT 65.130 121.065 65.510 121.445 ;
        RECT 65.750 121.060 66.580 121.230 ;
        RECT 62.140 120.725 63.350 120.895 ;
        RECT 60.090 119.805 60.890 120.135 ;
        RECT 59.740 119.075 59.995 119.605 ;
        RECT 60.175 118.895 60.460 119.355 ;
        RECT 60.640 119.155 60.890 119.805 ;
        RECT 61.090 120.555 61.410 120.575 ;
        RECT 61.090 120.385 63.010 120.555 ;
        RECT 61.090 119.490 61.280 120.385 ;
        RECT 63.180 120.215 63.350 120.725 ;
        RECT 63.520 120.465 64.040 120.775 ;
        RECT 61.450 120.045 63.350 120.215 ;
        RECT 61.450 119.985 61.780 120.045 ;
        RECT 61.930 119.815 62.260 119.875 ;
        RECT 61.600 119.545 62.260 119.815 ;
        RECT 61.090 119.160 61.410 119.490 ;
        RECT 61.590 118.895 62.250 119.375 ;
        RECT 62.450 119.285 62.620 120.045 ;
        RECT 63.520 119.875 63.700 120.285 ;
        RECT 62.790 119.705 63.120 119.825 ;
        RECT 63.870 119.705 64.040 120.465 ;
        RECT 62.790 119.535 64.040 119.705 ;
        RECT 64.210 120.645 65.580 120.895 ;
        RECT 64.210 119.875 64.400 120.645 ;
        RECT 65.330 120.385 65.580 120.645 ;
        RECT 64.570 120.215 64.820 120.375 ;
        RECT 65.750 120.215 65.920 121.060 ;
        RECT 66.815 120.775 66.985 121.275 ;
        RECT 67.155 120.945 67.485 121.445 ;
        RECT 66.090 120.385 66.590 120.765 ;
        RECT 66.815 120.605 67.510 120.775 ;
        RECT 64.570 120.045 65.920 120.215 ;
        RECT 65.500 120.005 65.920 120.045 ;
        RECT 64.210 119.535 64.630 119.875 ;
        RECT 64.920 119.545 65.330 119.875 ;
        RECT 62.450 119.115 63.300 119.285 ;
        RECT 63.860 118.895 64.180 119.355 ;
        RECT 64.380 119.105 64.630 119.535 ;
        RECT 64.920 118.895 65.330 119.335 ;
        RECT 65.500 119.275 65.670 120.005 ;
        RECT 65.840 119.455 66.190 119.825 ;
        RECT 66.370 119.515 66.590 120.385 ;
        RECT 66.760 119.815 67.170 120.435 ;
        RECT 67.340 119.635 67.510 120.605 ;
        RECT 66.815 119.445 67.510 119.635 ;
        RECT 65.500 119.075 66.515 119.275 ;
        RECT 66.815 119.115 66.985 119.445 ;
        RECT 67.155 118.895 67.485 119.275 ;
        RECT 67.700 119.155 67.925 121.275 ;
        RECT 68.095 120.945 68.425 121.445 ;
        RECT 68.595 120.775 68.765 121.275 ;
        RECT 68.100 120.605 68.765 120.775 ;
        RECT 68.100 119.615 68.330 120.605 ;
        RECT 68.500 119.785 68.850 120.435 ;
        RECT 69.025 120.370 69.295 121.275 ;
        RECT 69.465 120.685 69.795 121.445 ;
        RECT 69.975 120.515 70.145 121.275 ;
        RECT 68.100 119.445 68.765 119.615 ;
        RECT 68.095 118.895 68.425 119.275 ;
        RECT 68.595 119.155 68.765 119.445 ;
        RECT 69.025 119.570 69.195 120.370 ;
        RECT 69.480 120.345 70.145 120.515 ;
        RECT 70.865 120.355 74.375 121.445 ;
        RECT 69.480 120.200 69.650 120.345 ;
        RECT 69.365 119.870 69.650 120.200 ;
        RECT 69.480 119.615 69.650 119.870 ;
        RECT 69.885 119.795 70.215 120.165 ;
        RECT 70.865 119.835 72.555 120.355 ;
        RECT 74.585 120.305 74.815 121.445 ;
        RECT 74.985 120.295 75.315 121.275 ;
        RECT 75.485 120.305 75.695 121.445 ;
        RECT 72.725 119.665 74.375 120.185 ;
        RECT 74.565 119.885 74.895 120.135 ;
        RECT 69.025 119.065 69.285 119.570 ;
        RECT 69.480 119.445 70.145 119.615 ;
        RECT 69.465 118.895 69.795 119.275 ;
        RECT 69.975 119.065 70.145 119.445 ;
        RECT 70.865 118.895 74.375 119.665 ;
        RECT 74.585 118.895 74.815 119.715 ;
        RECT 75.065 119.695 75.315 120.295 ;
        RECT 75.925 120.280 76.215 121.445 ;
        RECT 76.845 120.685 77.360 121.095 ;
        RECT 77.595 120.685 77.765 121.445 ;
        RECT 77.935 121.105 79.965 121.275 ;
        RECT 76.845 119.875 77.185 120.685 ;
        RECT 77.935 120.440 78.105 121.105 ;
        RECT 78.500 120.765 79.625 120.935 ;
        RECT 77.355 120.250 78.105 120.440 ;
        RECT 78.275 120.425 79.285 120.595 ;
        RECT 74.985 119.065 75.315 119.695 ;
        RECT 75.485 118.895 75.695 119.715 ;
        RECT 76.845 119.705 78.075 119.875 ;
        RECT 75.925 118.895 76.215 119.620 ;
        RECT 77.120 119.100 77.365 119.705 ;
        RECT 77.585 118.895 78.095 119.430 ;
        RECT 78.275 119.065 78.465 120.425 ;
        RECT 78.635 119.405 78.910 120.225 ;
        RECT 79.115 119.625 79.285 120.425 ;
        RECT 79.455 119.635 79.625 120.765 ;
        RECT 79.795 120.135 79.965 121.105 ;
        RECT 80.135 120.305 80.305 121.445 ;
        RECT 80.475 120.305 80.810 121.275 ;
        RECT 79.795 119.805 79.990 120.135 ;
        RECT 80.215 119.805 80.470 120.135 ;
        RECT 80.215 119.635 80.385 119.805 ;
        RECT 80.640 119.635 80.810 120.305 ;
        RECT 79.455 119.465 80.385 119.635 ;
        RECT 79.455 119.430 79.630 119.465 ;
        RECT 78.635 119.235 78.915 119.405 ;
        RECT 78.635 119.065 78.910 119.235 ;
        RECT 79.100 119.065 79.630 119.430 ;
        RECT 80.055 118.895 80.385 119.295 ;
        RECT 80.555 119.065 80.810 119.635 ;
        RECT 80.985 120.370 81.255 121.275 ;
        RECT 81.425 120.685 81.755 121.445 ;
        RECT 81.935 120.515 82.105 121.275 ;
        RECT 80.985 119.570 81.155 120.370 ;
        RECT 81.440 120.345 82.105 120.515 ;
        RECT 81.440 120.200 81.610 120.345 ;
        RECT 82.425 120.305 82.635 121.445 ;
        RECT 81.325 119.870 81.610 120.200 ;
        RECT 82.805 120.295 83.135 121.275 ;
        RECT 83.305 120.305 83.535 121.445 ;
        RECT 84.295 120.515 84.465 121.275 ;
        RECT 84.645 120.685 84.975 121.445 ;
        RECT 84.295 120.345 84.960 120.515 ;
        RECT 85.145 120.370 85.415 121.275 ;
        RECT 85.590 121.010 90.935 121.445 ;
        RECT 81.440 119.615 81.610 119.870 ;
        RECT 81.845 119.795 82.175 120.165 ;
        RECT 80.985 119.065 81.245 119.570 ;
        RECT 81.440 119.445 82.105 119.615 ;
        RECT 81.425 118.895 81.755 119.275 ;
        RECT 81.935 119.065 82.105 119.445 ;
        RECT 82.425 118.895 82.635 119.715 ;
        RECT 82.805 119.695 83.055 120.295 ;
        RECT 84.790 120.200 84.960 120.345 ;
        RECT 83.225 119.885 83.555 120.135 ;
        RECT 84.225 119.795 84.555 120.165 ;
        RECT 84.790 119.870 85.075 120.200 ;
        RECT 82.805 119.065 83.135 119.695 ;
        RECT 83.305 118.895 83.535 119.715 ;
        RECT 84.790 119.615 84.960 119.870 ;
        RECT 84.295 119.445 84.960 119.615 ;
        RECT 85.245 119.570 85.415 120.370 ;
        RECT 87.180 119.760 87.530 121.010 ;
        RECT 91.110 120.305 91.445 121.275 ;
        RECT 91.615 120.305 91.785 121.445 ;
        RECT 91.955 121.105 93.985 121.275 ;
        RECT 84.295 119.065 84.465 119.445 ;
        RECT 84.645 118.895 84.975 119.275 ;
        RECT 85.155 119.065 85.415 119.570 ;
        RECT 89.010 119.440 89.350 120.270 ;
        RECT 91.110 119.635 91.280 120.305 ;
        RECT 91.955 120.135 92.125 121.105 ;
        RECT 91.450 119.805 91.705 120.135 ;
        RECT 91.930 119.805 92.125 120.135 ;
        RECT 92.295 120.765 93.420 120.935 ;
        RECT 91.535 119.635 91.705 119.805 ;
        RECT 92.295 119.635 92.465 120.765 ;
        RECT 85.590 118.895 90.935 119.440 ;
        RECT 91.110 119.065 91.365 119.635 ;
        RECT 91.535 119.465 92.465 119.635 ;
        RECT 92.635 120.425 93.645 120.595 ;
        RECT 92.635 119.625 92.805 120.425 ;
        RECT 92.290 119.430 92.465 119.465 ;
        RECT 91.535 118.895 91.865 119.295 ;
        RECT 92.290 119.065 92.820 119.430 ;
        RECT 93.010 119.405 93.285 120.225 ;
        RECT 93.005 119.235 93.285 119.405 ;
        RECT 93.010 119.065 93.285 119.235 ;
        RECT 93.455 119.065 93.645 120.425 ;
        RECT 93.815 120.440 93.985 121.105 ;
        RECT 94.155 120.685 94.325 121.445 ;
        RECT 94.560 120.685 95.075 121.095 ;
        RECT 93.815 120.250 94.565 120.440 ;
        RECT 94.735 119.875 95.075 120.685 ;
        RECT 93.845 119.705 95.075 119.875 ;
        RECT 95.705 120.355 97.375 121.445 ;
        RECT 97.545 120.685 98.060 121.095 ;
        RECT 98.295 120.685 98.465 121.445 ;
        RECT 98.635 121.105 100.665 121.275 ;
        RECT 95.705 119.835 96.455 120.355 ;
        RECT 93.825 118.895 94.335 119.430 ;
        RECT 94.555 119.100 94.800 119.705 ;
        RECT 96.625 119.665 97.375 120.185 ;
        RECT 97.545 119.875 97.885 120.685 ;
        RECT 98.635 120.440 98.805 121.105 ;
        RECT 99.200 120.765 100.325 120.935 ;
        RECT 98.055 120.250 98.805 120.440 ;
        RECT 98.975 120.425 99.985 120.595 ;
        RECT 97.545 119.705 98.775 119.875 ;
        RECT 95.705 118.895 97.375 119.665 ;
        RECT 97.820 119.100 98.065 119.705 ;
        RECT 98.285 118.895 98.795 119.430 ;
        RECT 98.975 119.065 99.165 120.425 ;
        RECT 99.335 120.085 99.610 120.225 ;
        RECT 99.335 119.915 99.615 120.085 ;
        RECT 99.335 119.065 99.610 119.915 ;
        RECT 99.815 119.625 99.985 120.425 ;
        RECT 100.155 119.635 100.325 120.765 ;
        RECT 100.495 120.135 100.665 121.105 ;
        RECT 100.835 120.305 101.005 121.445 ;
        RECT 101.175 120.305 101.510 121.275 ;
        RECT 100.495 119.805 100.690 120.135 ;
        RECT 100.915 119.805 101.170 120.135 ;
        RECT 100.915 119.635 101.085 119.805 ;
        RECT 101.340 119.635 101.510 120.305 ;
        RECT 101.685 120.280 101.975 121.445 ;
        RECT 102.145 120.355 103.355 121.445 ;
        RECT 102.145 119.815 102.665 120.355 ;
        RECT 103.565 120.305 103.795 121.445 ;
        RECT 103.965 120.295 104.295 121.275 ;
        RECT 104.465 120.305 104.675 121.445 ;
        RECT 104.905 120.685 105.420 121.095 ;
        RECT 105.655 120.685 105.825 121.445 ;
        RECT 105.995 121.105 108.025 121.275 ;
        RECT 102.835 119.645 103.355 120.185 ;
        RECT 103.545 119.885 103.875 120.135 ;
        RECT 100.155 119.465 101.085 119.635 ;
        RECT 100.155 119.430 100.330 119.465 ;
        RECT 99.800 119.065 100.330 119.430 ;
        RECT 100.755 118.895 101.085 119.295 ;
        RECT 101.255 119.065 101.510 119.635 ;
        RECT 101.685 118.895 101.975 119.620 ;
        RECT 102.145 118.895 103.355 119.645 ;
        RECT 103.565 118.895 103.795 119.715 ;
        RECT 104.045 119.695 104.295 120.295 ;
        RECT 104.905 119.875 105.245 120.685 ;
        RECT 105.995 120.440 106.165 121.105 ;
        RECT 106.560 120.765 107.685 120.935 ;
        RECT 105.415 120.250 106.165 120.440 ;
        RECT 106.335 120.425 107.345 120.595 ;
        RECT 103.965 119.065 104.295 119.695 ;
        RECT 104.465 118.895 104.675 119.715 ;
        RECT 104.905 119.705 106.135 119.875 ;
        RECT 105.180 119.100 105.425 119.705 ;
        RECT 105.645 118.895 106.155 119.430 ;
        RECT 106.335 119.065 106.525 120.425 ;
        RECT 106.695 119.745 106.970 120.225 ;
        RECT 106.695 119.575 106.975 119.745 ;
        RECT 107.175 119.625 107.345 120.425 ;
        RECT 107.515 119.635 107.685 120.765 ;
        RECT 107.855 120.135 108.025 121.105 ;
        RECT 108.195 120.305 108.365 121.445 ;
        RECT 108.535 120.305 108.870 121.275 ;
        RECT 109.420 120.465 109.675 121.135 ;
        RECT 109.855 120.645 110.140 121.445 ;
        RECT 110.320 120.725 110.650 121.235 ;
        RECT 109.420 120.425 109.600 120.465 ;
        RECT 107.855 119.805 108.050 120.135 ;
        RECT 108.275 119.805 108.530 120.135 ;
        RECT 108.275 119.635 108.445 119.805 ;
        RECT 108.700 119.635 108.870 120.305 ;
        RECT 109.335 120.255 109.600 120.425 ;
        RECT 106.695 119.065 106.970 119.575 ;
        RECT 107.515 119.465 108.445 119.635 ;
        RECT 107.515 119.430 107.690 119.465 ;
        RECT 107.160 119.065 107.690 119.430 ;
        RECT 108.115 118.895 108.445 119.295 ;
        RECT 108.615 119.065 108.870 119.635 ;
        RECT 109.420 119.605 109.600 120.255 ;
        RECT 110.320 120.135 110.570 120.725 ;
        RECT 110.920 120.575 111.090 121.185 ;
        RECT 111.260 120.755 111.590 121.445 ;
        RECT 111.820 120.895 112.060 121.185 ;
        RECT 112.260 121.065 112.680 121.445 ;
        RECT 112.860 120.975 113.490 121.225 ;
        RECT 113.960 121.065 114.290 121.445 ;
        RECT 112.860 120.895 113.030 120.975 ;
        RECT 114.460 120.895 114.630 121.185 ;
        RECT 114.810 121.065 115.190 121.445 ;
        RECT 115.430 121.060 116.260 121.230 ;
        RECT 111.820 120.725 113.030 120.895 ;
        RECT 109.770 119.805 110.570 120.135 ;
        RECT 109.420 119.075 109.675 119.605 ;
        RECT 109.855 118.895 110.140 119.355 ;
        RECT 110.320 119.155 110.570 119.805 ;
        RECT 110.770 120.555 111.090 120.575 ;
        RECT 110.770 120.385 112.690 120.555 ;
        RECT 110.770 119.490 110.960 120.385 ;
        RECT 112.860 120.215 113.030 120.725 ;
        RECT 113.200 120.465 113.720 120.775 ;
        RECT 111.130 120.045 113.030 120.215 ;
        RECT 111.130 119.985 111.460 120.045 ;
        RECT 111.610 119.815 111.940 119.875 ;
        RECT 111.280 119.545 111.940 119.815 ;
        RECT 110.770 119.160 111.090 119.490 ;
        RECT 111.270 118.895 111.930 119.375 ;
        RECT 112.130 119.285 112.300 120.045 ;
        RECT 113.200 119.875 113.380 120.285 ;
        RECT 112.470 119.705 112.800 119.825 ;
        RECT 113.550 119.705 113.720 120.465 ;
        RECT 112.470 119.535 113.720 119.705 ;
        RECT 113.890 120.645 115.260 120.895 ;
        RECT 113.890 119.875 114.080 120.645 ;
        RECT 115.010 120.385 115.260 120.645 ;
        RECT 114.250 120.215 114.500 120.375 ;
        RECT 115.430 120.215 115.600 121.060 ;
        RECT 116.495 120.775 116.665 121.275 ;
        RECT 116.835 120.945 117.165 121.445 ;
        RECT 115.770 120.385 116.270 120.765 ;
        RECT 116.495 120.605 117.190 120.775 ;
        RECT 114.250 120.045 115.600 120.215 ;
        RECT 115.180 120.005 115.600 120.045 ;
        RECT 113.890 119.535 114.310 119.875 ;
        RECT 114.600 119.545 115.010 119.875 ;
        RECT 112.130 119.115 112.980 119.285 ;
        RECT 113.540 118.895 113.860 119.355 ;
        RECT 114.060 119.105 114.310 119.535 ;
        RECT 114.600 118.895 115.010 119.335 ;
        RECT 115.180 119.275 115.350 120.005 ;
        RECT 115.520 119.455 115.870 119.825 ;
        RECT 116.050 119.515 116.270 120.385 ;
        RECT 116.440 119.815 116.850 120.435 ;
        RECT 117.020 119.635 117.190 120.605 ;
        RECT 116.495 119.445 117.190 119.635 ;
        RECT 115.180 119.075 116.195 119.275 ;
        RECT 116.495 119.115 116.665 119.445 ;
        RECT 116.835 118.895 117.165 119.275 ;
        RECT 117.380 119.155 117.605 121.275 ;
        RECT 117.775 120.945 118.105 121.445 ;
        RECT 118.275 120.775 118.445 121.275 ;
        RECT 117.780 120.605 118.445 120.775 ;
        RECT 117.780 119.615 118.010 120.605 ;
        RECT 118.180 119.785 118.530 120.435 ;
        RECT 118.745 120.305 118.975 121.445 ;
        RECT 119.145 120.295 119.475 121.275 ;
        RECT 119.645 120.305 119.855 121.445 ;
        RECT 120.635 120.515 120.805 121.275 ;
        RECT 120.985 120.685 121.315 121.445 ;
        RECT 120.635 120.345 121.300 120.515 ;
        RECT 121.485 120.370 121.755 121.275 ;
        RECT 118.725 119.885 119.055 120.135 ;
        RECT 117.780 119.445 118.445 119.615 ;
        RECT 117.775 118.895 118.105 119.275 ;
        RECT 118.275 119.155 118.445 119.445 ;
        RECT 118.745 118.895 118.975 119.715 ;
        RECT 119.225 119.695 119.475 120.295 ;
        RECT 121.130 120.200 121.300 120.345 ;
        RECT 120.565 119.795 120.895 120.165 ;
        RECT 121.130 119.870 121.415 120.200 ;
        RECT 119.145 119.065 119.475 119.695 ;
        RECT 119.645 118.895 119.855 119.715 ;
        RECT 121.130 119.615 121.300 119.870 ;
        RECT 120.635 119.445 121.300 119.615 ;
        RECT 121.585 119.570 121.755 120.370 ;
        RECT 122.845 120.355 126.355 121.445 ;
        RECT 126.525 120.355 127.735 121.445 ;
        RECT 122.845 119.835 124.535 120.355 ;
        RECT 124.705 119.665 126.355 120.185 ;
        RECT 126.525 119.815 127.045 120.355 ;
        RECT 120.635 119.065 120.805 119.445 ;
        RECT 120.985 118.895 121.315 119.275 ;
        RECT 121.495 119.065 121.755 119.570 ;
        RECT 122.845 118.895 126.355 119.665 ;
        RECT 127.215 119.645 127.735 120.185 ;
        RECT 126.525 118.895 127.735 119.645 ;
        RECT 14.660 118.725 127.820 118.895 ;
        RECT 14.745 117.975 15.955 118.725 ;
        RECT 14.745 117.435 15.265 117.975 ;
        RECT 16.645 117.905 16.855 118.725 ;
        RECT 17.025 117.925 17.355 118.555 ;
        RECT 15.435 117.265 15.955 117.805 ;
        RECT 17.025 117.325 17.275 117.925 ;
        RECT 17.525 117.905 17.755 118.725 ;
        RECT 18.340 118.385 18.595 118.545 ;
        RECT 18.255 118.215 18.595 118.385 ;
        RECT 18.775 118.265 19.060 118.725 ;
        RECT 18.340 118.015 18.595 118.215 ;
        RECT 17.445 117.485 17.775 117.735 ;
        RECT 14.745 116.175 15.955 117.265 ;
        RECT 16.645 116.175 16.855 117.315 ;
        RECT 17.025 116.345 17.355 117.325 ;
        RECT 17.525 116.175 17.755 117.315 ;
        RECT 18.340 117.155 18.520 118.015 ;
        RECT 19.240 117.815 19.490 118.465 ;
        RECT 18.690 117.485 19.490 117.815 ;
        RECT 18.340 116.485 18.595 117.155 ;
        RECT 18.775 116.175 19.060 116.975 ;
        RECT 19.240 116.895 19.490 117.485 ;
        RECT 19.690 118.130 20.010 118.460 ;
        RECT 20.190 118.245 20.850 118.725 ;
        RECT 21.050 118.335 21.900 118.505 ;
        RECT 19.690 117.235 19.880 118.130 ;
        RECT 20.200 117.805 20.860 118.075 ;
        RECT 20.530 117.745 20.860 117.805 ;
        RECT 20.050 117.575 20.380 117.635 ;
        RECT 21.050 117.575 21.220 118.335 ;
        RECT 22.460 118.265 22.780 118.725 ;
        RECT 22.980 118.085 23.230 118.515 ;
        RECT 23.520 118.285 23.930 118.725 ;
        RECT 24.100 118.345 25.115 118.545 ;
        RECT 21.390 117.915 22.640 118.085 ;
        RECT 21.390 117.795 21.720 117.915 ;
        RECT 20.050 117.405 21.950 117.575 ;
        RECT 19.690 117.065 21.610 117.235 ;
        RECT 19.690 117.045 20.010 117.065 ;
        RECT 19.240 116.385 19.570 116.895 ;
        RECT 19.840 116.435 20.010 117.045 ;
        RECT 21.780 116.895 21.950 117.405 ;
        RECT 22.120 117.335 22.300 117.745 ;
        RECT 22.470 117.155 22.640 117.915 ;
        RECT 20.180 116.175 20.510 116.865 ;
        RECT 20.740 116.725 21.950 116.895 ;
        RECT 22.120 116.845 22.640 117.155 ;
        RECT 22.810 117.745 23.230 118.085 ;
        RECT 23.520 117.745 23.930 118.075 ;
        RECT 22.810 116.975 23.000 117.745 ;
        RECT 24.100 117.615 24.270 118.345 ;
        RECT 25.415 118.175 25.585 118.505 ;
        RECT 25.755 118.345 26.085 118.725 ;
        RECT 24.440 117.795 24.790 118.165 ;
        RECT 24.100 117.575 24.520 117.615 ;
        RECT 23.170 117.405 24.520 117.575 ;
        RECT 23.170 117.245 23.420 117.405 ;
        RECT 23.930 116.975 24.180 117.235 ;
        RECT 22.810 116.725 24.180 116.975 ;
        RECT 20.740 116.435 20.980 116.725 ;
        RECT 21.780 116.645 21.950 116.725 ;
        RECT 21.180 116.175 21.600 116.555 ;
        RECT 21.780 116.395 22.410 116.645 ;
        RECT 22.880 116.175 23.210 116.555 ;
        RECT 23.380 116.435 23.550 116.725 ;
        RECT 24.350 116.560 24.520 117.405 ;
        RECT 24.970 117.235 25.190 118.105 ;
        RECT 25.415 117.985 26.110 118.175 ;
        RECT 24.690 116.855 25.190 117.235 ;
        RECT 25.360 117.185 25.770 117.805 ;
        RECT 25.940 117.015 26.110 117.985 ;
        RECT 25.415 116.845 26.110 117.015 ;
        RECT 23.730 116.175 24.110 116.555 ;
        RECT 24.350 116.390 25.180 116.560 ;
        RECT 25.415 116.345 25.585 116.845 ;
        RECT 25.755 116.175 26.085 116.675 ;
        RECT 26.300 116.345 26.525 118.465 ;
        RECT 26.695 118.345 27.025 118.725 ;
        RECT 27.195 118.175 27.365 118.465 ;
        RECT 26.700 118.005 27.365 118.175 ;
        RECT 27.715 118.175 27.885 118.465 ;
        RECT 28.055 118.345 28.385 118.725 ;
        RECT 27.715 118.005 28.380 118.175 ;
        RECT 26.700 117.015 26.930 118.005 ;
        RECT 27.100 117.185 27.450 117.835 ;
        RECT 27.630 117.185 27.980 117.835 ;
        RECT 28.150 117.015 28.380 118.005 ;
        RECT 26.700 116.845 27.365 117.015 ;
        RECT 26.695 116.175 27.025 116.675 ;
        RECT 27.195 116.345 27.365 116.845 ;
        RECT 27.715 116.845 28.380 117.015 ;
        RECT 27.715 116.345 27.885 116.845 ;
        RECT 28.055 116.175 28.385 116.675 ;
        RECT 28.555 116.345 28.780 118.465 ;
        RECT 28.995 118.345 29.325 118.725 ;
        RECT 29.495 118.175 29.665 118.505 ;
        RECT 29.965 118.345 30.980 118.545 ;
        RECT 28.970 117.985 29.665 118.175 ;
        RECT 28.970 117.015 29.140 117.985 ;
        RECT 29.310 117.185 29.720 117.805 ;
        RECT 29.890 117.235 30.110 118.105 ;
        RECT 30.290 117.795 30.640 118.165 ;
        RECT 30.810 117.615 30.980 118.345 ;
        RECT 31.150 118.285 31.560 118.725 ;
        RECT 31.850 118.085 32.100 118.515 ;
        RECT 32.300 118.265 32.620 118.725 ;
        RECT 33.180 118.335 34.030 118.505 ;
        RECT 31.150 117.745 31.560 118.075 ;
        RECT 31.850 117.745 32.270 118.085 ;
        RECT 30.560 117.575 30.980 117.615 ;
        RECT 30.560 117.405 31.910 117.575 ;
        RECT 28.970 116.845 29.665 117.015 ;
        RECT 29.890 116.855 30.390 117.235 ;
        RECT 28.995 116.175 29.325 116.675 ;
        RECT 29.495 116.345 29.665 116.845 ;
        RECT 30.560 116.560 30.730 117.405 ;
        RECT 31.660 117.245 31.910 117.405 ;
        RECT 30.900 116.975 31.150 117.235 ;
        RECT 32.080 116.975 32.270 117.745 ;
        RECT 30.900 116.725 32.270 116.975 ;
        RECT 32.440 117.915 33.690 118.085 ;
        RECT 32.440 117.155 32.610 117.915 ;
        RECT 33.360 117.795 33.690 117.915 ;
        RECT 32.780 117.335 32.960 117.745 ;
        RECT 33.860 117.575 34.030 118.335 ;
        RECT 34.230 118.245 34.890 118.725 ;
        RECT 35.070 118.130 35.390 118.460 ;
        RECT 34.220 117.805 34.880 118.075 ;
        RECT 34.220 117.745 34.550 117.805 ;
        RECT 34.700 117.575 35.030 117.635 ;
        RECT 33.130 117.405 35.030 117.575 ;
        RECT 32.440 116.845 32.960 117.155 ;
        RECT 33.130 116.895 33.300 117.405 ;
        RECT 35.200 117.235 35.390 118.130 ;
        RECT 33.470 117.065 35.390 117.235 ;
        RECT 35.070 117.045 35.390 117.065 ;
        RECT 35.590 117.815 35.840 118.465 ;
        RECT 36.020 118.265 36.305 118.725 ;
        RECT 36.485 118.385 36.740 118.545 ;
        RECT 36.485 118.215 36.825 118.385 ;
        RECT 36.485 118.015 36.740 118.215 ;
        RECT 35.590 117.485 36.390 117.815 ;
        RECT 33.130 116.725 34.340 116.895 ;
        RECT 29.900 116.390 30.730 116.560 ;
        RECT 30.970 116.175 31.350 116.555 ;
        RECT 31.530 116.435 31.700 116.725 ;
        RECT 33.130 116.645 33.300 116.725 ;
        RECT 31.870 116.175 32.200 116.555 ;
        RECT 32.670 116.395 33.300 116.645 ;
        RECT 33.480 116.175 33.900 116.555 ;
        RECT 34.100 116.435 34.340 116.725 ;
        RECT 34.570 116.175 34.900 116.865 ;
        RECT 35.070 116.435 35.240 117.045 ;
        RECT 35.590 116.895 35.840 117.485 ;
        RECT 36.560 117.155 36.740 118.015 ;
        RECT 37.285 118.000 37.575 118.725 ;
        RECT 38.120 118.385 38.375 118.545 ;
        RECT 38.035 118.215 38.375 118.385 ;
        RECT 38.555 118.265 38.840 118.725 ;
        RECT 38.120 118.015 38.375 118.215 ;
        RECT 35.510 116.385 35.840 116.895 ;
        RECT 36.020 116.175 36.305 116.975 ;
        RECT 36.485 116.485 36.740 117.155 ;
        RECT 37.285 116.175 37.575 117.340 ;
        RECT 38.120 117.155 38.300 118.015 ;
        RECT 39.020 117.815 39.270 118.465 ;
        RECT 38.470 117.485 39.270 117.815 ;
        RECT 38.120 116.485 38.375 117.155 ;
        RECT 38.555 116.175 38.840 116.975 ;
        RECT 39.020 116.895 39.270 117.485 ;
        RECT 39.470 118.130 39.790 118.460 ;
        RECT 39.970 118.245 40.630 118.725 ;
        RECT 40.830 118.335 41.680 118.505 ;
        RECT 39.470 117.235 39.660 118.130 ;
        RECT 39.980 117.805 40.640 118.075 ;
        RECT 40.310 117.745 40.640 117.805 ;
        RECT 39.830 117.575 40.160 117.635 ;
        RECT 40.830 117.575 41.000 118.335 ;
        RECT 42.240 118.265 42.560 118.725 ;
        RECT 42.760 118.085 43.010 118.515 ;
        RECT 43.300 118.285 43.710 118.725 ;
        RECT 43.880 118.345 44.895 118.545 ;
        RECT 41.170 117.915 42.420 118.085 ;
        RECT 41.170 117.795 41.500 117.915 ;
        RECT 39.830 117.405 41.730 117.575 ;
        RECT 39.470 117.065 41.390 117.235 ;
        RECT 39.470 117.045 39.790 117.065 ;
        RECT 39.020 116.385 39.350 116.895 ;
        RECT 39.620 116.435 39.790 117.045 ;
        RECT 41.560 116.895 41.730 117.405 ;
        RECT 41.900 117.335 42.080 117.745 ;
        RECT 42.250 117.155 42.420 117.915 ;
        RECT 39.960 116.175 40.290 116.865 ;
        RECT 40.520 116.725 41.730 116.895 ;
        RECT 41.900 116.845 42.420 117.155 ;
        RECT 42.590 117.745 43.010 118.085 ;
        RECT 43.300 117.745 43.710 118.075 ;
        RECT 42.590 116.975 42.780 117.745 ;
        RECT 43.880 117.615 44.050 118.345 ;
        RECT 45.195 118.175 45.365 118.505 ;
        RECT 45.535 118.345 45.865 118.725 ;
        RECT 44.220 117.795 44.570 118.165 ;
        RECT 43.880 117.575 44.300 117.615 ;
        RECT 42.950 117.405 44.300 117.575 ;
        RECT 42.950 117.245 43.200 117.405 ;
        RECT 43.710 116.975 43.960 117.235 ;
        RECT 42.590 116.725 43.960 116.975 ;
        RECT 40.520 116.435 40.760 116.725 ;
        RECT 41.560 116.645 41.730 116.725 ;
        RECT 40.960 116.175 41.380 116.555 ;
        RECT 41.560 116.395 42.190 116.645 ;
        RECT 42.660 116.175 42.990 116.555 ;
        RECT 43.160 116.435 43.330 116.725 ;
        RECT 44.130 116.560 44.300 117.405 ;
        RECT 44.750 117.235 44.970 118.105 ;
        RECT 45.195 117.985 45.890 118.175 ;
        RECT 44.470 116.855 44.970 117.235 ;
        RECT 45.140 117.185 45.550 117.805 ;
        RECT 45.720 117.015 45.890 117.985 ;
        RECT 45.195 116.845 45.890 117.015 ;
        RECT 43.510 116.175 43.890 116.555 ;
        RECT 44.130 116.390 44.960 116.560 ;
        RECT 45.195 116.345 45.365 116.845 ;
        RECT 45.535 116.175 45.865 116.675 ;
        RECT 46.080 116.345 46.305 118.465 ;
        RECT 46.475 118.345 46.805 118.725 ;
        RECT 46.975 118.175 47.145 118.465 ;
        RECT 46.480 118.005 47.145 118.175 ;
        RECT 47.780 118.015 48.035 118.545 ;
        RECT 48.215 118.265 48.500 118.725 ;
        RECT 46.480 117.015 46.710 118.005 ;
        RECT 46.880 117.185 47.230 117.835 ;
        RECT 47.780 117.155 47.960 118.015 ;
        RECT 48.680 117.815 48.930 118.465 ;
        RECT 48.130 117.485 48.930 117.815 ;
        RECT 46.480 116.845 47.145 117.015 ;
        RECT 46.475 116.175 46.805 116.675 ;
        RECT 46.975 116.345 47.145 116.845 ;
        RECT 47.780 116.685 48.035 117.155 ;
        RECT 47.695 116.515 48.035 116.685 ;
        RECT 47.780 116.485 48.035 116.515 ;
        RECT 48.215 116.175 48.500 116.975 ;
        RECT 48.680 116.895 48.930 117.485 ;
        RECT 49.130 118.130 49.450 118.460 ;
        RECT 49.630 118.245 50.290 118.725 ;
        RECT 50.490 118.335 51.340 118.505 ;
        RECT 49.130 117.235 49.320 118.130 ;
        RECT 49.640 117.805 50.300 118.075 ;
        RECT 49.970 117.745 50.300 117.805 ;
        RECT 49.490 117.575 49.820 117.635 ;
        RECT 50.490 117.575 50.660 118.335 ;
        RECT 51.900 118.265 52.220 118.725 ;
        RECT 52.420 118.085 52.670 118.515 ;
        RECT 52.960 118.285 53.370 118.725 ;
        RECT 53.540 118.345 54.555 118.545 ;
        RECT 50.830 117.915 52.080 118.085 ;
        RECT 50.830 117.795 51.160 117.915 ;
        RECT 49.490 117.405 51.390 117.575 ;
        RECT 49.130 117.065 51.050 117.235 ;
        RECT 49.130 117.045 49.450 117.065 ;
        RECT 48.680 116.385 49.010 116.895 ;
        RECT 49.280 116.435 49.450 117.045 ;
        RECT 51.220 116.895 51.390 117.405 ;
        RECT 51.560 117.335 51.740 117.745 ;
        RECT 51.910 117.155 52.080 117.915 ;
        RECT 49.620 116.175 49.950 116.865 ;
        RECT 50.180 116.725 51.390 116.895 ;
        RECT 51.560 116.845 52.080 117.155 ;
        RECT 52.250 117.745 52.670 118.085 ;
        RECT 52.960 117.745 53.370 118.075 ;
        RECT 52.250 116.975 52.440 117.745 ;
        RECT 53.540 117.615 53.710 118.345 ;
        RECT 54.855 118.175 55.025 118.505 ;
        RECT 55.195 118.345 55.525 118.725 ;
        RECT 53.880 117.795 54.230 118.165 ;
        RECT 53.540 117.575 53.960 117.615 ;
        RECT 52.610 117.405 53.960 117.575 ;
        RECT 52.610 117.245 52.860 117.405 ;
        RECT 53.370 116.975 53.620 117.235 ;
        RECT 52.250 116.725 53.620 116.975 ;
        RECT 50.180 116.435 50.420 116.725 ;
        RECT 51.220 116.645 51.390 116.725 ;
        RECT 50.620 116.175 51.040 116.555 ;
        RECT 51.220 116.395 51.850 116.645 ;
        RECT 52.320 116.175 52.650 116.555 ;
        RECT 52.820 116.435 52.990 116.725 ;
        RECT 53.790 116.560 53.960 117.405 ;
        RECT 54.410 117.235 54.630 118.105 ;
        RECT 54.855 117.985 55.550 118.175 ;
        RECT 54.130 116.855 54.630 117.235 ;
        RECT 54.800 117.185 55.210 117.805 ;
        RECT 55.380 117.015 55.550 117.985 ;
        RECT 54.855 116.845 55.550 117.015 ;
        RECT 53.170 116.175 53.550 116.555 ;
        RECT 53.790 116.390 54.620 116.560 ;
        RECT 54.855 116.345 55.025 116.845 ;
        RECT 55.195 116.175 55.525 116.675 ;
        RECT 55.740 116.345 55.965 118.465 ;
        RECT 56.135 118.345 56.465 118.725 ;
        RECT 56.635 118.175 56.805 118.465 ;
        RECT 56.140 118.005 56.805 118.175 ;
        RECT 56.140 117.015 56.370 118.005 ;
        RECT 57.985 117.955 61.495 118.725 ;
        RECT 56.540 117.185 56.890 117.835 ;
        RECT 57.985 117.265 59.675 117.785 ;
        RECT 59.845 117.435 61.495 117.955 ;
        RECT 61.705 117.905 61.935 118.725 ;
        RECT 62.105 117.925 62.435 118.555 ;
        RECT 61.685 117.485 62.015 117.735 ;
        RECT 62.185 117.325 62.435 117.925 ;
        RECT 62.605 117.905 62.815 118.725 ;
        RECT 63.045 118.000 63.335 118.725 ;
        RECT 63.880 118.385 64.135 118.545 ;
        RECT 63.795 118.215 64.135 118.385 ;
        RECT 64.315 118.265 64.600 118.725 ;
        RECT 63.880 118.015 64.135 118.215 ;
        RECT 56.140 116.845 56.805 117.015 ;
        RECT 56.135 116.175 56.465 116.675 ;
        RECT 56.635 116.345 56.805 116.845 ;
        RECT 57.985 116.175 61.495 117.265 ;
        RECT 61.705 116.175 61.935 117.315 ;
        RECT 62.105 116.345 62.435 117.325 ;
        RECT 62.605 116.175 62.815 117.315 ;
        RECT 63.045 116.175 63.335 117.340 ;
        RECT 63.880 117.155 64.060 118.015 ;
        RECT 64.780 117.815 65.030 118.465 ;
        RECT 64.230 117.485 65.030 117.815 ;
        RECT 63.880 116.485 64.135 117.155 ;
        RECT 64.315 116.175 64.600 116.975 ;
        RECT 64.780 116.895 65.030 117.485 ;
        RECT 65.230 118.130 65.550 118.460 ;
        RECT 65.730 118.245 66.390 118.725 ;
        RECT 66.590 118.335 67.440 118.505 ;
        RECT 65.230 117.235 65.420 118.130 ;
        RECT 65.740 117.805 66.400 118.075 ;
        RECT 66.070 117.745 66.400 117.805 ;
        RECT 65.590 117.575 65.920 117.635 ;
        RECT 66.590 117.575 66.760 118.335 ;
        RECT 68.000 118.265 68.320 118.725 ;
        RECT 68.520 118.085 68.770 118.515 ;
        RECT 69.060 118.285 69.470 118.725 ;
        RECT 69.640 118.345 70.655 118.545 ;
        RECT 66.930 117.915 68.180 118.085 ;
        RECT 66.930 117.795 67.260 117.915 ;
        RECT 65.590 117.405 67.490 117.575 ;
        RECT 65.230 117.065 67.150 117.235 ;
        RECT 65.230 117.045 65.550 117.065 ;
        RECT 64.780 116.385 65.110 116.895 ;
        RECT 65.380 116.435 65.550 117.045 ;
        RECT 67.320 116.895 67.490 117.405 ;
        RECT 67.660 117.335 67.840 117.745 ;
        RECT 68.010 117.155 68.180 117.915 ;
        RECT 65.720 116.175 66.050 116.865 ;
        RECT 66.280 116.725 67.490 116.895 ;
        RECT 67.660 116.845 68.180 117.155 ;
        RECT 68.350 117.745 68.770 118.085 ;
        RECT 69.060 117.745 69.470 118.075 ;
        RECT 68.350 116.975 68.540 117.745 ;
        RECT 69.640 117.615 69.810 118.345 ;
        RECT 70.955 118.175 71.125 118.505 ;
        RECT 71.295 118.345 71.625 118.725 ;
        RECT 69.980 117.795 70.330 118.165 ;
        RECT 69.640 117.575 70.060 117.615 ;
        RECT 68.710 117.405 70.060 117.575 ;
        RECT 68.710 117.245 68.960 117.405 ;
        RECT 69.470 116.975 69.720 117.235 ;
        RECT 68.350 116.725 69.720 116.975 ;
        RECT 66.280 116.435 66.520 116.725 ;
        RECT 67.320 116.645 67.490 116.725 ;
        RECT 66.720 116.175 67.140 116.555 ;
        RECT 67.320 116.395 67.950 116.645 ;
        RECT 68.420 116.175 68.750 116.555 ;
        RECT 68.920 116.435 69.090 116.725 ;
        RECT 69.890 116.560 70.060 117.405 ;
        RECT 70.510 117.235 70.730 118.105 ;
        RECT 70.955 117.985 71.650 118.175 ;
        RECT 70.230 116.855 70.730 117.235 ;
        RECT 70.900 117.185 71.310 117.805 ;
        RECT 71.480 117.015 71.650 117.985 ;
        RECT 70.955 116.845 71.650 117.015 ;
        RECT 69.270 116.175 69.650 116.555 ;
        RECT 69.890 116.390 70.720 116.560 ;
        RECT 70.955 116.345 71.125 116.845 ;
        RECT 71.295 116.175 71.625 116.675 ;
        RECT 71.840 116.345 72.065 118.465 ;
        RECT 72.235 118.345 72.565 118.725 ;
        RECT 72.735 118.175 72.905 118.465 ;
        RECT 73.540 118.385 73.795 118.545 ;
        RECT 73.455 118.215 73.795 118.385 ;
        RECT 73.975 118.265 74.260 118.725 ;
        RECT 72.240 118.005 72.905 118.175 ;
        RECT 73.540 118.015 73.795 118.215 ;
        RECT 72.240 117.015 72.470 118.005 ;
        RECT 72.640 117.185 72.990 117.835 ;
        RECT 73.540 117.155 73.720 118.015 ;
        RECT 74.440 117.815 74.690 118.465 ;
        RECT 73.890 117.485 74.690 117.815 ;
        RECT 72.240 116.845 72.905 117.015 ;
        RECT 72.235 116.175 72.565 116.675 ;
        RECT 72.735 116.345 72.905 116.845 ;
        RECT 73.540 116.485 73.795 117.155 ;
        RECT 73.975 116.175 74.260 116.975 ;
        RECT 74.440 116.895 74.690 117.485 ;
        RECT 74.890 118.130 75.210 118.460 ;
        RECT 75.390 118.245 76.050 118.725 ;
        RECT 76.250 118.335 77.100 118.505 ;
        RECT 74.890 117.235 75.080 118.130 ;
        RECT 75.400 117.805 76.060 118.075 ;
        RECT 75.730 117.745 76.060 117.805 ;
        RECT 75.250 117.575 75.580 117.635 ;
        RECT 76.250 117.575 76.420 118.335 ;
        RECT 77.660 118.265 77.980 118.725 ;
        RECT 78.180 118.085 78.430 118.515 ;
        RECT 78.720 118.285 79.130 118.725 ;
        RECT 79.300 118.345 80.315 118.545 ;
        RECT 76.590 117.915 77.840 118.085 ;
        RECT 76.590 117.795 76.920 117.915 ;
        RECT 75.250 117.405 77.150 117.575 ;
        RECT 74.890 117.065 76.810 117.235 ;
        RECT 74.890 117.045 75.210 117.065 ;
        RECT 74.440 116.385 74.770 116.895 ;
        RECT 75.040 116.435 75.210 117.045 ;
        RECT 76.980 116.895 77.150 117.405 ;
        RECT 77.320 117.335 77.500 117.745 ;
        RECT 77.670 117.155 77.840 117.915 ;
        RECT 75.380 116.175 75.710 116.865 ;
        RECT 75.940 116.725 77.150 116.895 ;
        RECT 77.320 116.845 77.840 117.155 ;
        RECT 78.010 117.745 78.430 118.085 ;
        RECT 78.720 117.745 79.130 118.075 ;
        RECT 78.010 116.975 78.200 117.745 ;
        RECT 79.300 117.615 79.470 118.345 ;
        RECT 80.615 118.175 80.785 118.505 ;
        RECT 80.955 118.345 81.285 118.725 ;
        RECT 79.640 117.795 79.990 118.165 ;
        RECT 79.300 117.575 79.720 117.615 ;
        RECT 78.370 117.405 79.720 117.575 ;
        RECT 78.370 117.245 78.620 117.405 ;
        RECT 79.130 116.975 79.380 117.235 ;
        RECT 78.010 116.725 79.380 116.975 ;
        RECT 75.940 116.435 76.180 116.725 ;
        RECT 76.980 116.645 77.150 116.725 ;
        RECT 76.380 116.175 76.800 116.555 ;
        RECT 76.980 116.395 77.610 116.645 ;
        RECT 78.080 116.175 78.410 116.555 ;
        RECT 78.580 116.435 78.750 116.725 ;
        RECT 79.550 116.560 79.720 117.405 ;
        RECT 80.170 117.235 80.390 118.105 ;
        RECT 80.615 117.985 81.310 118.175 ;
        RECT 79.890 116.855 80.390 117.235 ;
        RECT 80.560 117.185 80.970 117.805 ;
        RECT 81.140 117.015 81.310 117.985 ;
        RECT 80.615 116.845 81.310 117.015 ;
        RECT 78.930 116.175 79.310 116.555 ;
        RECT 79.550 116.390 80.380 116.560 ;
        RECT 80.615 116.345 80.785 116.845 ;
        RECT 80.955 116.175 81.285 116.675 ;
        RECT 81.500 116.345 81.725 118.465 ;
        RECT 81.895 118.345 82.225 118.725 ;
        RECT 82.395 118.175 82.565 118.465 ;
        RECT 81.900 118.005 82.565 118.175 ;
        RECT 81.900 117.015 82.130 118.005 ;
        RECT 82.830 117.985 83.085 118.555 ;
        RECT 83.255 118.325 83.585 118.725 ;
        RECT 84.010 118.190 84.540 118.555 ;
        RECT 84.010 118.155 84.185 118.190 ;
        RECT 83.255 117.985 84.185 118.155 ;
        RECT 82.300 117.185 82.650 117.835 ;
        RECT 82.830 117.315 83.000 117.985 ;
        RECT 83.255 117.815 83.425 117.985 ;
        RECT 83.170 117.485 83.425 117.815 ;
        RECT 83.650 117.485 83.845 117.815 ;
        RECT 81.900 116.845 82.565 117.015 ;
        RECT 81.895 116.175 82.225 116.675 ;
        RECT 82.395 116.345 82.565 116.845 ;
        RECT 82.830 116.345 83.165 117.315 ;
        RECT 83.335 116.175 83.505 117.315 ;
        RECT 83.675 116.515 83.845 117.485 ;
        RECT 84.015 116.855 84.185 117.985 ;
        RECT 84.355 117.195 84.525 117.995 ;
        RECT 84.730 117.705 85.005 118.555 ;
        RECT 84.725 117.535 85.005 117.705 ;
        RECT 84.730 117.395 85.005 117.535 ;
        RECT 85.175 117.195 85.365 118.555 ;
        RECT 85.545 118.190 86.055 118.725 ;
        RECT 86.275 117.915 86.520 118.520 ;
        RECT 87.515 118.175 87.685 118.555 ;
        RECT 87.865 118.345 88.195 118.725 ;
        RECT 87.515 118.005 88.180 118.175 ;
        RECT 88.375 118.050 88.635 118.555 ;
        RECT 85.565 117.745 86.795 117.915 ;
        RECT 84.355 117.025 85.365 117.195 ;
        RECT 85.535 117.180 86.285 117.370 ;
        RECT 84.015 116.685 85.140 116.855 ;
        RECT 85.535 116.515 85.705 117.180 ;
        RECT 86.455 116.935 86.795 117.745 ;
        RECT 87.445 117.455 87.775 117.825 ;
        RECT 88.010 117.750 88.180 118.005 ;
        RECT 88.010 117.420 88.295 117.750 ;
        RECT 88.010 117.275 88.180 117.420 ;
        RECT 83.675 116.345 85.705 116.515 ;
        RECT 85.875 116.175 86.045 116.935 ;
        RECT 86.280 116.525 86.795 116.935 ;
        RECT 87.515 117.105 88.180 117.275 ;
        RECT 88.465 117.250 88.635 118.050 ;
        RECT 88.805 118.000 89.095 118.725 ;
        RECT 89.305 117.905 89.535 118.725 ;
        RECT 89.705 117.925 90.035 118.555 ;
        RECT 89.285 117.485 89.615 117.735 ;
        RECT 87.515 116.345 87.685 117.105 ;
        RECT 87.865 116.175 88.195 116.935 ;
        RECT 88.365 116.345 88.635 117.250 ;
        RECT 88.805 116.175 89.095 117.340 ;
        RECT 89.785 117.325 90.035 117.925 ;
        RECT 90.205 117.905 90.415 118.725 ;
        RECT 90.685 117.905 90.915 118.725 ;
        RECT 91.085 117.925 91.415 118.555 ;
        RECT 90.665 117.485 90.995 117.735 ;
        RECT 91.165 117.325 91.415 117.925 ;
        RECT 91.585 117.905 91.795 118.725 ;
        RECT 93.320 118.385 93.575 118.545 ;
        RECT 93.235 118.215 93.575 118.385 ;
        RECT 93.755 118.265 94.040 118.725 ;
        RECT 93.320 118.015 93.575 118.215 ;
        RECT 89.305 116.175 89.535 117.315 ;
        RECT 89.705 116.345 90.035 117.325 ;
        RECT 90.205 116.175 90.415 117.315 ;
        RECT 90.685 116.175 90.915 117.315 ;
        RECT 91.085 116.345 91.415 117.325 ;
        RECT 91.585 116.175 91.795 117.315 ;
        RECT 93.320 117.155 93.500 118.015 ;
        RECT 94.220 117.815 94.470 118.465 ;
        RECT 93.670 117.485 94.470 117.815 ;
        RECT 93.320 116.485 93.575 117.155 ;
        RECT 93.755 116.175 94.040 116.975 ;
        RECT 94.220 116.895 94.470 117.485 ;
        RECT 94.670 118.130 94.990 118.460 ;
        RECT 95.170 118.245 95.830 118.725 ;
        RECT 96.030 118.335 96.880 118.505 ;
        RECT 94.670 117.235 94.860 118.130 ;
        RECT 95.180 117.805 95.840 118.075 ;
        RECT 95.510 117.745 95.840 117.805 ;
        RECT 95.030 117.575 95.360 117.635 ;
        RECT 96.030 117.575 96.200 118.335 ;
        RECT 97.440 118.265 97.760 118.725 ;
        RECT 97.960 118.085 98.210 118.515 ;
        RECT 98.500 118.285 98.910 118.725 ;
        RECT 99.080 118.345 100.095 118.545 ;
        RECT 96.370 117.915 97.620 118.085 ;
        RECT 96.370 117.795 96.700 117.915 ;
        RECT 95.030 117.405 96.930 117.575 ;
        RECT 94.670 117.065 96.590 117.235 ;
        RECT 94.670 117.045 94.990 117.065 ;
        RECT 94.220 116.385 94.550 116.895 ;
        RECT 94.820 116.435 94.990 117.045 ;
        RECT 96.760 116.895 96.930 117.405 ;
        RECT 97.100 117.335 97.280 117.745 ;
        RECT 97.450 117.155 97.620 117.915 ;
        RECT 95.160 116.175 95.490 116.865 ;
        RECT 95.720 116.725 96.930 116.895 ;
        RECT 97.100 116.845 97.620 117.155 ;
        RECT 97.790 117.745 98.210 118.085 ;
        RECT 98.500 117.745 98.910 118.075 ;
        RECT 97.790 116.975 97.980 117.745 ;
        RECT 99.080 117.615 99.250 118.345 ;
        RECT 100.395 118.175 100.565 118.505 ;
        RECT 100.735 118.345 101.065 118.725 ;
        RECT 99.420 117.795 99.770 118.165 ;
        RECT 99.080 117.575 99.500 117.615 ;
        RECT 98.150 117.405 99.500 117.575 ;
        RECT 98.150 117.245 98.400 117.405 ;
        RECT 98.910 116.975 99.160 117.235 ;
        RECT 97.790 116.725 99.160 116.975 ;
        RECT 95.720 116.435 95.960 116.725 ;
        RECT 96.760 116.645 96.930 116.725 ;
        RECT 96.160 116.175 96.580 116.555 ;
        RECT 96.760 116.395 97.390 116.645 ;
        RECT 97.860 116.175 98.190 116.555 ;
        RECT 98.360 116.435 98.530 116.725 ;
        RECT 99.330 116.560 99.500 117.405 ;
        RECT 99.950 117.235 100.170 118.105 ;
        RECT 100.395 117.985 101.090 118.175 ;
        RECT 99.670 116.855 100.170 117.235 ;
        RECT 100.340 117.185 100.750 117.805 ;
        RECT 100.920 117.015 101.090 117.985 ;
        RECT 100.395 116.845 101.090 117.015 ;
        RECT 98.710 116.175 99.090 116.555 ;
        RECT 99.330 116.390 100.160 116.560 ;
        RECT 100.395 116.345 100.565 116.845 ;
        RECT 100.735 116.175 101.065 116.675 ;
        RECT 101.280 116.345 101.505 118.465 ;
        RECT 101.675 118.345 102.005 118.725 ;
        RECT 102.175 118.175 102.345 118.465 ;
        RECT 102.980 118.385 103.235 118.545 ;
        RECT 102.895 118.215 103.235 118.385 ;
        RECT 103.415 118.265 103.700 118.725 ;
        RECT 101.680 118.005 102.345 118.175 ;
        RECT 102.980 118.015 103.235 118.215 ;
        RECT 101.680 117.015 101.910 118.005 ;
        RECT 102.080 117.185 102.430 117.835 ;
        RECT 102.980 117.155 103.160 118.015 ;
        RECT 103.880 117.815 104.130 118.465 ;
        RECT 103.330 117.485 104.130 117.815 ;
        RECT 101.680 116.845 102.345 117.015 ;
        RECT 101.675 116.175 102.005 116.675 ;
        RECT 102.175 116.345 102.345 116.845 ;
        RECT 102.980 116.485 103.235 117.155 ;
        RECT 103.415 116.175 103.700 116.975 ;
        RECT 103.880 116.895 104.130 117.485 ;
        RECT 104.330 118.130 104.650 118.460 ;
        RECT 104.830 118.245 105.490 118.725 ;
        RECT 105.690 118.335 106.540 118.505 ;
        RECT 104.330 117.235 104.520 118.130 ;
        RECT 104.840 117.805 105.500 118.075 ;
        RECT 105.170 117.745 105.500 117.805 ;
        RECT 104.690 117.575 105.020 117.635 ;
        RECT 105.690 117.575 105.860 118.335 ;
        RECT 107.100 118.265 107.420 118.725 ;
        RECT 107.620 118.085 107.870 118.515 ;
        RECT 108.160 118.285 108.570 118.725 ;
        RECT 108.740 118.345 109.755 118.545 ;
        RECT 106.030 117.915 107.280 118.085 ;
        RECT 106.030 117.795 106.360 117.915 ;
        RECT 104.690 117.405 106.590 117.575 ;
        RECT 104.330 117.065 106.250 117.235 ;
        RECT 104.330 117.045 104.650 117.065 ;
        RECT 103.880 116.385 104.210 116.895 ;
        RECT 104.480 116.435 104.650 117.045 ;
        RECT 106.420 116.895 106.590 117.405 ;
        RECT 106.760 117.335 106.940 117.745 ;
        RECT 107.110 117.155 107.280 117.915 ;
        RECT 104.820 116.175 105.150 116.865 ;
        RECT 105.380 116.725 106.590 116.895 ;
        RECT 106.760 116.845 107.280 117.155 ;
        RECT 107.450 117.745 107.870 118.085 ;
        RECT 108.160 117.745 108.570 118.075 ;
        RECT 107.450 116.975 107.640 117.745 ;
        RECT 108.740 117.615 108.910 118.345 ;
        RECT 110.055 118.175 110.225 118.505 ;
        RECT 110.395 118.345 110.725 118.725 ;
        RECT 109.080 117.795 109.430 118.165 ;
        RECT 108.740 117.575 109.160 117.615 ;
        RECT 107.810 117.405 109.160 117.575 ;
        RECT 107.810 117.245 108.060 117.405 ;
        RECT 108.570 116.975 108.820 117.235 ;
        RECT 107.450 116.725 108.820 116.975 ;
        RECT 105.380 116.435 105.620 116.725 ;
        RECT 106.420 116.645 106.590 116.725 ;
        RECT 105.820 116.175 106.240 116.555 ;
        RECT 106.420 116.395 107.050 116.645 ;
        RECT 107.520 116.175 107.850 116.555 ;
        RECT 108.020 116.435 108.190 116.725 ;
        RECT 108.990 116.560 109.160 117.405 ;
        RECT 109.610 117.235 109.830 118.105 ;
        RECT 110.055 117.985 110.750 118.175 ;
        RECT 109.330 116.855 109.830 117.235 ;
        RECT 110.000 117.185 110.410 117.805 ;
        RECT 110.580 117.015 110.750 117.985 ;
        RECT 110.055 116.845 110.750 117.015 ;
        RECT 108.370 116.175 108.750 116.555 ;
        RECT 108.990 116.390 109.820 116.560 ;
        RECT 110.055 116.345 110.225 116.845 ;
        RECT 110.395 116.175 110.725 116.675 ;
        RECT 110.940 116.345 111.165 118.465 ;
        RECT 111.335 118.345 111.665 118.725 ;
        RECT 111.835 118.175 112.005 118.465 ;
        RECT 111.340 118.005 112.005 118.175 ;
        RECT 111.340 117.015 111.570 118.005 ;
        RECT 113.245 117.905 113.455 118.725 ;
        RECT 113.625 117.925 113.955 118.555 ;
        RECT 111.740 117.185 112.090 117.835 ;
        RECT 113.625 117.325 113.875 117.925 ;
        RECT 114.125 117.905 114.355 118.725 ;
        RECT 114.565 118.000 114.855 118.725 ;
        RECT 115.575 118.175 115.745 118.555 ;
        RECT 115.925 118.345 116.255 118.725 ;
        RECT 115.575 118.005 116.240 118.175 ;
        RECT 116.435 118.050 116.695 118.555 ;
        RECT 114.045 117.485 114.375 117.735 ;
        RECT 115.505 117.455 115.835 117.825 ;
        RECT 116.070 117.750 116.240 118.005 ;
        RECT 116.070 117.420 116.355 117.750 ;
        RECT 111.340 116.845 112.005 117.015 ;
        RECT 111.335 116.175 111.665 116.675 ;
        RECT 111.835 116.345 112.005 116.845 ;
        RECT 113.245 116.175 113.455 117.315 ;
        RECT 113.625 116.345 113.955 117.325 ;
        RECT 114.125 116.175 114.355 117.315 ;
        RECT 114.565 116.175 114.855 117.340 ;
        RECT 116.070 117.275 116.240 117.420 ;
        RECT 115.575 117.105 116.240 117.275 ;
        RECT 116.525 117.250 116.695 118.050 ;
        RECT 117.325 117.955 120.835 118.725 ;
        RECT 121.010 118.180 126.355 118.725 ;
        RECT 115.575 116.345 115.745 117.105 ;
        RECT 115.925 116.175 116.255 116.935 ;
        RECT 116.425 116.345 116.695 117.250 ;
        RECT 117.325 117.265 119.015 117.785 ;
        RECT 119.185 117.435 120.835 117.955 ;
        RECT 117.325 116.175 120.835 117.265 ;
        RECT 122.600 116.610 122.950 117.860 ;
        RECT 124.430 117.350 124.770 118.180 ;
        RECT 126.525 117.975 127.735 118.725 ;
        RECT 126.525 117.265 127.045 117.805 ;
        RECT 127.215 117.435 127.735 117.975 ;
        RECT 121.010 116.175 126.355 116.610 ;
        RECT 126.525 116.175 127.735 117.265 ;
        RECT 14.660 116.005 127.820 116.175 ;
        RECT 14.745 114.915 15.955 116.005 ;
        RECT 14.745 114.205 15.265 114.745 ;
        RECT 15.435 114.375 15.955 114.915 ;
        RECT 16.125 114.915 17.335 116.005 ;
        RECT 17.505 114.915 21.015 116.005 ;
        RECT 21.275 115.075 21.445 115.835 ;
        RECT 21.625 115.245 21.955 116.005 ;
        RECT 16.125 114.375 16.645 114.915 ;
        RECT 16.815 114.205 17.335 114.745 ;
        RECT 17.505 114.395 19.195 114.915 ;
        RECT 21.275 114.905 21.940 115.075 ;
        RECT 22.125 114.930 22.395 115.835 ;
        RECT 21.770 114.760 21.940 114.905 ;
        RECT 19.365 114.225 21.015 114.745 ;
        RECT 21.205 114.355 21.535 114.725 ;
        RECT 21.770 114.430 22.055 114.760 ;
        RECT 14.745 113.455 15.955 114.205 ;
        RECT 16.125 113.455 17.335 114.205 ;
        RECT 17.505 113.455 21.015 114.225 ;
        RECT 21.770 114.175 21.940 114.430 ;
        RECT 21.275 114.005 21.940 114.175 ;
        RECT 22.225 114.130 22.395 114.930 ;
        RECT 22.625 114.865 22.835 116.005 ;
        RECT 23.005 114.855 23.335 115.835 ;
        RECT 23.505 114.865 23.735 116.005 ;
        RECT 21.275 113.625 21.445 114.005 ;
        RECT 21.625 113.455 21.955 113.835 ;
        RECT 22.135 113.625 22.395 114.130 ;
        RECT 22.625 113.455 22.835 114.275 ;
        RECT 23.005 114.255 23.255 114.855 ;
        RECT 24.405 114.840 24.695 116.005 ;
        RECT 24.955 115.335 25.125 115.835 ;
        RECT 25.295 115.505 25.625 116.005 ;
        RECT 24.955 115.165 25.620 115.335 ;
        RECT 23.425 114.445 23.755 114.695 ;
        RECT 24.870 114.345 25.220 114.995 ;
        RECT 23.005 113.625 23.335 114.255 ;
        RECT 23.505 113.455 23.735 114.275 ;
        RECT 24.405 113.455 24.695 114.180 ;
        RECT 25.390 114.175 25.620 115.165 ;
        RECT 24.955 114.005 25.620 114.175 ;
        RECT 24.955 113.715 25.125 114.005 ;
        RECT 25.295 113.455 25.625 113.835 ;
        RECT 25.795 113.715 26.020 115.835 ;
        RECT 26.235 115.505 26.565 116.005 ;
        RECT 26.735 115.335 26.905 115.835 ;
        RECT 27.140 115.620 27.970 115.790 ;
        RECT 28.210 115.625 28.590 116.005 ;
        RECT 26.210 115.165 26.905 115.335 ;
        RECT 26.210 114.195 26.380 115.165 ;
        RECT 26.550 114.375 26.960 114.995 ;
        RECT 27.130 114.945 27.630 115.325 ;
        RECT 26.210 114.005 26.905 114.195 ;
        RECT 27.130 114.075 27.350 114.945 ;
        RECT 27.800 114.775 27.970 115.620 ;
        RECT 28.770 115.455 28.940 115.745 ;
        RECT 29.110 115.625 29.440 116.005 ;
        RECT 29.910 115.535 30.540 115.785 ;
        RECT 30.720 115.625 31.140 116.005 ;
        RECT 30.370 115.455 30.540 115.535 ;
        RECT 31.340 115.455 31.580 115.745 ;
        RECT 28.140 115.205 29.510 115.455 ;
        RECT 28.140 114.945 28.390 115.205 ;
        RECT 28.900 114.775 29.150 114.935 ;
        RECT 27.800 114.605 29.150 114.775 ;
        RECT 27.800 114.565 28.220 114.605 ;
        RECT 27.530 114.015 27.880 114.385 ;
        RECT 26.235 113.455 26.565 113.835 ;
        RECT 26.735 113.675 26.905 114.005 ;
        RECT 28.050 113.835 28.220 114.565 ;
        RECT 29.320 114.435 29.510 115.205 ;
        RECT 28.390 114.105 28.800 114.435 ;
        RECT 29.090 114.095 29.510 114.435 ;
        RECT 29.680 115.025 30.200 115.335 ;
        RECT 30.370 115.285 31.580 115.455 ;
        RECT 31.810 115.315 32.140 116.005 ;
        RECT 29.680 114.265 29.850 115.025 ;
        RECT 30.020 114.435 30.200 114.845 ;
        RECT 30.370 114.775 30.540 115.285 ;
        RECT 32.310 115.135 32.480 115.745 ;
        RECT 32.750 115.285 33.080 115.795 ;
        RECT 32.310 115.115 32.630 115.135 ;
        RECT 30.710 114.945 32.630 115.115 ;
        RECT 30.370 114.605 32.270 114.775 ;
        RECT 30.600 114.265 30.930 114.385 ;
        RECT 29.680 114.095 30.930 114.265 ;
        RECT 27.205 113.635 28.220 113.835 ;
        RECT 28.390 113.455 28.800 113.895 ;
        RECT 29.090 113.665 29.340 114.095 ;
        RECT 29.540 113.455 29.860 113.915 ;
        RECT 31.100 113.845 31.270 114.605 ;
        RECT 31.940 114.545 32.270 114.605 ;
        RECT 31.460 114.375 31.790 114.435 ;
        RECT 31.460 114.105 32.120 114.375 ;
        RECT 32.440 114.050 32.630 114.945 ;
        RECT 30.420 113.675 31.270 113.845 ;
        RECT 31.470 113.455 32.130 113.935 ;
        RECT 32.310 113.720 32.630 114.050 ;
        RECT 32.830 114.695 33.080 115.285 ;
        RECT 33.260 115.205 33.545 116.005 ;
        RECT 33.725 115.665 33.980 115.695 ;
        RECT 33.725 115.495 34.065 115.665 ;
        RECT 33.725 115.025 33.980 115.495 ;
        RECT 32.830 114.365 33.630 114.695 ;
        RECT 32.830 113.715 33.080 114.365 ;
        RECT 33.800 114.165 33.980 115.025 ;
        RECT 35.045 114.865 35.255 116.005 ;
        RECT 35.425 114.855 35.755 115.835 ;
        RECT 35.925 114.865 36.155 116.005 ;
        RECT 36.915 115.075 37.085 115.835 ;
        RECT 37.265 115.245 37.595 116.005 ;
        RECT 36.915 114.905 37.580 115.075 ;
        RECT 37.765 114.930 38.035 115.835 ;
        RECT 33.260 113.455 33.545 113.915 ;
        RECT 33.725 113.635 33.980 114.165 ;
        RECT 35.045 113.455 35.255 114.275 ;
        RECT 35.425 114.255 35.675 114.855 ;
        RECT 37.410 114.760 37.580 114.905 ;
        RECT 35.845 114.445 36.175 114.695 ;
        RECT 36.845 114.355 37.175 114.725 ;
        RECT 37.410 114.430 37.695 114.760 ;
        RECT 35.425 113.625 35.755 114.255 ;
        RECT 35.925 113.455 36.155 114.275 ;
        RECT 37.410 114.175 37.580 114.430 ;
        RECT 36.915 114.005 37.580 114.175 ;
        RECT 37.865 114.130 38.035 114.930 ;
        RECT 36.915 113.625 37.085 114.005 ;
        RECT 37.265 113.455 37.595 113.835 ;
        RECT 37.775 113.625 38.035 114.130 ;
        RECT 39.125 114.930 39.395 115.835 ;
        RECT 39.565 115.245 39.895 116.005 ;
        RECT 40.075 115.075 40.245 115.835 ;
        RECT 39.125 114.130 39.295 114.930 ;
        RECT 39.580 114.905 40.245 115.075 ;
        RECT 40.505 114.915 44.015 116.005 ;
        RECT 39.580 114.760 39.750 114.905 ;
        RECT 39.465 114.430 39.750 114.760 ;
        RECT 39.580 114.175 39.750 114.430 ;
        RECT 39.985 114.355 40.315 114.725 ;
        RECT 40.505 114.395 42.195 114.915 ;
        RECT 44.245 114.865 44.455 116.005 ;
        RECT 44.625 114.855 44.955 115.835 ;
        RECT 45.125 114.865 45.355 116.005 ;
        RECT 45.570 114.865 45.905 115.835 ;
        RECT 46.075 114.865 46.245 116.005 ;
        RECT 46.415 115.665 48.445 115.835 ;
        RECT 42.365 114.225 44.015 114.745 ;
        RECT 39.125 113.625 39.385 114.130 ;
        RECT 39.580 114.005 40.245 114.175 ;
        RECT 39.565 113.455 39.895 113.835 ;
        RECT 40.075 113.625 40.245 114.005 ;
        RECT 40.505 113.455 44.015 114.225 ;
        RECT 44.245 113.455 44.455 114.275 ;
        RECT 44.625 114.255 44.875 114.855 ;
        RECT 45.045 114.445 45.375 114.695 ;
        RECT 44.625 113.625 44.955 114.255 ;
        RECT 45.125 113.455 45.355 114.275 ;
        RECT 45.570 114.195 45.740 114.865 ;
        RECT 46.415 114.695 46.585 115.665 ;
        RECT 45.910 114.365 46.165 114.695 ;
        RECT 46.390 114.365 46.585 114.695 ;
        RECT 46.755 115.325 47.880 115.495 ;
        RECT 45.995 114.195 46.165 114.365 ;
        RECT 46.755 114.195 46.925 115.325 ;
        RECT 45.570 113.625 45.825 114.195 ;
        RECT 45.995 114.025 46.925 114.195 ;
        RECT 47.095 114.985 48.105 115.155 ;
        RECT 47.095 114.185 47.265 114.985 ;
        RECT 47.470 114.305 47.745 114.785 ;
        RECT 47.465 114.135 47.745 114.305 ;
        RECT 46.750 113.990 46.925 114.025 ;
        RECT 45.995 113.455 46.325 113.855 ;
        RECT 46.750 113.625 47.280 113.990 ;
        RECT 47.470 113.625 47.745 114.135 ;
        RECT 47.915 113.625 48.105 114.985 ;
        RECT 48.275 115.000 48.445 115.665 ;
        RECT 48.615 115.245 48.785 116.005 ;
        RECT 49.020 115.245 49.535 115.655 ;
        RECT 48.275 114.810 49.025 115.000 ;
        RECT 49.195 114.435 49.535 115.245 ;
        RECT 50.165 114.840 50.455 116.005 ;
        RECT 50.625 114.915 52.295 116.005 ;
        RECT 52.555 115.075 52.725 115.835 ;
        RECT 52.905 115.245 53.235 116.005 ;
        RECT 48.305 114.265 49.535 114.435 ;
        RECT 50.625 114.395 51.375 114.915 ;
        RECT 52.555 114.905 53.220 115.075 ;
        RECT 53.405 114.930 53.675 115.835 ;
        RECT 53.050 114.760 53.220 114.905 ;
        RECT 48.285 113.455 48.795 113.990 ;
        RECT 49.015 113.660 49.260 114.265 ;
        RECT 51.545 114.225 52.295 114.745 ;
        RECT 52.485 114.355 52.815 114.725 ;
        RECT 53.050 114.430 53.335 114.760 ;
        RECT 50.165 113.455 50.455 114.180 ;
        RECT 50.625 113.455 52.295 114.225 ;
        RECT 53.050 114.175 53.220 114.430 ;
        RECT 52.555 114.005 53.220 114.175 ;
        RECT 53.505 114.130 53.675 114.930 ;
        RECT 53.845 114.915 55.055 116.005 ;
        RECT 55.230 115.570 60.575 116.005 ;
        RECT 60.750 115.570 66.095 116.005 ;
        RECT 53.845 114.375 54.365 114.915 ;
        RECT 54.535 114.205 55.055 114.745 ;
        RECT 56.820 114.320 57.170 115.570 ;
        RECT 52.555 113.625 52.725 114.005 ;
        RECT 52.905 113.455 53.235 113.835 ;
        RECT 53.415 113.625 53.675 114.130 ;
        RECT 53.845 113.455 55.055 114.205 ;
        RECT 58.650 114.000 58.990 114.830 ;
        RECT 62.340 114.320 62.690 115.570 ;
        RECT 66.305 114.865 66.535 116.005 ;
        RECT 66.705 114.855 67.035 115.835 ;
        RECT 67.205 114.865 67.415 116.005 ;
        RECT 68.195 115.075 68.365 115.835 ;
        RECT 68.545 115.245 68.875 116.005 ;
        RECT 68.195 114.905 68.860 115.075 ;
        RECT 69.045 114.930 69.315 115.835 ;
        RECT 70.410 115.570 75.755 116.005 ;
        RECT 64.170 114.000 64.510 114.830 ;
        RECT 66.285 114.445 66.615 114.695 ;
        RECT 55.230 113.455 60.575 114.000 ;
        RECT 60.750 113.455 66.095 114.000 ;
        RECT 66.305 113.455 66.535 114.275 ;
        RECT 66.785 114.255 67.035 114.855 ;
        RECT 68.690 114.760 68.860 114.905 ;
        RECT 68.125 114.355 68.455 114.725 ;
        RECT 68.690 114.430 68.975 114.760 ;
        RECT 66.705 113.625 67.035 114.255 ;
        RECT 67.205 113.455 67.415 114.275 ;
        RECT 68.690 114.175 68.860 114.430 ;
        RECT 68.195 114.005 68.860 114.175 ;
        RECT 69.145 114.130 69.315 114.930 ;
        RECT 72.000 114.320 72.350 115.570 ;
        RECT 75.925 114.840 76.215 116.005 ;
        RECT 77.680 115.665 77.935 115.695 ;
        RECT 77.595 115.495 77.935 115.665 ;
        RECT 77.680 115.025 77.935 115.495 ;
        RECT 78.115 115.205 78.400 116.005 ;
        RECT 78.580 115.285 78.910 115.795 ;
        RECT 68.195 113.625 68.365 114.005 ;
        RECT 68.545 113.455 68.875 113.835 ;
        RECT 69.055 113.625 69.315 114.130 ;
        RECT 73.830 114.000 74.170 114.830 ;
        RECT 70.410 113.455 75.755 114.000 ;
        RECT 75.925 113.455 76.215 114.180 ;
        RECT 77.680 114.165 77.860 115.025 ;
        RECT 78.580 114.695 78.830 115.285 ;
        RECT 79.180 115.135 79.350 115.745 ;
        RECT 79.520 115.315 79.850 116.005 ;
        RECT 80.080 115.455 80.320 115.745 ;
        RECT 80.520 115.625 80.940 116.005 ;
        RECT 81.120 115.535 81.750 115.785 ;
        RECT 82.220 115.625 82.550 116.005 ;
        RECT 81.120 115.455 81.290 115.535 ;
        RECT 82.720 115.455 82.890 115.745 ;
        RECT 83.070 115.625 83.450 116.005 ;
        RECT 83.690 115.620 84.520 115.790 ;
        RECT 80.080 115.285 81.290 115.455 ;
        RECT 78.030 114.365 78.830 114.695 ;
        RECT 77.680 113.635 77.935 114.165 ;
        RECT 78.115 113.455 78.400 113.915 ;
        RECT 78.580 113.715 78.830 114.365 ;
        RECT 79.030 115.115 79.350 115.135 ;
        RECT 79.030 114.945 80.950 115.115 ;
        RECT 79.030 114.050 79.220 114.945 ;
        RECT 81.120 114.775 81.290 115.285 ;
        RECT 81.460 115.025 81.980 115.335 ;
        RECT 79.390 114.605 81.290 114.775 ;
        RECT 79.390 114.545 79.720 114.605 ;
        RECT 79.870 114.375 80.200 114.435 ;
        RECT 79.540 114.105 80.200 114.375 ;
        RECT 79.030 113.720 79.350 114.050 ;
        RECT 79.530 113.455 80.190 113.935 ;
        RECT 80.390 113.845 80.560 114.605 ;
        RECT 81.460 114.435 81.640 114.845 ;
        RECT 80.730 114.265 81.060 114.385 ;
        RECT 81.810 114.265 81.980 115.025 ;
        RECT 80.730 114.095 81.980 114.265 ;
        RECT 82.150 115.205 83.520 115.455 ;
        RECT 82.150 114.435 82.340 115.205 ;
        RECT 83.270 114.945 83.520 115.205 ;
        RECT 82.510 114.775 82.760 114.935 ;
        RECT 83.690 114.775 83.860 115.620 ;
        RECT 84.755 115.335 84.925 115.835 ;
        RECT 85.095 115.505 85.425 116.005 ;
        RECT 84.030 114.945 84.530 115.325 ;
        RECT 84.755 115.165 85.450 115.335 ;
        RECT 82.510 114.605 83.860 114.775 ;
        RECT 83.440 114.565 83.860 114.605 ;
        RECT 82.150 114.095 82.570 114.435 ;
        RECT 82.860 114.105 83.270 114.435 ;
        RECT 80.390 113.675 81.240 113.845 ;
        RECT 81.800 113.455 82.120 113.915 ;
        RECT 82.320 113.665 82.570 114.095 ;
        RECT 82.860 113.455 83.270 113.895 ;
        RECT 83.440 113.835 83.610 114.565 ;
        RECT 83.780 114.015 84.130 114.385 ;
        RECT 84.310 114.075 84.530 114.945 ;
        RECT 84.700 114.375 85.110 114.995 ;
        RECT 85.280 114.195 85.450 115.165 ;
        RECT 84.755 114.005 85.450 114.195 ;
        RECT 83.440 113.635 84.455 113.835 ;
        RECT 84.755 113.675 84.925 114.005 ;
        RECT 85.095 113.455 85.425 113.835 ;
        RECT 85.640 113.715 85.865 115.835 ;
        RECT 86.035 115.505 86.365 116.005 ;
        RECT 86.535 115.335 86.705 115.835 ;
        RECT 86.040 115.165 86.705 115.335 ;
        RECT 87.515 115.335 87.685 115.835 ;
        RECT 87.855 115.505 88.185 116.005 ;
        RECT 87.515 115.165 88.180 115.335 ;
        RECT 86.040 114.175 86.270 115.165 ;
        RECT 86.440 114.345 86.790 114.995 ;
        RECT 87.430 114.345 87.780 114.995 ;
        RECT 87.950 114.175 88.180 115.165 ;
        RECT 86.040 114.005 86.705 114.175 ;
        RECT 86.035 113.455 86.365 113.835 ;
        RECT 86.535 113.715 86.705 114.005 ;
        RECT 87.515 114.005 88.180 114.175 ;
        RECT 87.515 113.715 87.685 114.005 ;
        RECT 87.855 113.455 88.185 113.835 ;
        RECT 88.355 113.715 88.580 115.835 ;
        RECT 88.795 115.505 89.125 116.005 ;
        RECT 89.295 115.335 89.465 115.835 ;
        RECT 89.700 115.620 90.530 115.790 ;
        RECT 90.770 115.625 91.150 116.005 ;
        RECT 88.770 115.165 89.465 115.335 ;
        RECT 88.770 114.195 88.940 115.165 ;
        RECT 89.110 114.375 89.520 114.995 ;
        RECT 89.690 114.945 90.190 115.325 ;
        RECT 88.770 114.005 89.465 114.195 ;
        RECT 89.690 114.075 89.910 114.945 ;
        RECT 90.360 114.775 90.530 115.620 ;
        RECT 91.330 115.455 91.500 115.745 ;
        RECT 91.670 115.625 92.000 116.005 ;
        RECT 92.470 115.535 93.100 115.785 ;
        RECT 93.280 115.625 93.700 116.005 ;
        RECT 92.930 115.455 93.100 115.535 ;
        RECT 93.900 115.455 94.140 115.745 ;
        RECT 90.700 115.205 92.070 115.455 ;
        RECT 90.700 114.945 90.950 115.205 ;
        RECT 91.460 114.775 91.710 114.935 ;
        RECT 90.360 114.605 91.710 114.775 ;
        RECT 90.360 114.565 90.780 114.605 ;
        RECT 90.090 114.015 90.440 114.385 ;
        RECT 88.795 113.455 89.125 113.835 ;
        RECT 89.295 113.675 89.465 114.005 ;
        RECT 90.610 113.835 90.780 114.565 ;
        RECT 91.880 114.435 92.070 115.205 ;
        RECT 90.950 114.105 91.360 114.435 ;
        RECT 91.650 114.095 92.070 114.435 ;
        RECT 92.240 115.025 92.760 115.335 ;
        RECT 92.930 115.285 94.140 115.455 ;
        RECT 94.370 115.315 94.700 116.005 ;
        RECT 92.240 114.265 92.410 115.025 ;
        RECT 92.580 114.435 92.760 114.845 ;
        RECT 92.930 114.775 93.100 115.285 ;
        RECT 94.870 115.135 95.040 115.745 ;
        RECT 95.310 115.285 95.640 115.795 ;
        RECT 94.870 115.115 95.190 115.135 ;
        RECT 93.270 114.945 95.190 115.115 ;
        RECT 92.930 114.605 94.830 114.775 ;
        RECT 93.160 114.265 93.490 114.385 ;
        RECT 92.240 114.095 93.490 114.265 ;
        RECT 89.765 113.635 90.780 113.835 ;
        RECT 90.950 113.455 91.360 113.895 ;
        RECT 91.650 113.665 91.900 114.095 ;
        RECT 92.100 113.455 92.420 113.915 ;
        RECT 93.660 113.845 93.830 114.605 ;
        RECT 94.500 114.545 94.830 114.605 ;
        RECT 94.020 114.375 94.350 114.435 ;
        RECT 94.020 114.105 94.680 114.375 ;
        RECT 95.000 114.050 95.190 114.945 ;
        RECT 92.980 113.675 93.830 113.845 ;
        RECT 94.030 113.455 94.690 113.935 ;
        RECT 94.870 113.720 95.190 114.050 ;
        RECT 95.390 114.695 95.640 115.285 ;
        RECT 95.820 115.205 96.105 116.005 ;
        RECT 96.285 115.665 96.540 115.695 ;
        RECT 96.285 115.495 96.625 115.665 ;
        RECT 96.285 115.025 96.540 115.495 ;
        RECT 95.390 114.365 96.190 114.695 ;
        RECT 95.390 113.715 95.640 114.365 ;
        RECT 96.360 114.165 96.540 115.025 ;
        RECT 97.545 114.915 100.135 116.005 ;
        RECT 100.305 114.930 100.575 115.835 ;
        RECT 100.745 115.245 101.075 116.005 ;
        RECT 101.255 115.075 101.425 115.835 ;
        RECT 97.545 114.395 98.755 114.915 ;
        RECT 98.925 114.225 100.135 114.745 ;
        RECT 95.820 113.455 96.105 113.915 ;
        RECT 96.285 113.635 96.540 114.165 ;
        RECT 97.545 113.455 100.135 114.225 ;
        RECT 100.305 114.130 100.475 114.930 ;
        RECT 100.760 114.905 101.425 115.075 ;
        RECT 100.760 114.760 100.930 114.905 ;
        RECT 101.685 114.840 101.975 116.005 ;
        RECT 102.610 115.570 107.955 116.005 ;
        RECT 100.645 114.430 100.930 114.760 ;
        RECT 100.760 114.175 100.930 114.430 ;
        RECT 101.165 114.355 101.495 114.725 ;
        RECT 104.200 114.320 104.550 115.570 ;
        RECT 108.215 115.075 108.385 115.835 ;
        RECT 108.565 115.245 108.895 116.005 ;
        RECT 108.215 114.905 108.880 115.075 ;
        RECT 109.065 114.930 109.335 115.835 ;
        RECT 100.305 113.625 100.565 114.130 ;
        RECT 100.760 114.005 101.425 114.175 ;
        RECT 100.745 113.455 101.075 113.835 ;
        RECT 101.255 113.625 101.425 114.005 ;
        RECT 101.685 113.455 101.975 114.180 ;
        RECT 106.030 114.000 106.370 114.830 ;
        RECT 108.710 114.760 108.880 114.905 ;
        RECT 108.145 114.355 108.475 114.725 ;
        RECT 108.710 114.430 108.995 114.760 ;
        RECT 108.710 114.175 108.880 114.430 ;
        RECT 108.215 114.005 108.880 114.175 ;
        RECT 109.165 114.130 109.335 114.930 ;
        RECT 109.505 114.915 111.175 116.005 ;
        RECT 111.345 115.245 111.860 115.655 ;
        RECT 112.095 115.245 112.265 116.005 ;
        RECT 112.435 115.665 114.465 115.835 ;
        RECT 109.505 114.395 110.255 114.915 ;
        RECT 110.425 114.225 111.175 114.745 ;
        RECT 111.345 114.435 111.685 115.245 ;
        RECT 112.435 115.000 112.605 115.665 ;
        RECT 113.000 115.325 114.125 115.495 ;
        RECT 111.855 114.810 112.605 115.000 ;
        RECT 112.775 114.985 113.785 115.155 ;
        RECT 111.345 114.265 112.575 114.435 ;
        RECT 102.610 113.455 107.955 114.000 ;
        RECT 108.215 113.625 108.385 114.005 ;
        RECT 108.565 113.455 108.895 113.835 ;
        RECT 109.075 113.625 109.335 114.130 ;
        RECT 109.505 113.455 111.175 114.225 ;
        RECT 111.620 113.660 111.865 114.265 ;
        RECT 112.085 113.455 112.595 113.990 ;
        RECT 112.775 113.625 112.965 114.985 ;
        RECT 113.135 114.645 113.410 114.785 ;
        RECT 113.135 114.475 113.415 114.645 ;
        RECT 113.135 113.625 113.410 114.475 ;
        RECT 113.615 114.185 113.785 114.985 ;
        RECT 113.955 114.195 114.125 115.325 ;
        RECT 114.295 114.695 114.465 115.665 ;
        RECT 114.635 114.865 114.805 116.005 ;
        RECT 114.975 114.865 115.310 115.835 ;
        RECT 115.490 115.570 120.835 116.005 ;
        RECT 121.010 115.570 126.355 116.005 ;
        RECT 114.295 114.365 114.490 114.695 ;
        RECT 114.715 114.365 114.970 114.695 ;
        RECT 114.715 114.195 114.885 114.365 ;
        RECT 115.140 114.195 115.310 114.865 ;
        RECT 117.080 114.320 117.430 115.570 ;
        RECT 113.955 114.025 114.885 114.195 ;
        RECT 113.955 113.990 114.130 114.025 ;
        RECT 113.600 113.625 114.130 113.990 ;
        RECT 114.555 113.455 114.885 113.855 ;
        RECT 115.055 113.625 115.310 114.195 ;
        RECT 118.910 114.000 119.250 114.830 ;
        RECT 122.600 114.320 122.950 115.570 ;
        RECT 126.525 114.915 127.735 116.005 ;
        RECT 124.430 114.000 124.770 114.830 ;
        RECT 126.525 114.375 127.045 114.915 ;
        RECT 127.215 114.205 127.735 114.745 ;
        RECT 115.490 113.455 120.835 114.000 ;
        RECT 121.010 113.455 126.355 114.000 ;
        RECT 126.525 113.455 127.735 114.205 ;
        RECT 14.660 113.285 127.820 113.455 ;
        RECT 14.745 112.535 15.955 113.285 ;
        RECT 16.435 112.815 16.605 113.285 ;
        RECT 16.775 112.635 17.105 113.115 ;
        RECT 17.275 112.815 17.445 113.285 ;
        RECT 17.615 112.635 17.945 113.115 ;
        RECT 14.745 111.995 15.265 112.535 ;
        RECT 16.180 112.465 17.945 112.635 ;
        RECT 18.115 112.475 18.285 113.285 ;
        RECT 18.485 112.905 19.555 113.075 ;
        RECT 18.485 112.550 18.805 112.905 ;
        RECT 15.435 111.825 15.955 112.365 ;
        RECT 14.745 110.735 15.955 111.825 ;
        RECT 16.180 111.915 16.590 112.465 ;
        RECT 18.480 112.295 18.805 112.550 ;
        RECT 16.775 112.085 18.805 112.295 ;
        RECT 18.460 112.075 18.805 112.085 ;
        RECT 18.975 112.335 19.215 112.735 ;
        RECT 19.385 112.675 19.555 112.905 ;
        RECT 19.725 112.845 19.915 113.285 ;
        RECT 20.085 112.835 21.035 113.115 ;
        RECT 21.255 112.925 21.605 113.095 ;
        RECT 19.385 112.505 19.915 112.675 ;
        RECT 16.180 111.745 17.905 111.915 ;
        RECT 16.435 110.735 16.605 111.575 ;
        RECT 16.815 110.905 17.065 111.745 ;
        RECT 17.275 110.735 17.445 111.575 ;
        RECT 17.615 110.905 17.905 111.745 ;
        RECT 18.115 110.735 18.285 111.795 ;
        RECT 18.460 111.455 18.630 112.075 ;
        RECT 18.975 111.965 19.515 112.335 ;
        RECT 19.695 112.225 19.915 112.505 ;
        RECT 20.085 112.055 20.255 112.835 ;
        RECT 19.850 111.885 20.255 112.055 ;
        RECT 20.425 112.045 20.775 112.665 ;
        RECT 19.850 111.795 20.020 111.885 ;
        RECT 20.945 111.875 21.155 112.665 ;
        RECT 18.800 111.625 20.020 111.795 ;
        RECT 20.480 111.715 21.155 111.875 ;
        RECT 18.460 111.285 19.260 111.455 ;
        RECT 18.580 110.735 18.910 111.115 ;
        RECT 19.090 110.995 19.260 111.285 ;
        RECT 19.850 111.245 20.020 111.625 ;
        RECT 20.190 111.705 21.155 111.715 ;
        RECT 21.345 112.535 21.605 112.925 ;
        RECT 21.815 112.825 22.145 113.285 ;
        RECT 23.020 112.895 23.875 113.065 ;
        RECT 24.080 112.895 24.575 113.065 ;
        RECT 24.745 112.925 25.075 113.285 ;
        RECT 21.345 111.845 21.515 112.535 ;
        RECT 21.685 112.185 21.855 112.365 ;
        RECT 22.025 112.355 22.815 112.605 ;
        RECT 23.020 112.185 23.190 112.895 ;
        RECT 23.360 112.385 23.715 112.605 ;
        RECT 21.685 112.015 23.375 112.185 ;
        RECT 20.190 111.415 20.650 111.705 ;
        RECT 21.345 111.675 22.845 111.845 ;
        RECT 21.345 111.535 21.515 111.675 ;
        RECT 20.955 111.365 21.515 111.535 ;
        RECT 19.430 110.735 19.680 111.195 ;
        RECT 19.850 110.905 20.720 111.245 ;
        RECT 20.955 110.905 21.125 111.365 ;
        RECT 21.960 111.335 23.035 111.505 ;
        RECT 21.295 110.735 21.665 111.195 ;
        RECT 21.960 110.995 22.130 111.335 ;
        RECT 22.300 110.735 22.630 111.165 ;
        RECT 22.865 110.995 23.035 111.335 ;
        RECT 23.205 111.235 23.375 112.015 ;
        RECT 23.545 111.795 23.715 112.385 ;
        RECT 23.885 111.985 24.235 112.605 ;
        RECT 23.545 111.405 24.010 111.795 ;
        RECT 24.405 111.535 24.575 112.895 ;
        RECT 24.745 111.705 25.205 112.755 ;
        RECT 24.180 111.365 24.575 111.535 ;
        RECT 24.180 111.235 24.350 111.365 ;
        RECT 23.205 110.905 23.885 111.235 ;
        RECT 24.100 110.905 24.350 111.235 ;
        RECT 24.520 110.735 24.770 111.195 ;
        RECT 24.940 110.920 25.265 111.705 ;
        RECT 25.435 110.905 25.605 113.025 ;
        RECT 25.775 112.905 26.105 113.285 ;
        RECT 26.275 112.735 26.530 113.025 ;
        RECT 25.780 112.565 26.530 112.735 ;
        RECT 25.780 111.575 26.010 112.565 ;
        RECT 26.705 112.515 28.375 113.285 ;
        RECT 28.550 112.740 33.895 113.285 ;
        RECT 26.180 111.745 26.530 112.395 ;
        RECT 26.705 111.825 27.455 112.345 ;
        RECT 27.625 111.995 28.375 112.515 ;
        RECT 25.780 111.405 26.530 111.575 ;
        RECT 25.775 110.735 26.105 111.235 ;
        RECT 26.275 110.905 26.530 111.405 ;
        RECT 26.705 110.735 28.375 111.825 ;
        RECT 30.140 111.170 30.490 112.420 ;
        RECT 31.970 111.910 32.310 112.740 ;
        RECT 34.125 112.465 34.335 113.285 ;
        RECT 34.505 112.485 34.835 113.115 ;
        RECT 34.505 111.885 34.755 112.485 ;
        RECT 35.005 112.465 35.235 113.285 ;
        RECT 35.445 112.515 37.115 113.285 ;
        RECT 37.285 112.560 37.575 113.285 ;
        RECT 38.295 112.805 38.595 113.285 ;
        RECT 38.765 112.635 39.025 113.090 ;
        RECT 39.195 112.805 39.455 113.285 ;
        RECT 39.635 112.635 39.895 113.090 ;
        RECT 40.065 112.805 40.315 113.285 ;
        RECT 40.495 112.635 40.755 113.090 ;
        RECT 40.925 112.805 41.175 113.285 ;
        RECT 41.355 112.635 41.615 113.090 ;
        RECT 41.785 112.805 42.030 113.285 ;
        RECT 42.200 112.635 42.475 113.090 ;
        RECT 42.645 112.805 42.890 113.285 ;
        RECT 43.060 112.635 43.320 113.090 ;
        RECT 43.490 112.805 43.750 113.285 ;
        RECT 43.920 112.635 44.180 113.090 ;
        RECT 44.350 112.805 44.610 113.285 ;
        RECT 44.780 112.635 45.040 113.090 ;
        RECT 45.210 112.725 45.470 113.285 ;
        RECT 34.925 112.045 35.255 112.295 ;
        RECT 28.550 110.735 33.895 111.170 ;
        RECT 34.125 110.735 34.335 111.875 ;
        RECT 34.505 110.905 34.835 111.885 ;
        RECT 35.005 110.735 35.235 111.875 ;
        RECT 35.445 111.825 36.195 112.345 ;
        RECT 36.365 111.995 37.115 112.515 ;
        RECT 38.295 112.465 45.040 112.635 ;
        RECT 35.445 110.735 37.115 111.825 ;
        RECT 37.285 110.735 37.575 111.900 ;
        RECT 38.295 111.875 39.460 112.465 ;
        RECT 45.640 112.295 45.890 113.105 ;
        RECT 46.070 112.760 46.330 113.285 ;
        RECT 46.500 112.295 46.750 113.105 ;
        RECT 46.930 112.775 47.235 113.285 ;
        RECT 39.630 112.045 46.750 112.295 ;
        RECT 46.920 112.045 47.235 112.605 ;
        RECT 48.325 112.515 51.835 113.285 ;
        RECT 52.010 112.740 57.355 113.285 ;
        RECT 57.530 112.740 62.875 113.285 ;
        RECT 38.295 111.650 45.040 111.875 ;
        RECT 38.295 110.735 38.565 111.480 ;
        RECT 38.735 110.910 39.025 111.650 ;
        RECT 39.635 111.635 45.040 111.650 ;
        RECT 39.195 110.740 39.450 111.465 ;
        RECT 39.635 110.910 39.895 111.635 ;
        RECT 40.065 110.740 40.310 111.465 ;
        RECT 40.495 110.910 40.755 111.635 ;
        RECT 40.925 110.740 41.170 111.465 ;
        RECT 41.355 110.910 41.615 111.635 ;
        RECT 41.785 110.740 42.030 111.465 ;
        RECT 42.200 110.910 42.460 111.635 ;
        RECT 42.630 110.740 42.890 111.465 ;
        RECT 43.060 110.910 43.320 111.635 ;
        RECT 43.490 110.740 43.750 111.465 ;
        RECT 43.920 110.910 44.180 111.635 ;
        RECT 44.350 110.740 44.610 111.465 ;
        RECT 44.780 110.910 45.040 111.635 ;
        RECT 45.210 110.740 45.470 111.535 ;
        RECT 45.640 110.910 45.890 112.045 ;
        RECT 39.195 110.735 45.470 110.740 ;
        RECT 46.070 110.735 46.330 111.545 ;
        RECT 46.505 110.905 46.750 112.045 ;
        RECT 48.325 111.825 50.015 112.345 ;
        RECT 50.185 111.995 51.835 112.515 ;
        RECT 46.930 110.735 47.225 111.545 ;
        RECT 48.325 110.735 51.835 111.825 ;
        RECT 53.600 111.170 53.950 112.420 ;
        RECT 55.430 111.910 55.770 112.740 ;
        RECT 59.120 111.170 59.470 112.420 ;
        RECT 60.950 111.910 61.290 112.740 ;
        RECT 63.045 112.560 63.335 113.285 ;
        RECT 63.970 112.740 69.315 113.285 ;
        RECT 69.490 112.740 74.835 113.285 ;
        RECT 75.010 112.740 80.355 113.285 ;
        RECT 52.010 110.735 57.355 111.170 ;
        RECT 57.530 110.735 62.875 111.170 ;
        RECT 63.045 110.735 63.335 111.900 ;
        RECT 65.560 111.170 65.910 112.420 ;
        RECT 67.390 111.910 67.730 112.740 ;
        RECT 71.080 111.170 71.430 112.420 ;
        RECT 72.910 111.910 73.250 112.740 ;
        RECT 76.600 111.170 76.950 112.420 ;
        RECT 78.430 111.910 78.770 112.740 ;
        RECT 80.585 112.465 80.795 113.285 ;
        RECT 80.965 112.485 81.295 113.115 ;
        RECT 80.965 111.885 81.215 112.485 ;
        RECT 81.465 112.465 81.695 113.285 ;
        RECT 81.905 112.535 83.115 113.285 ;
        RECT 83.290 112.740 88.635 113.285 ;
        RECT 81.385 112.045 81.715 112.295 ;
        RECT 63.970 110.735 69.315 111.170 ;
        RECT 69.490 110.735 74.835 111.170 ;
        RECT 75.010 110.735 80.355 111.170 ;
        RECT 80.585 110.735 80.795 111.875 ;
        RECT 80.965 110.905 81.295 111.885 ;
        RECT 81.465 110.735 81.695 111.875 ;
        RECT 81.905 111.825 82.425 112.365 ;
        RECT 82.595 111.995 83.115 112.535 ;
        RECT 81.905 110.735 83.115 111.825 ;
        RECT 84.880 111.170 85.230 112.420 ;
        RECT 86.710 111.910 87.050 112.740 ;
        RECT 88.805 112.560 89.095 113.285 ;
        RECT 89.265 112.515 92.775 113.285 ;
        RECT 92.945 112.775 93.250 113.285 ;
        RECT 83.290 110.735 88.635 111.170 ;
        RECT 88.805 110.735 89.095 111.900 ;
        RECT 89.265 111.825 90.955 112.345 ;
        RECT 91.125 111.995 92.775 112.515 ;
        RECT 92.945 112.045 93.260 112.605 ;
        RECT 93.430 112.295 93.680 113.105 ;
        RECT 93.850 112.760 94.110 113.285 ;
        RECT 94.290 112.295 94.540 113.105 ;
        RECT 94.710 112.725 94.970 113.285 ;
        RECT 95.140 112.635 95.400 113.090 ;
        RECT 95.570 112.805 95.830 113.285 ;
        RECT 96.000 112.635 96.260 113.090 ;
        RECT 96.430 112.805 96.690 113.285 ;
        RECT 96.860 112.635 97.120 113.090 ;
        RECT 97.290 112.805 97.535 113.285 ;
        RECT 97.705 112.635 97.980 113.090 ;
        RECT 98.150 112.805 98.395 113.285 ;
        RECT 98.565 112.635 98.825 113.090 ;
        RECT 99.005 112.805 99.255 113.285 ;
        RECT 99.425 112.635 99.685 113.090 ;
        RECT 99.865 112.805 100.115 113.285 ;
        RECT 100.285 112.635 100.545 113.090 ;
        RECT 100.725 112.805 100.985 113.285 ;
        RECT 101.155 112.635 101.415 113.090 ;
        RECT 101.585 112.805 101.885 113.285 ;
        RECT 102.145 112.780 102.430 113.285 ;
        RECT 95.140 112.605 101.885 112.635 ;
        RECT 102.600 112.610 102.925 113.115 ;
        RECT 95.140 112.465 101.915 112.605 ;
        RECT 100.720 112.435 101.915 112.465 ;
        RECT 93.430 112.045 100.550 112.295 ;
        RECT 89.265 110.735 92.775 111.825 ;
        RECT 92.955 110.735 93.250 111.545 ;
        RECT 93.430 110.905 93.675 112.045 ;
        RECT 93.850 110.735 94.110 111.545 ;
        RECT 94.290 110.910 94.540 112.045 ;
        RECT 100.720 111.875 101.885 112.435 ;
        RECT 102.145 112.080 102.925 112.610 ;
        RECT 95.140 111.650 101.885 111.875 ;
        RECT 95.140 111.635 100.545 111.650 ;
        RECT 94.710 110.740 94.970 111.535 ;
        RECT 95.140 110.910 95.400 111.635 ;
        RECT 95.570 110.740 95.830 111.465 ;
        RECT 96.000 110.910 96.260 111.635 ;
        RECT 96.430 110.740 96.690 111.465 ;
        RECT 96.860 110.910 97.120 111.635 ;
        RECT 97.290 110.740 97.550 111.465 ;
        RECT 97.720 110.910 97.980 111.635 ;
        RECT 98.150 110.740 98.395 111.465 ;
        RECT 98.565 110.910 98.825 111.635 ;
        RECT 99.010 110.740 99.255 111.465 ;
        RECT 99.425 110.910 99.685 111.635 ;
        RECT 99.870 110.740 100.115 111.465 ;
        RECT 100.285 110.910 100.545 111.635 ;
        RECT 100.730 110.740 100.985 111.465 ;
        RECT 101.155 110.910 101.445 111.650 ;
        RECT 94.710 110.735 100.985 110.740 ;
        RECT 101.615 110.735 101.885 111.480 ;
        RECT 102.145 110.735 102.425 111.705 ;
        RECT 102.595 110.905 102.925 112.080 ;
        RECT 103.115 112.045 103.355 112.995 ;
        RECT 103.530 112.740 108.875 113.285 ;
        RECT 109.050 112.740 114.395 113.285 ;
        RECT 103.095 110.735 103.355 111.705 ;
        RECT 105.120 111.170 105.470 112.420 ;
        RECT 106.950 111.910 107.290 112.740 ;
        RECT 110.640 111.170 110.990 112.420 ;
        RECT 112.470 111.910 112.810 112.740 ;
        RECT 114.565 112.560 114.855 113.285 ;
        RECT 115.945 112.515 119.455 113.285 ;
        RECT 103.530 110.735 108.875 111.170 ;
        RECT 109.050 110.735 114.395 111.170 ;
        RECT 114.565 110.735 114.855 111.900 ;
        RECT 115.945 111.825 117.635 112.345 ;
        RECT 117.805 111.995 119.455 112.515 ;
        RECT 119.665 112.465 119.895 113.285 ;
        RECT 120.065 112.485 120.395 113.115 ;
        RECT 119.645 112.045 119.975 112.295 ;
        RECT 120.145 111.885 120.395 112.485 ;
        RECT 120.565 112.465 120.775 113.285 ;
        RECT 121.005 112.610 121.265 113.115 ;
        RECT 121.445 112.905 121.775 113.285 ;
        RECT 121.955 112.735 122.125 113.115 ;
        RECT 115.945 110.735 119.455 111.825 ;
        RECT 119.665 110.735 119.895 111.875 ;
        RECT 120.065 110.905 120.395 111.885 ;
        RECT 120.565 110.735 120.775 111.875 ;
        RECT 121.005 111.810 121.175 112.610 ;
        RECT 121.460 112.565 122.125 112.735 ;
        RECT 122.385 112.610 122.645 113.115 ;
        RECT 122.825 112.905 123.155 113.285 ;
        RECT 123.335 112.735 123.505 113.115 ;
        RECT 121.460 112.310 121.630 112.565 ;
        RECT 121.345 111.980 121.630 112.310 ;
        RECT 121.865 112.015 122.195 112.385 ;
        RECT 121.460 111.835 121.630 111.980 ;
        RECT 121.005 110.905 121.275 111.810 ;
        RECT 121.460 111.665 122.125 111.835 ;
        RECT 121.445 110.735 121.775 111.495 ;
        RECT 121.955 110.905 122.125 111.665 ;
        RECT 122.385 111.810 122.555 112.610 ;
        RECT 122.840 112.565 123.505 112.735 ;
        RECT 122.840 112.310 123.010 112.565 ;
        RECT 123.765 112.515 126.355 113.285 ;
        RECT 126.525 112.535 127.735 113.285 ;
        RECT 122.725 111.980 123.010 112.310 ;
        RECT 123.245 112.015 123.575 112.385 ;
        RECT 122.840 111.835 123.010 111.980 ;
        RECT 122.385 110.905 122.655 111.810 ;
        RECT 122.840 111.665 123.505 111.835 ;
        RECT 122.825 110.735 123.155 111.495 ;
        RECT 123.335 110.905 123.505 111.665 ;
        RECT 123.765 111.825 124.975 112.345 ;
        RECT 125.145 111.995 126.355 112.515 ;
        RECT 126.525 111.825 127.045 112.365 ;
        RECT 127.215 111.995 127.735 112.535 ;
        RECT 123.765 110.735 126.355 111.825 ;
        RECT 126.525 110.735 127.735 111.825 ;
        RECT 14.660 110.565 127.820 110.735 ;
        RECT 14.745 109.475 15.955 110.565 ;
        RECT 14.745 108.765 15.265 109.305 ;
        RECT 15.435 108.935 15.955 109.475 ;
        RECT 17.045 109.475 20.555 110.565 ;
        RECT 17.045 108.955 18.735 109.475 ;
        RECT 20.785 109.425 20.995 110.565 ;
        RECT 21.165 109.415 21.495 110.395 ;
        RECT 21.665 109.425 21.895 110.565 ;
        RECT 23.085 109.425 23.295 110.565 ;
        RECT 23.465 109.415 23.795 110.395 ;
        RECT 23.965 109.425 24.195 110.565 ;
        RECT 18.905 108.785 20.555 109.305 ;
        RECT 14.745 108.015 15.955 108.765 ;
        RECT 17.045 108.015 20.555 108.785 ;
        RECT 20.785 108.015 20.995 108.835 ;
        RECT 21.165 108.815 21.415 109.415 ;
        RECT 21.585 109.005 21.915 109.255 ;
        RECT 21.165 108.185 21.495 108.815 ;
        RECT 21.665 108.015 21.895 108.835 ;
        RECT 23.085 108.015 23.295 108.835 ;
        RECT 23.465 108.815 23.715 109.415 ;
        RECT 24.405 109.400 24.695 110.565 ;
        RECT 24.865 109.475 27.455 110.565 ;
        RECT 27.625 109.490 27.895 110.395 ;
        RECT 28.065 109.805 28.395 110.565 ;
        RECT 28.575 109.635 28.745 110.395 ;
        RECT 23.885 109.005 24.215 109.255 ;
        RECT 24.865 108.955 26.075 109.475 ;
        RECT 23.465 108.185 23.795 108.815 ;
        RECT 23.965 108.015 24.195 108.835 ;
        RECT 26.245 108.785 27.455 109.305 ;
        RECT 24.405 108.015 24.695 108.740 ;
        RECT 24.865 108.015 27.455 108.785 ;
        RECT 27.625 108.690 27.795 109.490 ;
        RECT 28.080 109.465 28.745 109.635 ;
        RECT 29.005 109.475 30.675 110.565 ;
        RECT 28.080 109.320 28.250 109.465 ;
        RECT 27.965 108.990 28.250 109.320 ;
        RECT 28.080 108.735 28.250 108.990 ;
        RECT 28.485 108.915 28.815 109.285 ;
        RECT 29.005 108.955 29.755 109.475 ;
        RECT 30.905 109.425 31.115 110.565 ;
        RECT 31.285 109.415 31.615 110.395 ;
        RECT 31.785 109.425 32.015 110.565 ;
        RECT 32.225 109.490 32.495 110.395 ;
        RECT 32.665 109.805 32.995 110.565 ;
        RECT 33.175 109.635 33.345 110.395 ;
        RECT 29.925 108.785 30.675 109.305 ;
        RECT 27.625 108.185 27.885 108.690 ;
        RECT 28.080 108.565 28.745 108.735 ;
        RECT 28.065 108.015 28.395 108.395 ;
        RECT 28.575 108.185 28.745 108.565 ;
        RECT 29.005 108.015 30.675 108.785 ;
        RECT 30.905 108.015 31.115 108.835 ;
        RECT 31.285 108.815 31.535 109.415 ;
        RECT 31.705 109.005 32.035 109.255 ;
        RECT 31.285 108.185 31.615 108.815 ;
        RECT 31.785 108.015 32.015 108.835 ;
        RECT 32.225 108.690 32.395 109.490 ;
        RECT 32.680 109.465 33.345 109.635 ;
        RECT 34.525 109.490 34.795 110.395 ;
        RECT 34.965 109.805 35.295 110.565 ;
        RECT 35.475 109.635 35.645 110.395 ;
        RECT 32.680 109.320 32.850 109.465 ;
        RECT 32.565 108.990 32.850 109.320 ;
        RECT 32.680 108.735 32.850 108.990 ;
        RECT 33.085 108.915 33.415 109.285 ;
        RECT 32.225 108.185 32.485 108.690 ;
        RECT 32.680 108.565 33.345 108.735 ;
        RECT 32.665 108.015 32.995 108.395 ;
        RECT 33.175 108.185 33.345 108.565 ;
        RECT 34.525 108.690 34.695 109.490 ;
        RECT 34.980 109.465 35.645 109.635 ;
        RECT 36.365 109.475 38.955 110.565 ;
        RECT 39.130 110.130 44.475 110.565 ;
        RECT 44.650 110.130 49.995 110.565 ;
        RECT 34.980 109.320 35.150 109.465 ;
        RECT 34.865 108.990 35.150 109.320 ;
        RECT 34.980 108.735 35.150 108.990 ;
        RECT 35.385 108.915 35.715 109.285 ;
        RECT 36.365 108.955 37.575 109.475 ;
        RECT 37.745 108.785 38.955 109.305 ;
        RECT 40.720 108.880 41.070 110.130 ;
        RECT 34.525 108.185 34.785 108.690 ;
        RECT 34.980 108.565 35.645 108.735 ;
        RECT 34.965 108.015 35.295 108.395 ;
        RECT 35.475 108.185 35.645 108.565 ;
        RECT 36.365 108.015 38.955 108.785 ;
        RECT 42.550 108.560 42.890 109.390 ;
        RECT 46.240 108.880 46.590 110.130 ;
        RECT 50.165 109.400 50.455 110.565 ;
        RECT 51.175 109.635 51.345 110.395 ;
        RECT 51.525 109.805 51.855 110.565 ;
        RECT 51.175 109.465 51.840 109.635 ;
        RECT 52.025 109.490 52.295 110.395 ;
        RECT 48.070 108.560 48.410 109.390 ;
        RECT 51.670 109.320 51.840 109.465 ;
        RECT 51.105 108.915 51.435 109.285 ;
        RECT 51.670 108.990 51.955 109.320 ;
        RECT 39.130 108.015 44.475 108.560 ;
        RECT 44.650 108.015 49.995 108.560 ;
        RECT 50.165 108.015 50.455 108.740 ;
        RECT 51.670 108.735 51.840 108.990 ;
        RECT 51.175 108.565 51.840 108.735 ;
        RECT 52.125 108.690 52.295 109.490 ;
        RECT 53.385 109.475 56.895 110.565 ;
        RECT 57.155 109.635 57.325 110.395 ;
        RECT 57.505 109.805 57.835 110.565 ;
        RECT 53.385 108.955 55.075 109.475 ;
        RECT 57.155 109.465 57.820 109.635 ;
        RECT 58.005 109.490 58.275 110.395 ;
        RECT 57.650 109.320 57.820 109.465 ;
        RECT 55.245 108.785 56.895 109.305 ;
        RECT 57.085 108.915 57.415 109.285 ;
        RECT 57.650 108.990 57.935 109.320 ;
        RECT 51.175 108.185 51.345 108.565 ;
        RECT 51.525 108.015 51.855 108.395 ;
        RECT 52.035 108.185 52.295 108.690 ;
        RECT 53.385 108.015 56.895 108.785 ;
        RECT 57.650 108.735 57.820 108.990 ;
        RECT 57.155 108.565 57.820 108.735 ;
        RECT 58.105 108.690 58.275 109.490 ;
        RECT 58.445 109.475 59.655 110.565 ;
        RECT 59.835 109.585 60.165 110.395 ;
        RECT 60.335 109.765 60.575 110.565 ;
        RECT 58.445 108.935 58.965 109.475 ;
        RECT 59.835 109.415 60.550 109.585 ;
        RECT 59.135 108.765 59.655 109.305 ;
        RECT 59.830 109.005 60.210 109.245 ;
        RECT 60.380 109.175 60.550 109.415 ;
        RECT 60.755 109.545 60.925 110.395 ;
        RECT 61.095 109.765 61.425 110.565 ;
        RECT 61.595 109.545 61.765 110.395 ;
        RECT 60.755 109.375 61.765 109.545 ;
        RECT 61.935 109.415 62.265 110.565 ;
        RECT 63.045 109.475 64.715 110.565 ;
        RECT 61.270 109.205 61.765 109.375 ;
        RECT 60.380 109.005 60.880 109.175 ;
        RECT 61.265 109.035 61.765 109.205 ;
        RECT 60.380 108.835 60.550 109.005 ;
        RECT 61.270 108.835 61.765 109.035 ;
        RECT 63.045 108.955 63.795 109.475 ;
        RECT 64.925 109.425 65.155 110.565 ;
        RECT 65.325 109.415 65.655 110.395 ;
        RECT 65.825 109.425 66.035 110.565 ;
        RECT 66.725 109.475 68.395 110.565 ;
        RECT 68.655 109.635 68.825 110.395 ;
        RECT 69.005 109.805 69.335 110.565 ;
        RECT 57.155 108.185 57.325 108.565 ;
        RECT 57.505 108.015 57.835 108.395 ;
        RECT 58.015 108.185 58.275 108.690 ;
        RECT 58.445 108.015 59.655 108.765 ;
        RECT 59.915 108.665 60.550 108.835 ;
        RECT 60.755 108.665 61.765 108.835 ;
        RECT 59.915 108.185 60.085 108.665 ;
        RECT 60.265 108.015 60.505 108.495 ;
        RECT 60.755 108.185 60.925 108.665 ;
        RECT 61.095 108.015 61.425 108.495 ;
        RECT 61.595 108.185 61.765 108.665 ;
        RECT 61.935 108.015 62.265 108.815 ;
        RECT 63.965 108.785 64.715 109.305 ;
        RECT 64.905 109.005 65.235 109.255 ;
        RECT 63.045 108.015 64.715 108.785 ;
        RECT 64.925 108.015 65.155 108.835 ;
        RECT 65.405 108.815 65.655 109.415 ;
        RECT 66.725 108.955 67.475 109.475 ;
        RECT 68.655 109.465 69.320 109.635 ;
        RECT 69.505 109.490 69.775 110.395 ;
        RECT 70.410 110.130 75.755 110.565 ;
        RECT 69.150 109.320 69.320 109.465 ;
        RECT 65.325 108.185 65.655 108.815 ;
        RECT 65.825 108.015 66.035 108.835 ;
        RECT 67.645 108.785 68.395 109.305 ;
        RECT 68.585 108.915 68.915 109.285 ;
        RECT 69.150 108.990 69.435 109.320 ;
        RECT 66.725 108.015 68.395 108.785 ;
        RECT 69.150 108.735 69.320 108.990 ;
        RECT 68.655 108.565 69.320 108.735 ;
        RECT 69.605 108.690 69.775 109.490 ;
        RECT 72.000 108.880 72.350 110.130 ;
        RECT 75.925 109.400 76.215 110.565 ;
        RECT 76.445 109.425 76.655 110.565 ;
        RECT 76.825 109.415 77.155 110.395 ;
        RECT 77.325 109.425 77.555 110.565 ;
        RECT 77.825 109.425 78.035 110.565 ;
        RECT 78.205 109.415 78.535 110.395 ;
        RECT 78.705 109.425 78.935 110.565 ;
        RECT 80.075 109.585 80.405 110.395 ;
        RECT 80.575 109.765 80.815 110.565 ;
        RECT 80.075 109.415 80.790 109.585 ;
        RECT 68.655 108.185 68.825 108.565 ;
        RECT 69.005 108.015 69.335 108.395 ;
        RECT 69.515 108.185 69.775 108.690 ;
        RECT 73.830 108.560 74.170 109.390 ;
        RECT 70.410 108.015 75.755 108.560 ;
        RECT 75.925 108.015 76.215 108.740 ;
        RECT 76.445 108.015 76.655 108.835 ;
        RECT 76.825 108.815 77.075 109.415 ;
        RECT 77.245 109.005 77.575 109.255 ;
        RECT 76.825 108.185 77.155 108.815 ;
        RECT 77.325 108.015 77.555 108.835 ;
        RECT 77.825 108.015 78.035 108.835 ;
        RECT 78.205 108.815 78.455 109.415 ;
        RECT 78.625 109.005 78.955 109.255 ;
        RECT 80.070 109.005 80.450 109.245 ;
        RECT 80.620 109.175 80.790 109.415 ;
        RECT 80.995 109.545 81.165 110.395 ;
        RECT 81.335 109.765 81.665 110.565 ;
        RECT 81.835 109.545 82.005 110.395 ;
        RECT 80.995 109.375 82.005 109.545 ;
        RECT 82.175 109.415 82.505 110.565 ;
        RECT 82.915 109.635 83.085 110.395 ;
        RECT 83.265 109.805 83.595 110.565 ;
        RECT 82.915 109.465 83.580 109.635 ;
        RECT 83.765 109.490 84.035 110.395 ;
        RECT 80.620 109.005 81.120 109.175 ;
        RECT 80.620 108.835 80.790 109.005 ;
        RECT 81.510 108.835 82.005 109.375 ;
        RECT 83.410 109.320 83.580 109.465 ;
        RECT 82.845 108.915 83.175 109.285 ;
        RECT 83.410 108.990 83.695 109.320 ;
        RECT 78.205 108.185 78.535 108.815 ;
        RECT 78.705 108.015 78.935 108.835 ;
        RECT 80.155 108.665 80.790 108.835 ;
        RECT 80.995 108.665 82.005 108.835 ;
        RECT 80.155 108.185 80.325 108.665 ;
        RECT 80.505 108.015 80.745 108.495 ;
        RECT 80.995 108.185 81.165 108.665 ;
        RECT 81.335 108.015 81.665 108.495 ;
        RECT 81.835 108.185 82.005 108.665 ;
        RECT 82.175 108.015 82.505 108.815 ;
        RECT 83.410 108.735 83.580 108.990 ;
        RECT 82.915 108.565 83.580 108.735 ;
        RECT 83.865 108.690 84.035 109.490 ;
        RECT 84.665 109.475 87.255 110.565 ;
        RECT 84.665 108.955 85.875 109.475 ;
        RECT 87.465 109.425 87.695 110.565 ;
        RECT 87.865 109.415 88.195 110.395 ;
        RECT 88.365 109.425 88.575 110.565 ;
        RECT 88.805 109.475 92.315 110.565 ;
        RECT 86.045 108.785 87.255 109.305 ;
        RECT 87.445 109.005 87.775 109.255 ;
        RECT 82.915 108.185 83.085 108.565 ;
        RECT 83.265 108.015 83.595 108.395 ;
        RECT 83.775 108.185 84.035 108.690 ;
        RECT 84.665 108.015 87.255 108.785 ;
        RECT 87.465 108.015 87.695 108.835 ;
        RECT 87.945 108.815 88.195 109.415 ;
        RECT 88.805 108.955 90.495 109.475 ;
        RECT 92.525 109.425 92.755 110.565 ;
        RECT 92.925 109.415 93.255 110.395 ;
        RECT 93.425 109.425 93.635 110.565 ;
        RECT 93.955 109.635 94.125 110.395 ;
        RECT 94.305 109.805 94.635 110.565 ;
        RECT 93.955 109.465 94.620 109.635 ;
        RECT 94.805 109.490 95.075 110.395 ;
        RECT 87.865 108.185 88.195 108.815 ;
        RECT 88.365 108.015 88.575 108.835 ;
        RECT 90.665 108.785 92.315 109.305 ;
        RECT 92.505 109.005 92.835 109.255 ;
        RECT 88.805 108.015 92.315 108.785 ;
        RECT 92.525 108.015 92.755 108.835 ;
        RECT 93.005 108.815 93.255 109.415 ;
        RECT 94.450 109.320 94.620 109.465 ;
        RECT 93.885 108.915 94.215 109.285 ;
        RECT 94.450 108.990 94.735 109.320 ;
        RECT 92.925 108.185 93.255 108.815 ;
        RECT 93.425 108.015 93.635 108.835 ;
        RECT 94.450 108.735 94.620 108.990 ;
        RECT 93.955 108.565 94.620 108.735 ;
        RECT 94.905 108.690 95.075 109.490 ;
        RECT 95.245 109.475 96.455 110.565 ;
        RECT 96.625 109.475 100.135 110.565 ;
        RECT 100.305 109.490 100.575 110.395 ;
        RECT 100.745 109.805 101.075 110.565 ;
        RECT 101.255 109.635 101.425 110.395 ;
        RECT 95.245 108.935 95.765 109.475 ;
        RECT 95.935 108.765 96.455 109.305 ;
        RECT 96.625 108.955 98.315 109.475 ;
        RECT 98.485 108.785 100.135 109.305 ;
        RECT 93.955 108.185 94.125 108.565 ;
        RECT 94.305 108.015 94.635 108.395 ;
        RECT 94.815 108.185 95.075 108.690 ;
        RECT 95.245 108.015 96.455 108.765 ;
        RECT 96.625 108.015 100.135 108.785 ;
        RECT 100.305 108.690 100.475 109.490 ;
        RECT 100.760 109.465 101.425 109.635 ;
        RECT 100.760 109.320 100.930 109.465 ;
        RECT 101.685 109.400 101.975 110.565 ;
        RECT 102.605 109.475 106.115 110.565 ;
        RECT 106.375 109.635 106.545 110.395 ;
        RECT 106.725 109.805 107.055 110.565 ;
        RECT 100.645 108.990 100.930 109.320 ;
        RECT 100.760 108.735 100.930 108.990 ;
        RECT 101.165 108.915 101.495 109.285 ;
        RECT 102.605 108.955 104.295 109.475 ;
        RECT 106.375 109.465 107.040 109.635 ;
        RECT 107.225 109.490 107.495 110.395 ;
        RECT 106.870 109.320 107.040 109.465 ;
        RECT 104.465 108.785 106.115 109.305 ;
        RECT 106.305 108.915 106.635 109.285 ;
        RECT 106.870 108.990 107.155 109.320 ;
        RECT 100.305 108.185 100.565 108.690 ;
        RECT 100.760 108.565 101.425 108.735 ;
        RECT 100.745 108.015 101.075 108.395 ;
        RECT 101.255 108.185 101.425 108.565 ;
        RECT 101.685 108.015 101.975 108.740 ;
        RECT 102.605 108.015 106.115 108.785 ;
        RECT 106.870 108.735 107.040 108.990 ;
        RECT 106.375 108.565 107.040 108.735 ;
        RECT 107.325 108.690 107.495 109.490 ;
        RECT 107.665 109.475 108.875 110.565 ;
        RECT 107.665 108.935 108.185 109.475 ;
        RECT 109.105 109.425 109.315 110.565 ;
        RECT 109.485 109.415 109.815 110.395 ;
        RECT 109.985 109.425 110.215 110.565 ;
        RECT 110.515 109.635 110.685 110.395 ;
        RECT 110.865 109.805 111.195 110.565 ;
        RECT 110.515 109.465 111.180 109.635 ;
        RECT 111.365 109.490 111.635 110.395 ;
        RECT 108.355 108.765 108.875 109.305 ;
        RECT 106.375 108.185 106.545 108.565 ;
        RECT 106.725 108.015 107.055 108.395 ;
        RECT 107.235 108.185 107.495 108.690 ;
        RECT 107.665 108.015 108.875 108.765 ;
        RECT 109.105 108.015 109.315 108.835 ;
        RECT 109.485 108.815 109.735 109.415 ;
        RECT 111.010 109.320 111.180 109.465 ;
        RECT 109.905 109.005 110.235 109.255 ;
        RECT 110.445 108.915 110.775 109.285 ;
        RECT 111.010 108.990 111.295 109.320 ;
        RECT 109.485 108.185 109.815 108.815 ;
        RECT 109.985 108.015 110.215 108.835 ;
        RECT 111.010 108.735 111.180 108.990 ;
        RECT 110.515 108.565 111.180 108.735 ;
        RECT 111.465 108.690 111.635 109.490 ;
        RECT 111.895 109.635 112.065 110.395 ;
        RECT 112.245 109.805 112.575 110.565 ;
        RECT 111.895 109.465 112.560 109.635 ;
        RECT 112.745 109.490 113.015 110.395 ;
        RECT 112.390 109.320 112.560 109.465 ;
        RECT 111.825 108.915 112.155 109.285 ;
        RECT 112.390 108.990 112.675 109.320 ;
        RECT 112.390 108.735 112.560 108.990 ;
        RECT 110.515 108.185 110.685 108.565 ;
        RECT 110.865 108.015 111.195 108.395 ;
        RECT 111.375 108.185 111.635 108.690 ;
        RECT 111.895 108.565 112.560 108.735 ;
        RECT 112.845 108.690 113.015 109.490 ;
        RECT 113.185 109.475 114.395 110.565 ;
        RECT 113.185 108.935 113.705 109.475 ;
        RECT 114.605 109.425 114.835 110.565 ;
        RECT 115.005 109.415 115.335 110.395 ;
        RECT 115.505 109.425 115.715 110.565 ;
        RECT 115.950 109.895 116.205 110.395 ;
        RECT 116.375 110.065 116.705 110.565 ;
        RECT 115.950 109.725 116.700 109.895 ;
        RECT 113.875 108.765 114.395 109.305 ;
        RECT 114.585 109.005 114.915 109.255 ;
        RECT 111.895 108.185 112.065 108.565 ;
        RECT 112.245 108.015 112.575 108.395 ;
        RECT 112.755 108.185 113.015 108.690 ;
        RECT 113.185 108.015 114.395 108.765 ;
        RECT 114.605 108.015 114.835 108.835 ;
        RECT 115.085 108.815 115.335 109.415 ;
        RECT 115.950 108.905 116.300 109.555 ;
        RECT 115.005 108.185 115.335 108.815 ;
        RECT 115.505 108.015 115.715 108.835 ;
        RECT 116.470 108.735 116.700 109.725 ;
        RECT 115.950 108.565 116.700 108.735 ;
        RECT 115.950 108.275 116.205 108.565 ;
        RECT 116.375 108.015 116.705 108.395 ;
        RECT 116.875 108.275 117.045 110.395 ;
        RECT 117.215 109.595 117.540 110.380 ;
        RECT 117.710 110.105 117.960 110.565 ;
        RECT 118.130 110.065 118.380 110.395 ;
        RECT 118.595 110.065 119.275 110.395 ;
        RECT 118.130 109.935 118.300 110.065 ;
        RECT 117.905 109.765 118.300 109.935 ;
        RECT 117.275 108.545 117.735 109.595 ;
        RECT 117.905 108.405 118.075 109.765 ;
        RECT 118.470 109.505 118.935 109.895 ;
        RECT 118.245 108.695 118.595 109.315 ;
        RECT 118.765 108.915 118.935 109.505 ;
        RECT 119.105 109.285 119.275 110.065 ;
        RECT 119.445 109.965 119.615 110.305 ;
        RECT 119.850 110.135 120.180 110.565 ;
        RECT 120.350 109.965 120.520 110.305 ;
        RECT 120.815 110.105 121.185 110.565 ;
        RECT 119.445 109.795 120.520 109.965 ;
        RECT 121.355 109.935 121.525 110.395 ;
        RECT 121.760 110.055 122.630 110.395 ;
        RECT 122.800 110.105 123.050 110.565 ;
        RECT 120.965 109.765 121.525 109.935 ;
        RECT 120.965 109.625 121.135 109.765 ;
        RECT 119.635 109.455 121.135 109.625 ;
        RECT 121.830 109.595 122.290 109.885 ;
        RECT 119.105 109.115 120.795 109.285 ;
        RECT 118.765 108.695 119.120 108.915 ;
        RECT 119.290 108.405 119.460 109.115 ;
        RECT 119.665 108.695 120.455 108.945 ;
        RECT 120.625 108.935 120.795 109.115 ;
        RECT 120.965 108.765 121.135 109.455 ;
        RECT 117.405 108.015 117.735 108.375 ;
        RECT 117.905 108.235 118.400 108.405 ;
        RECT 118.605 108.235 119.460 108.405 ;
        RECT 120.335 108.015 120.665 108.475 ;
        RECT 120.875 108.375 121.135 108.765 ;
        RECT 121.325 109.585 122.290 109.595 ;
        RECT 122.460 109.675 122.630 110.055 ;
        RECT 123.220 110.015 123.390 110.305 ;
        RECT 123.570 110.185 123.900 110.565 ;
        RECT 123.220 109.845 124.020 110.015 ;
        RECT 121.325 109.425 122.000 109.585 ;
        RECT 122.460 109.505 123.680 109.675 ;
        RECT 121.325 108.635 121.535 109.425 ;
        RECT 122.460 109.415 122.630 109.505 ;
        RECT 121.705 108.635 122.055 109.255 ;
        RECT 122.225 109.245 122.630 109.415 ;
        RECT 122.225 108.465 122.395 109.245 ;
        RECT 122.565 108.795 122.785 109.075 ;
        RECT 122.965 108.965 123.505 109.335 ;
        RECT 123.850 109.225 124.020 109.845 ;
        RECT 124.195 109.505 124.365 110.565 ;
        RECT 124.575 109.555 124.865 110.395 ;
        RECT 125.035 109.725 125.205 110.565 ;
        RECT 125.415 109.555 125.665 110.395 ;
        RECT 125.875 109.725 126.045 110.565 ;
        RECT 124.575 109.385 126.300 109.555 ;
        RECT 122.565 108.625 123.095 108.795 ;
        RECT 120.875 108.205 121.225 108.375 ;
        RECT 121.445 108.185 122.395 108.465 ;
        RECT 122.565 108.015 122.755 108.455 ;
        RECT 122.925 108.395 123.095 108.625 ;
        RECT 123.265 108.565 123.505 108.965 ;
        RECT 123.675 109.215 124.020 109.225 ;
        RECT 123.675 109.005 125.705 109.215 ;
        RECT 123.675 108.750 124.000 109.005 ;
        RECT 125.890 108.835 126.300 109.385 ;
        RECT 126.525 109.475 127.735 110.565 ;
        RECT 126.525 108.935 127.045 109.475 ;
        RECT 123.675 108.395 123.995 108.750 ;
        RECT 122.925 108.225 123.995 108.395 ;
        RECT 124.195 108.015 124.365 108.825 ;
        RECT 124.535 108.665 126.300 108.835 ;
        RECT 127.215 108.765 127.735 109.305 ;
        RECT 124.535 108.185 124.865 108.665 ;
        RECT 125.035 108.015 125.205 108.485 ;
        RECT 125.375 108.185 125.705 108.665 ;
        RECT 125.875 108.015 126.045 108.485 ;
        RECT 126.525 108.015 127.735 108.765 ;
        RECT 14.660 107.845 127.820 108.015 ;
        RECT 14.745 107.095 15.955 107.845 ;
        RECT 16.435 107.375 16.605 107.845 ;
        RECT 16.775 107.195 17.105 107.675 ;
        RECT 17.275 107.375 17.445 107.845 ;
        RECT 17.615 107.195 17.945 107.675 ;
        RECT 14.745 106.555 15.265 107.095 ;
        RECT 16.180 107.025 17.945 107.195 ;
        RECT 18.115 107.035 18.285 107.845 ;
        RECT 18.485 107.465 19.555 107.635 ;
        RECT 18.485 107.110 18.805 107.465 ;
        RECT 15.435 106.385 15.955 106.925 ;
        RECT 14.745 105.295 15.955 106.385 ;
        RECT 16.180 106.475 16.590 107.025 ;
        RECT 18.480 106.855 18.805 107.110 ;
        RECT 16.775 106.645 18.805 106.855 ;
        RECT 18.460 106.635 18.805 106.645 ;
        RECT 18.975 106.895 19.215 107.295 ;
        RECT 19.385 107.235 19.555 107.465 ;
        RECT 19.725 107.405 19.915 107.845 ;
        RECT 20.085 107.395 21.035 107.675 ;
        RECT 21.255 107.485 21.605 107.655 ;
        RECT 19.385 107.065 19.915 107.235 ;
        RECT 16.180 106.305 17.905 106.475 ;
        RECT 16.435 105.295 16.605 106.135 ;
        RECT 16.815 105.465 17.065 106.305 ;
        RECT 17.275 105.295 17.445 106.135 ;
        RECT 17.615 105.465 17.905 106.305 ;
        RECT 18.115 105.295 18.285 106.355 ;
        RECT 18.460 106.015 18.630 106.635 ;
        RECT 18.975 106.525 19.515 106.895 ;
        RECT 19.695 106.785 19.915 107.065 ;
        RECT 20.085 106.615 20.255 107.395 ;
        RECT 19.850 106.445 20.255 106.615 ;
        RECT 20.425 106.605 20.775 107.225 ;
        RECT 19.850 106.355 20.020 106.445 ;
        RECT 20.945 106.435 21.155 107.225 ;
        RECT 18.800 106.185 20.020 106.355 ;
        RECT 20.480 106.275 21.155 106.435 ;
        RECT 18.460 105.845 19.260 106.015 ;
        RECT 18.580 105.295 18.910 105.675 ;
        RECT 19.090 105.555 19.260 105.845 ;
        RECT 19.850 105.805 20.020 106.185 ;
        RECT 20.190 106.265 21.155 106.275 ;
        RECT 21.345 107.095 21.605 107.485 ;
        RECT 21.815 107.385 22.145 107.845 ;
        RECT 23.020 107.455 23.875 107.625 ;
        RECT 24.080 107.455 24.575 107.625 ;
        RECT 24.745 107.485 25.075 107.845 ;
        RECT 21.345 106.405 21.515 107.095 ;
        RECT 21.685 106.745 21.855 106.925 ;
        RECT 22.025 106.915 22.815 107.165 ;
        RECT 23.020 106.745 23.190 107.455 ;
        RECT 23.360 106.945 23.715 107.165 ;
        RECT 21.685 106.575 23.375 106.745 ;
        RECT 20.190 105.975 20.650 106.265 ;
        RECT 21.345 106.235 22.845 106.405 ;
        RECT 21.345 106.095 21.515 106.235 ;
        RECT 20.955 105.925 21.515 106.095 ;
        RECT 19.430 105.295 19.680 105.755 ;
        RECT 19.850 105.465 20.720 105.805 ;
        RECT 20.955 105.465 21.125 105.925 ;
        RECT 21.960 105.895 23.035 106.065 ;
        RECT 21.295 105.295 21.665 105.755 ;
        RECT 21.960 105.555 22.130 105.895 ;
        RECT 22.300 105.295 22.630 105.725 ;
        RECT 22.865 105.555 23.035 105.895 ;
        RECT 23.205 105.795 23.375 106.575 ;
        RECT 23.545 106.355 23.715 106.945 ;
        RECT 23.885 106.545 24.235 107.165 ;
        RECT 23.545 105.965 24.010 106.355 ;
        RECT 24.405 106.095 24.575 107.455 ;
        RECT 24.745 106.265 25.205 107.315 ;
        RECT 24.180 105.925 24.575 106.095 ;
        RECT 24.180 105.795 24.350 105.925 ;
        RECT 23.205 105.465 23.885 105.795 ;
        RECT 24.100 105.465 24.350 105.795 ;
        RECT 24.520 105.295 24.770 105.755 ;
        RECT 24.940 105.480 25.265 106.265 ;
        RECT 25.435 105.465 25.605 107.585 ;
        RECT 25.775 107.465 26.105 107.845 ;
        RECT 26.275 107.295 26.530 107.585 ;
        RECT 27.015 107.375 27.185 107.845 ;
        RECT 25.780 107.125 26.530 107.295 ;
        RECT 27.355 107.195 27.685 107.675 ;
        RECT 27.855 107.375 28.025 107.845 ;
        RECT 28.195 107.195 28.525 107.675 ;
        RECT 25.780 106.135 26.010 107.125 ;
        RECT 26.760 107.025 28.525 107.195 ;
        RECT 28.695 107.035 28.865 107.845 ;
        RECT 29.065 107.465 30.135 107.635 ;
        RECT 29.065 107.110 29.385 107.465 ;
        RECT 26.180 106.305 26.530 106.955 ;
        RECT 26.760 106.475 27.170 107.025 ;
        RECT 29.060 106.855 29.385 107.110 ;
        RECT 27.355 106.645 29.385 106.855 ;
        RECT 29.040 106.635 29.385 106.645 ;
        RECT 29.555 106.895 29.795 107.295 ;
        RECT 29.965 107.235 30.135 107.465 ;
        RECT 30.305 107.405 30.495 107.845 ;
        RECT 30.665 107.395 31.615 107.675 ;
        RECT 31.835 107.485 32.185 107.655 ;
        RECT 29.965 107.065 30.495 107.235 ;
        RECT 26.760 106.305 28.485 106.475 ;
        RECT 25.780 105.965 26.530 106.135 ;
        RECT 25.775 105.295 26.105 105.795 ;
        RECT 26.275 105.465 26.530 105.965 ;
        RECT 27.015 105.295 27.185 106.135 ;
        RECT 27.395 105.465 27.645 106.305 ;
        RECT 27.855 105.295 28.025 106.135 ;
        RECT 28.195 105.465 28.485 106.305 ;
        RECT 28.695 105.295 28.865 106.355 ;
        RECT 29.040 106.015 29.210 106.635 ;
        RECT 29.555 106.525 30.095 106.895 ;
        RECT 30.275 106.785 30.495 107.065 ;
        RECT 30.665 106.615 30.835 107.395 ;
        RECT 30.430 106.445 30.835 106.615 ;
        RECT 31.005 106.605 31.355 107.225 ;
        RECT 30.430 106.355 30.600 106.445 ;
        RECT 31.525 106.435 31.735 107.225 ;
        RECT 29.380 106.185 30.600 106.355 ;
        RECT 31.060 106.275 31.735 106.435 ;
        RECT 29.040 105.845 29.840 106.015 ;
        RECT 29.160 105.295 29.490 105.675 ;
        RECT 29.670 105.555 29.840 105.845 ;
        RECT 30.430 105.805 30.600 106.185 ;
        RECT 30.770 106.265 31.735 106.275 ;
        RECT 31.925 107.095 32.185 107.485 ;
        RECT 32.395 107.385 32.725 107.845 ;
        RECT 33.600 107.455 34.455 107.625 ;
        RECT 34.660 107.455 35.155 107.625 ;
        RECT 35.325 107.485 35.655 107.845 ;
        RECT 31.925 106.405 32.095 107.095 ;
        RECT 32.265 106.745 32.435 106.925 ;
        RECT 32.605 106.915 33.395 107.165 ;
        RECT 33.600 106.745 33.770 107.455 ;
        RECT 33.940 106.945 34.295 107.165 ;
        RECT 32.265 106.575 33.955 106.745 ;
        RECT 30.770 105.975 31.230 106.265 ;
        RECT 31.925 106.235 33.425 106.405 ;
        RECT 31.925 106.095 32.095 106.235 ;
        RECT 31.535 105.925 32.095 106.095 ;
        RECT 30.010 105.295 30.260 105.755 ;
        RECT 30.430 105.465 31.300 105.805 ;
        RECT 31.535 105.465 31.705 105.925 ;
        RECT 32.540 105.895 33.615 106.065 ;
        RECT 31.875 105.295 32.245 105.755 ;
        RECT 32.540 105.555 32.710 105.895 ;
        RECT 32.880 105.295 33.210 105.725 ;
        RECT 33.445 105.555 33.615 105.895 ;
        RECT 33.785 105.795 33.955 106.575 ;
        RECT 34.125 106.355 34.295 106.945 ;
        RECT 34.465 106.545 34.815 107.165 ;
        RECT 34.125 105.965 34.590 106.355 ;
        RECT 34.985 106.095 35.155 107.455 ;
        RECT 35.325 106.265 35.785 107.315 ;
        RECT 34.760 105.925 35.155 106.095 ;
        RECT 34.760 105.795 34.930 105.925 ;
        RECT 33.785 105.465 34.465 105.795 ;
        RECT 34.680 105.465 34.930 105.795 ;
        RECT 35.100 105.295 35.350 105.755 ;
        RECT 35.520 105.480 35.845 106.265 ;
        RECT 36.015 105.465 36.185 107.585 ;
        RECT 36.355 107.465 36.685 107.845 ;
        RECT 36.855 107.295 37.110 107.585 ;
        RECT 36.360 107.125 37.110 107.295 ;
        RECT 36.360 106.135 36.590 107.125 ;
        RECT 37.285 107.120 37.575 107.845 ;
        RECT 37.745 107.170 38.005 107.675 ;
        RECT 38.185 107.465 38.515 107.845 ;
        RECT 38.695 107.295 38.865 107.675 ;
        RECT 36.760 106.305 37.110 106.955 ;
        RECT 36.360 105.965 37.110 106.135 ;
        RECT 36.355 105.295 36.685 105.795 ;
        RECT 36.855 105.465 37.110 105.965 ;
        RECT 37.285 105.295 37.575 106.460 ;
        RECT 37.745 106.370 37.915 107.170 ;
        RECT 38.200 107.125 38.865 107.295 ;
        RECT 38.200 106.870 38.370 107.125 ;
        RECT 39.645 107.025 39.855 107.845 ;
        RECT 40.025 107.045 40.355 107.675 ;
        RECT 38.085 106.540 38.370 106.870 ;
        RECT 38.605 106.575 38.935 106.945 ;
        RECT 38.200 106.395 38.370 106.540 ;
        RECT 40.025 106.445 40.275 107.045 ;
        RECT 40.525 107.025 40.755 107.845 ;
        RECT 40.965 107.095 42.175 107.845 ;
        RECT 40.445 106.605 40.775 106.855 ;
        RECT 37.745 105.465 38.015 106.370 ;
        RECT 38.200 106.225 38.865 106.395 ;
        RECT 38.185 105.295 38.515 106.055 ;
        RECT 38.695 105.465 38.865 106.225 ;
        RECT 39.645 105.295 39.855 106.435 ;
        RECT 40.025 105.465 40.355 106.445 ;
        RECT 40.525 105.295 40.755 106.435 ;
        RECT 40.965 106.385 41.485 106.925 ;
        RECT 41.655 106.555 42.175 107.095 ;
        RECT 42.345 107.170 42.605 107.675 ;
        RECT 42.785 107.465 43.115 107.845 ;
        RECT 43.295 107.295 43.465 107.675 ;
        RECT 40.965 105.295 42.175 106.385 ;
        RECT 42.345 106.370 42.515 107.170 ;
        RECT 42.800 107.125 43.465 107.295 ;
        RECT 42.800 106.870 42.970 107.125 ;
        RECT 44.245 107.025 44.455 107.845 ;
        RECT 44.625 107.045 44.955 107.675 ;
        RECT 42.685 106.540 42.970 106.870 ;
        RECT 43.205 106.575 43.535 106.945 ;
        RECT 42.800 106.395 42.970 106.540 ;
        RECT 44.625 106.445 44.875 107.045 ;
        RECT 45.125 107.025 45.355 107.845 ;
        RECT 45.655 107.295 45.825 107.675 ;
        RECT 46.005 107.465 46.335 107.845 ;
        RECT 45.655 107.125 46.320 107.295 ;
        RECT 46.515 107.170 46.775 107.675 ;
        RECT 47.255 107.375 47.425 107.845 ;
        RECT 47.595 107.195 47.925 107.675 ;
        RECT 48.095 107.375 48.265 107.845 ;
        RECT 48.435 107.195 48.765 107.675 ;
        RECT 45.045 106.605 45.375 106.855 ;
        RECT 45.585 106.575 45.915 106.945 ;
        RECT 46.150 106.870 46.320 107.125 ;
        RECT 46.150 106.540 46.435 106.870 ;
        RECT 42.345 105.465 42.615 106.370 ;
        RECT 42.800 106.225 43.465 106.395 ;
        RECT 42.785 105.295 43.115 106.055 ;
        RECT 43.295 105.465 43.465 106.225 ;
        RECT 44.245 105.295 44.455 106.435 ;
        RECT 44.625 105.465 44.955 106.445 ;
        RECT 45.125 105.295 45.355 106.435 ;
        RECT 46.150 106.395 46.320 106.540 ;
        RECT 45.655 106.225 46.320 106.395 ;
        RECT 46.605 106.370 46.775 107.170 ;
        RECT 45.655 105.465 45.825 106.225 ;
        RECT 46.005 105.295 46.335 106.055 ;
        RECT 46.505 105.465 46.775 106.370 ;
        RECT 47.000 107.025 48.765 107.195 ;
        RECT 48.935 107.035 49.105 107.845 ;
        RECT 49.305 107.465 50.375 107.635 ;
        RECT 49.305 107.110 49.625 107.465 ;
        RECT 47.000 106.475 47.410 107.025 ;
        RECT 49.300 106.855 49.625 107.110 ;
        RECT 47.595 106.645 49.625 106.855 ;
        RECT 49.280 106.635 49.625 106.645 ;
        RECT 49.795 106.895 50.035 107.295 ;
        RECT 50.205 107.235 50.375 107.465 ;
        RECT 50.545 107.405 50.735 107.845 ;
        RECT 50.905 107.395 51.855 107.675 ;
        RECT 52.075 107.485 52.425 107.655 ;
        RECT 50.205 107.065 50.735 107.235 ;
        RECT 47.000 106.305 48.725 106.475 ;
        RECT 47.255 105.295 47.425 106.135 ;
        RECT 47.635 105.465 47.885 106.305 ;
        RECT 48.095 105.295 48.265 106.135 ;
        RECT 48.435 105.465 48.725 106.305 ;
        RECT 48.935 105.295 49.105 106.355 ;
        RECT 49.280 106.015 49.450 106.635 ;
        RECT 49.795 106.525 50.335 106.895 ;
        RECT 50.515 106.785 50.735 107.065 ;
        RECT 50.905 106.615 51.075 107.395 ;
        RECT 50.670 106.445 51.075 106.615 ;
        RECT 51.245 106.605 51.595 107.225 ;
        RECT 50.670 106.355 50.840 106.445 ;
        RECT 51.765 106.435 51.975 107.225 ;
        RECT 49.620 106.185 50.840 106.355 ;
        RECT 51.300 106.275 51.975 106.435 ;
        RECT 49.280 105.845 50.080 106.015 ;
        RECT 49.400 105.295 49.730 105.675 ;
        RECT 49.910 105.555 50.080 105.845 ;
        RECT 50.670 105.805 50.840 106.185 ;
        RECT 51.010 106.265 51.975 106.275 ;
        RECT 52.165 107.095 52.425 107.485 ;
        RECT 52.635 107.385 52.965 107.845 ;
        RECT 53.840 107.455 54.695 107.625 ;
        RECT 54.900 107.455 55.395 107.625 ;
        RECT 55.565 107.485 55.895 107.845 ;
        RECT 52.165 106.405 52.335 107.095 ;
        RECT 52.505 106.745 52.675 106.925 ;
        RECT 52.845 106.915 53.635 107.165 ;
        RECT 53.840 106.745 54.010 107.455 ;
        RECT 54.180 106.945 54.535 107.165 ;
        RECT 52.505 106.575 54.195 106.745 ;
        RECT 51.010 105.975 51.470 106.265 ;
        RECT 52.165 106.235 53.665 106.405 ;
        RECT 52.165 106.095 52.335 106.235 ;
        RECT 51.775 105.925 52.335 106.095 ;
        RECT 50.250 105.295 50.500 105.755 ;
        RECT 50.670 105.465 51.540 105.805 ;
        RECT 51.775 105.465 51.945 105.925 ;
        RECT 52.780 105.895 53.855 106.065 ;
        RECT 52.115 105.295 52.485 105.755 ;
        RECT 52.780 105.555 52.950 105.895 ;
        RECT 53.120 105.295 53.450 105.725 ;
        RECT 53.685 105.555 53.855 105.895 ;
        RECT 54.025 105.795 54.195 106.575 ;
        RECT 54.365 106.355 54.535 106.945 ;
        RECT 54.705 106.545 55.055 107.165 ;
        RECT 54.365 105.965 54.830 106.355 ;
        RECT 55.225 106.095 55.395 107.455 ;
        RECT 55.565 106.265 56.025 107.315 ;
        RECT 55.000 105.925 55.395 106.095 ;
        RECT 55.000 105.795 55.170 105.925 ;
        RECT 54.025 105.465 54.705 105.795 ;
        RECT 54.920 105.465 55.170 105.795 ;
        RECT 55.340 105.295 55.590 105.755 ;
        RECT 55.760 105.480 56.085 106.265 ;
        RECT 56.255 105.465 56.425 107.585 ;
        RECT 56.595 107.465 56.925 107.845 ;
        RECT 57.095 107.295 57.350 107.585 ;
        RECT 56.600 107.125 57.350 107.295 ;
        RECT 56.600 106.135 56.830 107.125 ;
        RECT 57.585 107.025 57.795 107.845 ;
        RECT 57.965 107.045 58.295 107.675 ;
        RECT 57.000 106.305 57.350 106.955 ;
        RECT 57.965 106.445 58.215 107.045 ;
        RECT 58.465 107.025 58.695 107.845 ;
        RECT 58.905 107.095 60.115 107.845 ;
        RECT 58.385 106.605 58.715 106.855 ;
        RECT 56.600 105.965 57.350 106.135 ;
        RECT 56.595 105.295 56.925 105.795 ;
        RECT 57.095 105.465 57.350 105.965 ;
        RECT 57.585 105.295 57.795 106.435 ;
        RECT 57.965 105.465 58.295 106.445 ;
        RECT 58.465 105.295 58.695 106.435 ;
        RECT 58.905 106.385 59.425 106.925 ;
        RECT 59.595 106.555 60.115 107.095 ;
        RECT 60.325 107.025 60.555 107.845 ;
        RECT 60.725 107.045 61.055 107.675 ;
        RECT 60.305 106.605 60.635 106.855 ;
        RECT 60.805 106.445 61.055 107.045 ;
        RECT 61.225 107.025 61.435 107.845 ;
        RECT 61.755 107.295 61.925 107.675 ;
        RECT 62.105 107.465 62.435 107.845 ;
        RECT 61.755 107.125 62.420 107.295 ;
        RECT 62.615 107.170 62.875 107.675 ;
        RECT 61.685 106.575 62.015 106.945 ;
        RECT 62.250 106.870 62.420 107.125 ;
        RECT 58.905 105.295 60.115 106.385 ;
        RECT 60.325 105.295 60.555 106.435 ;
        RECT 60.725 105.465 61.055 106.445 ;
        RECT 62.250 106.540 62.535 106.870 ;
        RECT 61.225 105.295 61.435 106.435 ;
        RECT 62.250 106.395 62.420 106.540 ;
        RECT 61.755 106.225 62.420 106.395 ;
        RECT 62.705 106.370 62.875 107.170 ;
        RECT 63.045 107.120 63.335 107.845 ;
        RECT 63.815 107.375 63.985 107.845 ;
        RECT 64.155 107.195 64.485 107.675 ;
        RECT 64.655 107.375 64.825 107.845 ;
        RECT 64.995 107.195 65.325 107.675 ;
        RECT 63.560 107.025 65.325 107.195 ;
        RECT 65.495 107.035 65.665 107.845 ;
        RECT 65.865 107.465 66.935 107.635 ;
        RECT 65.865 107.110 66.185 107.465 ;
        RECT 63.560 106.475 63.970 107.025 ;
        RECT 65.860 106.855 66.185 107.110 ;
        RECT 64.155 106.645 66.185 106.855 ;
        RECT 65.840 106.635 66.185 106.645 ;
        RECT 66.355 106.895 66.595 107.295 ;
        RECT 66.765 107.235 66.935 107.465 ;
        RECT 67.105 107.405 67.295 107.845 ;
        RECT 67.465 107.395 68.415 107.675 ;
        RECT 68.635 107.485 68.985 107.655 ;
        RECT 66.765 107.065 67.295 107.235 ;
        RECT 61.755 105.465 61.925 106.225 ;
        RECT 62.105 105.295 62.435 106.055 ;
        RECT 62.605 105.465 62.875 106.370 ;
        RECT 63.045 105.295 63.335 106.460 ;
        RECT 63.560 106.305 65.285 106.475 ;
        RECT 63.815 105.295 63.985 106.135 ;
        RECT 64.195 105.465 64.445 106.305 ;
        RECT 64.655 105.295 64.825 106.135 ;
        RECT 64.995 105.465 65.285 106.305 ;
        RECT 65.495 105.295 65.665 106.355 ;
        RECT 65.840 106.015 66.010 106.635 ;
        RECT 66.355 106.525 66.895 106.895 ;
        RECT 67.075 106.785 67.295 107.065 ;
        RECT 67.465 106.615 67.635 107.395 ;
        RECT 67.230 106.445 67.635 106.615 ;
        RECT 67.805 106.605 68.155 107.225 ;
        RECT 67.230 106.355 67.400 106.445 ;
        RECT 68.325 106.435 68.535 107.225 ;
        RECT 66.180 106.185 67.400 106.355 ;
        RECT 67.860 106.275 68.535 106.435 ;
        RECT 65.840 105.845 66.640 106.015 ;
        RECT 65.960 105.295 66.290 105.675 ;
        RECT 66.470 105.555 66.640 105.845 ;
        RECT 67.230 105.805 67.400 106.185 ;
        RECT 67.570 106.265 68.535 106.275 ;
        RECT 68.725 107.095 68.985 107.485 ;
        RECT 69.195 107.385 69.525 107.845 ;
        RECT 70.400 107.455 71.255 107.625 ;
        RECT 71.460 107.455 71.955 107.625 ;
        RECT 72.125 107.485 72.455 107.845 ;
        RECT 68.725 106.405 68.895 107.095 ;
        RECT 69.065 106.745 69.235 106.925 ;
        RECT 69.405 106.915 70.195 107.165 ;
        RECT 70.400 106.745 70.570 107.455 ;
        RECT 70.740 106.945 71.095 107.165 ;
        RECT 69.065 106.575 70.755 106.745 ;
        RECT 67.570 105.975 68.030 106.265 ;
        RECT 68.725 106.235 70.225 106.405 ;
        RECT 68.725 106.095 68.895 106.235 ;
        RECT 68.335 105.925 68.895 106.095 ;
        RECT 66.810 105.295 67.060 105.755 ;
        RECT 67.230 105.465 68.100 105.805 ;
        RECT 68.335 105.465 68.505 105.925 ;
        RECT 69.340 105.895 70.415 106.065 ;
        RECT 68.675 105.295 69.045 105.755 ;
        RECT 69.340 105.555 69.510 105.895 ;
        RECT 69.680 105.295 70.010 105.725 ;
        RECT 70.245 105.555 70.415 105.895 ;
        RECT 70.585 105.795 70.755 106.575 ;
        RECT 70.925 106.355 71.095 106.945 ;
        RECT 71.265 106.545 71.615 107.165 ;
        RECT 70.925 105.965 71.390 106.355 ;
        RECT 71.785 106.095 71.955 107.455 ;
        RECT 72.125 106.265 72.585 107.315 ;
        RECT 71.560 105.925 71.955 106.095 ;
        RECT 71.560 105.795 71.730 105.925 ;
        RECT 70.585 105.465 71.265 105.795 ;
        RECT 71.480 105.465 71.730 105.795 ;
        RECT 71.900 105.295 72.150 105.755 ;
        RECT 72.320 105.480 72.645 106.265 ;
        RECT 72.815 105.465 72.985 107.585 ;
        RECT 73.155 107.465 73.485 107.845 ;
        RECT 73.655 107.295 73.910 107.585 ;
        RECT 73.160 107.125 73.910 107.295 ;
        RECT 75.095 107.295 75.265 107.675 ;
        RECT 75.445 107.465 75.775 107.845 ;
        RECT 75.095 107.125 75.760 107.295 ;
        RECT 75.955 107.170 76.215 107.675 ;
        RECT 76.695 107.375 76.865 107.845 ;
        RECT 77.035 107.195 77.365 107.675 ;
        RECT 77.535 107.375 77.705 107.845 ;
        RECT 77.875 107.195 78.205 107.675 ;
        RECT 73.160 106.135 73.390 107.125 ;
        RECT 73.560 106.305 73.910 106.955 ;
        RECT 75.025 106.575 75.355 106.945 ;
        RECT 75.590 106.870 75.760 107.125 ;
        RECT 75.590 106.540 75.875 106.870 ;
        RECT 75.590 106.395 75.760 106.540 ;
        RECT 75.095 106.225 75.760 106.395 ;
        RECT 76.045 106.370 76.215 107.170 ;
        RECT 73.160 105.965 73.910 106.135 ;
        RECT 73.155 105.295 73.485 105.795 ;
        RECT 73.655 105.465 73.910 105.965 ;
        RECT 75.095 105.465 75.265 106.225 ;
        RECT 75.445 105.295 75.775 106.055 ;
        RECT 75.945 105.465 76.215 106.370 ;
        RECT 76.440 107.025 78.205 107.195 ;
        RECT 78.375 107.035 78.545 107.845 ;
        RECT 78.745 107.465 79.815 107.635 ;
        RECT 78.745 107.110 79.065 107.465 ;
        RECT 76.440 106.475 76.850 107.025 ;
        RECT 78.740 106.855 79.065 107.110 ;
        RECT 77.035 106.645 79.065 106.855 ;
        RECT 78.720 106.635 79.065 106.645 ;
        RECT 79.235 106.895 79.475 107.295 ;
        RECT 79.645 107.235 79.815 107.465 ;
        RECT 79.985 107.405 80.175 107.845 ;
        RECT 80.345 107.395 81.295 107.675 ;
        RECT 81.515 107.485 81.865 107.655 ;
        RECT 79.645 107.065 80.175 107.235 ;
        RECT 76.440 106.305 78.165 106.475 ;
        RECT 76.695 105.295 76.865 106.135 ;
        RECT 77.075 105.465 77.325 106.305 ;
        RECT 77.535 105.295 77.705 106.135 ;
        RECT 77.875 105.465 78.165 106.305 ;
        RECT 78.375 105.295 78.545 106.355 ;
        RECT 78.720 106.015 78.890 106.635 ;
        RECT 79.235 106.525 79.775 106.895 ;
        RECT 79.955 106.785 80.175 107.065 ;
        RECT 80.345 106.615 80.515 107.395 ;
        RECT 80.110 106.445 80.515 106.615 ;
        RECT 80.685 106.605 81.035 107.225 ;
        RECT 80.110 106.355 80.280 106.445 ;
        RECT 81.205 106.435 81.415 107.225 ;
        RECT 79.060 106.185 80.280 106.355 ;
        RECT 80.740 106.275 81.415 106.435 ;
        RECT 78.720 105.845 79.520 106.015 ;
        RECT 78.840 105.295 79.170 105.675 ;
        RECT 79.350 105.555 79.520 105.845 ;
        RECT 80.110 105.805 80.280 106.185 ;
        RECT 80.450 106.265 81.415 106.275 ;
        RECT 81.605 107.095 81.865 107.485 ;
        RECT 82.075 107.385 82.405 107.845 ;
        RECT 83.280 107.455 84.135 107.625 ;
        RECT 84.340 107.455 84.835 107.625 ;
        RECT 85.005 107.485 85.335 107.845 ;
        RECT 81.605 106.405 81.775 107.095 ;
        RECT 81.945 106.745 82.115 106.925 ;
        RECT 82.285 106.915 83.075 107.165 ;
        RECT 83.280 106.745 83.450 107.455 ;
        RECT 83.620 106.945 83.975 107.165 ;
        RECT 81.945 106.575 83.635 106.745 ;
        RECT 80.450 105.975 80.910 106.265 ;
        RECT 81.605 106.235 83.105 106.405 ;
        RECT 81.605 106.095 81.775 106.235 ;
        RECT 81.215 105.925 81.775 106.095 ;
        RECT 79.690 105.295 79.940 105.755 ;
        RECT 80.110 105.465 80.980 105.805 ;
        RECT 81.215 105.465 81.385 105.925 ;
        RECT 82.220 105.895 83.295 106.065 ;
        RECT 81.555 105.295 81.925 105.755 ;
        RECT 82.220 105.555 82.390 105.895 ;
        RECT 82.560 105.295 82.890 105.725 ;
        RECT 83.125 105.555 83.295 105.895 ;
        RECT 83.465 105.795 83.635 106.575 ;
        RECT 83.805 106.355 83.975 106.945 ;
        RECT 84.145 106.545 84.495 107.165 ;
        RECT 83.805 105.965 84.270 106.355 ;
        RECT 84.665 106.095 84.835 107.455 ;
        RECT 85.005 106.265 85.465 107.315 ;
        RECT 84.440 105.925 84.835 106.095 ;
        RECT 84.440 105.795 84.610 105.925 ;
        RECT 83.465 105.465 84.145 105.795 ;
        RECT 84.360 105.465 84.610 105.795 ;
        RECT 84.780 105.295 85.030 105.755 ;
        RECT 85.200 105.480 85.525 106.265 ;
        RECT 85.695 105.465 85.865 107.585 ;
        RECT 86.035 107.465 86.365 107.845 ;
        RECT 86.535 107.295 86.790 107.585 ;
        RECT 86.040 107.125 86.790 107.295 ;
        RECT 87.515 107.295 87.685 107.675 ;
        RECT 87.865 107.465 88.195 107.845 ;
        RECT 87.515 107.125 88.180 107.295 ;
        RECT 88.375 107.170 88.635 107.675 ;
        RECT 86.040 106.135 86.270 107.125 ;
        RECT 86.440 106.305 86.790 106.955 ;
        RECT 87.445 106.575 87.775 106.945 ;
        RECT 88.010 106.870 88.180 107.125 ;
        RECT 88.010 106.540 88.295 106.870 ;
        RECT 88.010 106.395 88.180 106.540 ;
        RECT 87.515 106.225 88.180 106.395 ;
        RECT 88.465 106.370 88.635 107.170 ;
        RECT 88.805 107.120 89.095 107.845 ;
        RECT 89.575 107.375 89.745 107.845 ;
        RECT 89.915 107.195 90.245 107.675 ;
        RECT 90.415 107.375 90.585 107.845 ;
        RECT 90.755 107.195 91.085 107.675 ;
        RECT 89.320 107.025 91.085 107.195 ;
        RECT 91.255 107.035 91.425 107.845 ;
        RECT 91.625 107.465 92.695 107.635 ;
        RECT 91.625 107.110 91.945 107.465 ;
        RECT 89.320 106.475 89.730 107.025 ;
        RECT 91.620 106.855 91.945 107.110 ;
        RECT 89.915 106.645 91.945 106.855 ;
        RECT 91.600 106.635 91.945 106.645 ;
        RECT 92.115 106.895 92.355 107.295 ;
        RECT 92.525 107.235 92.695 107.465 ;
        RECT 92.865 107.405 93.055 107.845 ;
        RECT 93.225 107.395 94.175 107.675 ;
        RECT 94.395 107.485 94.745 107.655 ;
        RECT 92.525 107.065 93.055 107.235 ;
        RECT 86.040 105.965 86.790 106.135 ;
        RECT 86.035 105.295 86.365 105.795 ;
        RECT 86.535 105.465 86.790 105.965 ;
        RECT 87.515 105.465 87.685 106.225 ;
        RECT 87.865 105.295 88.195 106.055 ;
        RECT 88.365 105.465 88.635 106.370 ;
        RECT 88.805 105.295 89.095 106.460 ;
        RECT 89.320 106.305 91.045 106.475 ;
        RECT 89.575 105.295 89.745 106.135 ;
        RECT 89.955 105.465 90.205 106.305 ;
        RECT 90.415 105.295 90.585 106.135 ;
        RECT 90.755 105.465 91.045 106.305 ;
        RECT 91.255 105.295 91.425 106.355 ;
        RECT 91.600 106.015 91.770 106.635 ;
        RECT 92.115 106.525 92.655 106.895 ;
        RECT 92.835 106.785 93.055 107.065 ;
        RECT 93.225 106.615 93.395 107.395 ;
        RECT 92.990 106.445 93.395 106.615 ;
        RECT 93.565 106.605 93.915 107.225 ;
        RECT 92.990 106.355 93.160 106.445 ;
        RECT 94.085 106.435 94.295 107.225 ;
        RECT 91.940 106.185 93.160 106.355 ;
        RECT 93.620 106.275 94.295 106.435 ;
        RECT 91.600 105.845 92.400 106.015 ;
        RECT 91.720 105.295 92.050 105.675 ;
        RECT 92.230 105.555 92.400 105.845 ;
        RECT 92.990 105.805 93.160 106.185 ;
        RECT 93.330 106.265 94.295 106.275 ;
        RECT 94.485 107.095 94.745 107.485 ;
        RECT 94.955 107.385 95.285 107.845 ;
        RECT 96.160 107.455 97.015 107.625 ;
        RECT 97.220 107.455 97.715 107.625 ;
        RECT 97.885 107.485 98.215 107.845 ;
        RECT 94.485 106.405 94.655 107.095 ;
        RECT 94.825 106.745 94.995 106.925 ;
        RECT 95.165 106.915 95.955 107.165 ;
        RECT 96.160 106.745 96.330 107.455 ;
        RECT 96.500 106.945 96.855 107.165 ;
        RECT 94.825 106.575 96.515 106.745 ;
        RECT 93.330 105.975 93.790 106.265 ;
        RECT 94.485 106.235 95.985 106.405 ;
        RECT 94.485 106.095 94.655 106.235 ;
        RECT 94.095 105.925 94.655 106.095 ;
        RECT 92.570 105.295 92.820 105.755 ;
        RECT 92.990 105.465 93.860 105.805 ;
        RECT 94.095 105.465 94.265 105.925 ;
        RECT 95.100 105.895 96.175 106.065 ;
        RECT 94.435 105.295 94.805 105.755 ;
        RECT 95.100 105.555 95.270 105.895 ;
        RECT 95.440 105.295 95.770 105.725 ;
        RECT 96.005 105.555 96.175 105.895 ;
        RECT 96.345 105.795 96.515 106.575 ;
        RECT 96.685 106.355 96.855 106.945 ;
        RECT 97.025 106.545 97.375 107.165 ;
        RECT 96.685 105.965 97.150 106.355 ;
        RECT 97.545 106.095 97.715 107.455 ;
        RECT 97.885 106.265 98.345 107.315 ;
        RECT 97.320 105.925 97.715 106.095 ;
        RECT 97.320 105.795 97.490 105.925 ;
        RECT 96.345 105.465 97.025 105.795 ;
        RECT 97.240 105.465 97.490 105.795 ;
        RECT 97.660 105.295 97.910 105.755 ;
        RECT 98.080 105.480 98.405 106.265 ;
        RECT 98.575 105.465 98.745 107.585 ;
        RECT 98.915 107.465 99.245 107.845 ;
        RECT 99.415 107.295 99.670 107.585 ;
        RECT 98.920 107.125 99.670 107.295 ;
        RECT 98.920 106.135 99.150 107.125 ;
        RECT 99.905 107.025 100.115 107.845 ;
        RECT 100.285 107.045 100.615 107.675 ;
        RECT 99.320 106.305 99.670 106.955 ;
        RECT 100.285 106.445 100.535 107.045 ;
        RECT 100.785 107.025 101.015 107.845 ;
        RECT 101.225 107.095 102.435 107.845 ;
        RECT 100.705 106.605 101.035 106.855 ;
        RECT 98.920 105.965 99.670 106.135 ;
        RECT 98.915 105.295 99.245 105.795 ;
        RECT 99.415 105.465 99.670 105.965 ;
        RECT 99.905 105.295 100.115 106.435 ;
        RECT 100.285 105.465 100.615 106.445 ;
        RECT 100.785 105.295 101.015 106.435 ;
        RECT 101.225 106.385 101.745 106.925 ;
        RECT 101.915 106.555 102.435 107.095 ;
        RECT 102.645 107.025 102.875 107.845 ;
        RECT 103.045 107.045 103.375 107.675 ;
        RECT 102.625 106.605 102.955 106.855 ;
        RECT 103.125 106.445 103.375 107.045 ;
        RECT 103.545 107.025 103.755 107.845 ;
        RECT 104.295 107.375 104.465 107.845 ;
        RECT 104.635 107.195 104.965 107.675 ;
        RECT 105.135 107.375 105.305 107.845 ;
        RECT 105.475 107.195 105.805 107.675 ;
        RECT 104.040 107.025 105.805 107.195 ;
        RECT 105.975 107.035 106.145 107.845 ;
        RECT 106.345 107.465 107.415 107.635 ;
        RECT 106.345 107.110 106.665 107.465 ;
        RECT 101.225 105.295 102.435 106.385 ;
        RECT 102.645 105.295 102.875 106.435 ;
        RECT 103.045 105.465 103.375 106.445 ;
        RECT 104.040 106.475 104.450 107.025 ;
        RECT 106.340 106.855 106.665 107.110 ;
        RECT 104.635 106.645 106.665 106.855 ;
        RECT 106.320 106.635 106.665 106.645 ;
        RECT 106.835 106.895 107.075 107.295 ;
        RECT 107.245 107.235 107.415 107.465 ;
        RECT 107.585 107.405 107.775 107.845 ;
        RECT 107.945 107.395 108.895 107.675 ;
        RECT 109.115 107.485 109.465 107.655 ;
        RECT 107.245 107.065 107.775 107.235 ;
        RECT 103.545 105.295 103.755 106.435 ;
        RECT 104.040 106.305 105.765 106.475 ;
        RECT 104.295 105.295 104.465 106.135 ;
        RECT 104.675 105.465 104.925 106.305 ;
        RECT 105.135 105.295 105.305 106.135 ;
        RECT 105.475 105.465 105.765 106.305 ;
        RECT 105.975 105.295 106.145 106.355 ;
        RECT 106.320 106.015 106.490 106.635 ;
        RECT 106.835 106.525 107.375 106.895 ;
        RECT 107.555 106.785 107.775 107.065 ;
        RECT 107.945 106.615 108.115 107.395 ;
        RECT 107.710 106.445 108.115 106.615 ;
        RECT 108.285 106.605 108.635 107.225 ;
        RECT 107.710 106.355 107.880 106.445 ;
        RECT 108.805 106.435 109.015 107.225 ;
        RECT 106.660 106.185 107.880 106.355 ;
        RECT 108.340 106.275 109.015 106.435 ;
        RECT 106.320 105.845 107.120 106.015 ;
        RECT 106.440 105.295 106.770 105.675 ;
        RECT 106.950 105.555 107.120 105.845 ;
        RECT 107.710 105.805 107.880 106.185 ;
        RECT 108.050 106.265 109.015 106.275 ;
        RECT 109.205 107.095 109.465 107.485 ;
        RECT 109.675 107.385 110.005 107.845 ;
        RECT 110.880 107.455 111.735 107.625 ;
        RECT 111.940 107.455 112.435 107.625 ;
        RECT 112.605 107.485 112.935 107.845 ;
        RECT 109.205 106.405 109.375 107.095 ;
        RECT 109.545 106.745 109.715 106.925 ;
        RECT 109.885 106.915 110.675 107.165 ;
        RECT 110.880 106.745 111.050 107.455 ;
        RECT 111.220 106.945 111.575 107.165 ;
        RECT 109.545 106.575 111.235 106.745 ;
        RECT 108.050 105.975 108.510 106.265 ;
        RECT 109.205 106.235 110.705 106.405 ;
        RECT 109.205 106.095 109.375 106.235 ;
        RECT 108.815 105.925 109.375 106.095 ;
        RECT 107.290 105.295 107.540 105.755 ;
        RECT 107.710 105.465 108.580 105.805 ;
        RECT 108.815 105.465 108.985 105.925 ;
        RECT 109.820 105.895 110.895 106.065 ;
        RECT 109.155 105.295 109.525 105.755 ;
        RECT 109.820 105.555 109.990 105.895 ;
        RECT 110.160 105.295 110.490 105.725 ;
        RECT 110.725 105.555 110.895 105.895 ;
        RECT 111.065 105.795 111.235 106.575 ;
        RECT 111.405 106.355 111.575 106.945 ;
        RECT 111.745 106.545 112.095 107.165 ;
        RECT 111.405 105.965 111.870 106.355 ;
        RECT 112.265 106.095 112.435 107.455 ;
        RECT 112.605 106.265 113.065 107.315 ;
        RECT 112.040 105.925 112.435 106.095 ;
        RECT 112.040 105.795 112.210 105.925 ;
        RECT 111.065 105.465 111.745 105.795 ;
        RECT 111.960 105.465 112.210 105.795 ;
        RECT 112.380 105.295 112.630 105.755 ;
        RECT 112.800 105.480 113.125 106.265 ;
        RECT 113.295 105.465 113.465 107.585 ;
        RECT 113.635 107.465 113.965 107.845 ;
        RECT 114.135 107.295 114.390 107.585 ;
        RECT 113.640 107.125 114.390 107.295 ;
        RECT 113.640 106.135 113.870 107.125 ;
        RECT 114.565 107.120 114.855 107.845 ;
        RECT 115.950 107.295 116.205 107.585 ;
        RECT 116.375 107.465 116.705 107.845 ;
        RECT 115.950 107.125 116.700 107.295 ;
        RECT 114.040 106.305 114.390 106.955 ;
        RECT 113.640 105.965 114.390 106.135 ;
        RECT 113.635 105.295 113.965 105.795 ;
        RECT 114.135 105.465 114.390 105.965 ;
        RECT 114.565 105.295 114.855 106.460 ;
        RECT 115.950 106.305 116.300 106.955 ;
        RECT 116.470 106.135 116.700 107.125 ;
        RECT 115.950 105.965 116.700 106.135 ;
        RECT 115.950 105.465 116.205 105.965 ;
        RECT 116.375 105.295 116.705 105.795 ;
        RECT 116.875 105.465 117.045 107.585 ;
        RECT 117.405 107.485 117.735 107.845 ;
        RECT 117.905 107.455 118.400 107.625 ;
        RECT 118.605 107.455 119.460 107.625 ;
        RECT 117.275 106.265 117.735 107.315 ;
        RECT 117.215 105.480 117.540 106.265 ;
        RECT 117.905 106.095 118.075 107.455 ;
        RECT 118.245 106.545 118.595 107.165 ;
        RECT 118.765 106.945 119.120 107.165 ;
        RECT 118.765 106.355 118.935 106.945 ;
        RECT 119.290 106.745 119.460 107.455 ;
        RECT 120.335 107.385 120.665 107.845 ;
        RECT 120.875 107.485 121.225 107.655 ;
        RECT 119.665 106.915 120.455 107.165 ;
        RECT 120.875 107.095 121.135 107.485 ;
        RECT 121.445 107.395 122.395 107.675 ;
        RECT 122.565 107.405 122.755 107.845 ;
        RECT 122.925 107.465 123.995 107.635 ;
        RECT 120.625 106.745 120.795 106.925 ;
        RECT 117.905 105.925 118.300 106.095 ;
        RECT 118.470 105.965 118.935 106.355 ;
        RECT 119.105 106.575 120.795 106.745 ;
        RECT 118.130 105.795 118.300 105.925 ;
        RECT 119.105 105.795 119.275 106.575 ;
        RECT 120.965 106.405 121.135 107.095 ;
        RECT 119.635 106.235 121.135 106.405 ;
        RECT 121.325 106.435 121.535 107.225 ;
        RECT 121.705 106.605 122.055 107.225 ;
        RECT 122.225 106.615 122.395 107.395 ;
        RECT 122.925 107.235 123.095 107.465 ;
        RECT 122.565 107.065 123.095 107.235 ;
        RECT 122.565 106.785 122.785 107.065 ;
        RECT 123.265 106.895 123.505 107.295 ;
        RECT 122.225 106.445 122.630 106.615 ;
        RECT 122.965 106.525 123.505 106.895 ;
        RECT 123.675 107.110 123.995 107.465 ;
        RECT 123.675 106.855 124.000 107.110 ;
        RECT 124.195 107.035 124.365 107.845 ;
        RECT 124.535 107.195 124.865 107.675 ;
        RECT 125.035 107.375 125.205 107.845 ;
        RECT 125.375 107.195 125.705 107.675 ;
        RECT 125.875 107.375 126.045 107.845 ;
        RECT 124.535 107.025 126.300 107.195 ;
        RECT 126.525 107.095 127.735 107.845 ;
        RECT 123.675 106.645 125.705 106.855 ;
        RECT 123.675 106.635 124.020 106.645 ;
        RECT 121.325 106.275 122.000 106.435 ;
        RECT 122.460 106.355 122.630 106.445 ;
        RECT 121.325 106.265 122.290 106.275 ;
        RECT 120.965 106.095 121.135 106.235 ;
        RECT 117.710 105.295 117.960 105.755 ;
        RECT 118.130 105.465 118.380 105.795 ;
        RECT 118.595 105.465 119.275 105.795 ;
        RECT 119.445 105.895 120.520 106.065 ;
        RECT 120.965 105.925 121.525 106.095 ;
        RECT 121.830 105.975 122.290 106.265 ;
        RECT 122.460 106.185 123.680 106.355 ;
        RECT 119.445 105.555 119.615 105.895 ;
        RECT 119.850 105.295 120.180 105.725 ;
        RECT 120.350 105.555 120.520 105.895 ;
        RECT 120.815 105.295 121.185 105.755 ;
        RECT 121.355 105.465 121.525 105.925 ;
        RECT 122.460 105.805 122.630 106.185 ;
        RECT 123.850 106.015 124.020 106.635 ;
        RECT 125.890 106.475 126.300 107.025 ;
        RECT 121.760 105.465 122.630 105.805 ;
        RECT 123.220 105.845 124.020 106.015 ;
        RECT 122.800 105.295 123.050 105.755 ;
        RECT 123.220 105.555 123.390 105.845 ;
        RECT 123.570 105.295 123.900 105.675 ;
        RECT 124.195 105.295 124.365 106.355 ;
        RECT 124.575 106.305 126.300 106.475 ;
        RECT 126.525 106.385 127.045 106.925 ;
        RECT 127.215 106.555 127.735 107.095 ;
        RECT 124.575 105.465 124.865 106.305 ;
        RECT 125.035 105.295 125.205 106.135 ;
        RECT 125.415 105.465 125.665 106.305 ;
        RECT 125.875 105.295 126.045 106.135 ;
        RECT 126.525 105.295 127.735 106.385 ;
        RECT 14.660 105.125 127.820 105.295 ;
        RECT 14.745 104.035 15.955 105.125 ;
        RECT 14.745 103.325 15.265 103.865 ;
        RECT 15.435 103.495 15.955 104.035 ;
        RECT 16.125 104.035 18.715 105.125 ;
        RECT 18.890 104.690 24.235 105.125 ;
        RECT 16.125 103.515 17.335 104.035 ;
        RECT 17.505 103.345 18.715 103.865 ;
        RECT 20.480 103.440 20.830 104.690 ;
        RECT 24.405 103.960 24.695 105.125 ;
        RECT 24.865 104.035 27.455 105.125 ;
        RECT 14.745 102.575 15.955 103.325 ;
        RECT 16.125 102.575 18.715 103.345 ;
        RECT 22.310 103.120 22.650 103.950 ;
        RECT 24.865 103.515 26.075 104.035 ;
        RECT 27.665 103.985 27.895 105.125 ;
        RECT 28.065 103.975 28.395 104.955 ;
        RECT 28.565 103.985 28.775 105.125 ;
        RECT 29.010 104.455 29.265 104.955 ;
        RECT 29.435 104.625 29.765 105.125 ;
        RECT 29.010 104.285 29.760 104.455 ;
        RECT 26.245 103.345 27.455 103.865 ;
        RECT 27.645 103.565 27.975 103.815 ;
        RECT 18.890 102.575 24.235 103.120 ;
        RECT 24.405 102.575 24.695 103.300 ;
        RECT 24.865 102.575 27.455 103.345 ;
        RECT 27.665 102.575 27.895 103.395 ;
        RECT 28.145 103.375 28.395 103.975 ;
        RECT 29.010 103.465 29.360 104.115 ;
        RECT 28.065 102.745 28.395 103.375 ;
        RECT 28.565 102.575 28.775 103.395 ;
        RECT 29.530 103.295 29.760 104.285 ;
        RECT 29.010 103.125 29.760 103.295 ;
        RECT 29.010 102.835 29.265 103.125 ;
        RECT 29.435 102.575 29.765 102.955 ;
        RECT 29.935 102.835 30.105 104.955 ;
        RECT 30.275 104.155 30.600 104.940 ;
        RECT 30.770 104.665 31.020 105.125 ;
        RECT 31.190 104.625 31.440 104.955 ;
        RECT 31.655 104.625 32.335 104.955 ;
        RECT 31.190 104.495 31.360 104.625 ;
        RECT 30.965 104.325 31.360 104.495 ;
        RECT 30.335 103.105 30.795 104.155 ;
        RECT 30.965 102.965 31.135 104.325 ;
        RECT 31.530 104.065 31.995 104.455 ;
        RECT 31.305 103.255 31.655 103.875 ;
        RECT 31.825 103.475 31.995 104.065 ;
        RECT 32.165 103.845 32.335 104.625 ;
        RECT 32.505 104.525 32.675 104.865 ;
        RECT 32.910 104.695 33.240 105.125 ;
        RECT 33.410 104.525 33.580 104.865 ;
        RECT 33.875 104.665 34.245 105.125 ;
        RECT 32.505 104.355 33.580 104.525 ;
        RECT 34.415 104.495 34.585 104.955 ;
        RECT 34.820 104.615 35.690 104.955 ;
        RECT 35.860 104.665 36.110 105.125 ;
        RECT 34.025 104.325 34.585 104.495 ;
        RECT 34.025 104.185 34.195 104.325 ;
        RECT 32.695 104.015 34.195 104.185 ;
        RECT 34.890 104.155 35.350 104.445 ;
        RECT 32.165 103.675 33.855 103.845 ;
        RECT 31.825 103.255 32.180 103.475 ;
        RECT 32.350 102.965 32.520 103.675 ;
        RECT 32.725 103.255 33.515 103.505 ;
        RECT 33.685 103.495 33.855 103.675 ;
        RECT 34.025 103.325 34.195 104.015 ;
        RECT 30.465 102.575 30.795 102.935 ;
        RECT 30.965 102.795 31.460 102.965 ;
        RECT 31.665 102.795 32.520 102.965 ;
        RECT 33.395 102.575 33.725 103.035 ;
        RECT 33.935 102.935 34.195 103.325 ;
        RECT 34.385 104.145 35.350 104.155 ;
        RECT 35.520 104.235 35.690 104.615 ;
        RECT 36.280 104.575 36.450 104.865 ;
        RECT 36.630 104.745 36.960 105.125 ;
        RECT 36.280 104.405 37.080 104.575 ;
        RECT 34.385 103.985 35.060 104.145 ;
        RECT 35.520 104.065 36.740 104.235 ;
        RECT 34.385 103.195 34.595 103.985 ;
        RECT 35.520 103.975 35.690 104.065 ;
        RECT 34.765 103.195 35.115 103.815 ;
        RECT 35.285 103.805 35.690 103.975 ;
        RECT 35.285 103.025 35.455 103.805 ;
        RECT 35.625 103.355 35.845 103.635 ;
        RECT 36.025 103.525 36.565 103.895 ;
        RECT 36.910 103.785 37.080 104.405 ;
        RECT 37.255 104.065 37.425 105.125 ;
        RECT 37.635 104.115 37.925 104.955 ;
        RECT 38.095 104.285 38.265 105.125 ;
        RECT 38.475 104.115 38.725 104.955 ;
        RECT 38.935 104.285 39.105 105.125 ;
        RECT 39.895 104.285 40.065 105.125 ;
        RECT 40.275 104.115 40.525 104.955 ;
        RECT 40.735 104.285 40.905 105.125 ;
        RECT 41.075 104.115 41.365 104.955 ;
        RECT 37.635 103.945 39.360 104.115 ;
        RECT 35.625 103.185 36.155 103.355 ;
        RECT 33.935 102.765 34.285 102.935 ;
        RECT 34.505 102.745 35.455 103.025 ;
        RECT 35.625 102.575 35.815 103.015 ;
        RECT 35.985 102.955 36.155 103.185 ;
        RECT 36.325 103.125 36.565 103.525 ;
        RECT 36.735 103.775 37.080 103.785 ;
        RECT 36.735 103.565 38.765 103.775 ;
        RECT 36.735 103.310 37.060 103.565 ;
        RECT 38.950 103.395 39.360 103.945 ;
        RECT 36.735 102.955 37.055 103.310 ;
        RECT 35.985 102.785 37.055 102.955 ;
        RECT 37.255 102.575 37.425 103.385 ;
        RECT 37.595 103.225 39.360 103.395 ;
        RECT 39.640 103.945 41.365 104.115 ;
        RECT 41.575 104.065 41.745 105.125 ;
        RECT 42.040 104.745 42.370 105.125 ;
        RECT 42.550 104.575 42.720 104.865 ;
        RECT 42.890 104.665 43.140 105.125 ;
        RECT 41.920 104.405 42.720 104.575 ;
        RECT 43.310 104.615 44.180 104.955 ;
        RECT 39.640 103.395 40.050 103.945 ;
        RECT 41.920 103.785 42.090 104.405 ;
        RECT 43.310 104.235 43.480 104.615 ;
        RECT 44.415 104.495 44.585 104.955 ;
        RECT 44.755 104.665 45.125 105.125 ;
        RECT 45.420 104.525 45.590 104.865 ;
        RECT 45.760 104.695 46.090 105.125 ;
        RECT 46.325 104.525 46.495 104.865 ;
        RECT 42.260 104.065 43.480 104.235 ;
        RECT 43.650 104.155 44.110 104.445 ;
        RECT 44.415 104.325 44.975 104.495 ;
        RECT 45.420 104.355 46.495 104.525 ;
        RECT 46.665 104.625 47.345 104.955 ;
        RECT 47.560 104.625 47.810 104.955 ;
        RECT 47.980 104.665 48.230 105.125 ;
        RECT 44.805 104.185 44.975 104.325 ;
        RECT 43.650 104.145 44.615 104.155 ;
        RECT 43.310 103.975 43.480 104.065 ;
        RECT 43.940 103.985 44.615 104.145 ;
        RECT 41.920 103.775 42.265 103.785 ;
        RECT 40.235 103.565 42.265 103.775 ;
        RECT 39.640 103.225 41.405 103.395 ;
        RECT 37.595 102.745 37.925 103.225 ;
        RECT 38.095 102.575 38.265 103.045 ;
        RECT 38.435 102.745 38.765 103.225 ;
        RECT 38.935 102.575 39.105 103.045 ;
        RECT 39.895 102.575 40.065 103.045 ;
        RECT 40.235 102.745 40.565 103.225 ;
        RECT 40.735 102.575 40.905 103.045 ;
        RECT 41.075 102.745 41.405 103.225 ;
        RECT 41.575 102.575 41.745 103.385 ;
        RECT 41.940 103.310 42.265 103.565 ;
        RECT 41.945 102.955 42.265 103.310 ;
        RECT 42.435 103.525 42.975 103.895 ;
        RECT 43.310 103.805 43.715 103.975 ;
        RECT 42.435 103.125 42.675 103.525 ;
        RECT 43.155 103.355 43.375 103.635 ;
        RECT 42.845 103.185 43.375 103.355 ;
        RECT 42.845 102.955 43.015 103.185 ;
        RECT 43.545 103.025 43.715 103.805 ;
        RECT 43.885 103.195 44.235 103.815 ;
        RECT 44.405 103.195 44.615 103.985 ;
        RECT 44.805 104.015 46.305 104.185 ;
        RECT 44.805 103.325 44.975 104.015 ;
        RECT 46.665 103.845 46.835 104.625 ;
        RECT 47.640 104.495 47.810 104.625 ;
        RECT 45.145 103.675 46.835 103.845 ;
        RECT 47.005 104.065 47.470 104.455 ;
        RECT 47.640 104.325 48.035 104.495 ;
        RECT 45.145 103.495 45.315 103.675 ;
        RECT 41.945 102.785 43.015 102.955 ;
        RECT 43.185 102.575 43.375 103.015 ;
        RECT 43.545 102.745 44.495 103.025 ;
        RECT 44.805 102.935 45.065 103.325 ;
        RECT 45.485 103.255 46.275 103.505 ;
        RECT 44.715 102.765 45.065 102.935 ;
        RECT 45.275 102.575 45.605 103.035 ;
        RECT 46.480 102.965 46.650 103.675 ;
        RECT 47.005 103.475 47.175 104.065 ;
        RECT 46.820 103.255 47.175 103.475 ;
        RECT 47.345 103.255 47.695 103.875 ;
        RECT 47.865 102.965 48.035 104.325 ;
        RECT 48.400 104.155 48.725 104.940 ;
        RECT 48.205 103.105 48.665 104.155 ;
        RECT 46.480 102.795 47.335 102.965 ;
        RECT 47.540 102.795 48.035 102.965 ;
        RECT 48.205 102.575 48.535 102.935 ;
        RECT 48.895 102.835 49.065 104.955 ;
        RECT 49.235 104.625 49.565 105.125 ;
        RECT 49.735 104.455 49.990 104.955 ;
        RECT 49.240 104.285 49.990 104.455 ;
        RECT 49.240 103.295 49.470 104.285 ;
        RECT 49.640 103.465 49.990 104.115 ;
        RECT 50.165 103.960 50.455 105.125 ;
        RECT 51.605 103.985 51.815 105.125 ;
        RECT 51.985 103.975 52.315 104.955 ;
        RECT 52.485 103.985 52.715 105.125 ;
        RECT 53.235 104.285 53.405 105.125 ;
        RECT 53.615 104.115 53.865 104.955 ;
        RECT 54.075 104.285 54.245 105.125 ;
        RECT 54.415 104.115 54.705 104.955 ;
        RECT 49.240 103.125 49.990 103.295 ;
        RECT 49.235 102.575 49.565 102.955 ;
        RECT 49.735 102.835 49.990 103.125 ;
        RECT 50.165 102.575 50.455 103.300 ;
        RECT 51.605 102.575 51.815 103.395 ;
        RECT 51.985 103.375 52.235 103.975 ;
        RECT 52.980 103.945 54.705 104.115 ;
        RECT 54.915 104.065 55.085 105.125 ;
        RECT 55.380 104.745 55.710 105.125 ;
        RECT 55.890 104.575 56.060 104.865 ;
        RECT 56.230 104.665 56.480 105.125 ;
        RECT 55.260 104.405 56.060 104.575 ;
        RECT 56.650 104.615 57.520 104.955 ;
        RECT 52.405 103.565 52.735 103.815 ;
        RECT 52.980 103.395 53.390 103.945 ;
        RECT 55.260 103.785 55.430 104.405 ;
        RECT 56.650 104.235 56.820 104.615 ;
        RECT 57.755 104.495 57.925 104.955 ;
        RECT 58.095 104.665 58.465 105.125 ;
        RECT 58.760 104.525 58.930 104.865 ;
        RECT 59.100 104.695 59.430 105.125 ;
        RECT 59.665 104.525 59.835 104.865 ;
        RECT 55.600 104.065 56.820 104.235 ;
        RECT 56.990 104.155 57.450 104.445 ;
        RECT 57.755 104.325 58.315 104.495 ;
        RECT 58.760 104.355 59.835 104.525 ;
        RECT 60.005 104.625 60.685 104.955 ;
        RECT 60.900 104.625 61.150 104.955 ;
        RECT 61.320 104.665 61.570 105.125 ;
        RECT 58.145 104.185 58.315 104.325 ;
        RECT 56.990 104.145 57.955 104.155 ;
        RECT 56.650 103.975 56.820 104.065 ;
        RECT 57.280 103.985 57.955 104.145 ;
        RECT 55.260 103.775 55.605 103.785 ;
        RECT 53.575 103.565 55.605 103.775 ;
        RECT 51.985 102.745 52.315 103.375 ;
        RECT 52.485 102.575 52.715 103.395 ;
        RECT 52.980 103.225 54.745 103.395 ;
        RECT 53.235 102.575 53.405 103.045 ;
        RECT 53.575 102.745 53.905 103.225 ;
        RECT 54.075 102.575 54.245 103.045 ;
        RECT 54.415 102.745 54.745 103.225 ;
        RECT 54.915 102.575 55.085 103.385 ;
        RECT 55.280 103.310 55.605 103.565 ;
        RECT 55.285 102.955 55.605 103.310 ;
        RECT 55.775 103.525 56.315 103.895 ;
        RECT 56.650 103.805 57.055 103.975 ;
        RECT 55.775 103.125 56.015 103.525 ;
        RECT 56.495 103.355 56.715 103.635 ;
        RECT 56.185 103.185 56.715 103.355 ;
        RECT 56.185 102.955 56.355 103.185 ;
        RECT 56.885 103.025 57.055 103.805 ;
        RECT 57.225 103.195 57.575 103.815 ;
        RECT 57.745 103.195 57.955 103.985 ;
        RECT 58.145 104.015 59.645 104.185 ;
        RECT 58.145 103.325 58.315 104.015 ;
        RECT 60.005 103.845 60.175 104.625 ;
        RECT 60.980 104.495 61.150 104.625 ;
        RECT 58.485 103.675 60.175 103.845 ;
        RECT 60.345 104.065 60.810 104.455 ;
        RECT 60.980 104.325 61.375 104.495 ;
        RECT 58.485 103.495 58.655 103.675 ;
        RECT 55.285 102.785 56.355 102.955 ;
        RECT 56.525 102.575 56.715 103.015 ;
        RECT 56.885 102.745 57.835 103.025 ;
        RECT 58.145 102.935 58.405 103.325 ;
        RECT 58.825 103.255 59.615 103.505 ;
        RECT 58.055 102.765 58.405 102.935 ;
        RECT 58.615 102.575 58.945 103.035 ;
        RECT 59.820 102.965 59.990 103.675 ;
        RECT 60.345 103.475 60.515 104.065 ;
        RECT 60.160 103.255 60.515 103.475 ;
        RECT 60.685 103.255 61.035 103.875 ;
        RECT 61.205 102.965 61.375 104.325 ;
        RECT 61.740 104.155 62.065 104.940 ;
        RECT 61.545 103.105 62.005 104.155 ;
        RECT 59.820 102.795 60.675 102.965 ;
        RECT 60.880 102.795 61.375 102.965 ;
        RECT 61.545 102.575 61.875 102.935 ;
        RECT 62.235 102.835 62.405 104.955 ;
        RECT 62.575 104.625 62.905 105.125 ;
        RECT 63.075 104.455 63.330 104.955 ;
        RECT 62.580 104.285 63.330 104.455 ;
        RECT 63.815 104.285 63.985 105.125 ;
        RECT 62.580 103.295 62.810 104.285 ;
        RECT 64.195 104.115 64.445 104.955 ;
        RECT 64.655 104.285 64.825 105.125 ;
        RECT 64.995 104.115 65.285 104.955 ;
        RECT 62.980 103.465 63.330 104.115 ;
        RECT 63.560 103.945 65.285 104.115 ;
        RECT 65.495 104.065 65.665 105.125 ;
        RECT 65.960 104.745 66.290 105.125 ;
        RECT 66.470 104.575 66.640 104.865 ;
        RECT 66.810 104.665 67.060 105.125 ;
        RECT 65.840 104.405 66.640 104.575 ;
        RECT 67.230 104.615 68.100 104.955 ;
        RECT 63.560 103.395 63.970 103.945 ;
        RECT 65.840 103.785 66.010 104.405 ;
        RECT 67.230 104.235 67.400 104.615 ;
        RECT 68.335 104.495 68.505 104.955 ;
        RECT 68.675 104.665 69.045 105.125 ;
        RECT 69.340 104.525 69.510 104.865 ;
        RECT 69.680 104.695 70.010 105.125 ;
        RECT 70.245 104.525 70.415 104.865 ;
        RECT 66.180 104.065 67.400 104.235 ;
        RECT 67.570 104.155 68.030 104.445 ;
        RECT 68.335 104.325 68.895 104.495 ;
        RECT 69.340 104.355 70.415 104.525 ;
        RECT 70.585 104.625 71.265 104.955 ;
        RECT 71.480 104.625 71.730 104.955 ;
        RECT 71.900 104.665 72.150 105.125 ;
        RECT 68.725 104.185 68.895 104.325 ;
        RECT 67.570 104.145 68.535 104.155 ;
        RECT 67.230 103.975 67.400 104.065 ;
        RECT 67.860 103.985 68.535 104.145 ;
        RECT 65.840 103.775 66.185 103.785 ;
        RECT 64.155 103.565 66.185 103.775 ;
        RECT 62.580 103.125 63.330 103.295 ;
        RECT 63.560 103.225 65.325 103.395 ;
        RECT 62.575 102.575 62.905 102.955 ;
        RECT 63.075 102.835 63.330 103.125 ;
        RECT 63.815 102.575 63.985 103.045 ;
        RECT 64.155 102.745 64.485 103.225 ;
        RECT 64.655 102.575 64.825 103.045 ;
        RECT 64.995 102.745 65.325 103.225 ;
        RECT 65.495 102.575 65.665 103.385 ;
        RECT 65.860 103.310 66.185 103.565 ;
        RECT 65.865 102.955 66.185 103.310 ;
        RECT 66.355 103.525 66.895 103.895 ;
        RECT 67.230 103.805 67.635 103.975 ;
        RECT 66.355 103.125 66.595 103.525 ;
        RECT 67.075 103.355 67.295 103.635 ;
        RECT 66.765 103.185 67.295 103.355 ;
        RECT 66.765 102.955 66.935 103.185 ;
        RECT 67.465 103.025 67.635 103.805 ;
        RECT 67.805 103.195 68.155 103.815 ;
        RECT 68.325 103.195 68.535 103.985 ;
        RECT 68.725 104.015 70.225 104.185 ;
        RECT 68.725 103.325 68.895 104.015 ;
        RECT 70.585 103.845 70.755 104.625 ;
        RECT 71.560 104.495 71.730 104.625 ;
        RECT 69.065 103.675 70.755 103.845 ;
        RECT 70.925 104.065 71.390 104.455 ;
        RECT 71.560 104.325 71.955 104.495 ;
        RECT 69.065 103.495 69.235 103.675 ;
        RECT 65.865 102.785 66.935 102.955 ;
        RECT 67.105 102.575 67.295 103.015 ;
        RECT 67.465 102.745 68.415 103.025 ;
        RECT 68.725 102.935 68.985 103.325 ;
        RECT 69.405 103.255 70.195 103.505 ;
        RECT 68.635 102.765 68.985 102.935 ;
        RECT 69.195 102.575 69.525 103.035 ;
        RECT 70.400 102.965 70.570 103.675 ;
        RECT 70.925 103.475 71.095 104.065 ;
        RECT 70.740 103.255 71.095 103.475 ;
        RECT 71.265 103.255 71.615 103.875 ;
        RECT 71.785 102.965 71.955 104.325 ;
        RECT 72.320 104.155 72.645 104.940 ;
        RECT 72.125 103.105 72.585 104.155 ;
        RECT 70.400 102.795 71.255 102.965 ;
        RECT 71.460 102.795 71.955 102.965 ;
        RECT 72.125 102.575 72.455 102.935 ;
        RECT 72.815 102.835 72.985 104.955 ;
        RECT 73.155 104.625 73.485 105.125 ;
        RECT 73.655 104.455 73.910 104.955 ;
        RECT 73.160 104.285 73.910 104.455 ;
        RECT 73.160 103.295 73.390 104.285 ;
        RECT 73.560 103.465 73.910 104.115 ;
        RECT 74.085 104.035 75.755 105.125 ;
        RECT 74.085 103.515 74.835 104.035 ;
        RECT 75.925 103.960 76.215 105.125 ;
        RECT 76.695 104.285 76.865 105.125 ;
        RECT 77.075 104.115 77.325 104.955 ;
        RECT 77.535 104.285 77.705 105.125 ;
        RECT 77.875 104.115 78.165 104.955 ;
        RECT 76.440 103.945 78.165 104.115 ;
        RECT 78.375 104.065 78.545 105.125 ;
        RECT 78.840 104.745 79.170 105.125 ;
        RECT 79.350 104.575 79.520 104.865 ;
        RECT 79.690 104.665 79.940 105.125 ;
        RECT 78.720 104.405 79.520 104.575 ;
        RECT 80.110 104.615 80.980 104.955 ;
        RECT 75.005 103.345 75.755 103.865 ;
        RECT 73.160 103.125 73.910 103.295 ;
        RECT 73.155 102.575 73.485 102.955 ;
        RECT 73.655 102.835 73.910 103.125 ;
        RECT 74.085 102.575 75.755 103.345 ;
        RECT 76.440 103.395 76.850 103.945 ;
        RECT 78.720 103.785 78.890 104.405 ;
        RECT 80.110 104.235 80.280 104.615 ;
        RECT 81.215 104.495 81.385 104.955 ;
        RECT 81.555 104.665 81.925 105.125 ;
        RECT 82.220 104.525 82.390 104.865 ;
        RECT 82.560 104.695 82.890 105.125 ;
        RECT 83.125 104.525 83.295 104.865 ;
        RECT 79.060 104.065 80.280 104.235 ;
        RECT 80.450 104.155 80.910 104.445 ;
        RECT 81.215 104.325 81.775 104.495 ;
        RECT 82.220 104.355 83.295 104.525 ;
        RECT 83.465 104.625 84.145 104.955 ;
        RECT 84.360 104.625 84.610 104.955 ;
        RECT 84.780 104.665 85.030 105.125 ;
        RECT 81.605 104.185 81.775 104.325 ;
        RECT 80.450 104.145 81.415 104.155 ;
        RECT 80.110 103.975 80.280 104.065 ;
        RECT 80.740 103.985 81.415 104.145 ;
        RECT 78.720 103.775 79.065 103.785 ;
        RECT 77.035 103.565 79.065 103.775 ;
        RECT 75.925 102.575 76.215 103.300 ;
        RECT 76.440 103.225 78.205 103.395 ;
        RECT 76.695 102.575 76.865 103.045 ;
        RECT 77.035 102.745 77.365 103.225 ;
        RECT 77.535 102.575 77.705 103.045 ;
        RECT 77.875 102.745 78.205 103.225 ;
        RECT 78.375 102.575 78.545 103.385 ;
        RECT 78.740 103.310 79.065 103.565 ;
        RECT 78.745 102.955 79.065 103.310 ;
        RECT 79.235 103.525 79.775 103.895 ;
        RECT 80.110 103.805 80.515 103.975 ;
        RECT 79.235 103.125 79.475 103.525 ;
        RECT 79.955 103.355 80.175 103.635 ;
        RECT 79.645 103.185 80.175 103.355 ;
        RECT 79.645 102.955 79.815 103.185 ;
        RECT 80.345 103.025 80.515 103.805 ;
        RECT 80.685 103.195 81.035 103.815 ;
        RECT 81.205 103.195 81.415 103.985 ;
        RECT 81.605 104.015 83.105 104.185 ;
        RECT 81.605 103.325 81.775 104.015 ;
        RECT 83.465 103.845 83.635 104.625 ;
        RECT 84.440 104.495 84.610 104.625 ;
        RECT 81.945 103.675 83.635 103.845 ;
        RECT 83.805 104.065 84.270 104.455 ;
        RECT 84.440 104.325 84.835 104.495 ;
        RECT 81.945 103.495 82.115 103.675 ;
        RECT 78.745 102.785 79.815 102.955 ;
        RECT 79.985 102.575 80.175 103.015 ;
        RECT 80.345 102.745 81.295 103.025 ;
        RECT 81.605 102.935 81.865 103.325 ;
        RECT 82.285 103.255 83.075 103.505 ;
        RECT 81.515 102.765 81.865 102.935 ;
        RECT 82.075 102.575 82.405 103.035 ;
        RECT 83.280 102.965 83.450 103.675 ;
        RECT 83.805 103.475 83.975 104.065 ;
        RECT 83.620 103.255 83.975 103.475 ;
        RECT 84.145 103.255 84.495 103.875 ;
        RECT 84.665 102.965 84.835 104.325 ;
        RECT 85.200 104.155 85.525 104.940 ;
        RECT 85.005 103.105 85.465 104.155 ;
        RECT 83.280 102.795 84.135 102.965 ;
        RECT 84.340 102.795 84.835 102.965 ;
        RECT 85.005 102.575 85.335 102.935 ;
        RECT 85.695 102.835 85.865 104.955 ;
        RECT 86.035 104.625 86.365 105.125 ;
        RECT 86.535 104.455 86.790 104.955 ;
        RECT 86.040 104.285 86.790 104.455 ;
        RECT 87.275 104.285 87.445 105.125 ;
        RECT 86.040 103.295 86.270 104.285 ;
        RECT 87.655 104.115 87.905 104.955 ;
        RECT 88.115 104.285 88.285 105.125 ;
        RECT 88.455 104.115 88.745 104.955 ;
        RECT 86.440 103.465 86.790 104.115 ;
        RECT 87.020 103.945 88.745 104.115 ;
        RECT 88.955 104.065 89.125 105.125 ;
        RECT 89.420 104.745 89.750 105.125 ;
        RECT 89.930 104.575 90.100 104.865 ;
        RECT 90.270 104.665 90.520 105.125 ;
        RECT 89.300 104.405 90.100 104.575 ;
        RECT 90.690 104.615 91.560 104.955 ;
        RECT 87.020 103.395 87.430 103.945 ;
        RECT 89.300 103.785 89.470 104.405 ;
        RECT 90.690 104.235 90.860 104.615 ;
        RECT 91.795 104.495 91.965 104.955 ;
        RECT 92.135 104.665 92.505 105.125 ;
        RECT 92.800 104.525 92.970 104.865 ;
        RECT 93.140 104.695 93.470 105.125 ;
        RECT 93.705 104.525 93.875 104.865 ;
        RECT 89.640 104.065 90.860 104.235 ;
        RECT 91.030 104.155 91.490 104.445 ;
        RECT 91.795 104.325 92.355 104.495 ;
        RECT 92.800 104.355 93.875 104.525 ;
        RECT 94.045 104.625 94.725 104.955 ;
        RECT 94.940 104.625 95.190 104.955 ;
        RECT 95.360 104.665 95.610 105.125 ;
        RECT 92.185 104.185 92.355 104.325 ;
        RECT 91.030 104.145 91.995 104.155 ;
        RECT 90.690 103.975 90.860 104.065 ;
        RECT 91.320 103.985 91.995 104.145 ;
        RECT 89.300 103.775 89.645 103.785 ;
        RECT 87.615 103.565 89.645 103.775 ;
        RECT 86.040 103.125 86.790 103.295 ;
        RECT 87.020 103.225 88.785 103.395 ;
        RECT 86.035 102.575 86.365 102.955 ;
        RECT 86.535 102.835 86.790 103.125 ;
        RECT 87.275 102.575 87.445 103.045 ;
        RECT 87.615 102.745 87.945 103.225 ;
        RECT 88.115 102.575 88.285 103.045 ;
        RECT 88.455 102.745 88.785 103.225 ;
        RECT 88.955 102.575 89.125 103.385 ;
        RECT 89.320 103.310 89.645 103.565 ;
        RECT 89.325 102.955 89.645 103.310 ;
        RECT 89.815 103.525 90.355 103.895 ;
        RECT 90.690 103.805 91.095 103.975 ;
        RECT 89.815 103.125 90.055 103.525 ;
        RECT 90.535 103.355 90.755 103.635 ;
        RECT 90.225 103.185 90.755 103.355 ;
        RECT 90.225 102.955 90.395 103.185 ;
        RECT 90.925 103.025 91.095 103.805 ;
        RECT 91.265 103.195 91.615 103.815 ;
        RECT 91.785 103.195 91.995 103.985 ;
        RECT 92.185 104.015 93.685 104.185 ;
        RECT 92.185 103.325 92.355 104.015 ;
        RECT 94.045 103.845 94.215 104.625 ;
        RECT 95.020 104.495 95.190 104.625 ;
        RECT 92.525 103.675 94.215 103.845 ;
        RECT 94.385 104.065 94.850 104.455 ;
        RECT 95.020 104.325 95.415 104.495 ;
        RECT 92.525 103.495 92.695 103.675 ;
        RECT 89.325 102.785 90.395 102.955 ;
        RECT 90.565 102.575 90.755 103.015 ;
        RECT 90.925 102.745 91.875 103.025 ;
        RECT 92.185 102.935 92.445 103.325 ;
        RECT 92.865 103.255 93.655 103.505 ;
        RECT 92.095 102.765 92.445 102.935 ;
        RECT 92.655 102.575 92.985 103.035 ;
        RECT 93.860 102.965 94.030 103.675 ;
        RECT 94.385 103.475 94.555 104.065 ;
        RECT 94.200 103.255 94.555 103.475 ;
        RECT 94.725 103.255 95.075 103.875 ;
        RECT 95.245 102.965 95.415 104.325 ;
        RECT 95.780 104.155 96.105 104.940 ;
        RECT 95.585 103.105 96.045 104.155 ;
        RECT 93.860 102.795 94.715 102.965 ;
        RECT 94.920 102.795 95.415 102.965 ;
        RECT 95.585 102.575 95.915 102.935 ;
        RECT 96.275 102.835 96.445 104.955 ;
        RECT 96.615 104.625 96.945 105.125 ;
        RECT 97.115 104.455 97.370 104.955 ;
        RECT 96.620 104.285 97.370 104.455 ;
        RECT 96.620 103.295 96.850 104.285 ;
        RECT 97.020 103.465 97.370 104.115 ;
        RECT 98.005 104.035 101.515 105.125 ;
        RECT 98.005 103.515 99.695 104.035 ;
        RECT 101.685 103.960 101.975 105.125 ;
        RECT 102.455 104.285 102.625 105.125 ;
        RECT 102.835 104.115 103.085 104.955 ;
        RECT 103.295 104.285 103.465 105.125 ;
        RECT 103.635 104.115 103.925 104.955 ;
        RECT 102.200 103.945 103.925 104.115 ;
        RECT 104.135 104.065 104.305 105.125 ;
        RECT 104.600 104.745 104.930 105.125 ;
        RECT 105.110 104.575 105.280 104.865 ;
        RECT 105.450 104.665 105.700 105.125 ;
        RECT 104.480 104.405 105.280 104.575 ;
        RECT 105.870 104.615 106.740 104.955 ;
        RECT 99.865 103.345 101.515 103.865 ;
        RECT 96.620 103.125 97.370 103.295 ;
        RECT 96.615 102.575 96.945 102.955 ;
        RECT 97.115 102.835 97.370 103.125 ;
        RECT 98.005 102.575 101.515 103.345 ;
        RECT 102.200 103.395 102.610 103.945 ;
        RECT 104.480 103.785 104.650 104.405 ;
        RECT 105.870 104.235 106.040 104.615 ;
        RECT 106.975 104.495 107.145 104.955 ;
        RECT 107.315 104.665 107.685 105.125 ;
        RECT 107.980 104.525 108.150 104.865 ;
        RECT 108.320 104.695 108.650 105.125 ;
        RECT 108.885 104.525 109.055 104.865 ;
        RECT 104.820 104.065 106.040 104.235 ;
        RECT 106.210 104.155 106.670 104.445 ;
        RECT 106.975 104.325 107.535 104.495 ;
        RECT 107.980 104.355 109.055 104.525 ;
        RECT 109.225 104.625 109.905 104.955 ;
        RECT 110.120 104.625 110.370 104.955 ;
        RECT 110.540 104.665 110.790 105.125 ;
        RECT 107.365 104.185 107.535 104.325 ;
        RECT 106.210 104.145 107.175 104.155 ;
        RECT 105.870 103.975 106.040 104.065 ;
        RECT 106.500 103.985 107.175 104.145 ;
        RECT 104.480 103.775 104.825 103.785 ;
        RECT 102.795 103.565 104.825 103.775 ;
        RECT 101.685 102.575 101.975 103.300 ;
        RECT 102.200 103.225 103.965 103.395 ;
        RECT 102.455 102.575 102.625 103.045 ;
        RECT 102.795 102.745 103.125 103.225 ;
        RECT 103.295 102.575 103.465 103.045 ;
        RECT 103.635 102.745 103.965 103.225 ;
        RECT 104.135 102.575 104.305 103.385 ;
        RECT 104.500 103.310 104.825 103.565 ;
        RECT 104.505 102.955 104.825 103.310 ;
        RECT 104.995 103.525 105.535 103.895 ;
        RECT 105.870 103.805 106.275 103.975 ;
        RECT 104.995 103.125 105.235 103.525 ;
        RECT 105.715 103.355 105.935 103.635 ;
        RECT 105.405 103.185 105.935 103.355 ;
        RECT 105.405 102.955 105.575 103.185 ;
        RECT 106.105 103.025 106.275 103.805 ;
        RECT 106.445 103.195 106.795 103.815 ;
        RECT 106.965 103.195 107.175 103.985 ;
        RECT 107.365 104.015 108.865 104.185 ;
        RECT 107.365 103.325 107.535 104.015 ;
        RECT 109.225 103.845 109.395 104.625 ;
        RECT 110.200 104.495 110.370 104.625 ;
        RECT 107.705 103.675 109.395 103.845 ;
        RECT 109.565 104.065 110.030 104.455 ;
        RECT 110.200 104.325 110.595 104.495 ;
        RECT 107.705 103.495 107.875 103.675 ;
        RECT 104.505 102.785 105.575 102.955 ;
        RECT 105.745 102.575 105.935 103.015 ;
        RECT 106.105 102.745 107.055 103.025 ;
        RECT 107.365 102.935 107.625 103.325 ;
        RECT 108.045 103.255 108.835 103.505 ;
        RECT 107.275 102.765 107.625 102.935 ;
        RECT 107.835 102.575 108.165 103.035 ;
        RECT 109.040 102.965 109.210 103.675 ;
        RECT 109.565 103.475 109.735 104.065 ;
        RECT 109.380 103.255 109.735 103.475 ;
        RECT 109.905 103.255 110.255 103.875 ;
        RECT 110.425 102.965 110.595 104.325 ;
        RECT 110.960 104.155 111.285 104.940 ;
        RECT 110.765 103.105 111.225 104.155 ;
        RECT 109.040 102.795 109.895 102.965 ;
        RECT 110.100 102.795 110.595 102.965 ;
        RECT 110.765 102.575 111.095 102.935 ;
        RECT 111.455 102.835 111.625 104.955 ;
        RECT 111.795 104.625 112.125 105.125 ;
        RECT 112.295 104.455 112.550 104.955 ;
        RECT 111.800 104.285 112.550 104.455 ;
        RECT 112.730 104.455 112.985 104.955 ;
        RECT 113.155 104.625 113.485 105.125 ;
        RECT 112.730 104.285 113.480 104.455 ;
        RECT 111.800 103.295 112.030 104.285 ;
        RECT 112.200 103.465 112.550 104.115 ;
        RECT 112.730 103.465 113.080 104.115 ;
        RECT 113.250 103.295 113.480 104.285 ;
        RECT 111.800 103.125 112.550 103.295 ;
        RECT 111.795 102.575 112.125 102.955 ;
        RECT 112.295 102.835 112.550 103.125 ;
        RECT 112.730 103.125 113.480 103.295 ;
        RECT 112.730 102.835 112.985 103.125 ;
        RECT 113.155 102.575 113.485 102.955 ;
        RECT 113.655 102.835 113.825 104.955 ;
        RECT 113.995 104.155 114.320 104.940 ;
        RECT 114.490 104.665 114.740 105.125 ;
        RECT 114.910 104.625 115.160 104.955 ;
        RECT 115.375 104.625 116.055 104.955 ;
        RECT 114.910 104.495 115.080 104.625 ;
        RECT 114.685 104.325 115.080 104.495 ;
        RECT 114.055 103.105 114.515 104.155 ;
        RECT 114.685 102.965 114.855 104.325 ;
        RECT 115.250 104.065 115.715 104.455 ;
        RECT 115.025 103.255 115.375 103.875 ;
        RECT 115.545 103.475 115.715 104.065 ;
        RECT 115.885 103.845 116.055 104.625 ;
        RECT 116.225 104.525 116.395 104.865 ;
        RECT 116.630 104.695 116.960 105.125 ;
        RECT 117.130 104.525 117.300 104.865 ;
        RECT 117.595 104.665 117.965 105.125 ;
        RECT 116.225 104.355 117.300 104.525 ;
        RECT 118.135 104.495 118.305 104.955 ;
        RECT 118.540 104.615 119.410 104.955 ;
        RECT 119.580 104.665 119.830 105.125 ;
        RECT 117.745 104.325 118.305 104.495 ;
        RECT 117.745 104.185 117.915 104.325 ;
        RECT 116.415 104.015 117.915 104.185 ;
        RECT 118.610 104.155 119.070 104.445 ;
        RECT 115.885 103.675 117.575 103.845 ;
        RECT 115.545 103.255 115.900 103.475 ;
        RECT 116.070 102.965 116.240 103.675 ;
        RECT 116.445 103.255 117.235 103.505 ;
        RECT 117.405 103.495 117.575 103.675 ;
        RECT 117.745 103.325 117.915 104.015 ;
        RECT 114.185 102.575 114.515 102.935 ;
        RECT 114.685 102.795 115.180 102.965 ;
        RECT 115.385 102.795 116.240 102.965 ;
        RECT 117.115 102.575 117.445 103.035 ;
        RECT 117.655 102.935 117.915 103.325 ;
        RECT 118.105 104.145 119.070 104.155 ;
        RECT 119.240 104.235 119.410 104.615 ;
        RECT 120.000 104.575 120.170 104.865 ;
        RECT 120.350 104.745 120.680 105.125 ;
        RECT 120.000 104.405 120.800 104.575 ;
        RECT 118.105 103.985 118.780 104.145 ;
        RECT 119.240 104.065 120.460 104.235 ;
        RECT 118.105 103.195 118.315 103.985 ;
        RECT 119.240 103.975 119.410 104.065 ;
        RECT 118.485 103.195 118.835 103.815 ;
        RECT 119.005 103.805 119.410 103.975 ;
        RECT 119.005 103.025 119.175 103.805 ;
        RECT 119.345 103.355 119.565 103.635 ;
        RECT 119.745 103.525 120.285 103.895 ;
        RECT 120.630 103.785 120.800 104.405 ;
        RECT 120.975 104.065 121.145 105.125 ;
        RECT 121.355 104.115 121.645 104.955 ;
        RECT 121.815 104.285 121.985 105.125 ;
        RECT 122.195 104.115 122.445 104.955 ;
        RECT 122.655 104.285 122.825 105.125 ;
        RECT 121.355 103.945 123.080 104.115 ;
        RECT 119.345 103.185 119.875 103.355 ;
        RECT 117.655 102.765 118.005 102.935 ;
        RECT 118.225 102.745 119.175 103.025 ;
        RECT 119.345 102.575 119.535 103.015 ;
        RECT 119.705 102.955 119.875 103.185 ;
        RECT 120.045 103.125 120.285 103.525 ;
        RECT 120.455 103.775 120.800 103.785 ;
        RECT 120.455 103.565 122.485 103.775 ;
        RECT 120.455 103.310 120.780 103.565 ;
        RECT 122.670 103.395 123.080 103.945 ;
        RECT 123.305 104.035 124.975 105.125 ;
        RECT 125.145 104.050 125.415 104.955 ;
        RECT 125.585 104.365 125.915 105.125 ;
        RECT 126.095 104.195 126.275 104.955 ;
        RECT 123.305 103.515 124.055 104.035 ;
        RECT 120.455 102.955 120.775 103.310 ;
        RECT 119.705 102.785 120.775 102.955 ;
        RECT 120.975 102.575 121.145 103.385 ;
        RECT 121.315 103.225 123.080 103.395 ;
        RECT 124.225 103.345 124.975 103.865 ;
        RECT 121.315 102.745 121.645 103.225 ;
        RECT 121.815 102.575 121.985 103.045 ;
        RECT 122.155 102.745 122.485 103.225 ;
        RECT 122.655 102.575 122.825 103.045 ;
        RECT 123.305 102.575 124.975 103.345 ;
        RECT 125.145 103.250 125.325 104.050 ;
        RECT 125.600 104.025 126.275 104.195 ;
        RECT 126.525 104.035 127.735 105.125 ;
        RECT 125.600 103.880 125.770 104.025 ;
        RECT 125.495 103.550 125.770 103.880 ;
        RECT 125.600 103.295 125.770 103.550 ;
        RECT 125.995 103.475 126.335 103.845 ;
        RECT 126.525 103.495 127.045 104.035 ;
        RECT 127.215 103.325 127.735 103.865 ;
        RECT 125.145 102.745 125.405 103.250 ;
        RECT 125.600 103.125 126.265 103.295 ;
        RECT 125.585 102.575 125.915 102.955 ;
        RECT 126.095 102.745 126.265 103.125 ;
        RECT 126.525 102.575 127.735 103.325 ;
        RECT 14.660 102.405 127.820 102.575 ;
        RECT 14.745 101.655 15.955 102.405 ;
        RECT 14.745 101.115 15.265 101.655 ;
        RECT 16.125 101.635 18.715 102.405 ;
        RECT 18.890 101.860 24.235 102.405 ;
        RECT 15.435 100.945 15.955 101.485 ;
        RECT 14.745 99.855 15.955 100.945 ;
        RECT 16.125 100.945 17.335 101.465 ;
        RECT 17.505 101.115 18.715 101.635 ;
        RECT 16.125 99.855 18.715 100.945 ;
        RECT 20.480 100.290 20.830 101.540 ;
        RECT 22.310 101.030 22.650 101.860 ;
        RECT 24.405 101.680 24.695 102.405 ;
        RECT 25.175 101.935 25.345 102.405 ;
        RECT 25.515 101.755 25.845 102.235 ;
        RECT 26.015 101.935 26.185 102.405 ;
        RECT 26.355 101.755 26.685 102.235 ;
        RECT 24.920 101.585 26.685 101.755 ;
        RECT 26.855 101.595 27.025 102.405 ;
        RECT 27.225 102.025 28.295 102.195 ;
        RECT 27.225 101.670 27.545 102.025 ;
        RECT 24.920 101.035 25.330 101.585 ;
        RECT 27.220 101.415 27.545 101.670 ;
        RECT 25.515 101.205 27.545 101.415 ;
        RECT 27.200 101.195 27.545 101.205 ;
        RECT 27.715 101.455 27.955 101.855 ;
        RECT 28.125 101.795 28.295 102.025 ;
        RECT 28.465 101.965 28.655 102.405 ;
        RECT 28.825 101.955 29.775 102.235 ;
        RECT 29.995 102.045 30.345 102.215 ;
        RECT 28.125 101.625 28.655 101.795 ;
        RECT 18.890 99.855 24.235 100.290 ;
        RECT 24.405 99.855 24.695 101.020 ;
        RECT 24.920 100.865 26.645 101.035 ;
        RECT 25.175 99.855 25.345 100.695 ;
        RECT 25.555 100.025 25.805 100.865 ;
        RECT 26.015 99.855 26.185 100.695 ;
        RECT 26.355 100.025 26.645 100.865 ;
        RECT 26.855 99.855 27.025 100.915 ;
        RECT 27.200 100.575 27.370 101.195 ;
        RECT 27.715 101.085 28.255 101.455 ;
        RECT 28.435 101.345 28.655 101.625 ;
        RECT 28.825 101.175 28.995 101.955 ;
        RECT 28.590 101.005 28.995 101.175 ;
        RECT 29.165 101.165 29.515 101.785 ;
        RECT 28.590 100.915 28.760 101.005 ;
        RECT 29.685 100.995 29.895 101.785 ;
        RECT 27.540 100.745 28.760 100.915 ;
        RECT 29.220 100.835 29.895 100.995 ;
        RECT 27.200 100.405 28.000 100.575 ;
        RECT 27.320 99.855 27.650 100.235 ;
        RECT 27.830 100.115 28.000 100.405 ;
        RECT 28.590 100.365 28.760 100.745 ;
        RECT 28.930 100.825 29.895 100.835 ;
        RECT 30.085 101.655 30.345 102.045 ;
        RECT 30.555 101.945 30.885 102.405 ;
        RECT 31.760 102.015 32.615 102.185 ;
        RECT 32.820 102.015 33.315 102.185 ;
        RECT 33.485 102.045 33.815 102.405 ;
        RECT 30.085 100.965 30.255 101.655 ;
        RECT 30.425 101.305 30.595 101.485 ;
        RECT 30.765 101.475 31.555 101.725 ;
        RECT 31.760 101.305 31.930 102.015 ;
        RECT 32.100 101.505 32.455 101.725 ;
        RECT 30.425 101.135 32.115 101.305 ;
        RECT 28.930 100.535 29.390 100.825 ;
        RECT 30.085 100.795 31.585 100.965 ;
        RECT 30.085 100.655 30.255 100.795 ;
        RECT 29.695 100.485 30.255 100.655 ;
        RECT 28.170 99.855 28.420 100.315 ;
        RECT 28.590 100.025 29.460 100.365 ;
        RECT 29.695 100.025 29.865 100.485 ;
        RECT 30.700 100.455 31.775 100.625 ;
        RECT 30.035 99.855 30.405 100.315 ;
        RECT 30.700 100.115 30.870 100.455 ;
        RECT 31.040 99.855 31.370 100.285 ;
        RECT 31.605 100.115 31.775 100.455 ;
        RECT 31.945 100.355 32.115 101.135 ;
        RECT 32.285 100.915 32.455 101.505 ;
        RECT 32.625 101.105 32.975 101.725 ;
        RECT 32.285 100.525 32.750 100.915 ;
        RECT 33.145 100.655 33.315 102.015 ;
        RECT 33.485 100.825 33.945 101.875 ;
        RECT 32.920 100.485 33.315 100.655 ;
        RECT 32.920 100.355 33.090 100.485 ;
        RECT 31.945 100.025 32.625 100.355 ;
        RECT 32.840 100.025 33.090 100.355 ;
        RECT 33.260 99.855 33.510 100.315 ;
        RECT 33.680 100.040 34.005 100.825 ;
        RECT 34.175 100.025 34.345 102.145 ;
        RECT 34.515 102.025 34.845 102.405 ;
        RECT 35.015 101.855 35.270 102.145 ;
        RECT 34.520 101.685 35.270 101.855 ;
        RECT 34.520 100.695 34.750 101.685 ;
        RECT 35.445 101.635 37.115 102.405 ;
        RECT 37.285 101.680 37.575 102.405 ;
        RECT 37.745 101.655 38.955 102.405 ;
        RECT 39.130 101.860 44.475 102.405 ;
        RECT 44.650 101.860 49.995 102.405 ;
        RECT 34.920 100.865 35.270 101.515 ;
        RECT 35.445 100.945 36.195 101.465 ;
        RECT 36.365 101.115 37.115 101.635 ;
        RECT 34.520 100.525 35.270 100.695 ;
        RECT 34.515 99.855 34.845 100.355 ;
        RECT 35.015 100.025 35.270 100.525 ;
        RECT 35.445 99.855 37.115 100.945 ;
        RECT 37.285 99.855 37.575 101.020 ;
        RECT 37.745 100.945 38.265 101.485 ;
        RECT 38.435 101.115 38.955 101.655 ;
        RECT 37.745 99.855 38.955 100.945 ;
        RECT 40.720 100.290 41.070 101.540 ;
        RECT 42.550 101.030 42.890 101.860 ;
        RECT 46.240 100.290 46.590 101.540 ;
        RECT 48.070 101.030 48.410 101.860 ;
        RECT 50.165 101.680 50.455 102.405 ;
        RECT 50.625 101.655 51.835 102.405 ;
        RECT 52.010 101.860 57.355 102.405 ;
        RECT 57.530 101.860 62.875 102.405 ;
        RECT 39.130 99.855 44.475 100.290 ;
        RECT 44.650 99.855 49.995 100.290 ;
        RECT 50.165 99.855 50.455 101.020 ;
        RECT 50.625 100.945 51.145 101.485 ;
        RECT 51.315 101.115 51.835 101.655 ;
        RECT 50.625 99.855 51.835 100.945 ;
        RECT 53.600 100.290 53.950 101.540 ;
        RECT 55.430 101.030 55.770 101.860 ;
        RECT 59.120 100.290 59.470 101.540 ;
        RECT 60.950 101.030 61.290 101.860 ;
        RECT 63.045 101.680 63.335 102.405 ;
        RECT 63.505 101.655 64.715 102.405 ;
        RECT 64.890 101.860 70.235 102.405 ;
        RECT 70.410 101.860 75.755 102.405 ;
        RECT 52.010 99.855 57.355 100.290 ;
        RECT 57.530 99.855 62.875 100.290 ;
        RECT 63.045 99.855 63.335 101.020 ;
        RECT 63.505 100.945 64.025 101.485 ;
        RECT 64.195 101.115 64.715 101.655 ;
        RECT 63.505 99.855 64.715 100.945 ;
        RECT 66.480 100.290 66.830 101.540 ;
        RECT 68.310 101.030 68.650 101.860 ;
        RECT 72.000 100.290 72.350 101.540 ;
        RECT 73.830 101.030 74.170 101.860 ;
        RECT 75.925 101.680 76.215 102.405 ;
        RECT 76.385 101.655 77.595 102.405 ;
        RECT 77.770 101.860 83.115 102.405 ;
        RECT 83.290 101.860 88.635 102.405 ;
        RECT 64.890 99.855 70.235 100.290 ;
        RECT 70.410 99.855 75.755 100.290 ;
        RECT 75.925 99.855 76.215 101.020 ;
        RECT 76.385 100.945 76.905 101.485 ;
        RECT 77.075 101.115 77.595 101.655 ;
        RECT 76.385 99.855 77.595 100.945 ;
        RECT 79.360 100.290 79.710 101.540 ;
        RECT 81.190 101.030 81.530 101.860 ;
        RECT 84.880 100.290 85.230 101.540 ;
        RECT 86.710 101.030 87.050 101.860 ;
        RECT 88.805 101.680 89.095 102.405 ;
        RECT 89.265 101.635 90.935 102.405 ;
        RECT 91.415 101.935 91.585 102.405 ;
        RECT 91.755 101.755 92.085 102.235 ;
        RECT 92.255 101.935 92.425 102.405 ;
        RECT 92.595 101.755 92.925 102.235 ;
        RECT 77.770 99.855 83.115 100.290 ;
        RECT 83.290 99.855 88.635 100.290 ;
        RECT 88.805 99.855 89.095 101.020 ;
        RECT 89.265 100.945 90.015 101.465 ;
        RECT 90.185 101.115 90.935 101.635 ;
        RECT 91.160 101.585 92.925 101.755 ;
        RECT 93.095 101.595 93.265 102.405 ;
        RECT 93.465 102.025 94.535 102.195 ;
        RECT 93.465 101.670 93.785 102.025 ;
        RECT 91.160 101.035 91.570 101.585 ;
        RECT 93.460 101.415 93.785 101.670 ;
        RECT 91.755 101.205 93.785 101.415 ;
        RECT 93.440 101.195 93.785 101.205 ;
        RECT 93.955 101.455 94.195 101.855 ;
        RECT 94.365 101.795 94.535 102.025 ;
        RECT 94.705 101.965 94.895 102.405 ;
        RECT 95.065 101.955 96.015 102.235 ;
        RECT 96.235 102.045 96.585 102.215 ;
        RECT 94.365 101.625 94.895 101.795 ;
        RECT 89.265 99.855 90.935 100.945 ;
        RECT 91.160 100.865 92.885 101.035 ;
        RECT 91.415 99.855 91.585 100.695 ;
        RECT 91.795 100.025 92.045 100.865 ;
        RECT 92.255 99.855 92.425 100.695 ;
        RECT 92.595 100.025 92.885 100.865 ;
        RECT 93.095 99.855 93.265 100.915 ;
        RECT 93.440 100.575 93.610 101.195 ;
        RECT 93.955 101.085 94.495 101.455 ;
        RECT 94.675 101.345 94.895 101.625 ;
        RECT 95.065 101.175 95.235 101.955 ;
        RECT 94.830 101.005 95.235 101.175 ;
        RECT 95.405 101.165 95.755 101.785 ;
        RECT 94.830 100.915 95.000 101.005 ;
        RECT 95.925 100.995 96.135 101.785 ;
        RECT 93.780 100.745 95.000 100.915 ;
        RECT 95.460 100.835 96.135 100.995 ;
        RECT 93.440 100.405 94.240 100.575 ;
        RECT 93.560 99.855 93.890 100.235 ;
        RECT 94.070 100.115 94.240 100.405 ;
        RECT 94.830 100.365 95.000 100.745 ;
        RECT 95.170 100.825 96.135 100.835 ;
        RECT 96.325 101.655 96.585 102.045 ;
        RECT 96.795 101.945 97.125 102.405 ;
        RECT 98.000 102.015 98.855 102.185 ;
        RECT 99.060 102.015 99.555 102.185 ;
        RECT 99.725 102.045 100.055 102.405 ;
        RECT 96.325 100.965 96.495 101.655 ;
        RECT 96.665 101.305 96.835 101.485 ;
        RECT 97.005 101.475 97.795 101.725 ;
        RECT 98.000 101.305 98.170 102.015 ;
        RECT 98.340 101.505 98.695 101.725 ;
        RECT 96.665 101.135 98.355 101.305 ;
        RECT 95.170 100.535 95.630 100.825 ;
        RECT 96.325 100.795 97.825 100.965 ;
        RECT 96.325 100.655 96.495 100.795 ;
        RECT 95.935 100.485 96.495 100.655 ;
        RECT 94.410 99.855 94.660 100.315 ;
        RECT 94.830 100.025 95.700 100.365 ;
        RECT 95.935 100.025 96.105 100.485 ;
        RECT 96.940 100.455 98.015 100.625 ;
        RECT 96.275 99.855 96.645 100.315 ;
        RECT 96.940 100.115 97.110 100.455 ;
        RECT 97.280 99.855 97.610 100.285 ;
        RECT 97.845 100.115 98.015 100.455 ;
        RECT 98.185 100.355 98.355 101.135 ;
        RECT 98.525 100.915 98.695 101.505 ;
        RECT 98.865 101.105 99.215 101.725 ;
        RECT 98.525 100.525 98.990 100.915 ;
        RECT 99.385 100.655 99.555 102.015 ;
        RECT 99.725 100.825 100.185 101.875 ;
        RECT 99.160 100.485 99.555 100.655 ;
        RECT 99.160 100.355 99.330 100.485 ;
        RECT 98.185 100.025 98.865 100.355 ;
        RECT 99.080 100.025 99.330 100.355 ;
        RECT 99.500 99.855 99.750 100.315 ;
        RECT 99.920 100.040 100.245 100.825 ;
        RECT 100.415 100.025 100.585 102.145 ;
        RECT 100.755 102.025 101.085 102.405 ;
        RECT 101.255 101.855 101.510 102.145 ;
        RECT 100.760 101.685 101.510 101.855 ;
        RECT 100.760 100.695 100.990 101.685 ;
        RECT 101.685 101.680 101.975 102.405 ;
        RECT 102.145 101.655 103.355 102.405 ;
        RECT 103.530 101.860 108.875 102.405 ;
        RECT 109.050 101.860 114.395 102.405 ;
        RECT 101.160 100.865 101.510 101.515 ;
        RECT 100.760 100.525 101.510 100.695 ;
        RECT 100.755 99.855 101.085 100.355 ;
        RECT 101.255 100.025 101.510 100.525 ;
        RECT 101.685 99.855 101.975 101.020 ;
        RECT 102.145 100.945 102.665 101.485 ;
        RECT 102.835 101.115 103.355 101.655 ;
        RECT 102.145 99.855 103.355 100.945 ;
        RECT 105.120 100.290 105.470 101.540 ;
        RECT 106.950 101.030 107.290 101.860 ;
        RECT 110.640 100.290 110.990 101.540 ;
        RECT 112.470 101.030 112.810 101.860 ;
        RECT 114.565 101.680 114.855 102.405 ;
        RECT 115.945 101.635 119.455 102.405 ;
        RECT 103.530 99.855 108.875 100.290 ;
        RECT 109.050 99.855 114.395 100.290 ;
        RECT 114.565 99.855 114.855 101.020 ;
        RECT 115.945 100.945 117.635 101.465 ;
        RECT 117.805 101.115 119.455 101.635 ;
        RECT 119.665 101.585 119.895 102.405 ;
        RECT 120.065 101.605 120.395 102.235 ;
        RECT 119.645 101.165 119.975 101.415 ;
        RECT 120.145 101.005 120.395 101.605 ;
        RECT 120.565 101.585 120.775 102.405 ;
        RECT 121.010 101.860 126.355 102.405 ;
        RECT 115.945 99.855 119.455 100.945 ;
        RECT 119.665 99.855 119.895 100.995 ;
        RECT 120.065 100.025 120.395 101.005 ;
        RECT 120.565 99.855 120.775 100.995 ;
        RECT 122.600 100.290 122.950 101.540 ;
        RECT 124.430 101.030 124.770 101.860 ;
        RECT 126.525 101.655 127.735 102.405 ;
        RECT 126.525 100.945 127.045 101.485 ;
        RECT 127.215 101.115 127.735 101.655 ;
        RECT 121.010 99.855 126.355 100.290 ;
        RECT 126.525 99.855 127.735 100.945 ;
        RECT 14.660 99.685 127.820 99.855 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 14.660 211.050 127.820 211.530 ;
        RECT 14.660 208.330 127.820 208.810 ;
        RECT 73.610 207.790 73.930 207.850 ;
        RECT 75.005 207.790 75.295 207.835 ;
        RECT 73.610 207.650 79.360 207.790 ;
        RECT 73.610 207.590 73.930 207.650 ;
        RECT 75.005 207.605 75.295 207.650 ;
        RECT 66.250 207.110 66.570 207.170 ;
        RECT 72.705 207.110 72.995 207.155 ;
        RECT 66.250 206.970 72.995 207.110 ;
        RECT 66.250 206.910 66.570 206.970 ;
        RECT 72.705 206.925 72.995 206.970 ;
        RECT 73.150 207.110 73.470 207.170 ;
        RECT 79.220 207.155 79.360 207.650 ;
        RECT 79.590 207.250 79.910 207.510 ;
        RECT 74.085 207.110 74.375 207.155 ;
        RECT 73.150 206.970 74.375 207.110 ;
        RECT 73.150 206.910 73.470 206.970 ;
        RECT 74.085 206.925 74.375 206.970 ;
        RECT 79.145 206.925 79.435 207.155 ;
        RECT 73.165 206.430 73.455 206.475 ;
        RECT 74.070 206.430 74.390 206.490 ;
        RECT 73.165 206.290 74.390 206.430 ;
        RECT 73.165 206.245 73.455 206.290 ;
        RECT 74.070 206.230 74.390 206.290 ;
        RECT 75.910 206.430 76.230 206.490 ;
        RECT 77.305 206.430 77.595 206.475 ;
        RECT 75.910 206.290 77.595 206.430 ;
        RECT 75.910 206.230 76.230 206.290 ;
        RECT 77.305 206.245 77.595 206.290 ;
        RECT 14.660 205.610 127.820 206.090 ;
        RECT 74.070 205.410 74.390 205.470 ;
        RECT 74.070 205.270 76.600 205.410 ;
        RECT 74.070 205.210 74.390 205.270 ;
        RECT 67.645 205.070 67.935 205.115 ;
        RECT 70.045 205.070 70.335 205.115 ;
        RECT 73.285 205.070 73.935 205.115 ;
        RECT 67.645 204.930 73.935 205.070 ;
        RECT 67.645 204.885 67.935 204.930 ;
        RECT 70.045 204.885 70.635 204.930 ;
        RECT 73.285 204.885 73.935 204.930 ;
        RECT 65.805 204.730 66.095 204.775 ;
        RECT 66.250 204.730 66.570 204.790 ;
        RECT 67.185 204.730 67.475 204.775 ;
        RECT 65.805 204.590 67.475 204.730 ;
        RECT 65.805 204.545 66.095 204.590 ;
        RECT 66.250 204.530 66.570 204.590 ;
        RECT 67.185 204.545 67.475 204.590 ;
        RECT 70.345 204.570 70.635 204.885 ;
        RECT 75.910 204.870 76.230 205.130 ;
        RECT 76.460 205.070 76.600 205.270 ;
        RECT 79.245 205.070 79.535 205.115 ;
        RECT 82.485 205.070 83.135 205.115 ;
        RECT 76.460 204.930 83.135 205.070 ;
        RECT 79.245 204.885 79.835 204.930 ;
        RECT 82.485 204.885 83.135 204.930 ;
        RECT 83.730 205.070 84.050 205.130 ;
        RECT 85.125 205.070 85.415 205.115 ;
        RECT 83.730 204.930 85.415 205.070 ;
        RECT 71.425 204.730 71.715 204.775 ;
        RECT 75.005 204.730 75.295 204.775 ;
        RECT 76.840 204.730 77.130 204.775 ;
        RECT 71.425 204.590 77.130 204.730 ;
        RECT 71.425 204.545 71.715 204.590 ;
        RECT 75.005 204.545 75.295 204.590 ;
        RECT 76.840 204.545 77.130 204.590 ;
        RECT 79.545 204.570 79.835 204.885 ;
        RECT 83.730 204.870 84.050 204.930 ;
        RECT 85.125 204.885 85.415 204.930 ;
        RECT 80.625 204.730 80.915 204.775 ;
        RECT 84.205 204.730 84.495 204.775 ;
        RECT 86.040 204.730 86.330 204.775 ;
        RECT 80.625 204.590 86.330 204.730 ;
        RECT 80.625 204.545 80.915 204.590 ;
        RECT 84.205 204.545 84.495 204.590 ;
        RECT 86.040 204.545 86.330 204.590 ;
        RECT 63.950 204.390 64.270 204.450 ;
        RECT 77.305 204.390 77.595 204.435 ;
        RECT 63.950 204.250 77.595 204.390 ;
        RECT 63.950 204.190 64.270 204.250 ;
        RECT 77.305 204.205 77.595 204.250 ;
        RECT 86.505 204.390 86.795 204.435 ;
        RECT 88.330 204.390 88.650 204.450 ;
        RECT 86.505 204.250 88.650 204.390 ;
        RECT 86.505 204.205 86.795 204.250 ;
        RECT 88.330 204.190 88.650 204.250 ;
        RECT 71.425 204.050 71.715 204.095 ;
        RECT 74.545 204.050 74.835 204.095 ;
        RECT 76.435 204.050 76.725 204.095 ;
        RECT 71.425 203.910 76.725 204.050 ;
        RECT 71.425 203.865 71.715 203.910 ;
        RECT 74.545 203.865 74.835 203.910 ;
        RECT 76.435 203.865 76.725 203.910 ;
        RECT 80.625 204.050 80.915 204.095 ;
        RECT 83.745 204.050 84.035 204.095 ;
        RECT 85.635 204.050 85.925 204.095 ;
        RECT 80.625 203.910 85.925 204.050 ;
        RECT 80.625 203.865 80.915 203.910 ;
        RECT 83.745 203.865 84.035 203.910 ;
        RECT 85.635 203.865 85.925 203.910 ;
        RECT 64.870 203.710 65.190 203.770 ;
        RECT 65.345 203.710 65.635 203.755 ;
        RECT 64.870 203.570 65.635 203.710 ;
        RECT 64.870 203.510 65.190 203.570 ;
        RECT 65.345 203.525 65.635 203.570 ;
        RECT 68.565 203.710 68.855 203.755 ;
        RECT 73.150 203.710 73.470 203.770 ;
        RECT 68.565 203.570 73.470 203.710 ;
        RECT 68.565 203.525 68.855 203.570 ;
        RECT 73.150 203.510 73.470 203.570 ;
        RECT 74.070 203.710 74.390 203.770 ;
        RECT 77.765 203.710 78.055 203.755 ;
        RECT 74.070 203.570 78.055 203.710 ;
        RECT 74.070 203.510 74.390 203.570 ;
        RECT 77.765 203.525 78.055 203.570 ;
        RECT 14.660 202.890 127.820 203.370 ;
        RECT 63.950 202.690 64.270 202.750 ;
        RECT 60.360 202.550 64.270 202.690 ;
        RECT 59.825 202.010 60.115 202.055 ;
        RECT 60.360 202.010 60.500 202.550 ;
        RECT 63.950 202.490 64.270 202.550 ;
        RECT 66.710 202.690 67.030 202.750 ;
        RECT 70.405 202.690 70.695 202.735 ;
        RECT 66.710 202.550 70.695 202.690 ;
        RECT 66.710 202.490 67.030 202.550 ;
        RECT 70.405 202.505 70.695 202.550 ;
        RECT 77.765 202.505 78.055 202.735 ;
        RECT 60.695 202.350 60.985 202.395 ;
        RECT 62.585 202.350 62.875 202.395 ;
        RECT 65.705 202.350 65.995 202.395 ;
        RECT 76.370 202.350 76.690 202.410 ;
        RECT 77.840 202.350 77.980 202.505 ;
        RECT 60.695 202.210 65.995 202.350 ;
        RECT 60.695 202.165 60.985 202.210 ;
        RECT 62.585 202.165 62.875 202.210 ;
        RECT 65.705 202.165 65.995 202.210 ;
        RECT 70.020 202.210 73.840 202.350 ;
        RECT 59.825 201.870 60.500 202.010 ;
        RECT 59.825 201.825 60.115 201.870 ;
        RECT 61.190 201.810 61.510 202.070 ;
        RECT 70.020 202.055 70.160 202.210 ;
        RECT 69.945 201.825 70.235 202.055 ;
        RECT 72.245 202.010 72.535 202.055 ;
        RECT 73.150 202.010 73.470 202.070 ;
        RECT 73.700 202.055 73.840 202.210 ;
        RECT 76.370 202.210 77.980 202.350 ;
        RECT 82.465 202.350 82.755 202.395 ;
        RECT 85.585 202.350 85.875 202.395 ;
        RECT 87.475 202.350 87.765 202.395 ;
        RECT 82.465 202.210 87.765 202.350 ;
        RECT 76.370 202.150 76.690 202.210 ;
        RECT 82.465 202.165 82.755 202.210 ;
        RECT 85.585 202.165 85.875 202.210 ;
        RECT 87.475 202.165 87.765 202.210 ;
        RECT 72.245 201.870 73.470 202.010 ;
        RECT 72.245 201.825 72.535 201.870 ;
        RECT 73.150 201.810 73.470 201.870 ;
        RECT 73.625 202.010 73.915 202.055 ;
        RECT 74.530 202.010 74.850 202.070 ;
        RECT 73.625 201.870 74.850 202.010 ;
        RECT 73.625 201.825 73.915 201.870 ;
        RECT 74.530 201.810 74.850 201.870 ;
        RECT 79.130 202.010 79.450 202.070 ;
        RECT 79.605 202.010 79.895 202.055 ;
        RECT 79.130 201.870 79.895 202.010 ;
        RECT 79.130 201.810 79.450 201.870 ;
        RECT 79.605 201.825 79.895 201.870 ;
        RECT 84.650 202.010 84.970 202.070 ;
        RECT 86.965 202.010 87.255 202.055 ;
        RECT 84.650 201.870 87.255 202.010 ;
        RECT 84.650 201.810 84.970 201.870 ;
        RECT 86.965 201.825 87.255 201.870 ;
        RECT 60.290 201.670 60.580 201.715 ;
        RECT 62.125 201.670 62.415 201.715 ;
        RECT 65.705 201.670 65.995 201.715 ;
        RECT 60.290 201.530 65.995 201.670 ;
        RECT 60.290 201.485 60.580 201.530 ;
        RECT 62.125 201.485 62.415 201.530 ;
        RECT 65.705 201.485 65.995 201.530 ;
        RECT 63.485 201.330 64.135 201.375 ;
        RECT 64.870 201.330 65.190 201.390 ;
        RECT 66.785 201.375 67.075 201.690 ;
        RECT 71.200 201.670 71.490 201.715 ;
        RECT 74.070 201.670 74.390 201.730 ;
        RECT 71.200 201.530 74.390 201.670 ;
        RECT 71.200 201.485 71.490 201.530 ;
        RECT 74.070 201.470 74.390 201.530 ;
        RECT 66.785 201.330 67.375 201.375 ;
        RECT 63.485 201.190 67.375 201.330 ;
        RECT 63.485 201.145 64.135 201.190 ;
        RECT 64.870 201.130 65.190 201.190 ;
        RECT 67.085 201.145 67.375 201.190 ;
        RECT 74.990 201.130 75.310 201.390 ;
        RECT 75.450 201.330 75.770 201.390 ;
        RECT 77.605 201.330 77.895 201.375 ;
        RECT 75.450 201.190 77.895 201.330 ;
        RECT 75.450 201.130 75.770 201.190 ;
        RECT 77.605 201.145 77.895 201.190 ;
        RECT 78.685 201.330 78.975 201.375 ;
        RECT 79.590 201.330 79.910 201.390 ;
        RECT 81.385 201.375 81.675 201.690 ;
        RECT 82.465 201.670 82.755 201.715 ;
        RECT 86.045 201.670 86.335 201.715 ;
        RECT 87.880 201.670 88.170 201.715 ;
        RECT 82.465 201.530 88.170 201.670 ;
        RECT 82.465 201.485 82.755 201.530 ;
        RECT 86.045 201.485 86.335 201.530 ;
        RECT 87.880 201.485 88.170 201.530 ;
        RECT 88.330 201.670 88.650 201.730 ;
        RECT 96.610 201.670 96.930 201.730 ;
        RECT 88.330 201.530 96.930 201.670 ;
        RECT 88.330 201.470 88.650 201.530 ;
        RECT 96.610 201.470 96.930 201.530 ;
        RECT 78.685 201.190 79.910 201.330 ;
        RECT 78.685 201.145 78.975 201.190 ;
        RECT 79.590 201.130 79.910 201.190 ;
        RECT 81.085 201.330 81.675 201.375 ;
        RECT 84.325 201.330 84.975 201.375 ;
        RECT 85.570 201.330 85.890 201.390 ;
        RECT 81.085 201.190 85.890 201.330 ;
        RECT 81.085 201.145 81.375 201.190 ;
        RECT 84.325 201.145 84.975 201.190 ;
        RECT 85.570 201.130 85.890 201.190 ;
        RECT 71.770 200.790 72.090 201.050 ;
        RECT 72.690 200.990 73.010 201.050 ;
        RECT 74.545 200.990 74.835 201.035 ;
        RECT 72.690 200.850 74.835 200.990 ;
        RECT 72.690 200.790 73.010 200.850 ;
        RECT 74.545 200.805 74.835 200.850 ;
        RECT 75.910 200.990 76.230 201.050 ;
        RECT 76.845 200.990 77.135 201.035 ;
        RECT 75.910 200.850 77.135 200.990 ;
        RECT 75.910 200.790 76.230 200.850 ;
        RECT 76.845 200.805 77.135 200.850 ;
        RECT 14.660 200.170 127.820 200.650 ;
        RECT 61.190 199.970 61.510 200.030 ;
        RECT 67.645 199.970 67.935 200.015 ;
        RECT 72.245 199.970 72.535 200.015 ;
        RECT 74.070 199.970 74.390 200.030 ;
        RECT 61.190 199.830 67.935 199.970 ;
        RECT 61.190 199.770 61.510 199.830 ;
        RECT 67.645 199.785 67.935 199.830 ;
        RECT 71.170 199.830 74.390 199.970 ;
        RECT 69.945 199.630 70.235 199.675 ;
        RECT 71.170 199.630 71.310 199.830 ;
        RECT 72.245 199.785 72.535 199.830 ;
        RECT 74.070 199.770 74.390 199.830 ;
        RECT 74.990 199.970 75.310 200.030 ;
        RECT 75.465 199.970 75.755 200.015 ;
        RECT 74.990 199.830 75.755 199.970 ;
        RECT 74.990 199.770 75.310 199.830 ;
        RECT 75.465 199.785 75.755 199.830 ;
        RECT 76.370 199.970 76.690 200.030 ;
        RECT 79.145 199.970 79.435 200.015 ;
        RECT 76.370 199.830 79.435 199.970 ;
        RECT 76.370 199.770 76.690 199.830 ;
        RECT 79.145 199.785 79.435 199.830 ;
        RECT 79.590 199.970 79.910 200.030 ;
        RECT 81.445 199.970 81.735 200.015 ;
        RECT 79.590 199.830 81.735 199.970 ;
        RECT 79.590 199.770 79.910 199.830 ;
        RECT 81.445 199.785 81.735 199.830 ;
        RECT 83.730 199.770 84.050 200.030 ;
        RECT 84.650 199.770 84.970 200.030 ;
        RECT 85.570 199.970 85.890 200.030 ;
        RECT 86.045 199.970 86.335 200.015 ;
        RECT 85.570 199.830 86.335 199.970 ;
        RECT 85.570 199.770 85.890 199.830 ;
        RECT 86.045 199.785 86.335 199.830 ;
        RECT 69.945 199.490 71.310 199.630 ;
        RECT 69.945 199.445 70.235 199.490 ;
        RECT 74.530 199.430 74.850 199.690 ;
        RECT 80.970 199.630 81.290 199.690 ;
        RECT 97.990 199.630 98.310 199.690 ;
        RECT 98.565 199.630 98.855 199.675 ;
        RECT 101.805 199.630 102.455 199.675 ;
        RECT 80.970 199.490 84.420 199.630 ;
        RECT 80.970 199.430 81.290 199.490 ;
        RECT 68.550 199.090 68.870 199.350 ;
        RECT 71.770 199.290 72.090 199.350 ;
        RECT 78.685 199.290 78.975 199.335 ;
        RECT 79.130 199.290 79.450 199.350 ;
        RECT 71.770 199.150 79.450 199.290 ;
        RECT 71.770 199.090 72.090 199.150 ;
        RECT 78.685 199.105 78.975 199.150 ;
        RECT 79.130 199.090 79.450 199.150 ;
        RECT 80.050 199.290 80.370 199.350 ;
        RECT 82.440 199.335 82.580 199.490 ;
        RECT 84.280 199.335 84.420 199.490 ;
        RECT 97.990 199.490 102.455 199.630 ;
        RECT 97.990 199.430 98.310 199.490 ;
        RECT 98.565 199.445 99.155 199.490 ;
        RECT 101.805 199.445 102.455 199.490 ;
        RECT 81.445 199.290 81.735 199.335 ;
        RECT 80.050 199.150 81.735 199.290 ;
        RECT 80.050 199.090 80.370 199.150 ;
        RECT 81.445 199.105 81.735 199.150 ;
        RECT 82.365 199.105 82.655 199.335 ;
        RECT 82.825 199.105 83.115 199.335 ;
        RECT 84.205 199.105 84.495 199.335 ;
        RECT 86.505 199.290 86.795 199.335 ;
        RECT 86.950 199.290 87.270 199.350 ;
        RECT 86.505 199.150 87.270 199.290 ;
        RECT 86.505 199.105 86.795 199.150 ;
        RECT 75.910 198.950 76.230 199.010 ;
        RECT 82.900 198.950 83.040 199.105 ;
        RECT 86.950 199.090 87.270 199.150 ;
        RECT 98.865 199.130 99.155 199.445 ;
        RECT 99.945 199.290 100.235 199.335 ;
        RECT 103.525 199.290 103.815 199.335 ;
        RECT 105.360 199.290 105.650 199.335 ;
        RECT 99.945 199.150 105.650 199.290 ;
        RECT 99.945 199.105 100.235 199.150 ;
        RECT 103.525 199.105 103.815 199.150 ;
        RECT 105.360 199.105 105.650 199.150 ;
        RECT 75.910 198.810 83.040 198.950 ;
        RECT 75.910 198.750 76.230 198.810 ;
        RECT 104.430 198.750 104.750 199.010 ;
        RECT 105.810 198.750 106.130 199.010 ;
        RECT 69.025 198.610 69.315 198.655 ;
        RECT 73.150 198.610 73.470 198.670 ;
        RECT 69.025 198.470 73.470 198.610 ;
        RECT 69.025 198.425 69.315 198.470 ;
        RECT 73.150 198.410 73.470 198.470 ;
        RECT 73.610 198.610 73.930 198.670 ;
        RECT 74.545 198.610 74.835 198.655 ;
        RECT 73.610 198.470 74.835 198.610 ;
        RECT 73.610 198.410 73.930 198.470 ;
        RECT 74.545 198.425 74.835 198.470 ;
        RECT 99.945 198.610 100.235 198.655 ;
        RECT 103.065 198.610 103.355 198.655 ;
        RECT 104.955 198.610 105.245 198.655 ;
        RECT 99.945 198.470 105.245 198.610 ;
        RECT 99.945 198.425 100.235 198.470 ;
        RECT 103.065 198.425 103.355 198.470 ;
        RECT 104.955 198.425 105.245 198.470 ;
        RECT 64.870 198.270 65.190 198.330 ;
        RECT 70.865 198.270 71.155 198.315 ;
        RECT 64.870 198.130 71.155 198.270 ;
        RECT 64.870 198.070 65.190 198.130 ;
        RECT 70.865 198.085 71.155 198.130 ;
        RECT 72.690 198.270 73.010 198.330 ;
        RECT 80.970 198.270 81.290 198.330 ;
        RECT 72.690 198.130 81.290 198.270 ;
        RECT 72.690 198.070 73.010 198.130 ;
        RECT 80.970 198.070 81.290 198.130 ;
        RECT 97.085 198.270 97.375 198.315 ;
        RECT 98.450 198.270 98.770 198.330 ;
        RECT 97.085 198.130 98.770 198.270 ;
        RECT 97.085 198.085 97.375 198.130 ;
        RECT 98.450 198.070 98.770 198.130 ;
        RECT 14.660 197.450 127.820 197.930 ;
        RECT 68.550 197.250 68.870 197.310 ;
        RECT 69.025 197.250 69.315 197.295 ;
        RECT 68.550 197.110 69.315 197.250 ;
        RECT 68.550 197.050 68.870 197.110 ;
        RECT 69.025 197.065 69.315 197.110 ;
        RECT 69.930 197.050 70.250 197.310 ;
        RECT 73.610 197.250 73.930 197.310 ;
        RECT 72.320 197.110 73.930 197.250 ;
        RECT 50.610 196.570 50.930 196.630 ;
        RECT 54.305 196.570 54.595 196.615 ;
        RECT 50.610 196.430 54.595 196.570 ;
        RECT 50.610 196.370 50.930 196.430 ;
        RECT 54.305 196.385 54.595 196.430 ;
        RECT 70.390 196.570 70.710 196.630 ;
        RECT 72.320 196.615 72.460 197.110 ;
        RECT 73.610 197.050 73.930 197.110 ;
        RECT 80.050 196.910 80.370 196.970 ;
        RECT 73.700 196.770 80.370 196.910 ;
        RECT 72.245 196.570 72.535 196.615 ;
        RECT 70.390 196.430 72.535 196.570 ;
        RECT 70.390 196.370 70.710 196.430 ;
        RECT 72.245 196.385 72.535 196.430 ;
        RECT 72.690 196.370 73.010 196.630 ;
        RECT 73.150 196.570 73.470 196.630 ;
        RECT 73.700 196.570 73.840 196.770 ;
        RECT 80.050 196.710 80.370 196.770 ;
        RECT 89.680 196.910 89.970 196.955 ;
        RECT 92.460 196.910 92.750 196.955 ;
        RECT 94.320 196.910 94.610 196.955 ;
        RECT 89.680 196.770 94.610 196.910 ;
        RECT 89.680 196.725 89.970 196.770 ;
        RECT 92.460 196.725 92.750 196.770 ;
        RECT 94.320 196.725 94.610 196.770 ;
        RECT 113.285 196.910 113.575 196.955 ;
        RECT 116.405 196.910 116.695 196.955 ;
        RECT 118.295 196.910 118.585 196.955 ;
        RECT 113.285 196.770 118.585 196.910 ;
        RECT 113.285 196.725 113.575 196.770 ;
        RECT 116.405 196.725 116.695 196.770 ;
        RECT 118.295 196.725 118.585 196.770 ;
        RECT 73.150 196.430 73.840 196.570 ;
        RECT 92.945 196.570 93.235 196.615 ;
        RECT 93.850 196.570 94.170 196.630 ;
        RECT 92.945 196.430 94.170 196.570 ;
        RECT 73.150 196.370 73.470 196.430 ;
        RECT 92.945 196.385 93.235 196.430 ;
        RECT 93.850 196.370 94.170 196.430 ;
        RECT 49.230 196.230 49.550 196.290 ;
        RECT 53.845 196.230 54.135 196.275 ;
        RECT 49.230 196.090 54.135 196.230 ;
        RECT 49.230 196.030 49.550 196.090 ;
        RECT 53.845 196.045 54.135 196.090 ;
        RECT 69.010 196.230 69.330 196.290 ;
        RECT 73.625 196.230 73.915 196.275 ;
        RECT 74.530 196.230 74.850 196.290 ;
        RECT 69.010 196.090 74.850 196.230 ;
        RECT 69.010 196.030 69.330 196.090 ;
        RECT 73.625 196.045 73.915 196.090 ;
        RECT 74.530 196.030 74.850 196.090 ;
        RECT 89.680 196.230 89.970 196.275 ;
        RECT 94.785 196.230 95.075 196.275 ;
        RECT 96.610 196.230 96.930 196.290 ;
        RECT 89.680 196.090 92.215 196.230 ;
        RECT 89.680 196.045 89.970 196.090 ;
        RECT 70.865 195.890 71.155 195.935 ;
        RECT 71.770 195.890 72.090 195.950 ;
        RECT 75.450 195.890 75.770 195.950 ;
        RECT 70.865 195.750 75.770 195.890 ;
        RECT 70.865 195.705 71.155 195.750 ;
        RECT 71.770 195.690 72.090 195.750 ;
        RECT 75.450 195.690 75.770 195.750 ;
        RECT 87.820 195.890 88.110 195.935 ;
        RECT 90.170 195.890 90.490 195.950 ;
        RECT 92.000 195.935 92.215 196.090 ;
        RECT 94.785 196.090 96.930 196.230 ;
        RECT 94.785 196.045 95.075 196.090 ;
        RECT 96.610 196.030 96.930 196.090 ;
        RECT 98.450 196.030 98.770 196.290 ;
        RECT 112.205 195.935 112.495 196.250 ;
        RECT 113.285 196.230 113.575 196.275 ;
        RECT 116.865 196.230 117.155 196.275 ;
        RECT 118.700 196.230 118.990 196.275 ;
        RECT 113.285 196.090 118.990 196.230 ;
        RECT 113.285 196.045 113.575 196.090 ;
        RECT 116.865 196.045 117.155 196.090 ;
        RECT 118.700 196.045 118.990 196.090 ;
        RECT 119.165 196.045 119.455 196.275 ;
        RECT 115.470 195.935 115.790 195.950 ;
        RECT 91.080 195.890 91.370 195.935 ;
        RECT 87.820 195.750 91.370 195.890 ;
        RECT 87.820 195.705 88.110 195.750 ;
        RECT 90.170 195.690 90.490 195.750 ;
        RECT 91.080 195.705 91.370 195.750 ;
        RECT 92.000 195.890 92.290 195.935 ;
        RECT 93.860 195.890 94.150 195.935 ;
        RECT 92.000 195.750 94.150 195.890 ;
        RECT 92.000 195.705 92.290 195.750 ;
        RECT 93.860 195.705 94.150 195.750 ;
        RECT 111.905 195.890 112.495 195.935 ;
        RECT 115.145 195.890 115.795 195.935 ;
        RECT 111.905 195.750 115.795 195.890 ;
        RECT 111.905 195.705 112.195 195.750 ;
        RECT 115.145 195.705 115.795 195.750 ;
        RECT 115.470 195.690 115.790 195.705 ;
        RECT 117.770 195.690 118.090 195.950 ;
        RECT 118.230 195.890 118.550 195.950 ;
        RECT 119.240 195.890 119.380 196.045 ;
        RECT 118.230 195.750 119.380 195.890 ;
        RECT 118.230 195.690 118.550 195.750 ;
        RECT 53.370 195.350 53.690 195.610 ;
        RECT 57.525 195.550 57.815 195.595 ;
        RECT 57.970 195.550 58.290 195.610 ;
        RECT 85.570 195.595 85.890 195.610 ;
        RECT 57.525 195.410 58.290 195.550 ;
        RECT 57.525 195.365 57.815 195.410 ;
        RECT 57.970 195.350 58.290 195.410 ;
        RECT 69.865 195.550 70.155 195.595 ;
        RECT 71.325 195.550 71.615 195.595 ;
        RECT 69.865 195.410 71.615 195.550 ;
        RECT 69.865 195.365 70.155 195.410 ;
        RECT 71.325 195.365 71.615 195.410 ;
        RECT 85.570 195.365 86.105 195.595 ;
        RECT 85.570 195.350 85.890 195.365 ;
        RECT 101.210 195.350 101.530 195.610 ;
        RECT 109.030 195.550 109.350 195.610 ;
        RECT 110.425 195.550 110.715 195.595 ;
        RECT 109.030 195.410 110.715 195.550 ;
        RECT 109.030 195.350 109.350 195.410 ;
        RECT 110.425 195.365 110.715 195.410 ;
        RECT 14.660 194.730 127.820 195.210 ;
        RECT 50.610 194.530 50.930 194.590 ;
        RECT 57.985 194.530 58.275 194.575 ;
        RECT 50.610 194.390 58.275 194.530 ;
        RECT 50.610 194.330 50.930 194.390 ;
        RECT 57.985 194.345 58.275 194.390 ;
        RECT 71.770 194.330 72.090 194.590 ;
        RECT 85.570 194.530 85.890 194.590 ;
        RECT 86.045 194.530 86.335 194.575 ;
        RECT 72.320 194.390 85.340 194.530 ;
        RECT 49.230 194.190 49.550 194.250 ;
        RECT 53.370 194.235 53.690 194.250 ;
        RECT 48.860 194.050 49.550 194.190 ;
        RECT 46.010 193.850 46.330 193.910 ;
        RECT 48.860 193.895 49.000 194.050 ;
        RECT 49.230 193.990 49.550 194.050 ;
        RECT 52.905 194.190 53.690 194.235 ;
        RECT 56.505 194.190 56.795 194.235 ;
        RECT 72.320 194.190 72.460 194.390 ;
        RECT 52.905 194.050 56.795 194.190 ;
        RECT 52.905 194.005 53.690 194.050 ;
        RECT 53.370 193.990 53.690 194.005 ;
        RECT 56.205 194.005 56.795 194.050 ;
        RECT 66.340 194.050 72.460 194.190 ;
        RECT 72.690 194.190 73.010 194.250 ;
        RECT 85.200 194.190 85.340 194.390 ;
        RECT 85.570 194.390 86.335 194.530 ;
        RECT 85.570 194.330 85.890 194.390 ;
        RECT 86.045 194.345 86.335 194.390 ;
        RECT 89.725 194.530 90.015 194.575 ;
        RECT 90.170 194.530 90.490 194.590 ;
        RECT 89.725 194.390 90.490 194.530 ;
        RECT 89.725 194.345 90.015 194.390 ;
        RECT 90.170 194.330 90.490 194.390 ;
        RECT 93.865 194.530 94.155 194.575 ;
        RECT 97.990 194.530 98.310 194.590 ;
        RECT 93.865 194.390 98.310 194.530 ;
        RECT 93.865 194.345 94.155 194.390 ;
        RECT 97.990 194.330 98.310 194.390 ;
        RECT 112.265 194.530 112.555 194.575 ;
        RECT 112.710 194.530 113.030 194.590 ;
        RECT 112.265 194.390 113.030 194.530 ;
        RECT 112.265 194.345 112.555 194.390 ;
        RECT 112.710 194.330 113.030 194.390 ;
        RECT 115.470 194.330 115.790 194.590 ;
        RECT 86.950 194.190 87.270 194.250 ;
        RECT 96.610 194.190 96.930 194.250 ;
        RECT 103.525 194.190 103.815 194.235 ;
        RECT 105.810 194.190 106.130 194.250 ;
        RECT 118.230 194.190 118.550 194.250 ;
        RECT 72.690 194.050 75.220 194.190 ;
        RECT 85.200 194.050 95.460 194.190 ;
        RECT 48.785 193.850 49.075 193.895 ;
        RECT 46.010 193.710 49.075 193.850 ;
        RECT 46.010 193.650 46.330 193.710 ;
        RECT 48.785 193.665 49.075 193.710 ;
        RECT 49.710 193.850 50.000 193.895 ;
        RECT 51.545 193.850 51.835 193.895 ;
        RECT 55.125 193.850 55.415 193.895 ;
        RECT 49.710 193.710 55.415 193.850 ;
        RECT 49.710 193.665 50.000 193.710 ;
        RECT 51.545 193.665 51.835 193.710 ;
        RECT 55.125 193.665 55.415 193.710 ;
        RECT 56.205 193.690 56.495 194.005 ;
        RECT 66.340 193.910 66.480 194.050 ;
        RECT 72.690 193.990 73.010 194.050 ;
        RECT 66.250 193.650 66.570 193.910 ;
        RECT 69.010 193.650 69.330 193.910 ;
        RECT 73.150 193.650 73.470 193.910 ;
        RECT 75.080 193.895 75.220 194.050 ;
        RECT 86.950 193.990 87.270 194.050 ;
        RECT 75.005 193.850 75.295 193.895 ;
        RECT 76.370 193.850 76.690 193.910 ;
        RECT 75.005 193.710 76.690 193.850 ;
        RECT 75.005 193.665 75.295 193.710 ;
        RECT 76.370 193.650 76.690 193.710 ;
        RECT 86.030 193.850 86.350 193.910 ;
        RECT 86.505 193.850 86.795 193.895 ;
        RECT 86.030 193.710 86.795 193.850 ;
        RECT 86.030 193.650 86.350 193.710 ;
        RECT 86.505 193.665 86.795 193.710 ;
        RECT 90.170 193.650 90.490 193.910 ;
        RECT 93.480 193.895 93.620 194.050 ;
        RECT 93.405 193.665 93.695 193.895 ;
        RECT 94.770 193.650 95.090 193.910 ;
        RECT 95.320 193.850 95.460 194.050 ;
        RECT 96.610 194.050 118.550 194.190 ;
        RECT 96.610 193.990 96.930 194.050 ;
        RECT 103.525 194.005 103.815 194.050 ;
        RECT 105.810 193.990 106.130 194.050 ;
        RECT 118.230 193.990 118.550 194.050 ;
        RECT 109.045 193.850 109.335 193.895 ;
        RECT 115.930 193.850 116.250 193.910 ;
        RECT 95.320 193.710 116.250 193.850 ;
        RECT 109.045 193.665 109.335 193.710 ;
        RECT 115.930 193.650 116.250 193.710 ;
        RECT 49.230 193.310 49.550 193.570 ;
        RECT 50.610 193.310 50.930 193.570 ;
        RECT 70.405 193.510 70.695 193.555 ;
        RECT 70.405 193.370 72.460 193.510 ;
        RECT 70.405 193.325 70.695 193.370 ;
        RECT 72.320 193.215 72.460 193.370 ;
        RECT 85.110 193.310 85.430 193.570 ;
        RECT 108.110 193.510 108.430 193.570 ;
        RECT 110.870 193.510 111.190 193.570 ;
        RECT 108.110 193.370 111.190 193.510 ;
        RECT 108.110 193.310 108.430 193.370 ;
        RECT 110.870 193.310 111.190 193.370 ;
        RECT 111.805 193.325 112.095 193.555 ;
        RECT 50.115 193.170 50.405 193.215 ;
        RECT 52.005 193.170 52.295 193.215 ;
        RECT 55.125 193.170 55.415 193.215 ;
        RECT 50.115 193.030 55.415 193.170 ;
        RECT 50.115 192.985 50.405 193.030 ;
        RECT 52.005 192.985 52.295 193.030 ;
        RECT 55.125 192.985 55.415 193.030 ;
        RECT 72.245 192.985 72.535 193.215 ;
        RECT 111.880 193.170 112.020 193.325 ;
        RECT 112.250 193.170 112.570 193.230 ;
        RECT 111.880 193.030 112.570 193.170 ;
        RECT 112.250 192.970 112.570 193.030 ;
        RECT 48.325 192.830 48.615 192.875 ;
        RECT 54.290 192.830 54.610 192.890 ;
        RECT 48.325 192.690 54.610 192.830 ;
        RECT 48.325 192.645 48.615 192.690 ;
        RECT 54.290 192.630 54.610 192.690 ;
        RECT 65.790 192.630 66.110 192.890 ;
        RECT 70.390 192.630 70.710 192.890 ;
        RECT 72.690 192.830 73.010 192.890 ;
        RECT 73.165 192.830 73.455 192.875 ;
        RECT 72.690 192.690 73.455 192.830 ;
        RECT 72.690 192.630 73.010 192.690 ;
        RECT 73.165 192.645 73.455 192.690 ;
        RECT 88.345 192.830 88.635 192.875 ;
        RECT 91.090 192.830 91.410 192.890 ;
        RECT 88.345 192.690 91.410 192.830 ;
        RECT 88.345 192.645 88.635 192.690 ;
        RECT 91.090 192.630 91.410 192.690 ;
        RECT 109.490 192.630 109.810 192.890 ;
        RECT 114.105 192.830 114.395 192.875 ;
        RECT 119.150 192.830 119.470 192.890 ;
        RECT 114.105 192.690 119.470 192.830 ;
        RECT 114.105 192.645 114.395 192.690 ;
        RECT 119.150 192.630 119.470 192.690 ;
        RECT 14.660 192.010 127.820 192.490 ;
        RECT 50.610 191.810 50.930 191.870 ;
        RECT 51.085 191.810 51.375 191.855 ;
        RECT 50.610 191.670 51.375 191.810 ;
        RECT 50.610 191.610 50.930 191.670 ;
        RECT 51.085 191.625 51.375 191.670 ;
        RECT 85.570 191.810 85.890 191.870 ;
        RECT 85.570 191.670 93.620 191.810 ;
        RECT 85.570 191.610 85.890 191.670 ;
        RECT 40.460 191.470 40.750 191.515 ;
        RECT 43.240 191.470 43.530 191.515 ;
        RECT 45.100 191.470 45.390 191.515 ;
        RECT 40.460 191.330 45.390 191.470 ;
        RECT 40.460 191.285 40.750 191.330 ;
        RECT 43.240 191.285 43.530 191.330 ;
        RECT 45.100 191.285 45.390 191.330 ;
        RECT 49.705 191.285 49.995 191.515 ;
        RECT 55.325 191.470 55.615 191.515 ;
        RECT 58.445 191.470 58.735 191.515 ;
        RECT 60.335 191.470 60.625 191.515 ;
        RECT 55.325 191.330 60.625 191.470 ;
        RECT 55.325 191.285 55.615 191.330 ;
        RECT 58.445 191.285 58.735 191.330 ;
        RECT 60.335 191.285 60.625 191.330 ;
        RECT 36.595 191.130 36.885 191.175 ;
        RECT 41.410 191.130 41.730 191.190 ;
        RECT 36.595 190.990 46.240 191.130 ;
        RECT 36.595 190.945 36.885 190.990 ;
        RECT 41.410 190.930 41.730 190.990 ;
        RECT 40.460 190.790 40.750 190.835 ;
        RECT 43.725 190.790 44.015 190.835 ;
        RECT 45.090 190.790 45.410 190.850 ;
        RECT 40.460 190.650 42.995 190.790 ;
        RECT 40.460 190.605 40.750 190.650 ;
        RECT 38.600 190.450 38.890 190.495 ;
        RECT 39.110 190.450 39.430 190.510 ;
        RECT 42.780 190.495 42.995 190.650 ;
        RECT 43.725 190.650 45.410 190.790 ;
        RECT 43.725 190.605 44.015 190.650 ;
        RECT 45.090 190.590 45.410 190.650 ;
        RECT 45.565 190.605 45.855 190.835 ;
        RECT 46.100 190.790 46.240 190.990 ;
        RECT 46.470 190.930 46.790 191.190 ;
        RECT 47.865 190.790 48.155 190.835 ;
        RECT 46.100 190.650 48.155 190.790 ;
        RECT 49.780 190.790 49.920 191.285 ;
        RECT 63.950 191.270 64.270 191.530 ;
        RECT 64.985 191.470 65.275 191.515 ;
        RECT 68.105 191.470 68.395 191.515 ;
        RECT 69.995 191.470 70.285 191.515 ;
        RECT 76.845 191.470 77.135 191.515 ;
        RECT 64.985 191.330 70.285 191.470 ;
        RECT 64.985 191.285 65.275 191.330 ;
        RECT 68.105 191.285 68.395 191.330 ;
        RECT 69.995 191.285 70.285 191.330 ;
        RECT 73.700 191.330 77.135 191.470 ;
        RECT 52.450 190.930 52.770 191.190 ;
        RECT 59.350 191.130 59.670 191.190 ;
        RECT 61.205 191.130 61.495 191.175 ;
        RECT 64.040 191.130 64.180 191.270 ;
        RECT 70.865 191.130 71.155 191.175 ;
        RECT 59.350 190.990 71.155 191.130 ;
        RECT 59.350 190.930 59.670 190.990 ;
        RECT 61.205 190.945 61.495 190.990 ;
        RECT 70.865 190.945 71.155 190.990 ;
        RECT 71.310 191.130 71.630 191.190 ;
        RECT 73.700 191.175 73.840 191.330 ;
        RECT 76.845 191.285 77.135 191.330 ;
        RECT 87.380 191.470 87.670 191.515 ;
        RECT 90.160 191.470 90.450 191.515 ;
        RECT 92.020 191.470 92.310 191.515 ;
        RECT 87.380 191.330 92.310 191.470 ;
        RECT 93.480 191.470 93.620 191.670 ;
        RECT 93.850 191.610 94.170 191.870 ;
        RECT 103.065 191.810 103.355 191.855 ;
        RECT 104.430 191.810 104.750 191.870 ;
        RECT 112.710 191.810 113.030 191.870 ;
        RECT 103.065 191.670 104.750 191.810 ;
        RECT 103.065 191.625 103.355 191.670 ;
        RECT 104.430 191.610 104.750 191.670 ;
        RECT 108.660 191.670 113.030 191.810 ;
        RECT 108.110 191.470 108.430 191.530 ;
        RECT 93.480 191.330 97.300 191.470 ;
        RECT 87.380 191.285 87.670 191.330 ;
        RECT 90.160 191.285 90.450 191.330 ;
        RECT 92.020 191.285 92.310 191.330 ;
        RECT 73.625 191.130 73.915 191.175 ;
        RECT 71.310 190.990 73.915 191.130 ;
        RECT 71.310 190.930 71.630 190.990 ;
        RECT 73.625 190.945 73.915 190.990 ;
        RECT 78.225 191.130 78.515 191.175 ;
        RECT 80.050 191.130 80.370 191.190 ;
        RECT 78.225 190.990 80.370 191.130 ;
        RECT 78.225 190.945 78.515 190.990 ;
        RECT 80.050 190.930 80.370 190.990 ;
        RECT 92.485 191.130 92.775 191.175 ;
        RECT 93.850 191.130 94.170 191.190 ;
        RECT 92.485 190.990 96.840 191.130 ;
        RECT 92.485 190.945 92.775 190.990 ;
        RECT 93.850 190.930 94.170 190.990 ;
        RECT 96.700 190.850 96.840 190.990 ;
        RECT 52.005 190.790 52.295 190.835 ;
        RECT 54.290 190.810 54.610 190.850 ;
        RECT 49.780 190.650 52.295 190.790 ;
        RECT 47.865 190.605 48.155 190.650 ;
        RECT 52.005 190.605 52.295 190.650 ;
        RECT 41.860 190.450 42.150 190.495 ;
        RECT 38.600 190.310 42.150 190.450 ;
        RECT 38.600 190.265 38.890 190.310 ;
        RECT 39.110 190.250 39.430 190.310 ;
        RECT 41.860 190.265 42.150 190.310 ;
        RECT 42.780 190.450 43.070 190.495 ;
        RECT 44.640 190.450 44.930 190.495 ;
        RECT 42.780 190.310 44.930 190.450 ;
        RECT 45.640 190.450 45.780 190.605 ;
        RECT 54.245 190.590 54.610 190.810 ;
        RECT 55.325 190.790 55.615 190.835 ;
        RECT 58.905 190.790 59.195 190.835 ;
        RECT 60.740 190.790 61.030 190.835 ;
        RECT 55.325 190.650 61.030 190.790 ;
        RECT 55.325 190.605 55.615 190.650 ;
        RECT 58.905 190.605 59.195 190.650 ;
        RECT 60.740 190.605 61.030 190.650 ;
        RECT 49.230 190.450 49.550 190.510 ;
        RECT 54.245 190.495 54.535 190.590 ;
        RECT 45.640 190.310 49.550 190.450 ;
        RECT 42.780 190.265 43.070 190.310 ;
        RECT 44.640 190.265 44.930 190.310 ;
        RECT 49.230 190.250 49.550 190.310 ;
        RECT 53.945 190.450 54.535 190.495 ;
        RECT 57.185 190.450 57.835 190.495 ;
        RECT 53.945 190.310 57.835 190.450 ;
        RECT 53.945 190.265 54.235 190.310 ;
        RECT 57.185 190.265 57.835 190.310 ;
        RECT 59.825 190.450 60.115 190.495 ;
        RECT 60.270 190.450 60.590 190.510 ;
        RECT 63.905 190.495 64.195 190.810 ;
        RECT 64.985 190.790 65.275 190.835 ;
        RECT 68.565 190.790 68.855 190.835 ;
        RECT 70.400 190.790 70.690 190.835 ;
        RECT 64.985 190.650 70.690 190.790 ;
        RECT 64.985 190.605 65.275 190.650 ;
        RECT 68.565 190.605 68.855 190.650 ;
        RECT 70.400 190.605 70.690 190.650 ;
        RECT 73.150 190.590 73.470 190.850 ;
        RECT 74.530 190.790 74.850 190.850 ;
        RECT 76.385 190.790 76.675 190.835 ;
        RECT 74.530 190.650 76.675 190.790 ;
        RECT 74.530 190.590 74.850 190.650 ;
        RECT 76.385 190.605 76.675 190.650 ;
        RECT 87.380 190.790 87.670 190.835 ;
        RECT 87.380 190.650 89.915 190.790 ;
        RECT 87.380 190.605 87.670 190.650 ;
        RECT 59.825 190.310 60.590 190.450 ;
        RECT 59.825 190.265 60.115 190.310 ;
        RECT 60.270 190.250 60.590 190.310 ;
        RECT 63.605 190.450 64.195 190.495 ;
        RECT 65.790 190.450 66.110 190.510 ;
        RECT 66.845 190.450 67.495 190.495 ;
        RECT 63.605 190.310 67.495 190.450 ;
        RECT 63.605 190.265 63.895 190.310 ;
        RECT 65.790 190.250 66.110 190.310 ;
        RECT 66.845 190.265 67.495 190.310 ;
        RECT 69.485 190.450 69.775 190.495 ;
        RECT 73.610 190.450 73.930 190.510 ;
        RECT 76.845 190.450 77.135 190.495 ;
        RECT 69.485 190.310 71.540 190.450 ;
        RECT 69.485 190.265 69.775 190.310 ;
        RECT 47.405 190.110 47.695 190.155 ;
        RECT 57.970 190.110 58.290 190.170 ;
        RECT 47.405 189.970 58.290 190.110 ;
        RECT 47.405 189.925 47.695 189.970 ;
        RECT 57.970 189.910 58.290 189.970 ;
        RECT 62.110 189.910 62.430 190.170 ;
        RECT 66.250 190.110 66.570 190.170 ;
        RECT 69.930 190.110 70.250 190.170 ;
        RECT 71.400 190.155 71.540 190.310 ;
        RECT 73.610 190.310 77.135 190.450 ;
        RECT 73.610 190.250 73.930 190.310 ;
        RECT 76.845 190.265 77.135 190.310 ;
        RECT 85.520 190.450 85.810 190.495 ;
        RECT 87.870 190.450 88.190 190.510 ;
        RECT 89.700 190.495 89.915 190.650 ;
        RECT 90.630 190.590 90.950 190.850 ;
        RECT 91.090 190.790 91.410 190.850 ;
        RECT 92.945 190.790 93.235 190.835 ;
        RECT 91.090 190.650 93.235 190.790 ;
        RECT 91.090 190.590 91.410 190.650 ;
        RECT 92.945 190.605 93.235 190.650 ;
        RECT 96.610 190.590 96.930 190.850 ;
        RECT 97.160 190.790 97.300 191.330 ;
        RECT 98.080 191.330 108.430 191.470 ;
        RECT 98.080 191.190 98.220 191.330 ;
        RECT 97.990 190.930 98.310 191.190 ;
        RECT 98.925 191.130 99.215 191.175 ;
        RECT 101.210 191.130 101.530 191.190 ;
        RECT 105.440 191.175 105.580 191.330 ;
        RECT 108.110 191.270 108.430 191.330 ;
        RECT 98.925 190.990 102.820 191.130 ;
        RECT 98.925 190.945 99.215 190.990 ;
        RECT 101.210 190.930 101.530 190.990 ;
        RECT 99.385 190.790 99.675 190.835 ;
        RECT 102.145 190.790 102.435 190.835 ;
        RECT 97.160 190.650 99.675 190.790 ;
        RECT 99.385 190.605 99.675 190.650 ;
        RECT 101.300 190.650 102.435 190.790 ;
        RECT 102.680 190.790 102.820 190.990 ;
        RECT 105.365 190.945 105.655 191.175 ;
        RECT 106.270 191.130 106.590 191.190 ;
        RECT 108.660 191.130 108.800 191.670 ;
        RECT 112.710 191.610 113.030 191.670 ;
        RECT 117.770 191.810 118.090 191.870 ;
        RECT 118.245 191.810 118.535 191.855 ;
        RECT 117.770 191.670 118.535 191.810 ;
        RECT 117.770 191.610 118.090 191.670 ;
        RECT 118.245 191.625 118.535 191.670 ;
        RECT 111.905 191.470 112.195 191.515 ;
        RECT 115.025 191.470 115.315 191.515 ;
        RECT 116.915 191.470 117.205 191.515 ;
        RECT 111.905 191.330 117.205 191.470 ;
        RECT 111.905 191.285 112.195 191.330 ;
        RECT 115.025 191.285 115.315 191.330 ;
        RECT 116.915 191.285 117.205 191.330 ;
        RECT 106.270 190.990 108.800 191.130 ;
        RECT 109.045 191.130 109.335 191.175 ;
        RECT 109.950 191.130 110.270 191.190 ;
        RECT 109.045 190.990 110.270 191.130 ;
        RECT 106.270 190.930 106.590 190.990 ;
        RECT 109.045 190.945 109.335 190.990 ;
        RECT 109.950 190.930 110.270 190.990 ;
        RECT 106.745 190.790 107.035 190.835 ;
        RECT 102.680 190.650 107.035 190.790 ;
        RECT 88.780 190.450 89.070 190.495 ;
        RECT 85.520 190.310 89.070 190.450 ;
        RECT 85.520 190.265 85.810 190.310 ;
        RECT 87.870 190.250 88.190 190.310 ;
        RECT 88.780 190.265 89.070 190.310 ;
        RECT 89.700 190.450 89.990 190.495 ;
        RECT 91.560 190.450 91.850 190.495 ;
        RECT 89.700 190.310 91.850 190.450 ;
        RECT 89.700 190.265 89.990 190.310 ;
        RECT 91.560 190.265 91.850 190.310 ;
        RECT 66.250 189.970 70.250 190.110 ;
        RECT 66.250 189.910 66.570 189.970 ;
        RECT 69.930 189.910 70.250 189.970 ;
        RECT 71.325 189.925 71.615 190.155 ;
        RECT 76.370 190.110 76.690 190.170 ;
        RECT 77.305 190.110 77.595 190.155 ;
        RECT 76.370 189.970 77.595 190.110 ;
        RECT 76.370 189.910 76.690 189.970 ;
        RECT 77.305 189.925 77.595 189.970 ;
        RECT 83.515 190.110 83.805 190.155 ;
        RECT 86.030 190.110 86.350 190.170 ;
        RECT 101.300 190.155 101.440 190.650 ;
        RECT 102.145 190.605 102.435 190.650 ;
        RECT 106.745 190.605 107.035 190.650 ;
        RECT 109.490 190.450 109.810 190.510 ;
        RECT 110.825 190.495 111.115 190.810 ;
        RECT 111.905 190.790 112.195 190.835 ;
        RECT 115.485 190.790 115.775 190.835 ;
        RECT 117.320 190.790 117.610 190.835 ;
        RECT 111.905 190.650 117.610 190.790 ;
        RECT 111.905 190.605 112.195 190.650 ;
        RECT 115.485 190.605 115.775 190.650 ;
        RECT 117.320 190.605 117.610 190.650 ;
        RECT 117.785 190.790 118.075 190.835 ;
        RECT 118.230 190.790 118.550 190.850 ;
        RECT 117.785 190.650 118.550 190.790 ;
        RECT 117.785 190.605 118.075 190.650 ;
        RECT 118.230 190.590 118.550 190.650 ;
        RECT 119.150 190.590 119.470 190.850 ;
        RECT 110.525 190.450 111.115 190.495 ;
        RECT 113.765 190.450 114.415 190.495 ;
        RECT 109.490 190.310 114.415 190.450 ;
        RECT 109.490 190.250 109.810 190.310 ;
        RECT 110.525 190.265 110.815 190.310 ;
        RECT 113.765 190.265 114.415 190.310 ;
        RECT 116.390 190.250 116.710 190.510 ;
        RECT 83.515 189.970 86.350 190.110 ;
        RECT 83.515 189.925 83.805 189.970 ;
        RECT 86.030 189.910 86.350 189.970 ;
        RECT 101.225 189.925 101.515 190.155 ;
        RECT 108.585 190.110 108.875 190.155 ;
        RECT 113.170 190.110 113.490 190.170 ;
        RECT 108.585 189.970 113.490 190.110 ;
        RECT 108.585 189.925 108.875 189.970 ;
        RECT 113.170 189.910 113.490 189.970 ;
        RECT 14.660 189.290 127.820 189.770 ;
        RECT 57.970 188.890 58.290 189.150 ;
        RECT 59.825 188.905 60.115 189.135 ;
        RECT 36.365 188.750 36.655 188.795 ;
        RECT 39.225 188.750 39.515 188.795 ;
        RECT 42.465 188.750 43.115 188.795 ;
        RECT 36.365 188.610 43.115 188.750 ;
        RECT 36.365 188.565 36.655 188.610 ;
        RECT 39.225 188.565 39.815 188.610 ;
        RECT 42.465 188.565 43.115 188.610 ;
        RECT 30.385 188.410 30.675 188.455 ;
        RECT 35.905 188.410 36.195 188.455 ;
        RECT 30.385 188.270 36.580 188.410 ;
        RECT 30.385 188.225 30.675 188.270 ;
        RECT 35.905 188.225 36.195 188.270 ;
        RECT 36.440 188.130 36.580 188.270 ;
        RECT 39.525 188.250 39.815 188.565 ;
        RECT 40.605 188.410 40.895 188.455 ;
        RECT 44.185 188.410 44.475 188.455 ;
        RECT 46.020 188.410 46.310 188.455 ;
        RECT 40.605 188.270 46.310 188.410 ;
        RECT 40.605 188.225 40.895 188.270 ;
        RECT 44.185 188.225 44.475 188.270 ;
        RECT 46.020 188.225 46.310 188.270 ;
        RECT 55.670 188.210 55.990 188.470 ;
        RECT 56.590 188.410 56.910 188.470 ;
        RECT 57.525 188.410 57.815 188.455 ;
        RECT 56.590 188.270 57.815 188.410 ;
        RECT 59.900 188.410 60.040 188.905 ;
        RECT 60.270 188.890 60.590 189.150 ;
        RECT 67.185 189.090 67.475 189.135 ;
        RECT 73.150 189.090 73.470 189.150 ;
        RECT 67.185 188.950 73.470 189.090 ;
        RECT 67.185 188.905 67.475 188.950 ;
        RECT 73.150 188.890 73.470 188.950 ;
        RECT 87.425 189.090 87.715 189.135 ;
        RECT 87.870 189.090 88.190 189.150 ;
        RECT 87.425 188.950 88.190 189.090 ;
        RECT 87.425 188.905 87.715 188.950 ;
        RECT 87.870 188.890 88.190 188.950 ;
        RECT 90.185 189.090 90.475 189.135 ;
        RECT 90.630 189.090 90.950 189.150 ;
        RECT 90.185 188.950 90.950 189.090 ;
        RECT 90.185 188.905 90.475 188.950 ;
        RECT 90.630 188.890 90.950 188.950 ;
        RECT 106.270 189.090 106.590 189.150 ;
        RECT 107.205 189.090 107.495 189.135 ;
        RECT 106.270 188.950 107.495 189.090 ;
        RECT 106.270 188.890 106.590 188.950 ;
        RECT 107.205 188.905 107.495 188.950 ;
        RECT 114.105 189.090 114.395 189.135 ;
        RECT 116.390 189.090 116.710 189.150 ;
        RECT 114.105 188.950 116.710 189.090 ;
        RECT 114.105 188.905 114.395 188.950 ;
        RECT 116.390 188.890 116.710 188.950 ;
        RECT 99.485 188.750 99.775 188.795 ;
        RECT 100.290 188.750 100.610 188.810 ;
        RECT 102.725 188.750 103.375 188.795 ;
        RECT 99.485 188.610 103.375 188.750 ;
        RECT 99.485 188.565 100.075 188.610 ;
        RECT 61.205 188.410 61.495 188.455 ;
        RECT 59.900 188.270 61.495 188.410 ;
        RECT 56.590 188.210 56.910 188.270 ;
        RECT 57.525 188.225 57.815 188.270 ;
        RECT 61.205 188.225 61.495 188.270 ;
        RECT 87.885 188.225 88.175 188.455 ;
        RECT 28.530 188.070 28.850 188.130 ;
        RECT 29.925 188.070 30.215 188.115 ;
        RECT 28.530 187.930 30.215 188.070 ;
        RECT 28.530 187.870 28.850 187.930 ;
        RECT 29.925 187.885 30.215 187.930 ;
        RECT 36.350 187.870 36.670 188.130 ;
        RECT 44.630 188.070 44.950 188.130 ;
        RECT 46.485 188.070 46.775 188.115 ;
        RECT 44.630 187.930 46.775 188.070 ;
        RECT 44.630 187.870 44.950 187.930 ;
        RECT 46.485 187.885 46.775 187.930 ;
        RECT 46.930 188.070 47.250 188.130 ;
        RECT 57.065 188.070 57.355 188.115 ;
        RECT 46.930 187.930 57.355 188.070 ;
        RECT 40.605 187.730 40.895 187.775 ;
        RECT 43.725 187.730 44.015 187.775 ;
        RECT 45.615 187.730 45.905 187.775 ;
        RECT 40.605 187.590 45.905 187.730 ;
        RECT 46.560 187.730 46.700 187.885 ;
        RECT 46.930 187.870 47.250 187.930 ;
        RECT 57.065 187.885 57.355 187.930 ;
        RECT 62.110 188.070 62.430 188.130 ;
        RECT 64.425 188.070 64.715 188.115 ;
        RECT 65.790 188.070 66.110 188.130 ;
        RECT 72.230 188.070 72.550 188.130 ;
        RECT 62.110 187.930 72.550 188.070 ;
        RECT 87.960 188.070 88.100 188.225 ;
        RECT 89.250 188.210 89.570 188.470 ;
        RECT 99.785 188.250 100.075 188.565 ;
        RECT 100.290 188.550 100.610 188.610 ;
        RECT 102.725 188.565 103.375 188.610 ;
        RECT 100.865 188.410 101.155 188.455 ;
        RECT 104.445 188.410 104.735 188.455 ;
        RECT 106.280 188.410 106.570 188.455 ;
        RECT 100.865 188.270 106.570 188.410 ;
        RECT 100.865 188.225 101.155 188.270 ;
        RECT 104.445 188.225 104.735 188.270 ;
        RECT 106.280 188.225 106.570 188.270 ;
        RECT 109.950 188.210 110.270 188.470 ;
        RECT 113.170 188.210 113.490 188.470 ;
        RECT 90.170 188.070 90.490 188.130 ;
        RECT 91.090 188.070 91.410 188.130 ;
        RECT 87.960 187.930 91.410 188.070 ;
        RECT 62.110 187.870 62.430 187.930 ;
        RECT 64.425 187.885 64.715 187.930 ;
        RECT 65.790 187.870 66.110 187.930 ;
        RECT 72.230 187.870 72.550 187.930 ;
        RECT 90.170 187.870 90.490 187.930 ;
        RECT 91.090 187.870 91.410 187.930 ;
        RECT 106.745 188.070 107.035 188.115 ;
        RECT 118.230 188.070 118.550 188.130 ;
        RECT 106.745 187.930 118.550 188.070 ;
        RECT 106.745 187.885 107.035 187.930 ;
        RECT 118.230 187.870 118.550 187.930 ;
        RECT 49.230 187.730 49.550 187.790 ;
        RECT 59.350 187.730 59.670 187.790 ;
        RECT 46.560 187.590 59.670 187.730 ;
        RECT 40.605 187.545 40.895 187.590 ;
        RECT 43.725 187.545 44.015 187.590 ;
        RECT 45.615 187.545 45.905 187.590 ;
        RECT 49.230 187.530 49.550 187.590 ;
        RECT 59.350 187.530 59.670 187.590 ;
        RECT 100.865 187.730 101.155 187.775 ;
        RECT 103.985 187.730 104.275 187.775 ;
        RECT 105.875 187.730 106.165 187.775 ;
        RECT 100.865 187.590 106.165 187.730 ;
        RECT 100.865 187.545 101.155 187.590 ;
        RECT 103.985 187.545 104.275 187.590 ;
        RECT 105.875 187.545 106.165 187.590 ;
        RECT 37.730 187.190 38.050 187.450 ;
        RECT 45.200 187.390 45.490 187.435 ;
        RECT 50.150 187.390 50.470 187.450 ;
        RECT 45.200 187.250 50.470 187.390 ;
        RECT 45.200 187.205 45.490 187.250 ;
        RECT 50.150 187.190 50.470 187.250 ;
        RECT 98.005 187.390 98.295 187.435 ;
        RECT 99.370 187.390 99.690 187.450 ;
        RECT 98.005 187.250 99.690 187.390 ;
        RECT 98.005 187.205 98.295 187.250 ;
        RECT 99.370 187.190 99.690 187.250 ;
        RECT 99.830 187.390 100.150 187.450 ;
        RECT 105.430 187.390 105.720 187.435 ;
        RECT 99.830 187.250 105.720 187.390 ;
        RECT 99.830 187.190 100.150 187.250 ;
        RECT 105.430 187.205 105.720 187.250 ;
        RECT 14.660 186.570 127.820 187.050 ;
        RECT 39.110 186.170 39.430 186.430 ;
        RECT 46.010 186.370 46.330 186.430 ;
        RECT 88.345 186.370 88.635 186.415 ;
        RECT 89.250 186.370 89.570 186.430 ;
        RECT 46.010 186.230 47.620 186.370 ;
        RECT 46.010 186.170 46.330 186.230 ;
        RECT 29.105 186.030 29.395 186.075 ;
        RECT 32.225 186.030 32.515 186.075 ;
        RECT 34.115 186.030 34.405 186.075 ;
        RECT 44.630 186.030 44.950 186.090 ;
        RECT 29.105 185.890 34.405 186.030 ;
        RECT 29.105 185.845 29.395 185.890 ;
        RECT 32.225 185.845 32.515 185.890 ;
        RECT 34.115 185.845 34.405 185.890 ;
        RECT 35.060 185.890 44.950 186.030 ;
        RECT 23.010 185.690 23.330 185.750 ;
        RECT 35.060 185.735 35.200 185.890 ;
        RECT 44.630 185.830 44.950 185.890 ;
        RECT 46.470 185.830 46.790 186.090 ;
        RECT 33.605 185.690 33.895 185.735 ;
        RECT 23.010 185.550 33.895 185.690 ;
        RECT 23.010 185.490 23.330 185.550 ;
        RECT 33.605 185.505 33.895 185.550 ;
        RECT 34.985 185.505 35.275 185.735 ;
        RECT 38.190 185.690 38.510 185.750 ;
        RECT 40.505 185.690 40.795 185.735 ;
        RECT 38.190 185.550 40.795 185.690 ;
        RECT 38.190 185.490 38.510 185.550 ;
        RECT 40.505 185.505 40.795 185.550 ;
        RECT 28.025 185.055 28.315 185.370 ;
        RECT 29.105 185.350 29.395 185.395 ;
        RECT 32.685 185.350 32.975 185.395 ;
        RECT 34.520 185.350 34.810 185.395 ;
        RECT 29.105 185.210 34.810 185.350 ;
        RECT 29.105 185.165 29.395 185.210 ;
        RECT 32.685 185.165 32.975 185.210 ;
        RECT 34.520 185.165 34.810 185.210 ;
        RECT 36.350 185.350 36.670 185.410 ;
        RECT 38.665 185.350 38.955 185.395 ;
        RECT 36.350 185.210 38.955 185.350 ;
        RECT 40.580 185.350 40.720 185.505 ;
        RECT 41.410 185.490 41.730 185.750 ;
        RECT 46.560 185.690 46.700 185.830 ;
        RECT 46.945 185.690 47.235 185.735 ;
        RECT 46.100 185.550 47.235 185.690 ;
        RECT 45.550 185.350 45.870 185.410 ;
        RECT 46.100 185.350 46.240 185.550 ;
        RECT 46.945 185.505 47.235 185.550 ;
        RECT 40.580 185.210 46.240 185.350 ;
        RECT 36.350 185.150 36.670 185.210 ;
        RECT 38.665 185.165 38.955 185.210 ;
        RECT 45.550 185.150 45.870 185.210 ;
        RECT 46.485 185.165 46.775 185.395 ;
        RECT 47.480 185.350 47.620 186.230 ;
        RECT 88.345 186.230 89.570 186.370 ;
        RECT 88.345 186.185 88.635 186.230 ;
        RECT 89.250 186.170 89.570 186.230 ;
        RECT 99.830 186.170 100.150 186.430 ;
        RECT 100.290 186.370 100.610 186.430 ;
        RECT 100.765 186.370 101.055 186.415 ;
        RECT 100.290 186.230 101.055 186.370 ;
        RECT 100.290 186.170 100.610 186.230 ;
        RECT 100.765 186.185 101.055 186.230 ;
        RECT 53.485 186.030 53.775 186.075 ;
        RECT 56.605 186.030 56.895 186.075 ;
        RECT 58.495 186.030 58.785 186.075 ;
        RECT 60.730 186.030 61.050 186.090 ;
        RECT 53.485 185.890 58.785 186.030 ;
        RECT 53.485 185.845 53.775 185.890 ;
        RECT 56.605 185.845 56.895 185.890 ;
        RECT 58.495 185.845 58.785 185.890 ;
        RECT 58.980 185.890 61.050 186.030 ;
        RECT 58.980 185.690 59.120 185.890 ;
        RECT 60.730 185.830 61.050 185.890 ;
        RECT 71.310 186.030 71.630 186.090 ;
        RECT 75.005 186.030 75.295 186.075 ;
        RECT 76.370 186.030 76.690 186.090 ;
        RECT 71.310 185.890 76.690 186.030 ;
        RECT 71.310 185.830 71.630 185.890 ;
        RECT 75.005 185.845 75.295 185.890 ;
        RECT 76.370 185.830 76.690 185.890 ;
        RECT 91.090 186.030 91.410 186.090 ;
        RECT 91.090 185.890 100.520 186.030 ;
        RECT 91.090 185.830 91.410 185.890 ;
        RECT 52.080 185.550 59.120 185.690 ;
        RECT 48.785 185.350 49.075 185.395 ;
        RECT 52.080 185.350 52.220 185.550 ;
        RECT 59.350 185.490 59.670 185.750 ;
        RECT 68.090 185.690 68.410 185.750 ;
        RECT 72.705 185.690 72.995 185.735 ;
        RECT 73.610 185.690 73.930 185.750 ;
        RECT 68.090 185.550 73.930 185.690 ;
        RECT 68.090 185.490 68.410 185.550 ;
        RECT 72.705 185.505 72.995 185.550 ;
        RECT 73.610 185.490 73.930 185.550 ;
        RECT 85.110 185.490 85.430 185.750 ;
        RECT 94.785 185.690 95.075 185.735 ;
        RECT 99.370 185.690 99.690 185.750 ;
        RECT 94.785 185.550 99.690 185.690 ;
        RECT 94.785 185.505 95.075 185.550 ;
        RECT 99.370 185.490 99.690 185.550 ;
        RECT 47.480 185.210 52.220 185.350 ;
        RECT 48.785 185.165 49.075 185.210 ;
        RECT 27.725 185.010 28.315 185.055 ;
        RECT 28.530 185.010 28.850 185.070 ;
        RECT 30.965 185.010 31.615 185.055 ;
        RECT 27.725 184.870 31.615 185.010 ;
        RECT 27.725 184.825 28.015 184.870 ;
        RECT 28.530 184.810 28.850 184.870 ;
        RECT 30.965 184.825 31.615 184.870 ;
        RECT 37.730 185.010 38.050 185.070 ;
        RECT 46.560 185.010 46.700 185.165 ;
        RECT 52.405 185.055 52.695 185.370 ;
        RECT 53.485 185.350 53.775 185.395 ;
        RECT 57.065 185.350 57.355 185.395 ;
        RECT 58.900 185.350 59.190 185.395 ;
        RECT 53.485 185.210 59.190 185.350 ;
        RECT 53.485 185.165 53.775 185.210 ;
        RECT 57.065 185.165 57.355 185.210 ;
        RECT 58.900 185.165 59.190 185.210 ;
        RECT 74.530 185.150 74.850 185.410 ;
        RECT 100.380 185.395 100.520 185.890 ;
        RECT 105.350 185.690 105.670 185.750 ;
        RECT 107.205 185.690 107.495 185.735 ;
        RECT 109.030 185.690 109.350 185.750 ;
        RECT 105.350 185.550 109.350 185.690 ;
        RECT 105.350 185.490 105.670 185.550 ;
        RECT 107.205 185.505 107.495 185.550 ;
        RECT 109.030 185.490 109.350 185.550 ;
        RECT 98.925 185.165 99.215 185.395 ;
        RECT 100.305 185.165 100.595 185.395 ;
        RECT 37.730 184.870 46.700 185.010 ;
        RECT 49.245 185.010 49.535 185.055 ;
        RECT 52.105 185.010 52.695 185.055 ;
        RECT 55.345 185.010 55.995 185.055 ;
        RECT 49.245 184.870 55.995 185.010 ;
        RECT 37.730 184.810 38.050 184.870 ;
        RECT 49.245 184.825 49.535 184.870 ;
        RECT 52.105 184.825 52.395 184.870 ;
        RECT 55.345 184.825 55.995 184.870 ;
        RECT 57.970 184.810 58.290 185.070 ;
        RECT 72.245 185.010 72.535 185.055 ;
        RECT 72.690 185.010 73.010 185.070 ;
        RECT 72.245 184.870 73.010 185.010 ;
        RECT 74.620 185.010 74.760 185.150 ;
        RECT 75.005 185.010 75.295 185.055 ;
        RECT 75.910 185.010 76.230 185.070 ;
        RECT 74.620 184.870 76.230 185.010 ;
        RECT 99.000 185.010 99.140 185.165 ;
        RECT 105.810 185.150 106.130 185.410 ;
        RECT 110.410 185.150 110.730 185.410 ;
        RECT 102.605 185.010 102.895 185.055 ;
        RECT 99.000 184.870 102.895 185.010 ;
        RECT 72.245 184.825 72.535 184.870 ;
        RECT 72.690 184.810 73.010 184.870 ;
        RECT 75.005 184.825 75.295 184.870 ;
        RECT 75.910 184.810 76.230 184.870 ;
        RECT 102.605 184.825 102.895 184.870 ;
        RECT 109.965 185.010 110.255 185.055 ;
        RECT 112.250 185.010 112.570 185.070 ;
        RECT 109.965 184.870 112.570 185.010 ;
        RECT 109.965 184.825 110.255 184.870 ;
        RECT 112.250 184.810 112.570 184.870 ;
        RECT 26.245 184.670 26.535 184.715 ;
        RECT 29.910 184.670 30.230 184.730 ;
        RECT 26.245 184.530 30.230 184.670 ;
        RECT 26.245 184.485 26.535 184.530 ;
        RECT 29.910 184.470 30.230 184.530 ;
        RECT 30.370 184.670 30.690 184.730 ;
        RECT 41.885 184.670 42.175 184.715 ;
        RECT 30.370 184.530 42.175 184.670 ;
        RECT 30.370 184.470 30.690 184.530 ;
        RECT 41.885 184.485 42.175 184.530 ;
        RECT 43.710 184.470 44.030 184.730 ;
        RECT 44.170 184.470 44.490 184.730 ;
        RECT 46.010 184.470 46.330 184.730 ;
        RECT 46.470 184.670 46.790 184.730 ;
        RECT 50.625 184.670 50.915 184.715 ;
        RECT 46.470 184.530 50.915 184.670 ;
        RECT 46.470 184.470 46.790 184.530 ;
        RECT 50.625 184.485 50.915 184.530 ;
        RECT 71.325 184.670 71.615 184.715 ;
        RECT 74.530 184.670 74.850 184.730 ;
        RECT 71.325 184.530 74.850 184.670 ;
        RECT 71.325 184.485 71.615 184.530 ;
        RECT 74.530 184.470 74.850 184.530 ;
        RECT 86.030 184.470 86.350 184.730 ;
        RECT 86.490 184.470 86.810 184.730 ;
        RECT 97.530 184.470 97.850 184.730 ;
        RECT 111.790 184.670 112.110 184.730 ;
        RECT 113.645 184.670 113.935 184.715 ;
        RECT 111.790 184.530 113.935 184.670 ;
        RECT 111.790 184.470 112.110 184.530 ;
        RECT 113.645 184.485 113.935 184.530 ;
        RECT 14.660 183.850 127.820 184.330 ;
        RECT 23.010 183.450 23.330 183.710 ;
        RECT 30.370 183.450 30.690 183.710 ;
        RECT 45.090 183.650 45.410 183.710 ;
        RECT 48.785 183.650 49.075 183.695 ;
        RECT 45.090 183.510 49.075 183.650 ;
        RECT 45.090 183.450 45.410 183.510 ;
        RECT 48.785 183.465 49.075 183.510 ;
        RECT 50.150 183.450 50.470 183.710 ;
        RECT 52.465 183.650 52.755 183.695 ;
        RECT 57.970 183.650 58.290 183.710 ;
        RECT 71.310 183.650 71.630 183.710 ;
        RECT 52.465 183.510 58.290 183.650 ;
        RECT 52.465 183.465 52.755 183.510 ;
        RECT 57.970 183.450 58.290 183.510 ;
        RECT 69.100 183.510 71.630 183.650 ;
        RECT 32.685 183.310 32.975 183.355 ;
        RECT 34.050 183.310 34.370 183.370 ;
        RECT 32.685 183.170 34.370 183.310 ;
        RECT 32.685 183.125 32.975 183.170 ;
        RECT 34.050 183.110 34.370 183.170 ;
        RECT 44.645 183.310 44.935 183.355 ;
        RECT 44.645 183.170 51.300 183.310 ;
        RECT 44.645 183.125 44.935 183.170 ;
        RECT 22.105 182.970 22.395 183.015 ;
        RECT 23.485 182.970 23.775 183.015 ;
        RECT 22.105 182.830 23.775 182.970 ;
        RECT 22.105 182.785 22.395 182.830 ;
        RECT 23.485 182.785 23.775 182.830 ;
        RECT 27.625 182.970 27.915 183.015 ;
        RECT 29.910 182.970 30.230 183.030 ;
        RECT 33.145 182.970 33.435 183.015 ;
        RECT 35.890 182.970 36.210 183.030 ;
        RECT 27.625 182.830 36.210 182.970 ;
        RECT 27.625 182.785 27.915 182.830 ;
        RECT 29.910 182.770 30.230 182.830 ;
        RECT 33.145 182.785 33.435 182.830 ;
        RECT 35.890 182.770 36.210 182.830 ;
        RECT 37.730 182.770 38.050 183.030 ;
        RECT 41.885 182.970 42.175 183.015 ;
        RECT 44.170 182.970 44.490 183.030 ;
        RECT 41.885 182.830 44.490 182.970 ;
        RECT 41.885 182.785 42.175 182.830 ;
        RECT 44.170 182.770 44.490 182.830 ;
        RECT 45.565 182.970 45.855 183.015 ;
        RECT 46.470 182.970 46.790 183.030 ;
        RECT 51.160 183.015 51.300 183.170 ;
        RECT 45.565 182.830 46.790 182.970 ;
        RECT 45.565 182.785 45.855 182.830 ;
        RECT 46.470 182.770 46.790 182.830 ;
        RECT 49.705 182.785 49.995 183.015 ;
        RECT 51.085 182.785 51.375 183.015 ;
        RECT 51.545 182.785 51.835 183.015 ;
        RECT 55.685 182.970 55.975 183.015 ;
        RECT 59.350 182.970 59.670 183.030 ;
        RECT 55.685 182.830 59.670 182.970 ;
        RECT 55.685 182.785 55.975 182.830 ;
        RECT 26.705 182.445 26.995 182.675 ;
        RECT 34.065 182.630 34.355 182.675 ;
        RECT 38.190 182.630 38.510 182.690 ;
        RECT 34.065 182.490 38.510 182.630 ;
        RECT 34.065 182.445 34.355 182.490 ;
        RECT 26.780 182.290 26.920 182.445 ;
        RECT 38.190 182.430 38.510 182.490 ;
        RECT 43.710 182.630 44.030 182.690 ;
        RECT 49.780 182.630 49.920 182.785 ;
        RECT 43.710 182.490 49.920 182.630 ;
        RECT 50.150 182.630 50.470 182.690 ;
        RECT 51.620 182.630 51.760 182.785 ;
        RECT 59.350 182.770 59.670 182.830 ;
        RECT 60.285 182.970 60.575 183.015 ;
        RECT 60.730 182.970 61.050 183.030 ;
        RECT 60.285 182.830 61.050 182.970 ;
        RECT 60.285 182.785 60.575 182.830 ;
        RECT 60.730 182.770 61.050 182.830 ;
        RECT 68.090 182.770 68.410 183.030 ;
        RECT 69.100 183.015 69.240 183.510 ;
        RECT 71.310 183.450 71.630 183.510 ;
        RECT 71.770 183.650 72.090 183.710 ;
        RECT 72.690 183.650 73.010 183.710 ;
        RECT 74.070 183.650 74.390 183.710 ;
        RECT 89.725 183.650 90.015 183.695 ;
        RECT 71.770 183.510 76.600 183.650 ;
        RECT 71.770 183.450 72.090 183.510 ;
        RECT 72.690 183.450 73.010 183.510 ;
        RECT 74.070 183.450 74.390 183.510 ;
        RECT 73.610 183.110 73.930 183.370 ;
        RECT 69.025 182.785 69.315 183.015 ;
        RECT 70.865 182.970 71.155 183.015 ;
        RECT 71.770 182.970 72.090 183.030 ;
        RECT 70.865 182.830 72.090 182.970 ;
        RECT 70.865 182.785 71.155 182.830 ;
        RECT 50.150 182.490 51.760 182.630 ;
        RECT 43.710 182.430 44.030 182.490 ;
        RECT 50.150 182.430 50.470 182.490 ;
        RECT 67.645 182.445 67.935 182.675 ;
        RECT 68.565 182.630 68.855 182.675 ;
        RECT 70.940 182.630 71.080 182.785 ;
        RECT 71.770 182.770 72.090 182.830 ;
        RECT 72.245 182.785 72.535 183.015 ;
        RECT 68.565 182.490 71.080 182.630 ;
        RECT 72.320 182.630 72.460 182.785 ;
        RECT 72.690 182.770 73.010 183.030 ;
        RECT 73.700 182.970 73.840 183.110 ;
        RECT 75.005 182.970 75.295 183.015 ;
        RECT 73.700 182.830 75.295 182.970 ;
        RECT 75.005 182.785 75.295 182.830 ;
        RECT 72.320 182.490 72.920 182.630 ;
        RECT 68.565 182.445 68.855 182.490 ;
        RECT 30.845 182.290 31.135 182.335 ;
        RECT 26.780 182.150 31.135 182.290 ;
        RECT 67.720 182.290 67.860 182.445 ;
        RECT 72.780 182.350 72.920 182.490 ;
        RECT 73.610 182.430 73.930 182.690 ;
        RECT 75.080 182.630 75.220 182.785 ;
        RECT 75.910 182.770 76.230 183.030 ;
        RECT 76.460 183.015 76.600 183.510 ;
        RECT 86.580 183.510 90.015 183.650 ;
        RECT 81.085 183.310 81.375 183.355 ;
        RECT 84.325 183.310 84.975 183.355 ;
        RECT 86.580 183.310 86.720 183.510 ;
        RECT 89.725 183.465 90.015 183.510 ;
        RECT 97.530 183.450 97.850 183.710 ;
        RECT 105.810 183.650 106.130 183.710 ;
        RECT 106.285 183.650 106.575 183.695 ;
        RECT 105.810 183.510 106.575 183.650 ;
        RECT 105.810 183.450 106.130 183.510 ;
        RECT 106.285 183.465 106.575 183.510 ;
        RECT 111.805 183.465 112.095 183.695 ;
        RECT 81.085 183.170 86.720 183.310 ;
        RECT 104.445 183.310 104.735 183.355 ;
        RECT 111.880 183.310 112.020 183.465 ;
        RECT 104.445 183.170 112.020 183.310 ;
        RECT 117.425 183.310 117.715 183.355 ;
        RECT 120.665 183.310 121.315 183.355 ;
        RECT 117.425 183.170 121.315 183.310 ;
        RECT 81.085 183.125 81.675 183.170 ;
        RECT 84.325 183.125 84.975 183.170 ;
        RECT 104.445 183.125 104.735 183.170 ;
        RECT 76.385 182.785 76.675 183.015 ;
        RECT 76.830 182.770 77.150 183.030 ;
        RECT 81.385 182.810 81.675 183.125 ;
        RECT 105.900 183.030 106.040 183.170 ;
        RECT 117.425 183.125 118.015 183.170 ;
        RECT 120.665 183.125 121.315 183.170 ;
        RECT 123.305 183.310 123.595 183.355 ;
        RECT 124.670 183.310 124.990 183.370 ;
        RECT 123.305 183.170 124.990 183.310 ;
        RECT 123.305 183.125 123.595 183.170 ;
        RECT 117.725 183.030 118.015 183.125 ;
        RECT 124.670 183.110 124.990 183.170 ;
        RECT 82.465 182.970 82.755 183.015 ;
        RECT 86.045 182.970 86.335 183.015 ;
        RECT 87.880 182.970 88.170 183.015 ;
        RECT 82.465 182.830 88.170 182.970 ;
        RECT 82.465 182.785 82.755 182.830 ;
        RECT 86.045 182.785 86.335 182.830 ;
        RECT 87.880 182.785 88.170 182.830 ;
        RECT 90.185 182.970 90.475 183.015 ;
        RECT 91.090 182.970 91.410 183.030 ;
        RECT 90.185 182.830 91.410 182.970 ;
        RECT 90.185 182.785 90.475 182.830 ;
        RECT 91.090 182.770 91.410 182.830 ;
        RECT 96.150 182.970 96.470 183.030 ;
        RECT 97.085 182.970 97.375 183.015 ;
        RECT 96.150 182.830 97.375 182.970 ;
        RECT 96.150 182.770 96.470 182.830 ;
        RECT 97.085 182.785 97.375 182.830 ;
        RECT 99.370 182.970 99.690 183.030 ;
        RECT 103.985 182.970 104.275 183.015 ;
        RECT 99.370 182.830 104.275 182.970 ;
        RECT 99.370 182.770 99.690 182.830 ;
        RECT 103.985 182.785 104.275 182.830 ;
        RECT 105.810 182.770 106.130 183.030 ;
        RECT 106.270 182.970 106.590 183.030 ;
        RECT 106.270 182.830 107.880 182.970 ;
        RECT 106.270 182.770 106.590 182.830 ;
        RECT 77.305 182.630 77.595 182.675 ;
        RECT 75.080 182.490 77.595 182.630 ;
        RECT 77.305 182.445 77.595 182.490 ;
        RECT 86.965 182.630 87.255 182.675 ;
        RECT 88.345 182.630 88.635 182.675 ;
        RECT 93.850 182.630 94.170 182.690 ;
        RECT 86.965 182.490 88.100 182.630 ;
        RECT 86.965 182.445 87.255 182.490 ;
        RECT 72.690 182.290 73.010 182.350 ;
        RECT 75.910 182.290 76.230 182.350 ;
        RECT 67.720 182.150 76.230 182.290 ;
        RECT 30.845 182.105 31.135 182.150 ;
        RECT 72.690 182.090 73.010 182.150 ;
        RECT 75.910 182.090 76.230 182.150 ;
        RECT 82.465 182.290 82.755 182.335 ;
        RECT 85.585 182.290 85.875 182.335 ;
        RECT 87.475 182.290 87.765 182.335 ;
        RECT 82.465 182.150 87.765 182.290 ;
        RECT 87.960 182.290 88.100 182.490 ;
        RECT 88.345 182.490 94.170 182.630 ;
        RECT 88.345 182.445 88.635 182.490 ;
        RECT 93.850 182.430 94.170 182.490 ;
        RECT 96.625 182.630 96.915 182.675 ;
        RECT 97.990 182.630 98.310 182.690 ;
        RECT 103.065 182.630 103.355 182.675 ;
        RECT 96.625 182.490 103.355 182.630 ;
        RECT 96.625 182.445 96.915 182.490 ;
        RECT 89.710 182.290 90.030 182.350 ;
        RECT 87.960 182.150 90.030 182.290 ;
        RECT 82.465 182.105 82.755 182.150 ;
        RECT 85.585 182.105 85.875 182.150 ;
        RECT 87.475 182.105 87.765 182.150 ;
        RECT 89.710 182.090 90.030 182.150 ;
        RECT 39.570 181.950 39.890 182.010 ;
        RECT 40.965 181.950 41.255 181.995 ;
        RECT 39.570 181.810 41.255 181.950 ;
        RECT 39.570 181.750 39.890 181.810 ;
        RECT 40.965 181.765 41.255 181.810 ;
        RECT 46.010 181.950 46.330 182.010 ;
        RECT 47.390 181.950 47.710 182.010 ;
        RECT 48.325 181.950 48.615 181.995 ;
        RECT 46.010 181.810 48.615 181.950 ;
        RECT 46.010 181.750 46.330 181.810 ;
        RECT 47.390 181.750 47.710 181.810 ;
        RECT 48.325 181.765 48.615 181.810 ;
        RECT 56.130 181.950 56.450 182.010 ;
        RECT 59.825 181.950 60.115 181.995 ;
        RECT 56.130 181.810 60.115 181.950 ;
        RECT 56.130 181.750 56.450 181.810 ;
        RECT 59.825 181.765 60.115 181.810 ;
        RECT 66.725 181.950 67.015 181.995 ;
        RECT 69.470 181.950 69.790 182.010 ;
        RECT 66.725 181.810 69.790 181.950 ;
        RECT 66.725 181.765 67.015 181.810 ;
        RECT 69.470 181.750 69.790 181.810 ;
        RECT 74.990 181.950 75.310 182.010 ;
        RECT 78.225 181.950 78.515 181.995 ;
        RECT 74.990 181.810 78.515 181.950 ;
        RECT 74.990 181.750 75.310 181.810 ;
        RECT 78.225 181.765 78.515 181.810 ;
        RECT 79.590 181.750 79.910 182.010 ;
        RECT 85.110 181.950 85.430 182.010 ;
        RECT 96.700 181.950 96.840 182.445 ;
        RECT 97.990 182.430 98.310 182.490 ;
        RECT 103.065 182.445 103.355 182.490 ;
        RECT 104.430 182.630 104.750 182.690 ;
        RECT 106.745 182.630 107.035 182.675 ;
        RECT 104.430 182.490 107.035 182.630 ;
        RECT 107.740 182.630 107.880 182.830 ;
        RECT 108.110 182.770 108.430 183.030 ;
        RECT 108.585 182.785 108.875 183.015 ;
        RECT 109.045 182.785 109.335 183.015 ;
        RECT 109.490 182.970 109.810 183.030 ;
        RECT 109.965 182.970 110.255 183.015 ;
        RECT 109.490 182.830 110.255 182.970 ;
        RECT 108.660 182.630 108.800 182.785 ;
        RECT 107.740 182.490 108.800 182.630 ;
        RECT 104.430 182.430 104.750 182.490 ;
        RECT 106.745 182.445 107.035 182.490 ;
        RECT 98.450 182.290 98.770 182.350 ;
        RECT 109.120 182.290 109.260 182.785 ;
        RECT 109.490 182.770 109.810 182.830 ;
        RECT 109.965 182.785 110.255 182.830 ;
        RECT 111.790 182.970 112.110 183.030 ;
        RECT 112.265 182.970 112.555 183.015 ;
        RECT 111.790 182.830 112.555 182.970 ;
        RECT 111.790 182.770 112.110 182.830 ;
        RECT 112.265 182.785 112.555 182.830 ;
        RECT 117.725 182.810 118.090 183.030 ;
        RECT 117.770 182.770 118.090 182.810 ;
        RECT 118.805 182.970 119.095 183.015 ;
        RECT 122.385 182.970 122.675 183.015 ;
        RECT 124.220 182.970 124.510 183.015 ;
        RECT 118.805 182.830 124.510 182.970 ;
        RECT 118.805 182.785 119.095 182.830 ;
        RECT 122.385 182.785 122.675 182.830 ;
        RECT 124.220 182.785 124.510 182.830 ;
        RECT 110.870 182.430 111.190 182.690 ;
        RECT 118.230 182.630 118.550 182.690 ;
        RECT 124.685 182.630 124.975 182.675 ;
        RECT 118.230 182.490 124.975 182.630 ;
        RECT 118.230 182.430 118.550 182.490 ;
        RECT 124.685 182.445 124.975 182.490 ;
        RECT 98.450 182.150 109.260 182.290 ;
        RECT 110.410 182.290 110.730 182.350 ;
        RECT 115.945 182.290 116.235 182.335 ;
        RECT 110.410 182.150 116.235 182.290 ;
        RECT 98.450 182.090 98.770 182.150 ;
        RECT 110.410 182.090 110.730 182.150 ;
        RECT 115.945 182.105 116.235 182.150 ;
        RECT 118.805 182.290 119.095 182.335 ;
        RECT 121.925 182.290 122.215 182.335 ;
        RECT 123.815 182.290 124.105 182.335 ;
        RECT 118.805 182.150 124.105 182.290 ;
        RECT 118.805 182.105 119.095 182.150 ;
        RECT 121.925 182.105 122.215 182.150 ;
        RECT 123.815 182.105 124.105 182.150 ;
        RECT 85.110 181.810 96.840 181.950 ;
        RECT 99.385 181.950 99.675 181.995 ;
        RECT 104.890 181.950 105.210 182.010 ;
        RECT 99.385 181.810 105.210 181.950 ;
        RECT 85.110 181.750 85.430 181.810 ;
        RECT 99.385 181.765 99.675 181.810 ;
        RECT 104.890 181.750 105.210 181.810 ;
        RECT 114.105 181.950 114.395 181.995 ;
        RECT 116.850 181.950 117.170 182.010 ;
        RECT 114.105 181.810 117.170 181.950 ;
        RECT 114.105 181.765 114.395 181.810 ;
        RECT 116.850 181.750 117.170 181.810 ;
        RECT 14.660 181.130 127.820 181.610 ;
        RECT 45.550 180.930 45.870 180.990 ;
        RECT 46.930 180.930 47.250 180.990 ;
        RECT 45.550 180.790 47.250 180.930 ;
        RECT 45.550 180.730 45.870 180.790 ;
        RECT 46.930 180.730 47.250 180.790 ;
        RECT 49.705 180.930 49.995 180.975 ;
        RECT 50.150 180.930 50.470 180.990 ;
        RECT 82.350 180.930 82.670 180.990 ;
        RECT 49.705 180.790 50.470 180.930 ;
        RECT 49.705 180.745 49.995 180.790 ;
        RECT 50.150 180.730 50.470 180.790 ;
        RECT 78.760 180.790 82.670 180.930 ;
        RECT 25.735 180.590 26.025 180.635 ;
        RECT 27.625 180.590 27.915 180.635 ;
        RECT 30.745 180.590 31.035 180.635 ;
        RECT 25.735 180.450 31.035 180.590 ;
        RECT 25.735 180.405 26.025 180.450 ;
        RECT 27.625 180.405 27.915 180.450 ;
        RECT 30.745 180.405 31.035 180.450 ;
        RECT 53.845 180.590 54.135 180.635 ;
        RECT 56.590 180.590 56.910 180.650 ;
        RECT 53.845 180.450 56.910 180.590 ;
        RECT 53.845 180.405 54.135 180.450 ;
        RECT 56.590 180.390 56.910 180.450 ;
        RECT 67.630 180.590 67.950 180.650 ;
        RECT 78.760 180.590 78.900 180.790 ;
        RECT 82.350 180.730 82.670 180.790 ;
        RECT 89.710 180.730 90.030 180.990 ;
        RECT 105.810 180.730 106.130 180.990 ;
        RECT 117.770 180.930 118.090 180.990 ;
        RECT 122.845 180.930 123.135 180.975 ;
        RECT 124.670 180.930 124.990 180.990 ;
        RECT 117.770 180.790 119.840 180.930 ;
        RECT 117.770 180.730 118.090 180.790 ;
        RECT 67.630 180.450 78.900 180.590 ;
        RECT 79.130 180.590 79.450 180.650 ;
        RECT 85.570 180.590 85.890 180.650 ;
        RECT 79.130 180.450 85.890 180.590 ;
        RECT 67.630 180.390 67.950 180.450 ;
        RECT 79.130 180.390 79.450 180.450 ;
        RECT 85.570 180.390 85.890 180.450 ;
        RECT 95.345 180.590 95.635 180.635 ;
        RECT 98.465 180.590 98.755 180.635 ;
        RECT 100.355 180.590 100.645 180.635 ;
        RECT 95.345 180.450 100.645 180.590 ;
        RECT 95.345 180.405 95.635 180.450 ;
        RECT 98.465 180.405 98.755 180.450 ;
        RECT 100.355 180.405 100.645 180.450 ;
        RECT 114.205 180.590 114.495 180.635 ;
        RECT 117.325 180.590 117.615 180.635 ;
        RECT 119.215 180.590 119.505 180.635 ;
        RECT 114.205 180.450 119.505 180.590 ;
        RECT 119.700 180.590 119.840 180.790 ;
        RECT 122.845 180.790 124.990 180.930 ;
        RECT 122.845 180.745 123.135 180.790 ;
        RECT 124.670 180.730 124.990 180.790 ;
        RECT 121.005 180.590 121.295 180.635 ;
        RECT 119.700 180.450 121.295 180.590 ;
        RECT 114.205 180.405 114.495 180.450 ;
        RECT 117.325 180.405 117.615 180.450 ;
        RECT 119.215 180.405 119.505 180.450 ;
        RECT 121.005 180.405 121.295 180.450 ;
        RECT 33.605 180.065 33.895 180.295 ;
        RECT 46.470 180.250 46.790 180.310 ;
        RECT 44.720 180.110 46.790 180.250 ;
        RECT 24.865 179.725 25.155 179.955 ;
        RECT 25.330 179.910 25.620 179.955 ;
        RECT 27.165 179.910 27.455 179.955 ;
        RECT 30.745 179.910 31.035 179.955 ;
        RECT 25.330 179.770 31.035 179.910 ;
        RECT 25.330 179.725 25.620 179.770 ;
        RECT 27.165 179.725 27.455 179.770 ;
        RECT 30.745 179.725 31.035 179.770 ;
        RECT 24.940 179.570 25.080 179.725 ;
        RECT 24.940 179.430 25.540 179.570 ;
        RECT 25.400 179.230 25.540 179.430 ;
        RECT 26.230 179.370 26.550 179.630 ;
        RECT 27.610 179.570 27.930 179.630 ;
        RECT 31.825 179.615 32.115 179.930 ;
        RECT 33.680 179.910 33.820 180.065 ;
        RECT 37.270 179.910 37.590 179.970 ;
        RECT 33.680 179.770 37.590 179.910 ;
        RECT 37.270 179.710 37.590 179.770 ;
        RECT 39.585 179.725 39.875 179.955 ;
        RECT 40.045 179.725 40.335 179.955 ;
        RECT 40.505 179.910 40.795 179.955 ;
        RECT 40.950 179.910 41.270 179.970 ;
        RECT 40.505 179.770 41.270 179.910 ;
        RECT 40.505 179.725 40.795 179.770 ;
        RECT 28.525 179.570 29.175 179.615 ;
        RECT 31.825 179.570 32.415 179.615 ;
        RECT 27.610 179.430 32.415 179.570 ;
        RECT 27.610 179.370 27.930 179.430 ;
        RECT 28.525 179.385 29.175 179.430 ;
        RECT 32.125 179.385 32.415 179.430 ;
        RECT 34.050 179.370 34.370 179.630 ;
        RECT 34.970 179.570 35.290 179.630 ;
        RECT 38.205 179.570 38.495 179.615 ;
        RECT 34.970 179.430 38.495 179.570 ;
        RECT 34.970 179.370 35.290 179.430 ;
        RECT 38.205 179.385 38.495 179.430 ;
        RECT 36.810 179.230 37.130 179.290 ;
        RECT 25.400 179.090 37.130 179.230 ;
        RECT 39.660 179.230 39.800 179.725 ;
        RECT 40.120 179.570 40.260 179.725 ;
        RECT 40.950 179.710 41.270 179.770 ;
        RECT 41.425 179.725 41.715 179.955 ;
        RECT 43.725 179.725 44.015 179.955 ;
        RECT 40.120 179.430 40.720 179.570 ;
        RECT 40.580 179.290 40.720 179.430 ;
        RECT 40.030 179.230 40.350 179.290 ;
        RECT 39.660 179.090 40.350 179.230 ;
        RECT 36.810 179.030 37.130 179.090 ;
        RECT 40.030 179.030 40.350 179.090 ;
        RECT 40.490 179.030 40.810 179.290 ;
        RECT 40.950 179.230 41.270 179.290 ;
        RECT 41.500 179.230 41.640 179.725 ;
        RECT 40.950 179.090 41.640 179.230 ;
        RECT 40.950 179.030 41.270 179.090 ;
        RECT 42.330 179.030 42.650 179.290 ;
        RECT 43.800 179.230 43.940 179.725 ;
        RECT 44.170 179.710 44.490 179.970 ;
        RECT 44.720 179.955 44.860 180.110 ;
        RECT 46.470 180.050 46.790 180.110 ;
        RECT 46.930 180.050 47.250 180.310 ;
        RECT 47.390 180.050 47.710 180.310 ;
        RECT 51.085 180.250 51.375 180.295 ;
        RECT 52.450 180.250 52.770 180.310 ;
        RECT 51.085 180.110 52.770 180.250 ;
        RECT 51.085 180.065 51.375 180.110 ;
        RECT 52.450 180.050 52.770 180.110 ;
        RECT 54.290 180.250 54.610 180.310 ;
        RECT 58.905 180.250 59.195 180.295 ;
        RECT 60.745 180.250 61.035 180.295 ;
        RECT 54.290 180.110 61.035 180.250 ;
        RECT 54.290 180.050 54.610 180.110 ;
        RECT 58.905 180.065 59.195 180.110 ;
        RECT 60.745 180.065 61.035 180.110 ;
        RECT 72.690 180.050 73.010 180.310 ;
        RECT 73.150 180.050 73.470 180.310 ;
        RECT 73.625 180.250 73.915 180.295 ;
        RECT 75.910 180.250 76.230 180.310 ;
        RECT 73.625 180.110 76.230 180.250 ;
        RECT 73.625 180.065 73.915 180.110 ;
        RECT 75.910 180.050 76.230 180.110 ;
        RECT 76.845 180.250 77.135 180.295 ;
        RECT 79.590 180.250 79.910 180.310 ;
        RECT 85.110 180.250 85.430 180.310 ;
        RECT 86.045 180.250 86.335 180.295 ;
        RECT 76.845 180.110 81.200 180.250 ;
        RECT 76.845 180.065 77.135 180.110 ;
        RECT 79.590 180.050 79.910 180.110 ;
        RECT 44.645 179.725 44.935 179.955 ;
        RECT 45.550 179.710 45.870 179.970 ;
        RECT 65.790 179.710 66.110 179.970 ;
        RECT 68.550 179.710 68.870 179.970 ;
        RECT 71.310 179.910 71.630 179.970 ;
        RECT 71.785 179.910 72.075 179.955 ;
        RECT 71.310 179.770 72.075 179.910 ;
        RECT 71.310 179.710 71.630 179.770 ;
        RECT 71.785 179.725 72.075 179.770 ;
        RECT 74.070 179.710 74.390 179.970 ;
        RECT 76.370 179.910 76.690 179.970 ;
        RECT 81.060 179.955 81.200 180.110 ;
        RECT 85.110 180.110 86.335 180.250 ;
        RECT 85.110 180.050 85.430 180.110 ;
        RECT 86.045 180.065 86.335 180.110 ;
        RECT 104.890 180.050 105.210 180.310 ;
        RECT 105.810 180.250 106.130 180.310 ;
        RECT 108.110 180.250 108.430 180.310 ;
        RECT 111.345 180.250 111.635 180.295 ;
        RECT 115.930 180.250 116.250 180.310 ;
        RECT 105.810 180.110 108.430 180.250 ;
        RECT 105.810 180.050 106.130 180.110 ;
        RECT 108.110 180.050 108.430 180.110 ;
        RECT 109.120 180.110 111.635 180.250 ;
        RECT 109.120 179.970 109.260 180.110 ;
        RECT 111.345 180.065 111.635 180.110 ;
        RECT 111.880 180.110 120.760 180.250 ;
        RECT 80.065 179.910 80.355 179.955 ;
        RECT 76.370 179.770 80.355 179.910 ;
        RECT 76.370 179.710 76.690 179.770 ;
        RECT 53.830 179.570 54.150 179.630 ;
        RECT 58.445 179.570 58.735 179.615 ;
        RECT 53.830 179.430 58.735 179.570 ;
        RECT 53.830 179.370 54.150 179.430 ;
        RECT 58.445 179.385 58.735 179.430 ;
        RECT 62.125 179.570 62.415 179.615 ;
        RECT 69.485 179.570 69.775 179.615 ;
        RECT 73.150 179.570 73.470 179.630 ;
        RECT 62.125 179.430 73.470 179.570 ;
        RECT 62.125 179.385 62.415 179.430 ;
        RECT 69.485 179.385 69.775 179.430 ;
        RECT 73.150 179.370 73.470 179.430 ;
        RECT 44.630 179.230 44.950 179.290 ;
        RECT 43.800 179.090 44.950 179.230 ;
        RECT 44.630 179.030 44.950 179.090 ;
        RECT 46.010 179.230 46.330 179.290 ;
        RECT 47.865 179.230 48.155 179.275 ;
        RECT 46.010 179.090 48.155 179.230 ;
        RECT 46.010 179.030 46.330 179.090 ;
        RECT 47.865 179.045 48.155 179.090 ;
        RECT 50.610 179.230 50.930 179.290 ;
        RECT 56.145 179.230 56.435 179.275 ;
        RECT 50.610 179.090 56.435 179.230 ;
        RECT 50.610 179.030 50.930 179.090 ;
        RECT 56.145 179.045 56.435 179.090 ;
        RECT 57.970 179.030 58.290 179.290 ;
        RECT 66.250 179.030 66.570 179.290 ;
        RECT 70.865 179.230 71.155 179.275 ;
        RECT 78.670 179.230 78.990 179.290 ;
        RECT 70.865 179.090 78.990 179.230 ;
        RECT 79.220 179.230 79.360 179.770 ;
        RECT 80.065 179.725 80.355 179.770 ;
        RECT 80.985 179.725 81.275 179.955 ;
        RECT 81.430 179.710 81.750 179.970 ;
        RECT 81.890 179.710 82.210 179.970 ;
        RECT 90.630 179.710 90.950 179.970 ;
        RECT 91.090 179.710 91.410 179.970 ;
        RECT 79.605 179.570 79.895 179.615 ;
        RECT 86.490 179.570 86.810 179.630 ;
        RECT 94.265 179.615 94.555 179.930 ;
        RECT 95.345 179.910 95.635 179.955 ;
        RECT 98.925 179.910 99.215 179.955 ;
        RECT 100.760 179.910 101.050 179.955 ;
        RECT 95.345 179.770 101.050 179.910 ;
        RECT 95.345 179.725 95.635 179.770 ;
        RECT 98.925 179.725 99.215 179.770 ;
        RECT 100.760 179.725 101.050 179.770 ;
        RECT 101.225 179.725 101.515 179.955 ;
        RECT 86.965 179.570 87.255 179.615 ;
        RECT 91.565 179.570 91.855 179.615 ;
        RECT 93.965 179.570 94.555 179.615 ;
        RECT 97.205 179.570 97.855 179.615 ;
        RECT 79.605 179.430 87.255 179.570 ;
        RECT 79.605 179.385 79.895 179.430 ;
        RECT 86.490 179.370 86.810 179.430 ;
        RECT 86.965 179.385 87.255 179.430 ;
        RECT 87.500 179.430 90.400 179.570 ;
        RECT 87.500 179.290 87.640 179.430 ;
        RECT 82.810 179.230 83.130 179.290 ;
        RECT 79.220 179.090 83.130 179.230 ;
        RECT 70.865 179.045 71.155 179.090 ;
        RECT 78.670 179.030 78.990 179.090 ;
        RECT 82.810 179.030 83.130 179.090 ;
        RECT 83.285 179.230 83.575 179.275 ;
        RECT 83.730 179.230 84.050 179.290 ;
        RECT 83.285 179.090 84.050 179.230 ;
        RECT 83.285 179.045 83.575 179.090 ;
        RECT 83.730 179.030 84.050 179.090 ;
        RECT 87.410 179.030 87.730 179.290 ;
        RECT 89.250 179.030 89.570 179.290 ;
        RECT 90.260 179.230 90.400 179.430 ;
        RECT 91.565 179.430 97.855 179.570 ;
        RECT 91.565 179.385 91.855 179.430 ;
        RECT 93.965 179.385 94.255 179.430 ;
        RECT 97.205 179.385 97.855 179.430 ;
        RECT 99.830 179.370 100.150 179.630 ;
        RECT 92.485 179.230 92.775 179.275 ;
        RECT 96.150 179.230 96.470 179.290 ;
        RECT 90.260 179.090 96.470 179.230 ;
        RECT 101.300 179.230 101.440 179.725 ;
        RECT 109.030 179.710 109.350 179.970 ;
        RECT 109.965 179.910 110.255 179.955 ;
        RECT 111.880 179.910 112.020 180.110 ;
        RECT 115.930 180.050 116.250 180.110 ;
        RECT 120.620 179.955 120.760 180.110 ;
        RECT 109.965 179.770 112.020 179.910 ;
        RECT 109.965 179.725 110.255 179.770 ;
        RECT 102.130 179.370 102.450 179.630 ;
        RECT 113.125 179.615 113.415 179.930 ;
        RECT 114.205 179.910 114.495 179.955 ;
        RECT 117.785 179.910 118.075 179.955 ;
        RECT 119.620 179.910 119.910 179.955 ;
        RECT 114.205 179.770 119.910 179.910 ;
        RECT 114.205 179.725 114.495 179.770 ;
        RECT 117.785 179.725 118.075 179.770 ;
        RECT 119.620 179.725 119.910 179.770 ;
        RECT 120.085 179.725 120.375 179.955 ;
        RECT 120.545 179.725 120.835 179.955 ;
        RECT 110.425 179.570 110.715 179.615 ;
        RECT 112.825 179.570 113.415 179.615 ;
        RECT 116.065 179.570 116.715 179.615 ;
        RECT 110.425 179.430 116.715 179.570 ;
        RECT 110.425 179.385 110.715 179.430 ;
        RECT 112.825 179.385 113.115 179.430 ;
        RECT 116.065 179.385 116.715 179.430 ;
        RECT 118.690 179.370 119.010 179.630 ;
        RECT 118.230 179.230 118.550 179.290 ;
        RECT 120.160 179.230 120.300 179.725 ;
        RECT 121.910 179.710 122.230 179.970 ;
        RECT 101.300 179.090 120.300 179.230 ;
        RECT 92.485 179.045 92.775 179.090 ;
        RECT 96.150 179.030 96.470 179.090 ;
        RECT 118.230 179.030 118.550 179.090 ;
        RECT 14.660 178.410 127.820 178.890 ;
        RECT 25.785 178.210 26.075 178.255 ;
        RECT 27.610 178.210 27.930 178.270 ;
        RECT 25.785 178.070 27.930 178.210 ;
        RECT 25.785 178.025 26.075 178.070 ;
        RECT 27.610 178.010 27.930 178.070 ;
        RECT 39.570 178.010 39.890 178.270 ;
        RECT 46.010 178.010 46.330 178.270 ;
        RECT 53.830 178.210 54.150 178.270 ;
        RECT 62.110 178.210 62.430 178.270 ;
        RECT 63.505 178.210 63.795 178.255 ;
        RECT 71.770 178.210 72.090 178.270 ;
        RECT 72.245 178.210 72.535 178.255 ;
        RECT 46.560 178.070 54.150 178.210 ;
        RECT 27.165 177.870 27.455 177.915 ;
        RECT 29.565 177.870 29.855 177.915 ;
        RECT 32.805 177.870 33.455 177.915 ;
        RECT 46.560 177.870 46.700 178.070 ;
        RECT 53.830 178.010 54.150 178.070 ;
        RECT 54.840 178.070 61.880 178.210 ;
        RECT 52.450 177.870 52.770 177.930 ;
        RECT 27.165 177.730 33.455 177.870 ;
        RECT 27.165 177.685 27.455 177.730 ;
        RECT 29.565 177.685 30.155 177.730 ;
        RECT 32.805 177.685 33.455 177.730 ;
        RECT 43.340 177.730 46.700 177.870 ;
        RECT 47.480 177.730 52.770 177.870 ;
        RECT 26.245 177.530 26.535 177.575 ;
        RECT 26.705 177.530 26.995 177.575 ;
        RECT 26.245 177.390 26.995 177.530 ;
        RECT 26.245 177.345 26.535 177.390 ;
        RECT 26.705 177.345 26.995 177.390 ;
        RECT 29.865 177.370 30.155 177.685 ;
        RECT 43.340 177.575 43.480 177.730 ;
        RECT 30.945 177.530 31.235 177.575 ;
        RECT 34.525 177.530 34.815 177.575 ;
        RECT 36.360 177.530 36.650 177.575 ;
        RECT 30.945 177.390 36.650 177.530 ;
        RECT 30.945 177.345 31.235 177.390 ;
        RECT 34.525 177.345 34.815 177.390 ;
        RECT 36.360 177.345 36.650 177.390 ;
        RECT 43.265 177.530 43.555 177.575 ;
        RECT 43.710 177.530 44.030 177.590 ;
        RECT 43.265 177.390 44.030 177.530 ;
        RECT 43.265 177.345 43.555 177.390 ;
        RECT 26.780 177.190 26.920 177.345 ;
        RECT 43.710 177.330 44.030 177.390 ;
        RECT 45.550 177.530 45.870 177.590 ;
        RECT 47.480 177.575 47.620 177.730 ;
        RECT 52.450 177.670 52.770 177.730 ;
        RECT 46.485 177.530 46.775 177.575 ;
        RECT 45.550 177.390 46.775 177.530 ;
        RECT 45.550 177.330 45.870 177.390 ;
        RECT 46.485 177.345 46.775 177.390 ;
        RECT 47.405 177.345 47.695 177.575 ;
        RECT 30.370 177.190 30.690 177.250 ;
        RECT 26.780 177.050 30.690 177.190 ;
        RECT 30.370 176.990 30.690 177.050 ;
        RECT 35.430 176.990 35.750 177.250 ;
        RECT 36.810 176.990 37.130 177.250 ;
        RECT 38.190 176.990 38.510 177.250 ;
        RECT 39.125 177.005 39.415 177.235 ;
        RECT 30.945 176.850 31.235 176.895 ;
        RECT 34.065 176.850 34.355 176.895 ;
        RECT 35.955 176.850 36.245 176.895 ;
        RECT 30.945 176.710 36.245 176.850 ;
        RECT 30.945 176.665 31.235 176.710 ;
        RECT 34.065 176.665 34.355 176.710 ;
        RECT 35.955 176.665 36.245 176.710 ;
        RECT 28.070 176.310 28.390 176.570 ;
        RECT 34.510 176.510 34.830 176.570 ;
        RECT 39.200 176.510 39.340 177.005 ;
        RECT 46.560 176.850 46.700 177.345 ;
        RECT 47.850 177.330 48.170 177.590 ;
        RECT 48.325 177.530 48.615 177.575 ;
        RECT 49.230 177.530 49.550 177.590 ;
        RECT 48.325 177.390 49.550 177.530 ;
        RECT 48.325 177.345 48.615 177.390 ;
        RECT 49.230 177.330 49.550 177.390 ;
        RECT 50.610 177.330 50.930 177.590 ;
        RECT 49.320 177.190 49.460 177.330 ;
        RECT 54.840 177.190 54.980 178.070 ;
        RECT 55.325 177.870 55.615 177.915 ;
        RECT 56.130 177.870 56.450 177.930 ;
        RECT 58.565 177.870 59.215 177.915 ;
        RECT 55.325 177.730 59.215 177.870 ;
        RECT 55.325 177.685 55.915 177.730 ;
        RECT 55.625 177.370 55.915 177.685 ;
        RECT 56.130 177.670 56.450 177.730 ;
        RECT 58.565 177.685 59.215 177.730 ;
        RECT 61.190 177.670 61.510 177.930 ;
        RECT 61.740 177.870 61.880 178.070 ;
        RECT 62.110 178.070 63.795 178.210 ;
        RECT 62.110 178.010 62.430 178.070 ;
        RECT 63.505 178.025 63.795 178.070 ;
        RECT 70.480 178.070 72.535 178.210 ;
        RECT 70.480 177.870 70.620 178.070 ;
        RECT 71.770 178.010 72.090 178.070 ;
        RECT 72.245 178.025 72.535 178.070 ;
        RECT 73.150 178.010 73.470 178.270 ;
        RECT 81.890 178.210 82.210 178.270 ;
        RECT 81.520 178.070 82.210 178.210 ;
        RECT 61.740 177.730 70.620 177.870 ;
        RECT 79.590 177.870 79.910 177.930 ;
        RECT 80.065 177.870 80.355 177.915 ;
        RECT 81.520 177.870 81.660 178.070 ;
        RECT 81.890 178.010 82.210 178.070 ;
        RECT 82.350 178.210 82.670 178.270 ;
        RECT 88.345 178.210 88.635 178.255 ;
        RECT 90.630 178.210 90.950 178.270 ;
        RECT 82.350 178.070 88.100 178.210 ;
        RECT 82.350 178.010 82.670 178.070 ;
        RECT 86.030 177.870 86.350 177.930 ;
        RECT 79.590 177.730 80.355 177.870 ;
        RECT 79.590 177.670 79.910 177.730 ;
        RECT 80.065 177.685 80.355 177.730 ;
        RECT 80.600 177.730 81.660 177.870 ;
        RECT 56.705 177.530 56.995 177.575 ;
        RECT 60.285 177.530 60.575 177.575 ;
        RECT 62.120 177.530 62.410 177.575 ;
        RECT 56.705 177.390 62.410 177.530 ;
        RECT 56.705 177.345 56.995 177.390 ;
        RECT 60.285 177.345 60.575 177.390 ;
        RECT 62.120 177.345 62.410 177.390 ;
        RECT 64.425 177.345 64.715 177.575 ;
        RECT 49.320 177.050 54.980 177.190 ;
        RECT 59.350 177.190 59.670 177.250 ;
        RECT 62.585 177.190 62.875 177.235 ;
        RECT 63.950 177.190 64.270 177.250 ;
        RECT 59.350 177.050 64.270 177.190 ;
        RECT 59.350 176.990 59.670 177.050 ;
        RECT 62.585 177.005 62.875 177.050 ;
        RECT 63.950 176.990 64.270 177.050 ;
        RECT 51.070 176.850 51.390 176.910 ;
        RECT 46.560 176.710 51.390 176.850 ;
        RECT 51.070 176.650 51.390 176.710 ;
        RECT 56.705 176.850 56.995 176.895 ;
        RECT 59.825 176.850 60.115 176.895 ;
        RECT 61.715 176.850 62.005 176.895 ;
        RECT 56.705 176.710 62.005 176.850 ;
        RECT 56.705 176.665 56.995 176.710 ;
        RECT 59.825 176.665 60.115 176.710 ;
        RECT 61.715 176.665 62.005 176.710 ;
        RECT 34.510 176.370 39.340 176.510 ;
        RECT 41.425 176.510 41.715 176.555 ;
        RECT 42.790 176.510 43.110 176.570 ;
        RECT 41.425 176.370 43.110 176.510 ;
        RECT 34.510 176.310 34.830 176.370 ;
        RECT 41.425 176.325 41.715 176.370 ;
        RECT 42.790 176.310 43.110 176.370 ;
        RECT 49.705 176.510 49.995 176.555 ;
        RECT 50.150 176.510 50.470 176.570 ;
        RECT 49.705 176.370 50.470 176.510 ;
        RECT 49.705 176.325 49.995 176.370 ;
        RECT 50.150 176.310 50.470 176.370 ;
        RECT 53.385 176.510 53.675 176.555 ;
        RECT 64.500 176.510 64.640 177.345 ;
        RECT 69.010 177.330 69.330 177.590 ;
        RECT 69.470 177.530 69.790 177.590 ;
        RECT 71.360 177.530 71.650 177.575 ;
        RECT 72.690 177.530 73.010 177.590 ;
        RECT 73.625 177.530 73.915 177.575 ;
        RECT 69.470 177.390 72.460 177.530 ;
        RECT 69.470 177.330 69.790 177.390 ;
        RECT 71.360 177.345 71.650 177.390 ;
        RECT 72.320 177.190 72.460 177.390 ;
        RECT 72.690 177.390 73.915 177.530 ;
        RECT 72.690 177.330 73.010 177.390 ;
        RECT 73.625 177.345 73.915 177.390 ;
        RECT 74.070 177.330 74.390 177.590 ;
        RECT 74.990 177.330 75.310 177.590 ;
        RECT 75.465 177.345 75.755 177.575 ;
        RECT 75.540 177.190 75.680 177.345 ;
        RECT 76.370 177.330 76.690 177.590 ;
        RECT 77.305 177.345 77.595 177.575 ;
        RECT 72.320 177.050 75.680 177.190 ;
        RECT 77.380 177.190 77.520 177.345 ;
        RECT 77.750 177.330 78.070 177.590 ;
        RECT 78.210 177.530 78.530 177.590 ;
        RECT 80.600 177.530 80.740 177.730 ;
        RECT 81.520 177.575 81.660 177.730 ;
        RECT 82.440 177.730 86.350 177.870 ;
        RECT 87.960 177.870 88.100 178.070 ;
        RECT 88.345 178.070 90.950 178.210 ;
        RECT 88.345 178.025 88.635 178.070 ;
        RECT 90.630 178.010 90.950 178.070 ;
        RECT 99.830 178.210 100.150 178.270 ;
        RECT 102.145 178.210 102.435 178.255 ;
        RECT 99.830 178.070 102.435 178.210 ;
        RECT 99.830 178.010 100.150 178.070 ;
        RECT 102.145 178.025 102.435 178.070 ;
        RECT 111.790 178.010 112.110 178.270 ;
        RECT 112.250 178.010 112.570 178.270 ;
        RECT 114.105 178.025 114.395 178.255 ;
        RECT 117.785 178.210 118.075 178.255 ;
        RECT 118.690 178.210 119.010 178.270 ;
        RECT 117.785 178.070 119.010 178.210 ;
        RECT 117.785 178.025 118.075 178.070 ;
        RECT 109.030 177.870 109.350 177.930 ;
        RECT 87.960 177.730 106.960 177.870 ;
        RECT 78.210 177.390 80.740 177.530 ;
        RECT 78.210 177.330 78.530 177.390 ;
        RECT 81.445 177.345 81.735 177.575 ;
        RECT 81.890 177.330 82.210 177.590 ;
        RECT 82.440 177.575 82.580 177.730 ;
        RECT 86.030 177.670 86.350 177.730 ;
        RECT 82.365 177.345 82.655 177.575 ;
        RECT 82.810 177.530 83.130 177.590 ;
        RECT 83.285 177.530 83.575 177.575 ;
        RECT 84.190 177.530 84.510 177.590 ;
        RECT 82.810 177.390 84.510 177.530 ;
        RECT 82.810 177.330 83.130 177.390 ;
        RECT 83.285 177.345 83.575 177.390 ;
        RECT 84.190 177.330 84.510 177.390 ;
        RECT 85.585 177.530 85.875 177.575 ;
        RECT 89.250 177.530 89.570 177.590 ;
        RECT 85.585 177.390 89.570 177.530 ;
        RECT 85.585 177.345 85.875 177.390 ;
        RECT 89.250 177.330 89.570 177.390 ;
        RECT 98.450 177.330 98.770 177.590 ;
        RECT 99.370 177.330 99.690 177.590 ;
        RECT 99.920 177.575 100.060 177.730 ;
        RECT 106.820 177.590 106.960 177.730 ;
        RECT 107.280 177.730 109.350 177.870 ;
        RECT 114.180 177.870 114.320 178.025 ;
        RECT 118.690 178.010 119.010 178.070 ;
        RECT 121.910 177.870 122.230 177.930 ;
        RECT 114.180 177.730 122.230 177.870 ;
        RECT 99.845 177.345 100.135 177.575 ;
        RECT 100.305 177.345 100.595 177.575 ;
        RECT 102.130 177.530 102.450 177.590 ;
        RECT 103.065 177.530 103.355 177.575 ;
        RECT 102.130 177.390 103.355 177.530 ;
        RECT 79.130 177.190 79.450 177.250 ;
        RECT 77.380 177.050 79.450 177.190 ;
        RECT 79.130 176.990 79.450 177.050 ;
        RECT 79.605 177.190 79.895 177.235 ;
        RECT 80.510 177.190 80.830 177.250 ;
        RECT 100.380 177.190 100.520 177.345 ;
        RECT 102.130 177.330 102.450 177.390 ;
        RECT 103.065 177.345 103.355 177.390 ;
        RECT 106.285 177.345 106.575 177.575 ;
        RECT 105.810 177.190 106.130 177.250 ;
        RECT 106.360 177.190 106.500 177.345 ;
        RECT 106.730 177.330 107.050 177.590 ;
        RECT 107.280 177.575 107.420 177.730 ;
        RECT 109.030 177.670 109.350 177.730 ;
        RECT 121.910 177.670 122.230 177.730 ;
        RECT 107.205 177.345 107.495 177.575 ;
        RECT 108.110 177.530 108.430 177.590 ;
        RECT 109.490 177.530 109.810 177.590 ;
        RECT 108.110 177.390 109.810 177.530 ;
        RECT 108.110 177.330 108.430 177.390 ;
        RECT 109.490 177.330 109.810 177.390 ;
        RECT 116.850 177.330 117.170 177.590 ;
        RECT 79.605 177.050 80.830 177.190 ;
        RECT 79.605 177.005 79.895 177.050 ;
        RECT 80.510 176.990 80.830 177.050 ;
        RECT 84.970 177.050 106.500 177.190 ;
        RECT 65.330 176.850 65.650 176.910 ;
        RECT 70.405 176.850 70.695 176.895 ;
        RECT 84.970 176.850 85.110 177.050 ;
        RECT 105.810 176.990 106.130 177.050 ;
        RECT 110.870 176.990 111.190 177.250 ;
        RECT 65.330 176.710 85.110 176.850 ;
        RECT 65.330 176.650 65.650 176.710 ;
        RECT 70.405 176.665 70.695 176.710 ;
        RECT 53.385 176.370 64.640 176.510 ;
        RECT 64.870 176.510 65.190 176.570 ;
        RECT 68.090 176.510 68.410 176.570 ;
        RECT 64.870 176.370 68.410 176.510 ;
        RECT 53.385 176.325 53.675 176.370 ;
        RECT 64.870 176.310 65.190 176.370 ;
        RECT 68.090 176.310 68.410 176.370 ;
        RECT 69.010 176.510 69.330 176.570 ;
        RECT 74.990 176.510 75.310 176.570 ;
        RECT 69.010 176.370 75.310 176.510 ;
        RECT 69.010 176.310 69.330 176.370 ;
        RECT 74.990 176.310 75.310 176.370 ;
        RECT 100.750 176.510 101.070 176.570 ;
        RECT 101.685 176.510 101.975 176.555 ;
        RECT 100.750 176.370 101.975 176.510 ;
        RECT 100.750 176.310 101.070 176.370 ;
        RECT 101.685 176.325 101.975 176.370 ;
        RECT 102.130 176.510 102.450 176.570 ;
        RECT 104.905 176.510 105.195 176.555 ;
        RECT 102.130 176.370 105.195 176.510 ;
        RECT 102.130 176.310 102.450 176.370 ;
        RECT 104.905 176.325 105.195 176.370 ;
        RECT 14.660 175.690 127.820 176.170 ;
        RECT 25.785 175.490 26.075 175.535 ;
        RECT 26.230 175.490 26.550 175.550 ;
        RECT 38.190 175.490 38.510 175.550 ;
        RECT 40.950 175.490 41.270 175.550 ;
        RECT 25.785 175.350 26.550 175.490 ;
        RECT 25.785 175.305 26.075 175.350 ;
        RECT 26.230 175.290 26.550 175.350 ;
        RECT 34.140 175.350 38.510 175.490 ;
        RECT 30.845 175.150 31.135 175.195 ;
        RECT 26.780 175.010 31.135 175.150 ;
        RECT 26.780 174.515 26.920 175.010 ;
        RECT 30.845 174.965 31.135 175.010 ;
        RECT 34.140 174.855 34.280 175.350 ;
        RECT 38.190 175.290 38.510 175.350 ;
        RECT 38.740 175.350 41.270 175.490 ;
        RECT 38.740 175.150 38.880 175.350 ;
        RECT 40.950 175.290 41.270 175.350 ;
        RECT 46.470 175.490 46.790 175.550 ;
        RECT 54.290 175.490 54.610 175.550 ;
        RECT 46.470 175.350 54.610 175.490 ;
        RECT 46.470 175.290 46.790 175.350 ;
        RECT 54.290 175.290 54.610 175.350 ;
        RECT 63.950 175.490 64.270 175.550 ;
        RECT 66.250 175.490 66.570 175.550 ;
        RECT 63.950 175.350 66.570 175.490 ;
        RECT 63.950 175.290 64.270 175.350 ;
        RECT 66.250 175.290 66.570 175.350 ;
        RECT 68.090 175.490 68.410 175.550 ;
        RECT 77.750 175.490 78.070 175.550 ;
        RECT 81.890 175.490 82.210 175.550 ;
        RECT 106.270 175.490 106.590 175.550 ;
        RECT 108.110 175.490 108.430 175.550 ;
        RECT 68.090 175.350 82.210 175.490 ;
        RECT 68.090 175.290 68.410 175.350 ;
        RECT 77.750 175.290 78.070 175.350 ;
        RECT 81.890 175.290 82.210 175.350 ;
        RECT 104.060 175.350 110.640 175.490 ;
        RECT 36.900 175.010 38.880 175.150 ;
        RECT 39.125 175.150 39.415 175.195 ;
        RECT 40.490 175.150 40.810 175.210 ;
        RECT 57.525 175.150 57.815 175.195 ;
        RECT 39.125 175.010 40.810 175.150 ;
        RECT 34.065 174.625 34.355 174.855 ;
        RECT 36.900 174.810 37.040 175.010 ;
        RECT 39.125 174.965 39.415 175.010 ;
        RECT 40.490 174.950 40.810 175.010 ;
        RECT 53.920 175.010 57.815 175.150 ;
        RECT 53.920 174.870 54.060 175.010 ;
        RECT 57.525 174.965 57.815 175.010 ;
        RECT 60.385 175.150 60.675 175.195 ;
        RECT 63.505 175.150 63.795 175.195 ;
        RECT 65.395 175.150 65.685 175.195 ;
        RECT 71.785 175.150 72.075 175.195 ;
        RECT 76.370 175.150 76.690 175.210 ;
        RECT 60.385 175.010 65.685 175.150 ;
        RECT 60.385 174.965 60.675 175.010 ;
        RECT 63.505 174.965 63.795 175.010 ;
        RECT 65.395 174.965 65.685 175.010 ;
        RECT 69.560 175.010 76.690 175.150 ;
        RECT 35.520 174.670 37.040 174.810 ;
        RECT 37.730 174.810 38.050 174.870 ;
        RECT 45.550 174.810 45.870 174.870 ;
        RECT 37.730 174.670 41.640 174.810 ;
        RECT 26.705 174.285 26.995 174.515 ;
        RECT 27.165 174.285 27.455 174.515 ;
        RECT 30.385 174.470 30.675 174.515 ;
        RECT 32.685 174.470 32.975 174.515 ;
        RECT 34.510 174.470 34.830 174.530 ;
        RECT 35.520 174.515 35.660 174.670 ;
        RECT 37.730 174.610 38.050 174.670 ;
        RECT 30.385 174.330 34.830 174.470 ;
        RECT 30.385 174.285 30.675 174.330 ;
        RECT 32.685 174.285 32.975 174.330 ;
        RECT 27.240 174.130 27.380 174.285 ;
        RECT 34.510 174.270 34.830 174.330 ;
        RECT 35.445 174.285 35.735 174.515 ;
        RECT 36.365 174.285 36.655 174.515 ;
        RECT 36.825 174.285 37.115 174.515 ;
        RECT 37.285 174.470 37.575 174.515 ;
        RECT 38.190 174.470 38.510 174.530 ;
        RECT 40.030 174.470 40.350 174.530 ;
        RECT 41.500 174.515 41.640 174.670 ;
        RECT 42.880 174.670 45.870 174.810 ;
        RECT 42.880 174.515 43.020 174.670 ;
        RECT 45.550 174.610 45.870 174.670 ;
        RECT 46.945 174.810 47.235 174.855 ;
        RECT 53.830 174.810 54.150 174.870 ;
        RECT 46.945 174.670 54.150 174.810 ;
        RECT 46.945 174.625 47.235 174.670 ;
        RECT 53.830 174.610 54.150 174.670 ;
        RECT 54.290 174.610 54.610 174.870 ;
        RECT 57.970 174.810 58.290 174.870 ;
        RECT 64.870 174.810 65.190 174.870 ;
        RECT 54.840 174.670 58.290 174.810 ;
        RECT 40.505 174.470 40.795 174.515 ;
        RECT 37.285 174.330 40.795 174.470 ;
        RECT 37.285 174.285 37.575 174.330 ;
        RECT 28.070 174.130 28.390 174.190 ;
        RECT 33.145 174.130 33.435 174.175 ;
        RECT 34.050 174.130 34.370 174.190 ;
        RECT 36.440 174.130 36.580 174.285 ;
        RECT 27.240 173.990 32.900 174.130 ;
        RECT 28.070 173.930 28.390 173.990 ;
        RECT 32.760 173.790 32.900 173.990 ;
        RECT 33.145 173.990 34.370 174.130 ;
        RECT 33.145 173.945 33.435 173.990 ;
        RECT 34.050 173.930 34.370 173.990 ;
        RECT 34.600 173.990 36.580 174.130 ;
        RECT 34.600 173.790 34.740 173.990 ;
        RECT 32.760 173.650 34.740 173.790 ;
        RECT 36.900 173.790 37.040 174.285 ;
        RECT 38.190 174.270 38.510 174.330 ;
        RECT 40.030 174.270 40.350 174.330 ;
        RECT 40.505 174.285 40.795 174.330 ;
        RECT 40.965 174.285 41.255 174.515 ;
        RECT 41.425 174.285 41.715 174.515 ;
        RECT 42.345 174.470 42.635 174.515 ;
        RECT 42.805 174.470 43.095 174.515 ;
        RECT 42.345 174.330 43.095 174.470 ;
        RECT 42.345 174.285 42.635 174.330 ;
        RECT 42.805 174.285 43.095 174.330 ;
        RECT 38.665 174.130 38.955 174.175 ;
        RECT 39.110 174.130 39.430 174.190 ;
        RECT 38.665 173.990 39.430 174.130 ;
        RECT 38.665 173.945 38.955 173.990 ;
        RECT 39.110 173.930 39.430 173.990 ;
        RECT 39.570 174.130 39.890 174.190 ;
        RECT 41.040 174.130 41.180 174.285 ;
        RECT 43.710 174.270 44.030 174.530 ;
        RECT 44.170 174.270 44.490 174.530 ;
        RECT 44.630 174.270 44.950 174.530 ;
        RECT 54.840 174.515 54.980 174.670 ;
        RECT 57.970 174.610 58.290 174.670 ;
        RECT 58.520 174.670 65.190 174.810 ;
        RECT 49.705 174.470 49.995 174.515 ;
        RECT 54.765 174.470 55.055 174.515 ;
        RECT 49.705 174.330 55.055 174.470 ;
        RECT 49.705 174.285 49.995 174.330 ;
        RECT 54.765 174.285 55.055 174.330 ;
        RECT 55.225 174.470 55.515 174.515 ;
        RECT 56.590 174.470 56.910 174.530 ;
        RECT 55.225 174.330 56.910 174.470 ;
        RECT 55.225 174.285 55.515 174.330 ;
        RECT 56.590 174.270 56.910 174.330 ;
        RECT 41.870 174.130 42.190 174.190 ;
        RECT 39.570 173.990 42.190 174.130 ;
        RECT 39.570 173.930 39.890 173.990 ;
        RECT 41.870 173.930 42.190 173.990 ;
        RECT 39.660 173.790 39.800 173.930 ;
        RECT 36.900 173.650 39.800 173.790 ;
        RECT 44.260 173.790 44.400 174.270 ;
        RECT 45.550 174.130 45.870 174.190 ;
        RECT 46.025 174.130 46.315 174.175 ;
        RECT 45.550 173.990 46.315 174.130 ;
        RECT 45.550 173.930 45.870 173.990 ;
        RECT 46.025 173.945 46.315 173.990 ;
        RECT 47.850 174.130 48.170 174.190 ;
        RECT 53.370 174.130 53.690 174.190 ;
        RECT 58.520 174.130 58.660 174.670 ;
        RECT 64.870 174.610 65.190 174.670 ;
        RECT 66.250 174.610 66.570 174.870 ;
        RECT 59.305 174.175 59.595 174.490 ;
        RECT 60.385 174.470 60.675 174.515 ;
        RECT 63.965 174.470 64.255 174.515 ;
        RECT 65.800 174.470 66.090 174.515 ;
        RECT 60.385 174.330 66.090 174.470 ;
        RECT 60.385 174.285 60.675 174.330 ;
        RECT 63.965 174.285 64.255 174.330 ;
        RECT 65.800 174.285 66.090 174.330 ;
        RECT 68.565 174.470 68.855 174.515 ;
        RECT 69.010 174.470 69.330 174.530 ;
        RECT 68.565 174.330 69.330 174.470 ;
        RECT 68.565 174.285 68.855 174.330 ;
        RECT 69.010 174.270 69.330 174.330 ;
        RECT 47.850 173.990 58.660 174.130 ;
        RECT 59.005 174.130 59.595 174.175 ;
        RECT 61.190 174.130 61.510 174.190 ;
        RECT 62.245 174.130 62.895 174.175 ;
        RECT 59.005 173.990 62.895 174.130 ;
        RECT 47.850 173.930 48.170 173.990 ;
        RECT 53.370 173.930 53.690 173.990 ;
        RECT 59.005 173.945 59.295 173.990 ;
        RECT 61.190 173.930 61.510 173.990 ;
        RECT 62.245 173.945 62.895 173.990 ;
        RECT 64.870 173.930 65.190 174.190 ;
        RECT 69.560 174.130 69.700 175.010 ;
        RECT 71.785 174.965 72.075 175.010 ;
        RECT 76.370 174.950 76.690 175.010 ;
        RECT 69.930 174.610 70.250 174.870 ;
        RECT 81.980 174.810 82.120 175.290 ;
        RECT 87.410 174.810 87.730 174.870 ;
        RECT 81.980 174.670 83.040 174.810 ;
        RECT 72.690 174.270 73.010 174.530 ;
        RECT 78.210 174.470 78.530 174.530 ;
        RECT 82.900 174.515 83.040 174.670 ;
        RECT 83.360 174.670 87.730 174.810 ;
        RECT 83.360 174.515 83.500 174.670 ;
        RECT 87.410 174.610 87.730 174.670 ;
        RECT 82.365 174.470 82.655 174.515 ;
        RECT 78.210 174.330 82.655 174.470 ;
        RECT 78.210 174.270 78.530 174.330 ;
        RECT 82.365 174.285 82.655 174.330 ;
        RECT 82.825 174.285 83.115 174.515 ;
        RECT 83.285 174.285 83.575 174.515 ;
        RECT 84.190 174.270 84.510 174.530 ;
        RECT 98.450 174.470 98.770 174.530 ;
        RECT 104.060 174.515 104.200 175.350 ;
        RECT 106.270 175.290 106.590 175.350 ;
        RECT 108.110 175.290 108.430 175.350 ;
        RECT 107.205 175.150 107.495 175.195 ;
        RECT 109.030 175.150 109.350 175.210 ;
        RECT 107.205 175.010 109.350 175.150 ;
        RECT 107.205 174.965 107.495 175.010 ;
        RECT 109.030 174.950 109.350 175.010 ;
        RECT 106.730 174.810 107.050 174.870 ;
        RECT 105.440 174.670 109.720 174.810 ;
        RECT 103.985 174.470 104.275 174.515 ;
        RECT 98.450 174.330 104.275 174.470 ;
        RECT 98.450 174.270 98.770 174.330 ;
        RECT 103.985 174.285 104.275 174.330 ;
        RECT 104.890 174.270 105.210 174.530 ;
        RECT 105.440 174.515 105.580 174.670 ;
        RECT 106.730 174.610 107.050 174.670 ;
        RECT 109.580 174.530 109.720 174.670 ;
        RECT 105.365 174.285 105.655 174.515 ;
        RECT 105.810 174.470 106.130 174.530 ;
        RECT 109.045 174.470 109.335 174.515 ;
        RECT 105.810 174.330 109.335 174.470 ;
        RECT 105.810 174.270 106.130 174.330 ;
        RECT 109.045 174.285 109.335 174.330 ;
        RECT 65.420 173.990 69.700 174.130 ;
        RECT 80.985 174.130 81.275 174.175 ;
        RECT 81.890 174.130 82.210 174.190 ;
        RECT 80.985 173.990 82.210 174.130 ;
        RECT 47.940 173.790 48.080 173.930 ;
        RECT 44.260 173.650 48.080 173.790 ;
        RECT 57.050 173.590 57.370 173.850 ;
        RECT 63.030 173.790 63.350 173.850 ;
        RECT 65.420 173.790 65.560 173.990 ;
        RECT 80.985 173.945 81.275 173.990 ;
        RECT 81.890 173.930 82.210 173.990 ;
        RECT 104.430 174.130 104.750 174.190 ;
        RECT 107.665 174.130 107.955 174.175 ;
        RECT 104.430 173.990 107.955 174.130 ;
        RECT 104.430 173.930 104.750 173.990 ;
        RECT 107.665 173.945 107.955 173.990 ;
        RECT 63.030 173.650 65.560 173.790 ;
        RECT 70.850 173.790 71.170 173.850 ;
        RECT 98.450 173.790 98.770 173.850 ;
        RECT 70.850 173.650 98.770 173.790 ;
        RECT 109.120 173.790 109.260 174.285 ;
        RECT 109.490 174.270 109.810 174.530 ;
        RECT 109.950 174.270 110.270 174.530 ;
        RECT 110.500 174.470 110.640 175.350 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 110.885 174.470 111.175 174.515 ;
        RECT 110.500 174.330 111.175 174.470 ;
        RECT 110.885 174.285 111.175 174.330 ;
        RECT 118.245 174.470 118.535 174.515 ;
        RECT 119.150 174.470 119.470 174.530 ;
        RECT 118.245 174.330 119.470 174.470 ;
        RECT 118.245 174.285 118.535 174.330 ;
        RECT 119.150 174.270 119.470 174.330 ;
        RECT 118.705 173.945 118.995 174.175 ;
        RECT 109.950 173.790 110.270 173.850 ;
        RECT 109.120 173.650 110.270 173.790 ;
        RECT 63.030 173.590 63.350 173.650 ;
        RECT 70.850 173.590 71.170 173.650 ;
        RECT 98.450 173.590 98.770 173.650 ;
        RECT 109.950 173.590 110.270 173.650 ;
        RECT 118.230 173.790 118.550 173.850 ;
        RECT 118.780 173.790 118.920 173.945 ;
        RECT 118.230 173.650 118.920 173.790 ;
        RECT 118.230 173.590 118.550 173.650 ;
        RECT 14.660 172.970 127.820 173.450 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 35.430 172.770 35.750 172.830 ;
        RECT 41.885 172.770 42.175 172.815 ;
        RECT 35.430 172.630 42.175 172.770 ;
        RECT 35.430 172.570 35.750 172.630 ;
        RECT 41.885 172.585 42.175 172.630 ;
        RECT 44.630 172.770 44.950 172.830 ;
        RECT 49.230 172.770 49.550 172.830 ;
        RECT 44.630 172.630 49.550 172.770 ;
        RECT 44.630 172.570 44.950 172.630 ;
        RECT 37.270 172.430 37.590 172.490 ;
        RECT 37.270 172.290 40.260 172.430 ;
        RECT 37.270 172.230 37.590 172.290 ;
        RECT 38.190 172.090 38.510 172.150 ;
        RECT 39.125 172.090 39.415 172.135 ;
        RECT 38.190 171.950 39.415 172.090 ;
        RECT 38.190 171.890 38.510 171.950 ;
        RECT 39.125 171.905 39.415 171.950 ;
        RECT 39.570 171.890 39.890 172.150 ;
        RECT 40.120 172.135 40.260 172.290 ;
        RECT 40.045 171.905 40.335 172.135 ;
        RECT 40.950 171.890 41.270 172.150 ;
        RECT 42.790 171.890 43.110 172.150 ;
        RECT 45.640 172.135 45.780 172.630 ;
        RECT 49.230 172.570 49.550 172.630 ;
        RECT 49.690 172.770 50.010 172.830 ;
        RECT 51.070 172.770 51.390 172.830 ;
        RECT 54.750 172.770 55.070 172.830 ;
        RECT 49.690 172.630 50.380 172.770 ;
        RECT 49.690 172.570 50.010 172.630 ;
        RECT 46.100 172.290 49.920 172.430 ;
        RECT 46.100 172.135 46.240 172.290 ;
        RECT 49.780 172.150 49.920 172.290 ;
        RECT 45.565 171.905 45.855 172.135 ;
        RECT 46.025 171.905 46.315 172.135 ;
        RECT 46.485 171.905 46.775 172.135 ;
        RECT 35.890 171.750 36.210 171.810 ;
        RECT 46.560 171.750 46.700 171.905 ;
        RECT 47.390 171.890 47.710 172.150 ;
        RECT 49.230 171.890 49.550 172.150 ;
        RECT 49.690 171.890 50.010 172.150 ;
        RECT 50.240 172.135 50.380 172.630 ;
        RECT 51.070 172.630 55.070 172.770 ;
        RECT 51.070 172.570 51.390 172.630 ;
        RECT 54.750 172.570 55.070 172.630 ;
        RECT 60.745 172.770 61.035 172.815 ;
        RECT 61.190 172.770 61.510 172.830 ;
        RECT 60.745 172.630 61.510 172.770 ;
        RECT 60.745 172.585 61.035 172.630 ;
        RECT 61.190 172.570 61.510 172.630 ;
        RECT 62.585 172.770 62.875 172.815 ;
        RECT 64.870 172.770 65.190 172.830 ;
        RECT 91.090 172.770 91.410 172.830 ;
        RECT 119.150 172.770 119.470 172.830 ;
        RECT 62.585 172.630 65.190 172.770 ;
        RECT 62.585 172.585 62.875 172.630 ;
        RECT 64.870 172.570 65.190 172.630 ;
        RECT 89.800 172.630 100.060 172.770 ;
        RECT 57.050 172.430 57.370 172.490 ;
        RECT 83.745 172.430 84.035 172.475 ;
        RECT 89.800 172.430 89.940 172.630 ;
        RECT 91.090 172.570 91.410 172.630 ;
        RECT 57.050 172.290 61.880 172.430 ;
        RECT 57.050 172.230 57.370 172.290 ;
        RECT 50.165 171.905 50.455 172.135 ;
        RECT 51.070 171.890 51.390 172.150 ;
        RECT 52.925 171.905 53.215 172.135 ;
        RECT 35.890 171.610 46.700 171.750 ;
        RECT 49.320 171.750 49.460 171.890 ;
        RECT 53.000 171.750 53.140 171.905 ;
        RECT 53.370 171.890 53.690 172.150 ;
        RECT 53.830 171.890 54.150 172.150 ;
        RECT 54.750 171.890 55.070 172.150 ;
        RECT 60.730 172.090 61.050 172.150 ;
        RECT 61.740 172.135 61.880 172.290 ;
        RECT 83.745 172.290 89.940 172.430 ;
        RECT 83.745 172.245 84.035 172.290 ;
        RECT 61.205 172.090 61.495 172.135 ;
        RECT 60.730 171.950 61.495 172.090 ;
        RECT 60.730 171.890 61.050 171.950 ;
        RECT 61.205 171.905 61.495 171.950 ;
        RECT 61.665 171.905 61.955 172.135 ;
        RECT 69.010 172.090 69.330 172.150 ;
        RECT 89.800 172.135 89.940 172.290 ;
        RECT 90.185 172.430 90.475 172.475 ;
        RECT 92.585 172.430 92.875 172.475 ;
        RECT 95.825 172.430 96.475 172.475 ;
        RECT 90.185 172.290 96.475 172.430 ;
        RECT 90.185 172.245 90.475 172.290 ;
        RECT 92.585 172.245 93.175 172.290 ;
        RECT 95.825 172.245 96.475 172.290 ;
        RECT 82.365 172.090 82.655 172.135 ;
        RECT 69.010 171.950 82.655 172.090 ;
        RECT 69.010 171.890 69.330 171.950 ;
        RECT 82.365 171.905 82.655 171.950 ;
        RECT 89.725 171.905 90.015 172.135 ;
        RECT 92.885 171.930 93.175 172.245 ;
        RECT 93.965 172.090 94.255 172.135 ;
        RECT 97.545 172.090 97.835 172.135 ;
        RECT 99.380 172.090 99.670 172.135 ;
        RECT 93.965 171.950 99.670 172.090 ;
        RECT 99.920 172.090 100.060 172.630 ;
        RECT 113.260 172.630 119.470 172.770 ;
        RECT 106.270 172.430 106.590 172.490 ;
        RECT 110.410 172.430 110.730 172.490 ;
        RECT 106.270 172.290 108.340 172.430 ;
        RECT 106.270 172.230 106.590 172.290 ;
        RECT 108.200 172.135 108.340 172.290 ;
        RECT 109.120 172.290 110.730 172.430 ;
        RECT 109.120 172.135 109.260 172.290 ;
        RECT 110.410 172.230 110.730 172.290 ;
        RECT 107.665 172.090 107.955 172.135 ;
        RECT 99.920 171.950 107.955 172.090 ;
        RECT 93.965 171.905 94.255 171.950 ;
        RECT 97.545 171.905 97.835 171.950 ;
        RECT 99.380 171.905 99.670 171.950 ;
        RECT 107.665 171.905 107.955 171.950 ;
        RECT 108.125 171.905 108.415 172.135 ;
        RECT 109.045 171.905 109.335 172.135 ;
        RECT 49.320 171.610 53.140 171.750 ;
        RECT 35.890 171.550 36.210 171.610 ;
        RECT 49.690 171.410 50.010 171.470 ;
        RECT 53.460 171.410 53.600 171.890 ;
        RECT 85.585 171.750 85.875 171.795 ;
        RECT 85.585 171.610 91.320 171.750 ;
        RECT 85.585 171.565 85.875 171.610 ;
        RECT 49.690 171.270 53.600 171.410 ;
        RECT 49.690 171.210 50.010 171.270 ;
        RECT 35.430 171.070 35.750 171.130 ;
        RECT 37.745 171.070 38.035 171.115 ;
        RECT 35.430 170.930 38.035 171.070 ;
        RECT 35.430 170.870 35.750 170.930 ;
        RECT 37.745 170.885 38.035 170.930 ;
        RECT 41.410 171.070 41.730 171.130 ;
        RECT 44.185 171.070 44.475 171.115 ;
        RECT 41.410 170.930 44.475 171.070 ;
        RECT 41.410 170.870 41.730 170.930 ;
        RECT 44.185 170.885 44.475 170.930 ;
        RECT 46.010 171.070 46.330 171.130 ;
        RECT 47.865 171.070 48.155 171.115 ;
        RECT 46.010 170.930 48.155 171.070 ;
        RECT 46.010 170.870 46.330 170.930 ;
        RECT 47.865 170.885 48.155 170.930 ;
        RECT 51.545 171.070 51.835 171.115 ;
        RECT 52.450 171.070 52.770 171.130 ;
        RECT 51.545 170.930 52.770 171.070 ;
        RECT 51.545 170.885 51.835 170.930 ;
        RECT 52.450 170.870 52.770 170.930 ;
        RECT 88.345 171.070 88.635 171.115 ;
        RECT 89.710 171.070 90.030 171.130 ;
        RECT 91.180 171.115 91.320 171.610 ;
        RECT 98.450 171.550 98.770 171.810 ;
        RECT 99.845 171.750 100.135 171.795 ;
        RECT 105.810 171.750 106.130 171.810 ;
        RECT 99.845 171.610 106.130 171.750 ;
        RECT 107.740 171.750 107.880 171.905 ;
        RECT 109.490 171.890 109.810 172.150 ;
        RECT 109.950 171.890 110.270 172.150 ;
        RECT 113.260 172.135 113.400 172.630 ;
        RECT 119.150 172.570 119.470 172.630 ;
        RECT 117.425 172.430 117.715 172.475 ;
        RECT 118.230 172.430 118.550 172.490 ;
        RECT 120.665 172.430 121.315 172.475 ;
        RECT 117.425 172.290 121.315 172.430 ;
        RECT 117.425 172.245 118.015 172.290 ;
        RECT 113.185 171.905 113.475 172.135 ;
        RECT 117.725 171.930 118.015 172.245 ;
        RECT 118.230 172.230 118.550 172.290 ;
        RECT 120.665 172.245 121.315 172.290 ;
        RECT 118.805 172.090 119.095 172.135 ;
        RECT 122.385 172.090 122.675 172.135 ;
        RECT 124.220 172.090 124.510 172.135 ;
        RECT 118.805 171.950 124.510 172.090 ;
        RECT 133.500 172.050 136.690 172.190 ;
        RECT 118.805 171.905 119.095 171.950 ;
        RECT 122.385 171.905 122.675 171.950 ;
        RECT 124.220 171.905 124.510 171.950 ;
        RECT 129.260 171.930 136.690 172.050 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 113.260 171.750 113.400 171.905 ;
        RECT 107.740 171.610 113.400 171.750 ;
        RECT 121.450 171.750 121.770 171.810 ;
        RECT 123.305 171.750 123.595 171.795 ;
        RECT 121.450 171.610 123.595 171.750 ;
        RECT 99.845 171.565 100.135 171.610 ;
        RECT 105.810 171.550 106.130 171.610 ;
        RECT 121.450 171.550 121.770 171.610 ;
        RECT 123.305 171.565 123.595 171.610 ;
        RECT 124.670 171.550 124.990 171.810 ;
        RECT 93.965 171.410 94.255 171.455 ;
        RECT 97.085 171.410 97.375 171.455 ;
        RECT 98.975 171.410 99.265 171.455 ;
        RECT 114.550 171.410 114.870 171.470 ;
        RECT 93.965 171.270 99.265 171.410 ;
        RECT 93.965 171.225 94.255 171.270 ;
        RECT 97.085 171.225 97.375 171.270 ;
        RECT 98.975 171.225 99.265 171.270 ;
        RECT 99.920 171.270 114.870 171.410 ;
        RECT 88.345 170.930 90.030 171.070 ;
        RECT 88.345 170.885 88.635 170.930 ;
        RECT 89.710 170.870 90.030 170.930 ;
        RECT 91.105 171.070 91.395 171.115 ;
        RECT 99.920 171.070 100.060 171.270 ;
        RECT 114.550 171.210 114.870 171.270 ;
        RECT 118.805 171.410 119.095 171.455 ;
        RECT 121.925 171.410 122.215 171.455 ;
        RECT 123.815 171.410 124.105 171.455 ;
        RECT 118.805 171.270 124.105 171.410 ;
        RECT 118.805 171.225 119.095 171.270 ;
        RECT 121.925 171.225 122.215 171.270 ;
        RECT 123.815 171.225 124.105 171.270 ;
        RECT 91.105 170.930 100.060 171.070 ;
        RECT 91.105 170.885 91.395 170.930 ;
        RECT 107.190 170.870 107.510 171.130 ;
        RECT 111.330 170.870 111.650 171.130 ;
        RECT 113.630 170.870 113.950 171.130 ;
        RECT 115.945 171.070 116.235 171.115 ;
        RECT 117.310 171.070 117.630 171.130 ;
        RECT 115.945 170.930 117.630 171.070 ;
        RECT 115.945 170.885 116.235 170.930 ;
        RECT 117.310 170.870 117.630 170.930 ;
        RECT 129.260 170.790 139.470 171.930 ;
        RECT 14.660 170.250 127.820 170.730 ;
        RECT 133.500 170.600 136.690 170.790 ;
        RECT 47.390 170.050 47.710 170.110 ;
        RECT 67.630 170.050 67.950 170.110 ;
        RECT 69.025 170.050 69.315 170.095 ;
        RECT 47.390 169.910 69.315 170.050 ;
        RECT 47.390 169.850 47.710 169.910 ;
        RECT 67.630 169.850 67.950 169.910 ;
        RECT 69.025 169.865 69.315 169.910 ;
        RECT 70.850 169.850 71.170 170.110 ;
        RECT 97.085 170.050 97.375 170.095 ;
        RECT 98.450 170.050 98.770 170.110 ;
        RECT 97.085 169.910 98.770 170.050 ;
        RECT 97.085 169.865 97.375 169.910 ;
        RECT 98.450 169.850 98.770 169.910 ;
        RECT 121.450 169.850 121.770 170.110 ;
        RECT 40.950 169.710 41.270 169.770 ;
        RECT 70.940 169.710 71.080 169.850 ;
        RECT 40.950 169.570 71.080 169.710 ;
        RECT 84.620 169.710 84.910 169.755 ;
        RECT 87.400 169.710 87.690 169.755 ;
        RECT 89.260 169.710 89.550 169.755 ;
        RECT 84.620 169.570 89.550 169.710 ;
        RECT 40.950 169.510 41.270 169.570 ;
        RECT 84.620 169.525 84.910 169.570 ;
        RECT 87.400 169.525 87.690 169.570 ;
        RECT 89.260 169.525 89.550 169.570 ;
        RECT 89.710 169.710 90.030 169.770 ;
        RECT 89.710 169.570 93.160 169.710 ;
        RECT 89.710 169.510 90.030 169.570 ;
        RECT 77.305 169.370 77.595 169.415 ;
        RECT 80.050 169.370 80.370 169.430 ;
        RECT 77.305 169.230 80.370 169.370 ;
        RECT 77.305 169.185 77.595 169.230 ;
        RECT 80.050 169.170 80.370 169.230 ;
        RECT 81.980 169.230 91.780 169.370 ;
        RECT 27.165 169.030 27.455 169.075 ;
        RECT 30.370 169.030 30.690 169.090 ;
        RECT 33.605 169.030 33.895 169.075 ;
        RECT 35.890 169.030 36.210 169.090 ;
        RECT 27.165 168.890 36.210 169.030 ;
        RECT 27.165 168.845 27.455 168.890 ;
        RECT 30.370 168.830 30.690 168.890 ;
        RECT 33.605 168.845 33.895 168.890 ;
        RECT 35.890 168.830 36.210 168.890 ;
        RECT 44.170 168.830 44.490 169.090 ;
        RECT 69.945 169.030 70.235 169.075 ;
        RECT 70.390 169.030 70.710 169.090 ;
        RECT 71.785 169.030 72.075 169.075 ;
        RECT 69.945 168.890 72.075 169.030 ;
        RECT 69.945 168.845 70.235 168.890 ;
        RECT 70.390 168.830 70.710 168.890 ;
        RECT 71.785 168.845 72.075 168.890 ;
        RECT 80.755 168.690 81.045 168.735 ;
        RECT 81.980 168.690 82.120 169.230 ;
        RECT 84.620 169.030 84.910 169.075 ;
        RECT 84.620 168.890 87.155 169.030 ;
        RECT 84.620 168.845 84.910 168.890 ;
        RECT 77.840 168.550 82.120 168.690 ;
        RECT 82.760 168.690 83.050 168.735 ;
        RECT 84.190 168.690 84.510 168.750 ;
        RECT 86.940 168.735 87.155 168.890 ;
        RECT 87.870 168.830 88.190 169.090 ;
        RECT 89.725 169.030 90.015 169.075 ;
        RECT 91.090 169.030 91.410 169.090 ;
        RECT 89.725 168.890 91.410 169.030 ;
        RECT 91.640 169.030 91.780 169.230 ;
        RECT 92.010 169.170 92.330 169.430 ;
        RECT 93.020 169.415 93.160 169.570 ;
        RECT 95.245 169.525 95.535 169.755 ;
        RECT 105.925 169.710 106.215 169.755 ;
        RECT 109.045 169.710 109.335 169.755 ;
        RECT 110.935 169.710 111.225 169.755 ;
        RECT 105.925 169.570 111.225 169.710 ;
        RECT 105.925 169.525 106.215 169.570 ;
        RECT 109.045 169.525 109.335 169.570 ;
        RECT 110.935 169.525 111.225 169.570 ;
        RECT 92.945 169.185 93.235 169.415 ;
        RECT 93.405 169.030 93.695 169.075 ;
        RECT 91.640 168.890 93.695 169.030 ;
        RECT 95.320 169.030 95.460 169.525 ;
        RECT 109.950 169.370 110.270 169.430 ;
        RECT 110.425 169.370 110.715 169.415 ;
        RECT 109.950 169.230 110.715 169.370 ;
        RECT 109.950 169.170 110.270 169.230 ;
        RECT 110.425 169.185 110.715 169.230 ;
        RECT 112.710 169.370 113.030 169.430 ;
        RECT 115.485 169.370 115.775 169.415 ;
        RECT 112.710 169.230 115.775 169.370 ;
        RECT 112.710 169.170 113.030 169.230 ;
        RECT 115.485 169.185 115.775 169.230 ;
        RECT 117.310 169.370 117.630 169.430 ;
        RECT 119.625 169.370 119.915 169.415 ;
        RECT 117.310 169.230 119.915 169.370 ;
        RECT 117.310 169.170 117.630 169.230 ;
        RECT 119.625 169.185 119.915 169.230 ;
        RECT 96.165 169.030 96.455 169.075 ;
        RECT 95.320 168.890 96.455 169.030 ;
        RECT 89.725 168.845 90.015 168.890 ;
        RECT 91.090 168.830 91.410 168.890 ;
        RECT 93.405 168.845 93.695 168.890 ;
        RECT 96.165 168.845 96.455 168.890 ;
        RECT 104.845 168.735 105.135 169.050 ;
        RECT 105.925 169.030 106.215 169.075 ;
        RECT 109.505 169.030 109.795 169.075 ;
        RECT 111.340 169.030 111.630 169.075 ;
        RECT 105.925 168.890 111.630 169.030 ;
        RECT 105.925 168.845 106.215 168.890 ;
        RECT 109.505 168.845 109.795 168.890 ;
        RECT 111.340 168.845 111.630 168.890 ;
        RECT 111.790 168.830 112.110 169.090 ;
        RECT 114.550 168.830 114.870 169.090 ;
        RECT 115.025 169.030 115.315 169.075 ;
        RECT 116.865 169.030 117.155 169.075 ;
        RECT 115.025 168.890 117.155 169.030 ;
        RECT 115.025 168.845 115.315 168.890 ;
        RECT 116.865 168.845 117.155 168.890 ;
        RECT 120.545 168.845 120.835 169.075 ;
        RECT 122.845 169.030 123.135 169.075 ;
        RECT 127.890 169.030 128.210 169.090 ;
        RECT 122.845 168.890 128.210 169.030 ;
        RECT 122.845 168.845 123.135 168.890 ;
        RECT 86.020 168.690 86.310 168.735 ;
        RECT 82.760 168.550 86.310 168.690 ;
        RECT 27.625 168.350 27.915 168.395 ;
        RECT 29.910 168.350 30.230 168.410 ;
        RECT 27.625 168.210 30.230 168.350 ;
        RECT 27.625 168.165 27.915 168.210 ;
        RECT 29.910 168.150 30.230 168.210 ;
        RECT 33.145 168.350 33.435 168.395 ;
        RECT 34.050 168.350 34.370 168.410 ;
        RECT 33.145 168.210 34.370 168.350 ;
        RECT 33.145 168.165 33.435 168.210 ;
        RECT 34.050 168.150 34.370 168.210 ;
        RECT 36.810 168.150 37.130 168.410 ;
        RECT 76.370 168.350 76.690 168.410 ;
        RECT 77.840 168.395 77.980 168.550 ;
        RECT 80.755 168.505 81.045 168.550 ;
        RECT 82.760 168.505 83.050 168.550 ;
        RECT 84.190 168.490 84.510 168.550 ;
        RECT 86.020 168.505 86.310 168.550 ;
        RECT 86.940 168.690 87.230 168.735 ;
        RECT 88.800 168.690 89.090 168.735 ;
        RECT 86.940 168.550 89.090 168.690 ;
        RECT 86.940 168.505 87.230 168.550 ;
        RECT 88.800 168.505 89.090 168.550 ;
        RECT 104.545 168.690 105.135 168.735 ;
        RECT 107.190 168.690 107.510 168.750 ;
        RECT 107.785 168.690 108.435 168.735 ;
        RECT 104.545 168.550 108.435 168.690 ;
        RECT 104.545 168.505 104.835 168.550 ;
        RECT 107.190 168.490 107.510 168.550 ;
        RECT 107.785 168.505 108.435 168.550 ;
        RECT 110.410 168.690 110.730 168.750 ;
        RECT 120.620 168.690 120.760 168.845 ;
        RECT 127.890 168.830 128.210 168.890 ;
        RECT 110.410 168.550 120.760 168.690 ;
        RECT 110.410 168.490 110.730 168.550 ;
        RECT 77.765 168.350 78.055 168.395 ;
        RECT 76.370 168.210 78.055 168.350 ;
        RECT 76.370 168.150 76.690 168.210 ;
        RECT 77.765 168.165 78.055 168.210 ;
        RECT 78.225 168.350 78.515 168.395 ;
        RECT 79.130 168.350 79.450 168.410 ;
        RECT 78.225 168.210 79.450 168.350 ;
        RECT 78.225 168.165 78.515 168.210 ;
        RECT 79.130 168.150 79.450 168.210 ;
        RECT 80.065 168.350 80.355 168.395 ;
        RECT 83.270 168.350 83.590 168.410 ;
        RECT 80.065 168.210 83.590 168.350 ;
        RECT 80.065 168.165 80.355 168.210 ;
        RECT 83.270 168.150 83.590 168.210 ;
        RECT 102.590 168.350 102.910 168.410 ;
        RECT 103.065 168.350 103.355 168.395 ;
        RECT 102.590 168.210 103.355 168.350 ;
        RECT 102.590 168.150 102.910 168.210 ;
        RECT 103.065 168.165 103.355 168.210 ;
        RECT 110.870 168.350 111.190 168.410 ;
        RECT 112.725 168.350 113.015 168.395 ;
        RECT 110.870 168.210 113.015 168.350 ;
        RECT 110.870 168.150 111.190 168.210 ;
        RECT 112.725 168.165 113.015 168.210 ;
        RECT 113.170 168.350 113.490 168.410 ;
        RECT 122.385 168.350 122.675 168.395 ;
        RECT 113.170 168.210 122.675 168.350 ;
        RECT 113.170 168.150 113.490 168.210 ;
        RECT 122.385 168.165 122.675 168.210 ;
        RECT 14.660 167.530 127.820 168.010 ;
        RECT 70.390 167.330 70.710 167.390 ;
        RECT 48.400 167.190 53.140 167.330 ;
        RECT 24.850 166.790 25.170 167.050 ;
        RECT 27.145 166.990 27.795 167.035 ;
        RECT 29.910 166.990 30.230 167.050 ;
        RECT 30.745 166.990 31.035 167.035 ;
        RECT 27.145 166.850 31.035 166.990 ;
        RECT 27.145 166.805 27.795 166.850 ;
        RECT 29.910 166.790 30.230 166.850 ;
        RECT 30.445 166.805 31.035 166.850 ;
        RECT 35.890 166.990 36.210 167.050 ;
        RECT 48.400 166.990 48.540 167.190 ;
        RECT 35.890 166.850 48.540 166.990 ;
        RECT 48.885 166.990 49.175 167.035 ;
        RECT 51.070 166.990 51.390 167.050 ;
        RECT 52.125 166.990 52.775 167.035 ;
        RECT 48.885 166.850 52.775 166.990 ;
        RECT 53.000 166.990 53.140 167.190 ;
        RECT 70.390 167.190 73.840 167.330 ;
        RECT 70.390 167.130 70.710 167.190 ;
        RECT 53.370 166.990 53.690 167.050 ;
        RECT 73.165 166.990 73.455 167.035 ;
        RECT 53.000 166.850 59.580 166.990 ;
        RECT 23.950 166.650 24.240 166.695 ;
        RECT 25.785 166.650 26.075 166.695 ;
        RECT 29.365 166.650 29.655 166.695 ;
        RECT 23.950 166.510 29.655 166.650 ;
        RECT 23.950 166.465 24.240 166.510 ;
        RECT 25.785 166.465 26.075 166.510 ;
        RECT 29.365 166.465 29.655 166.510 ;
        RECT 30.445 166.490 30.735 166.805 ;
        RECT 35.890 166.790 36.210 166.850 ;
        RECT 33.605 166.650 33.895 166.695 ;
        RECT 34.510 166.650 34.830 166.710 ;
        RECT 33.605 166.510 34.830 166.650 ;
        RECT 33.605 166.465 33.895 166.510 ;
        RECT 34.510 166.450 34.830 166.510 ;
        RECT 36.365 166.650 36.655 166.695 ;
        RECT 36.810 166.650 37.130 166.710 ;
        RECT 37.820 166.695 37.960 166.850 ;
        RECT 48.885 166.805 49.475 166.850 ;
        RECT 36.365 166.510 37.130 166.650 ;
        RECT 36.365 166.465 36.655 166.510 ;
        RECT 36.810 166.450 37.130 166.510 ;
        RECT 37.745 166.465 38.035 166.695 ;
        RECT 45.640 166.510 49.000 166.650 ;
        RECT 23.485 166.310 23.775 166.355 ;
        RECT 27.150 166.310 27.470 166.370 ;
        RECT 23.485 166.170 27.470 166.310 ;
        RECT 23.485 166.125 23.775 166.170 ;
        RECT 27.150 166.110 27.470 166.170 ;
        RECT 32.225 166.310 32.515 166.355 ;
        RECT 39.585 166.310 39.875 166.355 ;
        RECT 43.250 166.310 43.570 166.370 ;
        RECT 32.225 166.170 43.570 166.310 ;
        RECT 32.225 166.125 32.515 166.170 ;
        RECT 39.585 166.125 39.875 166.170 ;
        RECT 43.250 166.110 43.570 166.170 ;
        RECT 24.355 165.970 24.645 166.015 ;
        RECT 26.245 165.970 26.535 166.015 ;
        RECT 29.365 165.970 29.655 166.015 ;
        RECT 24.355 165.830 29.655 165.970 ;
        RECT 24.355 165.785 24.645 165.830 ;
        RECT 26.245 165.785 26.535 165.830 ;
        RECT 29.365 165.785 29.655 165.830 ;
        RECT 29.910 165.970 30.230 166.030 ;
        RECT 42.345 165.970 42.635 166.015 ;
        RECT 45.640 165.970 45.780 166.510 ;
        RECT 46.025 166.310 46.315 166.355 ;
        RECT 48.860 166.310 49.000 166.510 ;
        RECT 49.185 166.490 49.475 166.805 ;
        RECT 51.070 166.790 51.390 166.850 ;
        RECT 52.125 166.805 52.775 166.850 ;
        RECT 53.370 166.790 53.690 166.850 ;
        RECT 59.440 166.695 59.580 166.850 ;
        RECT 68.640 166.850 73.455 166.990 ;
        RECT 68.640 166.710 68.780 166.850 ;
        RECT 73.165 166.805 73.455 166.850 ;
        RECT 50.265 166.650 50.555 166.695 ;
        RECT 53.845 166.650 54.135 166.695 ;
        RECT 55.680 166.650 55.970 166.695 ;
        RECT 50.265 166.510 55.970 166.650 ;
        RECT 50.265 166.465 50.555 166.510 ;
        RECT 53.845 166.465 54.135 166.510 ;
        RECT 55.680 166.465 55.970 166.510 ;
        RECT 59.365 166.650 59.655 166.695 ;
        RECT 61.205 166.650 61.495 166.695 ;
        RECT 59.365 166.510 61.495 166.650 ;
        RECT 59.365 166.465 59.655 166.510 ;
        RECT 61.205 166.465 61.495 166.510 ;
        RECT 61.650 166.650 61.970 166.710 ;
        RECT 62.585 166.650 62.875 166.695 ;
        RECT 67.185 166.650 67.475 166.695 ;
        RECT 61.650 166.510 67.475 166.650 ;
        RECT 61.650 166.450 61.970 166.510 ;
        RECT 62.585 166.465 62.875 166.510 ;
        RECT 67.185 166.465 67.475 166.510 ;
        RECT 68.550 166.450 68.870 166.710 ;
        RECT 70.850 166.450 71.170 166.710 ;
        RECT 72.705 166.650 72.995 166.695 ;
        RECT 73.700 166.650 73.840 167.190 ;
        RECT 110.410 167.130 110.730 167.390 ;
        RECT 77.700 166.990 77.990 167.035 ;
        RECT 80.960 166.990 81.250 167.035 ;
        RECT 77.700 166.850 81.250 166.990 ;
        RECT 77.700 166.805 77.990 166.850 ;
        RECT 72.705 166.510 73.840 166.650 ;
        RECT 72.705 166.465 72.995 166.510 ;
        RECT 54.290 166.310 54.610 166.370 ;
        RECT 46.025 166.170 47.620 166.310 ;
        RECT 48.860 166.170 54.610 166.310 ;
        RECT 46.025 166.125 46.315 166.170 ;
        RECT 29.910 165.830 45.780 165.970 ;
        RECT 29.910 165.770 30.230 165.830 ;
        RECT 42.345 165.785 42.635 165.830 ;
        RECT 28.530 165.630 28.850 165.690 ;
        RECT 32.685 165.630 32.975 165.675 ;
        RECT 28.530 165.490 32.975 165.630 ;
        RECT 28.530 165.430 28.850 165.490 ;
        RECT 32.685 165.445 32.975 165.490 ;
        RECT 38.190 165.430 38.510 165.690 ;
        RECT 42.790 165.430 43.110 165.690 ;
        RECT 47.480 165.675 47.620 166.170 ;
        RECT 54.290 166.110 54.610 166.170 ;
        RECT 54.750 166.110 55.070 166.370 ;
        RECT 56.145 166.310 56.435 166.355 ;
        RECT 57.510 166.310 57.830 166.370 ;
        RECT 63.950 166.310 64.270 166.370 ;
        RECT 56.145 166.170 64.270 166.310 ;
        RECT 56.145 166.125 56.435 166.170 ;
        RECT 57.510 166.110 57.830 166.170 ;
        RECT 63.950 166.110 64.270 166.170 ;
        RECT 66.710 166.310 67.030 166.370 ;
        RECT 71.325 166.310 71.615 166.355 ;
        RECT 66.710 166.170 71.615 166.310 ;
        RECT 66.710 166.110 67.030 166.170 ;
        RECT 71.325 166.125 71.615 166.170 ;
        RECT 72.245 166.310 72.535 166.355 ;
        RECT 74.070 166.310 74.390 166.370 ;
        RECT 74.990 166.310 75.310 166.370 ;
        RECT 72.245 166.170 75.310 166.310 ;
        RECT 79.220 166.310 79.360 166.850 ;
        RECT 80.960 166.805 81.250 166.850 ;
        RECT 81.880 166.990 82.170 167.035 ;
        RECT 83.740 166.990 84.030 167.035 ;
        RECT 81.880 166.850 84.030 166.990 ;
        RECT 81.880 166.805 82.170 166.850 ;
        RECT 83.740 166.805 84.030 166.850 ;
        RECT 84.190 166.990 84.510 167.050 ;
        RECT 86.965 166.990 87.255 167.035 ;
        RECT 84.190 166.850 87.255 166.990 ;
        RECT 79.560 166.650 79.850 166.695 ;
        RECT 81.880 166.650 82.095 166.805 ;
        RECT 84.190 166.790 84.510 166.850 ;
        RECT 86.965 166.805 87.255 166.850 ;
        RECT 99.780 166.990 100.070 167.035 ;
        RECT 100.290 166.990 100.610 167.050 ;
        RECT 103.040 166.990 103.330 167.035 ;
        RECT 99.780 166.850 103.330 166.990 ;
        RECT 99.780 166.805 100.070 166.850 ;
        RECT 100.290 166.790 100.610 166.850 ;
        RECT 103.040 166.805 103.330 166.850 ;
        RECT 103.960 166.990 104.250 167.035 ;
        RECT 105.820 166.990 106.110 167.035 ;
        RECT 103.960 166.850 106.110 166.990 ;
        RECT 103.960 166.805 104.250 166.850 ;
        RECT 105.820 166.805 106.110 166.850 ;
        RECT 117.425 166.990 117.715 167.035 ;
        RECT 119.610 166.990 119.930 167.050 ;
        RECT 120.665 166.990 121.315 167.035 ;
        RECT 117.425 166.850 121.315 166.990 ;
        RECT 117.425 166.805 118.015 166.850 ;
        RECT 85.585 166.650 85.875 166.695 ;
        RECT 79.560 166.510 82.095 166.650 ;
        RECT 82.440 166.510 85.875 166.650 ;
        RECT 79.560 166.465 79.850 166.510 ;
        RECT 82.440 166.310 82.580 166.510 ;
        RECT 85.585 166.465 85.875 166.510 ;
        RECT 86.045 166.650 86.335 166.695 ;
        RECT 87.425 166.650 87.715 166.695 ;
        RECT 88.790 166.650 89.110 166.710 ;
        RECT 86.045 166.510 89.110 166.650 ;
        RECT 86.045 166.465 86.335 166.510 ;
        RECT 87.425 166.465 87.715 166.510 ;
        RECT 88.790 166.450 89.110 166.510 ;
        RECT 95.245 166.465 95.535 166.695 ;
        RECT 101.640 166.650 101.930 166.695 ;
        RECT 103.960 166.650 104.175 166.805 ;
        RECT 101.640 166.510 104.175 166.650 ;
        RECT 107.665 166.650 107.955 166.695 ;
        RECT 110.870 166.650 111.190 166.710 ;
        RECT 107.665 166.510 111.190 166.650 ;
        RECT 101.640 166.465 101.930 166.510 ;
        RECT 107.665 166.465 107.955 166.510 ;
        RECT 79.220 166.170 82.580 166.310 ;
        RECT 72.245 166.125 72.535 166.170 ;
        RECT 74.070 166.110 74.390 166.170 ;
        RECT 74.990 166.110 75.310 166.170 ;
        RECT 82.810 166.110 83.130 166.370 ;
        RECT 84.665 166.310 84.955 166.355 ;
        RECT 91.090 166.310 91.410 166.370 ;
        RECT 84.665 166.170 91.410 166.310 ;
        RECT 84.665 166.125 84.955 166.170 ;
        RECT 91.090 166.110 91.410 166.170 ;
        RECT 92.010 166.310 92.330 166.370 ;
        RECT 93.850 166.310 94.170 166.370 ;
        RECT 92.010 166.170 94.170 166.310 ;
        RECT 92.010 166.110 92.330 166.170 ;
        RECT 93.850 166.110 94.170 166.170 ;
        RECT 94.770 166.110 95.090 166.370 ;
        RECT 95.320 166.310 95.460 166.465 ;
        RECT 110.870 166.450 111.190 166.510 ;
        RECT 111.345 166.650 111.635 166.695 ;
        RECT 112.250 166.650 112.570 166.710 ;
        RECT 111.345 166.510 112.570 166.650 ;
        RECT 111.345 166.465 111.635 166.510 ;
        RECT 112.250 166.450 112.570 166.510 ;
        RECT 117.725 166.490 118.015 166.805 ;
        RECT 119.610 166.790 119.930 166.850 ;
        RECT 120.665 166.805 121.315 166.850 ;
        RECT 118.805 166.650 119.095 166.695 ;
        RECT 122.385 166.650 122.675 166.695 ;
        RECT 124.220 166.650 124.510 166.695 ;
        RECT 118.805 166.510 124.510 166.650 ;
        RECT 118.805 166.465 119.095 166.510 ;
        RECT 122.385 166.465 122.675 166.510 ;
        RECT 124.220 166.465 124.510 166.510 ;
        RECT 124.670 166.450 124.990 166.710 ;
        RECT 97.775 166.310 98.065 166.355 ;
        RECT 98.450 166.310 98.770 166.370 ;
        RECT 95.320 166.170 98.770 166.310 ;
        RECT 97.775 166.125 98.065 166.170 ;
        RECT 98.450 166.110 98.770 166.170 ;
        RECT 104.890 166.110 105.210 166.370 ;
        RECT 105.810 166.310 106.130 166.370 ;
        RECT 106.745 166.310 107.035 166.355 ;
        RECT 111.790 166.310 112.110 166.370 ;
        RECT 124.760 166.310 124.900 166.450 ;
        RECT 105.810 166.170 124.900 166.310 ;
        RECT 105.810 166.110 106.130 166.170 ;
        RECT 106.745 166.125 107.035 166.170 ;
        RECT 111.790 166.110 112.110 166.170 ;
        RECT 50.265 165.970 50.555 166.015 ;
        RECT 53.385 165.970 53.675 166.015 ;
        RECT 55.275 165.970 55.565 166.015 ;
        RECT 50.265 165.830 55.565 165.970 ;
        RECT 50.265 165.785 50.555 165.830 ;
        RECT 53.385 165.785 53.675 165.830 ;
        RECT 55.275 165.785 55.565 165.830 ;
        RECT 69.945 165.970 70.235 166.015 ;
        RECT 78.670 165.970 78.990 166.030 ;
        RECT 69.945 165.830 78.990 165.970 ;
        RECT 69.945 165.785 70.235 165.830 ;
        RECT 78.670 165.770 78.990 165.830 ;
        RECT 79.560 165.970 79.850 166.015 ;
        RECT 82.340 165.970 82.630 166.015 ;
        RECT 84.200 165.970 84.490 166.015 ;
        RECT 79.560 165.830 84.490 165.970 ;
        RECT 79.560 165.785 79.850 165.830 ;
        RECT 82.340 165.785 82.630 165.830 ;
        RECT 84.200 165.785 84.490 165.830 ;
        RECT 101.640 165.970 101.930 166.015 ;
        RECT 104.420 165.970 104.710 166.015 ;
        RECT 106.280 165.970 106.570 166.015 ;
        RECT 101.640 165.830 106.570 165.970 ;
        RECT 101.640 165.785 101.930 165.830 ;
        RECT 104.420 165.785 104.710 165.830 ;
        RECT 106.280 165.785 106.570 165.830 ;
        RECT 109.030 165.970 109.350 166.030 ;
        RECT 110.870 165.970 111.190 166.030 ;
        RECT 109.030 165.830 111.190 165.970 ;
        RECT 109.030 165.770 109.350 165.830 ;
        RECT 110.870 165.770 111.190 165.830 ;
        RECT 112.250 165.970 112.570 166.030 ;
        RECT 115.945 165.970 116.235 166.015 ;
        RECT 112.250 165.830 116.235 165.970 ;
        RECT 112.250 165.770 112.570 165.830 ;
        RECT 115.945 165.785 116.235 165.830 ;
        RECT 118.805 165.970 119.095 166.015 ;
        RECT 121.925 165.970 122.215 166.015 ;
        RECT 123.815 165.970 124.105 166.015 ;
        RECT 118.805 165.830 124.105 165.970 ;
        RECT 118.805 165.785 119.095 165.830 ;
        RECT 121.925 165.785 122.215 165.830 ;
        RECT 123.815 165.785 124.105 165.830 ;
        RECT 47.405 165.630 47.695 165.675 ;
        RECT 49.690 165.630 50.010 165.690 ;
        RECT 47.405 165.490 50.010 165.630 ;
        RECT 47.405 165.445 47.695 165.490 ;
        RECT 49.690 165.430 50.010 165.490 ;
        RECT 58.890 165.430 59.210 165.690 ;
        RECT 66.725 165.630 67.015 165.675 ;
        RECT 69.010 165.630 69.330 165.690 ;
        RECT 66.725 165.490 69.330 165.630 ;
        RECT 66.725 165.445 67.015 165.490 ;
        RECT 69.010 165.430 69.330 165.490 ;
        RECT 73.150 165.630 73.470 165.690 ;
        RECT 75.695 165.630 75.985 165.675 ;
        RECT 73.150 165.490 75.985 165.630 ;
        RECT 78.760 165.630 78.900 165.770 ;
        RECT 80.050 165.630 80.370 165.690 ;
        RECT 92.010 165.630 92.330 165.690 ;
        RECT 78.760 165.490 92.330 165.630 ;
        RECT 73.150 165.430 73.470 165.490 ;
        RECT 75.695 165.445 75.985 165.490 ;
        RECT 80.050 165.430 80.370 165.490 ;
        RECT 92.010 165.430 92.330 165.490 ;
        RECT 96.610 165.630 96.930 165.690 ;
        RECT 97.085 165.630 97.375 165.675 ;
        RECT 96.610 165.490 97.375 165.630 ;
        RECT 96.610 165.430 96.930 165.490 ;
        RECT 97.085 165.445 97.375 165.490 ;
        RECT 114.090 165.430 114.410 165.690 ;
        RECT 121.450 165.630 121.770 165.690 ;
        RECT 123.370 165.630 123.660 165.675 ;
        RECT 121.450 165.490 123.660 165.630 ;
        RECT 121.450 165.430 121.770 165.490 ;
        RECT 123.370 165.445 123.660 165.490 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 14.660 164.810 127.820 165.290 ;
        RECT 24.850 164.610 25.170 164.670 ;
        RECT 25.785 164.610 26.075 164.655 ;
        RECT 24.850 164.470 26.075 164.610 ;
        RECT 24.850 164.410 25.170 164.470 ;
        RECT 25.785 164.425 26.075 164.470 ;
        RECT 51.070 164.410 51.390 164.670 ;
        RECT 54.750 164.410 55.070 164.670 ;
        RECT 61.650 164.610 61.970 164.670 ;
        RECT 82.810 164.610 83.130 164.670 ;
        RECT 83.285 164.610 83.575 164.655 ;
        RECT 61.650 164.470 71.310 164.610 ;
        RECT 61.650 164.410 61.970 164.470 ;
        RECT 28.035 164.270 28.325 164.315 ;
        RECT 29.925 164.270 30.215 164.315 ;
        RECT 33.045 164.270 33.335 164.315 ;
        RECT 28.035 164.130 33.335 164.270 ;
        RECT 28.035 164.085 28.325 164.130 ;
        RECT 29.925 164.085 30.215 164.130 ;
        RECT 33.045 164.085 33.335 164.130 ;
        RECT 39.225 164.270 39.515 164.315 ;
        RECT 42.345 164.270 42.635 164.315 ;
        RECT 44.235 164.270 44.525 164.315 ;
        RECT 57.510 164.270 57.830 164.330 ;
        RECT 39.225 164.130 44.525 164.270 ;
        RECT 39.225 164.085 39.515 164.130 ;
        RECT 42.345 164.085 42.635 164.130 ;
        RECT 44.235 164.085 44.525 164.130 ;
        RECT 45.180 164.130 57.830 164.270 ;
        RECT 28.530 163.730 28.850 163.990 ;
        RECT 28.990 163.930 29.310 163.990 ;
        RECT 36.810 163.930 37.130 163.990 ;
        RECT 45.180 163.975 45.320 164.130 ;
        RECT 57.510 164.070 57.830 164.130 ;
        RECT 58.085 164.270 58.375 164.315 ;
        RECT 61.205 164.270 61.495 164.315 ;
        RECT 63.095 164.270 63.385 164.315 ;
        RECT 58.085 164.130 63.385 164.270 ;
        RECT 58.085 164.085 58.375 164.130 ;
        RECT 61.205 164.085 61.495 164.130 ;
        RECT 63.095 164.085 63.385 164.130 ;
        RECT 45.105 163.930 45.395 163.975 ;
        RECT 28.990 163.790 45.395 163.930 ;
        RECT 28.990 163.730 29.310 163.790 ;
        RECT 36.810 163.730 37.130 163.790 ;
        RECT 45.105 163.745 45.395 163.790 ;
        RECT 49.705 163.930 49.995 163.975 ;
        RECT 60.730 163.930 61.050 163.990 ;
        RECT 49.705 163.790 54.060 163.930 ;
        RECT 49.705 163.745 49.995 163.790 ;
        RECT 26.690 163.390 27.010 163.650 ;
        RECT 27.150 163.390 27.470 163.650 ;
        RECT 27.630 163.590 27.920 163.635 ;
        RECT 29.465 163.590 29.755 163.635 ;
        RECT 33.045 163.590 33.335 163.635 ;
        RECT 27.630 163.450 33.335 163.590 ;
        RECT 27.630 163.405 27.920 163.450 ;
        RECT 29.465 163.405 29.755 163.450 ;
        RECT 33.045 163.405 33.335 163.450 ;
        RECT 34.050 163.610 34.370 163.650 ;
        RECT 38.190 163.610 38.510 163.650 ;
        RECT 34.050 163.390 34.415 163.610 ;
        RECT 27.240 163.250 27.380 163.390 ;
        RECT 28.990 163.250 29.310 163.310 ;
        RECT 34.125 163.295 34.415 163.390 ;
        RECT 38.145 163.390 38.510 163.610 ;
        RECT 39.225 163.590 39.515 163.635 ;
        RECT 42.805 163.590 43.095 163.635 ;
        RECT 44.640 163.590 44.930 163.635 ;
        RECT 39.225 163.450 44.930 163.590 ;
        RECT 39.225 163.405 39.515 163.450 ;
        RECT 42.805 163.405 43.095 163.450 ;
        RECT 44.640 163.405 44.930 163.450 ;
        RECT 46.945 163.590 47.235 163.635 ;
        RECT 49.230 163.590 49.550 163.650 ;
        RECT 46.945 163.450 49.550 163.590 ;
        RECT 46.945 163.405 47.235 163.450 ;
        RECT 49.230 163.390 49.550 163.450 ;
        RECT 51.545 163.590 51.835 163.635 ;
        RECT 53.370 163.590 53.690 163.650 ;
        RECT 53.920 163.635 54.060 163.790 ;
        RECT 60.730 163.790 65.560 163.930 ;
        RECT 60.730 163.730 61.050 163.790 ;
        RECT 51.545 163.450 53.690 163.590 ;
        RECT 51.545 163.405 51.835 163.450 ;
        RECT 53.370 163.390 53.690 163.450 ;
        RECT 53.845 163.405 54.135 163.635 ;
        RECT 38.145 163.295 38.435 163.390 ;
        RECT 27.240 163.110 29.310 163.250 ;
        RECT 28.990 163.050 29.310 163.110 ;
        RECT 30.825 163.250 31.475 163.295 ;
        RECT 34.125 163.250 34.715 163.295 ;
        RECT 30.825 163.110 34.715 163.250 ;
        RECT 30.825 163.065 31.475 163.110 ;
        RECT 34.425 163.065 34.715 163.110 ;
        RECT 37.845 163.250 38.435 163.295 ;
        RECT 41.085 163.250 41.735 163.295 ;
        RECT 37.845 163.110 41.735 163.250 ;
        RECT 37.845 163.065 38.135 163.110 ;
        RECT 41.085 163.065 41.735 163.110 ;
        RECT 43.725 163.250 44.015 163.295 ;
        RECT 46.470 163.250 46.790 163.310 ;
        RECT 57.005 163.295 57.295 163.610 ;
        RECT 58.085 163.590 58.375 163.635 ;
        RECT 61.665 163.590 61.955 163.635 ;
        RECT 63.500 163.590 63.790 163.635 ;
        RECT 58.085 163.450 63.790 163.590 ;
        RECT 58.085 163.405 58.375 163.450 ;
        RECT 61.665 163.405 61.955 163.450 ;
        RECT 63.500 163.405 63.790 163.450 ;
        RECT 63.950 163.390 64.270 163.650 ;
        RECT 43.725 163.110 46.790 163.250 ;
        RECT 43.725 163.065 44.015 163.110 ;
        RECT 46.470 163.050 46.790 163.110 ;
        RECT 56.705 163.250 57.295 163.295 ;
        RECT 58.890 163.250 59.210 163.310 ;
        RECT 59.945 163.250 60.595 163.295 ;
        RECT 56.705 163.110 60.595 163.250 ;
        RECT 56.705 163.065 56.995 163.110 ;
        RECT 58.890 163.050 59.210 163.110 ;
        RECT 59.945 163.065 60.595 163.110 ;
        RECT 62.570 163.050 62.890 163.310 ;
        RECT 65.420 163.295 65.560 163.790 ;
        RECT 65.880 163.590 66.020 164.470 ;
        RECT 71.170 164.270 71.310 164.470 ;
        RECT 82.810 164.470 83.575 164.610 ;
        RECT 82.810 164.410 83.130 164.470 ;
        RECT 83.285 164.425 83.575 164.470 ;
        RECT 86.505 164.610 86.795 164.655 ;
        RECT 87.870 164.610 88.190 164.670 ;
        RECT 113.170 164.610 113.490 164.670 ;
        RECT 86.505 164.470 88.190 164.610 ;
        RECT 86.505 164.425 86.795 164.470 ;
        RECT 87.870 164.410 88.190 164.470 ;
        RECT 105.900 164.470 113.490 164.610 ;
        RECT 105.900 164.270 106.040 164.470 ;
        RECT 113.170 164.410 113.490 164.470 ;
        RECT 71.170 164.130 106.040 164.270 ;
        RECT 106.745 164.270 107.035 164.315 ;
        RECT 109.030 164.270 109.350 164.330 ;
        RECT 106.745 164.130 109.350 164.270 ;
        RECT 106.745 164.085 107.035 164.130 ;
        RECT 109.030 164.070 109.350 164.130 ;
        RECT 116.505 164.270 116.795 164.315 ;
        RECT 119.625 164.270 119.915 164.315 ;
        RECT 121.515 164.270 121.805 164.315 ;
        RECT 116.505 164.130 121.805 164.270 ;
        RECT 116.505 164.085 116.795 164.130 ;
        RECT 119.625 164.085 119.915 164.130 ;
        RECT 121.515 164.085 121.805 164.130 ;
        RECT 78.670 163.730 78.990 163.990 ;
        RECT 93.850 163.930 94.170 163.990 ;
        RECT 102.605 163.930 102.895 163.975 ;
        RECT 109.505 163.930 109.795 163.975 ;
        RECT 93.850 163.790 109.795 163.930 ;
        RECT 93.850 163.730 94.170 163.790 ;
        RECT 102.605 163.745 102.895 163.790 ;
        RECT 109.505 163.745 109.795 163.790 ;
        RECT 110.410 163.930 110.730 163.990 ;
        RECT 113.645 163.930 113.935 163.975 ;
        RECT 110.410 163.790 113.935 163.930 ;
        RECT 66.725 163.590 67.015 163.635 ;
        RECT 65.880 163.450 67.015 163.590 ;
        RECT 66.725 163.405 67.015 163.450 ;
        RECT 68.550 163.590 68.870 163.650 ;
        RECT 69.025 163.590 69.315 163.635 ;
        RECT 68.550 163.450 69.315 163.590 ;
        RECT 68.550 163.390 68.870 163.450 ;
        RECT 69.025 163.405 69.315 163.450 ;
        RECT 73.150 163.590 73.470 163.650 ;
        RECT 79.605 163.590 79.895 163.635 ;
        RECT 82.365 163.590 82.655 163.635 ;
        RECT 73.150 163.450 79.895 163.590 ;
        RECT 73.150 163.390 73.470 163.450 ;
        RECT 79.220 163.310 79.360 163.450 ;
        RECT 79.605 163.405 79.895 163.450 ;
        RECT 81.980 163.450 82.655 163.590 ;
        RECT 65.345 163.250 65.635 163.295 ;
        RECT 75.450 163.250 75.770 163.310 ;
        RECT 65.345 163.110 75.770 163.250 ;
        RECT 65.345 163.065 65.635 163.110 ;
        RECT 75.450 163.050 75.770 163.110 ;
        RECT 79.130 163.050 79.450 163.310 ;
        RECT 35.890 162.710 36.210 162.970 ;
        RECT 36.350 162.710 36.670 162.970 ;
        RECT 52.910 162.910 53.230 162.970 ;
        RECT 55.225 162.910 55.515 162.955 ;
        RECT 52.910 162.770 55.515 162.910 ;
        RECT 52.910 162.710 53.230 162.770 ;
        RECT 55.225 162.725 55.515 162.770 ;
        RECT 67.170 162.910 67.490 162.970 ;
        RECT 67.645 162.910 67.935 162.955 ;
        RECT 67.170 162.770 67.935 162.910 ;
        RECT 67.170 162.710 67.490 162.770 ;
        RECT 67.645 162.725 67.935 162.770 ;
        RECT 80.065 162.910 80.355 162.955 ;
        RECT 80.970 162.910 81.290 162.970 ;
        RECT 81.980 162.955 82.120 163.450 ;
        RECT 82.365 163.405 82.655 163.450 ;
        RECT 83.270 163.590 83.590 163.650 ;
        RECT 85.585 163.590 85.875 163.635 ;
        RECT 83.270 163.450 85.875 163.590 ;
        RECT 83.270 163.390 83.590 163.450 ;
        RECT 85.585 163.405 85.875 163.450 ;
        RECT 101.210 163.390 101.530 163.650 ;
        RECT 109.580 163.590 109.720 163.745 ;
        RECT 110.410 163.730 110.730 163.790 ;
        RECT 113.645 163.745 113.935 163.790 ;
        RECT 122.385 163.930 122.675 163.975 ;
        RECT 124.670 163.930 124.990 163.990 ;
        RECT 122.385 163.790 124.990 163.930 ;
        RECT 122.385 163.745 122.675 163.790 ;
        RECT 124.670 163.730 124.990 163.790 ;
        RECT 112.710 163.590 113.030 163.650 ;
        RECT 109.580 163.450 113.030 163.590 ;
        RECT 112.710 163.390 113.030 163.450 ;
        RECT 113.170 163.390 113.490 163.650 ;
        RECT 98.450 163.250 98.770 163.310 ;
        RECT 103.525 163.250 103.815 163.295 ;
        RECT 98.450 163.110 103.815 163.250 ;
        RECT 98.450 163.050 98.770 163.110 ;
        RECT 103.525 163.065 103.815 163.110 ;
        RECT 103.985 163.250 104.275 163.295 ;
        RECT 106.270 163.250 106.590 163.310 ;
        RECT 109.045 163.250 109.335 163.295 ;
        RECT 103.985 163.110 109.335 163.250 ;
        RECT 103.985 163.065 104.275 163.110 ;
        RECT 106.270 163.050 106.590 163.110 ;
        RECT 109.045 163.065 109.335 163.110 ;
        RECT 111.790 163.050 112.110 163.310 ;
        RECT 113.630 163.250 113.950 163.310 ;
        RECT 115.425 163.295 115.715 163.610 ;
        RECT 116.505 163.590 116.795 163.635 ;
        RECT 120.085 163.590 120.375 163.635 ;
        RECT 121.920 163.590 122.210 163.635 ;
        RECT 116.505 163.450 122.210 163.590 ;
        RECT 116.505 163.405 116.795 163.450 ;
        RECT 120.085 163.405 120.375 163.450 ;
        RECT 121.920 163.405 122.210 163.450 ;
        RECT 123.750 163.390 124.070 163.650 ;
        RECT 115.125 163.250 115.715 163.295 ;
        RECT 118.365 163.250 119.015 163.295 ;
        RECT 113.630 163.110 119.015 163.250 ;
        RECT 113.630 163.050 113.950 163.110 ;
        RECT 115.125 163.065 115.415 163.110 ;
        RECT 118.365 163.065 119.015 163.110 ;
        RECT 121.005 163.065 121.295 163.295 ;
        RECT 80.065 162.770 81.290 162.910 ;
        RECT 80.065 162.725 80.355 162.770 ;
        RECT 80.970 162.710 81.290 162.770 ;
        RECT 81.905 162.725 82.195 162.955 ;
        RECT 91.090 162.910 91.410 162.970 ;
        RECT 94.785 162.910 95.075 162.955 ;
        RECT 97.530 162.910 97.850 162.970 ;
        RECT 91.090 162.770 97.850 162.910 ;
        RECT 91.090 162.710 91.410 162.770 ;
        RECT 94.785 162.725 95.075 162.770 ;
        RECT 97.530 162.710 97.850 162.770 ;
        RECT 105.350 162.910 105.670 162.970 ;
        RECT 105.825 162.910 106.115 162.955 ;
        RECT 105.350 162.770 106.115 162.910 ;
        RECT 105.350 162.710 105.670 162.770 ;
        RECT 105.825 162.725 106.115 162.770 ;
        RECT 108.585 162.910 108.875 162.955 ;
        RECT 109.950 162.910 110.270 162.970 ;
        RECT 108.585 162.770 110.270 162.910 ;
        RECT 121.080 162.910 121.220 163.065 ;
        RECT 122.845 162.910 123.135 162.955 ;
        RECT 121.080 162.770 123.135 162.910 ;
        RECT 108.585 162.725 108.875 162.770 ;
        RECT 109.950 162.710 110.270 162.770 ;
        RECT 122.845 162.725 123.135 162.770 ;
        RECT 14.660 162.090 127.820 162.570 ;
        RECT 26.690 161.890 27.010 161.950 ;
        RECT 27.625 161.890 27.915 161.935 ;
        RECT 26.690 161.750 27.915 161.890 ;
        RECT 26.690 161.690 27.010 161.750 ;
        RECT 27.625 161.705 27.915 161.750 ;
        RECT 29.910 161.690 30.230 161.950 ;
        RECT 33.145 161.890 33.435 161.935 ;
        RECT 34.510 161.890 34.830 161.950 ;
        RECT 33.145 161.750 34.830 161.890 ;
        RECT 33.145 161.705 33.435 161.750 ;
        RECT 34.510 161.690 34.830 161.750 ;
        RECT 42.790 161.890 43.110 161.950 ;
        RECT 45.565 161.890 45.855 161.935 ;
        RECT 42.790 161.750 45.855 161.890 ;
        RECT 42.790 161.690 43.110 161.750 ;
        RECT 45.565 161.705 45.855 161.750 ;
        RECT 46.470 161.890 46.790 161.950 ;
        RECT 47.865 161.890 48.155 161.935 ;
        RECT 46.470 161.750 48.155 161.890 ;
        RECT 46.470 161.690 46.790 161.750 ;
        RECT 47.865 161.705 48.155 161.750 ;
        RECT 49.230 161.690 49.550 161.950 ;
        RECT 49.690 161.690 50.010 161.950 ;
        RECT 54.290 161.890 54.610 161.950 ;
        RECT 55.225 161.890 55.515 161.935 ;
        RECT 54.290 161.750 55.515 161.890 ;
        RECT 54.290 161.690 54.610 161.750 ;
        RECT 55.225 161.705 55.515 161.750 ;
        RECT 57.065 161.705 57.355 161.935 ;
        RECT 60.745 161.890 61.035 161.935 ;
        RECT 62.570 161.890 62.890 161.950 ;
        RECT 60.745 161.750 62.890 161.890 ;
        RECT 60.745 161.705 61.035 161.750 ;
        RECT 18.870 161.550 19.190 161.610 ;
        RECT 20.200 161.550 20.490 161.595 ;
        RECT 23.460 161.550 23.750 161.595 ;
        RECT 18.870 161.410 23.750 161.550 ;
        RECT 18.870 161.350 19.190 161.410 ;
        RECT 20.200 161.365 20.490 161.410 ;
        RECT 23.460 161.365 23.750 161.410 ;
        RECT 24.380 161.550 24.670 161.595 ;
        RECT 26.240 161.550 26.530 161.595 ;
        RECT 24.380 161.410 26.530 161.550 ;
        RECT 24.380 161.365 24.670 161.410 ;
        RECT 26.240 161.365 26.530 161.410 ;
        RECT 29.465 161.365 29.755 161.595 ;
        RECT 31.290 161.550 31.610 161.610 ;
        RECT 34.985 161.550 35.275 161.595 ;
        RECT 31.290 161.410 35.275 161.550 ;
        RECT 22.060 161.210 22.350 161.255 ;
        RECT 24.380 161.210 24.595 161.365 ;
        RECT 22.060 161.070 24.595 161.210 ;
        RECT 27.150 161.210 27.470 161.270 ;
        RECT 28.990 161.210 29.310 161.270 ;
        RECT 27.150 161.070 29.310 161.210 ;
        RECT 22.060 161.025 22.350 161.070 ;
        RECT 27.150 161.010 27.470 161.070 ;
        RECT 28.990 161.010 29.310 161.070 ;
        RECT 25.325 160.870 25.615 160.915 ;
        RECT 25.770 160.870 26.090 160.930 ;
        RECT 25.325 160.730 26.090 160.870 ;
        RECT 25.325 160.685 25.615 160.730 ;
        RECT 25.770 160.670 26.090 160.730 ;
        RECT 22.060 160.530 22.350 160.575 ;
        RECT 24.840 160.530 25.130 160.575 ;
        RECT 26.700 160.530 26.990 160.575 ;
        RECT 22.060 160.390 26.990 160.530 ;
        RECT 22.060 160.345 22.350 160.390 ;
        RECT 24.840 160.345 25.130 160.390 ;
        RECT 26.700 160.345 26.990 160.390 ;
        RECT 29.540 160.530 29.680 161.365 ;
        RECT 31.290 161.350 31.610 161.410 ;
        RECT 34.985 161.365 35.275 161.410 ;
        RECT 35.445 161.365 35.735 161.595 ;
        RECT 36.350 161.550 36.670 161.610 ;
        RECT 46.025 161.550 46.315 161.595 ;
        RECT 49.780 161.550 49.920 161.690 ;
        RECT 36.350 161.410 46.315 161.550 ;
        RECT 34.050 161.210 34.370 161.270 ;
        RECT 35.520 161.210 35.660 161.365 ;
        RECT 36.350 161.350 36.670 161.410 ;
        RECT 46.025 161.365 46.315 161.410 ;
        RECT 49.320 161.410 49.920 161.550 ;
        RECT 43.265 161.210 43.555 161.255 ;
        RECT 48.785 161.210 49.075 161.255 ;
        RECT 34.050 161.070 35.660 161.210 ;
        RECT 40.120 161.070 41.180 161.210 ;
        RECT 34.050 161.010 34.370 161.070 ;
        RECT 30.830 160.870 31.150 160.930 ;
        RECT 36.365 160.870 36.655 160.915 ;
        RECT 40.120 160.870 40.260 161.070 ;
        RECT 30.830 160.730 40.260 160.870 ;
        RECT 30.830 160.670 31.150 160.730 ;
        RECT 36.365 160.685 36.655 160.730 ;
        RECT 40.505 160.685 40.795 160.915 ;
        RECT 41.040 160.870 41.180 161.070 ;
        RECT 43.265 161.070 49.075 161.210 ;
        RECT 43.265 161.025 43.555 161.070 ;
        RECT 48.785 161.025 49.075 161.070 ;
        RECT 49.320 160.930 49.460 161.410 ;
        RECT 49.690 161.210 50.010 161.270 ;
        RECT 51.085 161.210 51.375 161.255 ;
        RECT 54.765 161.210 55.055 161.255 ;
        RECT 49.690 161.070 55.055 161.210 ;
        RECT 57.140 161.210 57.280 161.705 ;
        RECT 62.570 161.690 62.890 161.750 ;
        RECT 82.810 161.890 83.130 161.950 ;
        RECT 89.955 161.890 90.245 161.935 ;
        RECT 94.770 161.890 95.090 161.950 ;
        RECT 82.810 161.750 84.420 161.890 ;
        RECT 82.810 161.690 83.130 161.750 ;
        RECT 84.280 161.595 84.420 161.750 ;
        RECT 87.960 161.750 95.090 161.890 ;
        RECT 84.205 161.550 84.495 161.595 ;
        RECT 87.960 161.550 88.100 161.750 ;
        RECT 89.955 161.705 90.245 161.750 ;
        RECT 94.770 161.690 95.090 161.750 ;
        RECT 105.825 161.890 106.115 161.935 ;
        RECT 106.270 161.890 106.590 161.950 ;
        RECT 105.825 161.750 106.590 161.890 ;
        RECT 105.825 161.705 106.115 161.750 ;
        RECT 106.270 161.690 106.590 161.750 ;
        RECT 109.950 161.890 110.270 161.950 ;
        RECT 111.805 161.890 112.095 161.935 ;
        RECT 109.950 161.750 112.095 161.890 ;
        RECT 109.950 161.690 110.270 161.750 ;
        RECT 111.805 161.705 112.095 161.750 ;
        RECT 114.105 161.705 114.395 161.935 ;
        RECT 116.390 161.890 116.710 161.950 ;
        RECT 116.865 161.890 117.155 161.935 ;
        RECT 117.310 161.890 117.630 161.950 ;
        RECT 116.390 161.750 117.630 161.890 ;
        RECT 68.180 161.410 70.620 161.550 ;
        RECT 59.825 161.210 60.115 161.255 ;
        RECT 57.140 161.070 60.115 161.210 ;
        RECT 49.690 161.010 50.010 161.070 ;
        RECT 51.085 161.025 51.375 161.070 ;
        RECT 54.765 161.025 55.055 161.070 ;
        RECT 59.825 161.025 60.115 161.070 ;
        RECT 66.265 161.210 66.555 161.255 ;
        RECT 66.710 161.210 67.030 161.270 ;
        RECT 68.180 161.255 68.320 161.410 ;
        RECT 70.480 161.255 70.620 161.410 ;
        RECT 84.205 161.410 88.100 161.550 ;
        RECT 91.960 161.550 92.250 161.595 ;
        RECT 94.310 161.550 94.630 161.610 ;
        RECT 95.220 161.550 95.510 161.595 ;
        RECT 91.960 161.410 95.510 161.550 ;
        RECT 84.205 161.365 84.495 161.410 ;
        RECT 91.960 161.365 92.250 161.410 ;
        RECT 94.310 161.350 94.630 161.410 ;
        RECT 95.220 161.365 95.510 161.410 ;
        RECT 96.140 161.550 96.430 161.595 ;
        RECT 98.000 161.550 98.290 161.595 ;
        RECT 96.140 161.410 98.290 161.550 ;
        RECT 114.180 161.550 114.320 161.705 ;
        RECT 116.390 161.690 116.710 161.750 ;
        RECT 116.865 161.705 117.155 161.750 ;
        RECT 117.310 161.690 117.630 161.750 ;
        RECT 119.610 161.690 119.930 161.950 ;
        RECT 121.450 161.890 121.770 161.950 ;
        RECT 121.925 161.890 122.215 161.935 ;
        RECT 121.450 161.750 122.215 161.890 ;
        RECT 121.450 161.690 121.770 161.750 ;
        RECT 121.925 161.705 122.215 161.750 ;
        RECT 123.750 161.550 124.070 161.610 ;
        RECT 114.180 161.410 124.070 161.550 ;
        RECT 96.140 161.365 96.430 161.410 ;
        RECT 98.000 161.365 98.290 161.410 ;
        RECT 66.265 161.070 67.860 161.210 ;
        RECT 66.265 161.025 66.555 161.070 ;
        RECT 66.710 161.010 67.030 161.070 ;
        RECT 46.945 160.870 47.235 160.915 ;
        RECT 41.040 160.730 47.235 160.870 ;
        RECT 46.945 160.685 47.235 160.730 ;
        RECT 49.230 160.870 49.550 160.930 ;
        RECT 51.545 160.870 51.835 160.915 ;
        RECT 49.230 160.730 51.835 160.870 ;
        RECT 37.730 160.530 38.050 160.590 ;
        RECT 29.540 160.390 38.050 160.530 ;
        RECT 40.580 160.530 40.720 160.685 ;
        RECT 43.725 160.530 44.015 160.575 ;
        RECT 40.580 160.390 44.015 160.530 ;
        RECT 47.020 160.530 47.160 160.685 ;
        RECT 49.230 160.670 49.550 160.730 ;
        RECT 51.545 160.685 51.835 160.730 ;
        RECT 52.465 160.870 52.755 160.915 ;
        RECT 54.305 160.870 54.595 160.915 ;
        RECT 67.170 160.870 67.490 160.930 ;
        RECT 52.465 160.730 67.490 160.870 ;
        RECT 67.720 160.870 67.860 161.070 ;
        RECT 68.105 161.025 68.395 161.255 ;
        RECT 68.565 161.025 68.855 161.255 ;
        RECT 70.405 161.210 70.695 161.255 ;
        RECT 71.310 161.210 71.630 161.270 ;
        RECT 70.405 161.070 71.630 161.210 ;
        RECT 70.405 161.025 70.695 161.070 ;
        RECT 68.640 160.870 68.780 161.025 ;
        RECT 71.310 161.010 71.630 161.070 ;
        RECT 81.905 161.210 82.195 161.255 ;
        RECT 86.505 161.210 86.795 161.255 ;
        RECT 81.905 161.070 85.800 161.210 ;
        RECT 81.905 161.025 82.195 161.070 ;
        RECT 67.720 160.730 68.780 160.870 ;
        RECT 80.050 160.870 80.370 160.930 ;
        RECT 82.825 160.870 83.115 160.915 ;
        RECT 80.050 160.730 83.115 160.870 ;
        RECT 52.465 160.685 52.755 160.730 ;
        RECT 54.305 160.685 54.595 160.730 ;
        RECT 52.540 160.530 52.680 160.685 ;
        RECT 67.170 160.670 67.490 160.730 ;
        RECT 80.050 160.670 80.370 160.730 ;
        RECT 82.825 160.685 83.115 160.730 ;
        RECT 83.745 160.685 84.035 160.915 ;
        RECT 47.020 160.390 52.680 160.530 ;
        RECT 53.370 160.530 53.690 160.590 ;
        RECT 65.345 160.530 65.635 160.575 ;
        RECT 70.850 160.530 71.170 160.590 ;
        RECT 53.370 160.390 71.170 160.530 ;
        RECT 18.195 160.190 18.485 160.235 ;
        RECT 21.630 160.190 21.950 160.250 ;
        RECT 29.540 160.190 29.680 160.390 ;
        RECT 37.730 160.330 38.050 160.390 ;
        RECT 43.725 160.345 44.015 160.390 ;
        RECT 53.370 160.330 53.690 160.390 ;
        RECT 65.345 160.345 65.635 160.390 ;
        RECT 70.850 160.330 71.170 160.390 ;
        RECT 80.970 160.530 81.290 160.590 ;
        RECT 83.820 160.530 83.960 160.685 ;
        RECT 80.970 160.390 83.960 160.530 ;
        RECT 80.970 160.330 81.290 160.390 ;
        RECT 18.195 160.050 29.680 160.190 ;
        RECT 34.050 160.190 34.370 160.250 ;
        RECT 34.970 160.190 35.290 160.250 ;
        RECT 34.050 160.050 35.290 160.190 ;
        RECT 18.195 160.005 18.485 160.050 ;
        RECT 21.630 159.990 21.950 160.050 ;
        RECT 34.050 159.990 34.370 160.050 ;
        RECT 34.970 159.990 35.290 160.050 ;
        RECT 67.170 159.990 67.490 160.250 ;
        RECT 69.485 160.190 69.775 160.235 ;
        RECT 69.930 160.190 70.250 160.250 ;
        RECT 69.485 160.050 70.250 160.190 ;
        RECT 69.485 160.005 69.775 160.050 ;
        RECT 69.930 159.990 70.250 160.050 ;
        RECT 71.325 160.190 71.615 160.235 ;
        RECT 74.070 160.190 74.390 160.250 ;
        RECT 71.325 160.050 74.390 160.190 ;
        RECT 71.325 160.005 71.615 160.050 ;
        RECT 74.070 159.990 74.390 160.050 ;
        RECT 81.445 160.190 81.735 160.235 ;
        RECT 83.270 160.190 83.590 160.250 ;
        RECT 81.445 160.050 83.590 160.190 ;
        RECT 85.660 160.190 85.800 161.070 ;
        RECT 86.120 161.070 86.795 161.210 ;
        RECT 86.120 160.575 86.260 161.070 ;
        RECT 86.505 161.025 86.795 161.070 ;
        RECT 93.820 161.210 94.110 161.255 ;
        RECT 96.140 161.210 96.355 161.365 ;
        RECT 123.750 161.350 124.070 161.410 ;
        RECT 93.820 161.070 96.355 161.210 ;
        RECT 97.530 161.210 97.850 161.270 ;
        RECT 98.925 161.210 99.215 161.255 ;
        RECT 102.145 161.210 102.435 161.255 ;
        RECT 97.530 161.070 102.435 161.210 ;
        RECT 93.820 161.025 94.110 161.070 ;
        RECT 97.530 161.010 97.850 161.070 ;
        RECT 98.925 161.025 99.215 161.070 ;
        RECT 102.145 161.025 102.435 161.070 ;
        RECT 97.070 160.670 97.390 160.930 ;
        RECT 102.220 160.870 102.360 161.025 ;
        RECT 102.590 161.010 102.910 161.270 ;
        RECT 107.205 161.210 107.495 161.255 ;
        RECT 110.410 161.210 110.730 161.270 ;
        RECT 107.205 161.070 110.730 161.210 ;
        RECT 107.205 161.025 107.495 161.070 ;
        RECT 110.410 161.010 110.730 161.070 ;
        RECT 112.265 161.210 112.555 161.255 ;
        RECT 114.090 161.210 114.410 161.270 ;
        RECT 116.405 161.210 116.695 161.255 ;
        RECT 112.265 161.070 116.695 161.210 ;
        RECT 112.265 161.025 112.555 161.070 ;
        RECT 114.090 161.010 114.410 161.070 ;
        RECT 116.405 161.025 116.695 161.070 ;
        RECT 119.150 161.010 119.470 161.270 ;
        RECT 120.990 161.010 121.310 161.270 ;
        RECT 105.810 160.870 106.130 160.930 ;
        RECT 102.220 160.730 106.130 160.870 ;
        RECT 105.810 160.670 106.130 160.730 ;
        RECT 86.045 160.345 86.335 160.575 ;
        RECT 88.790 160.530 89.110 160.590 ;
        RECT 86.580 160.390 89.110 160.530 ;
        RECT 86.580 160.190 86.720 160.390 ;
        RECT 88.790 160.330 89.110 160.390 ;
        RECT 93.820 160.530 94.110 160.575 ;
        RECT 96.600 160.530 96.890 160.575 ;
        RECT 98.460 160.530 98.750 160.575 ;
        RECT 93.820 160.390 98.750 160.530 ;
        RECT 93.820 160.345 94.110 160.390 ;
        RECT 96.600 160.345 96.890 160.390 ;
        RECT 98.460 160.345 98.750 160.390 ;
        RECT 85.660 160.050 86.720 160.190 ;
        RECT 87.425 160.190 87.715 160.235 ;
        RECT 88.330 160.190 88.650 160.250 ;
        RECT 87.425 160.050 88.650 160.190 ;
        RECT 110.500 160.190 110.640 161.010 ;
        RECT 111.345 160.870 111.635 160.915 ;
        RECT 112.710 160.870 113.030 160.930 ;
        RECT 115.485 160.870 115.775 160.915 ;
        RECT 111.345 160.730 115.775 160.870 ;
        RECT 111.345 160.685 111.635 160.730 ;
        RECT 112.710 160.670 113.030 160.730 ;
        RECT 115.485 160.685 115.775 160.730 ;
        RECT 110.870 160.190 111.190 160.250 ;
        RECT 110.500 160.050 111.190 160.190 ;
        RECT 81.445 160.005 81.735 160.050 ;
        RECT 83.270 159.990 83.590 160.050 ;
        RECT 87.425 160.005 87.715 160.050 ;
        RECT 88.330 159.990 88.650 160.050 ;
        RECT 110.870 159.990 111.190 160.050 ;
        RECT 116.850 160.190 117.170 160.250 ;
        RECT 118.705 160.190 118.995 160.235 ;
        RECT 116.850 160.050 118.995 160.190 ;
        RECT 116.850 159.990 117.170 160.050 ;
        RECT 118.705 160.005 118.995 160.050 ;
        RECT 14.660 159.370 127.820 159.850 ;
        RECT 17.965 159.170 18.255 159.215 ;
        RECT 18.870 159.170 19.190 159.230 ;
        RECT 17.965 159.030 19.190 159.170 ;
        RECT 17.965 158.985 18.255 159.030 ;
        RECT 18.870 158.970 19.190 159.030 ;
        RECT 25.770 158.970 26.090 159.230 ;
        RECT 31.290 158.970 31.610 159.230 ;
        RECT 49.690 158.970 50.010 159.230 ;
        RECT 50.610 159.170 50.930 159.230 ;
        RECT 52.910 159.170 53.230 159.230 ;
        RECT 50.610 159.030 53.230 159.170 ;
        RECT 50.610 158.970 50.930 159.030 ;
        RECT 52.910 158.970 53.230 159.030 ;
        RECT 71.325 159.170 71.615 159.215 ;
        RECT 71.770 159.170 72.090 159.230 ;
        RECT 71.325 159.030 72.090 159.170 ;
        RECT 71.325 158.985 71.615 159.030 ;
        RECT 71.770 158.970 72.090 159.030 ;
        RECT 80.050 158.970 80.370 159.230 ;
        RECT 80.970 159.215 81.290 159.230 ;
        RECT 80.970 158.985 81.505 159.215 ;
        RECT 93.405 159.170 93.695 159.215 ;
        RECT 94.310 159.170 94.630 159.230 ;
        RECT 93.405 159.030 94.630 159.170 ;
        RECT 93.405 158.985 93.695 159.030 ;
        RECT 80.970 158.970 81.290 158.985 ;
        RECT 94.310 158.970 94.630 159.030 ;
        RECT 97.070 159.170 97.390 159.230 ;
        RECT 97.545 159.170 97.835 159.215 ;
        RECT 97.070 159.030 97.835 159.170 ;
        RECT 97.070 158.970 97.390 159.030 ;
        RECT 97.545 158.985 97.835 159.030 ;
        RECT 100.290 158.970 100.610 159.230 ;
        RECT 104.445 159.170 104.735 159.215 ;
        RECT 104.890 159.170 105.210 159.230 ;
        RECT 112.250 159.170 112.570 159.230 ;
        RECT 104.445 159.030 105.210 159.170 ;
        RECT 104.445 158.985 104.735 159.030 ;
        RECT 104.890 158.970 105.210 159.030 ;
        RECT 110.500 159.030 112.570 159.170 ;
        RECT 30.830 158.830 31.150 158.890 ;
        RECT 21.260 158.690 31.150 158.830 ;
        RECT 21.260 158.550 21.400 158.690 ;
        RECT 30.830 158.630 31.150 158.690 ;
        RECT 42.650 158.690 54.060 158.830 ;
        RECT 21.170 158.290 21.490 158.550 ;
        RECT 21.630 158.290 21.950 158.550 ;
        RECT 29.910 158.490 30.230 158.550 ;
        RECT 42.650 158.490 42.790 158.690 ;
        RECT 22.870 158.350 30.230 158.490 ;
        RECT 18.425 158.150 18.715 158.195 ;
        RECT 18.885 158.150 19.175 158.195 ;
        RECT 22.870 158.150 23.010 158.350 ;
        RECT 29.910 158.290 30.230 158.350 ;
        RECT 39.200 158.350 42.790 158.490 ;
        RECT 24.865 158.150 25.155 158.195 ;
        RECT 18.425 158.010 23.010 158.150 ;
        RECT 24.020 158.010 25.155 158.150 ;
        RECT 18.425 157.965 18.715 158.010 ;
        RECT 18.885 157.965 19.175 158.010 ;
        RECT 19.330 157.270 19.650 157.530 ;
        RECT 22.090 157.270 22.410 157.530 ;
        RECT 24.020 157.515 24.160 158.010 ;
        RECT 24.865 157.965 25.155 158.010 ;
        RECT 28.545 157.965 28.835 158.195 ;
        RECT 32.210 158.150 32.530 158.210 ;
        RECT 35.890 158.150 36.210 158.210 ;
        RECT 39.200 158.195 39.340 158.350 ;
        RECT 32.210 158.010 36.210 158.150 ;
        RECT 28.620 157.810 28.760 157.965 ;
        RECT 32.210 157.950 32.530 158.010 ;
        RECT 35.890 157.950 36.210 158.010 ;
        RECT 39.125 157.965 39.415 158.195 ;
        RECT 40.045 157.965 40.335 158.195 ;
        RECT 40.505 157.965 40.795 158.195 ;
        RECT 40.965 158.150 41.255 158.195 ;
        RECT 41.870 158.150 42.190 158.210 ;
        RECT 40.965 158.010 42.190 158.150 ;
        RECT 42.650 158.195 42.790 158.350 ;
        RECT 46.945 158.490 47.235 158.535 ;
        RECT 50.610 158.490 50.930 158.550 ;
        RECT 53.920 158.490 54.060 158.690 ;
        RECT 69.485 158.645 69.775 158.875 ;
        RECT 70.850 158.830 71.170 158.890 ;
        RECT 85.080 158.830 85.370 158.875 ;
        RECT 87.860 158.830 88.150 158.875 ;
        RECT 89.720 158.830 90.010 158.875 ;
        RECT 70.850 158.690 78.440 158.830 ;
        RECT 69.560 158.490 69.700 158.645 ;
        RECT 70.850 158.630 71.170 158.690 ;
        RECT 46.945 158.350 50.930 158.490 ;
        RECT 46.945 158.305 47.235 158.350 ;
        RECT 50.610 158.290 50.930 158.350 ;
        RECT 52.080 158.350 53.600 158.490 ;
        RECT 42.650 158.010 43.035 158.195 ;
        RECT 40.965 157.965 41.255 158.010 ;
        RECT 36.350 157.810 36.670 157.870 ;
        RECT 40.120 157.810 40.260 157.965 ;
        RECT 28.620 157.670 40.260 157.810 ;
        RECT 40.580 157.810 40.720 157.965 ;
        RECT 41.870 157.950 42.190 158.010 ;
        RECT 42.745 157.965 43.035 158.010 ;
        RECT 43.250 158.150 43.570 158.210 ;
        RECT 43.725 158.150 44.015 158.195 ;
        RECT 43.250 158.010 44.015 158.150 ;
        RECT 43.250 157.950 43.570 158.010 ;
        RECT 43.725 157.965 44.015 158.010 ;
        RECT 44.185 157.965 44.475 158.195 ;
        RECT 44.645 158.150 44.935 158.195 ;
        RECT 45.090 158.150 45.410 158.210 ;
        RECT 52.080 158.195 52.220 158.350 ;
        RECT 52.005 158.150 52.295 158.195 ;
        RECT 44.645 158.010 52.295 158.150 ;
        RECT 44.645 157.965 44.935 158.010 ;
        RECT 44.260 157.810 44.400 157.965 ;
        RECT 45.090 157.950 45.410 158.010 ;
        RECT 52.005 157.965 52.295 158.010 ;
        RECT 52.465 157.965 52.755 158.195 ;
        RECT 52.540 157.810 52.680 157.965 ;
        RECT 52.910 157.950 53.230 158.210 ;
        RECT 40.580 157.670 52.680 157.810 ;
        RECT 53.460 157.810 53.600 158.350 ;
        RECT 53.920 158.350 72.460 158.490 ;
        RECT 53.920 158.210 54.060 158.350 ;
        RECT 53.830 157.950 54.150 158.210 ;
        RECT 57.050 158.150 57.370 158.210 ;
        RECT 61.205 158.150 61.495 158.195 ;
        RECT 62.585 158.150 62.875 158.195 ;
        RECT 57.050 158.010 62.875 158.150 ;
        RECT 57.050 157.950 57.370 158.010 ;
        RECT 61.205 157.965 61.495 158.010 ;
        RECT 62.585 157.965 62.875 158.010 ;
        RECT 63.030 158.150 63.350 158.210 ;
        RECT 63.965 158.150 64.255 158.195 ;
        RECT 63.030 158.010 64.255 158.150 ;
        RECT 63.030 157.950 63.350 158.010 ;
        RECT 63.965 157.965 64.255 158.010 ;
        RECT 68.565 158.150 68.855 158.195 ;
        RECT 69.470 158.150 69.790 158.210 ;
        RECT 70.390 158.150 70.710 158.210 ;
        RECT 72.320 158.195 72.460 158.350 ;
        RECT 68.565 158.010 70.710 158.150 ;
        RECT 68.565 157.965 68.855 158.010 ;
        RECT 69.470 157.950 69.790 158.010 ;
        RECT 70.390 157.950 70.710 158.010 ;
        RECT 72.245 157.965 72.535 158.195 ;
        RECT 72.320 157.810 72.460 157.965 ;
        RECT 73.150 157.950 73.470 158.210 ;
        RECT 73.700 158.195 73.840 158.690 ;
        RECT 76.370 158.490 76.690 158.550 ;
        RECT 76.370 158.350 77.980 158.490 ;
        RECT 76.370 158.290 76.690 158.350 ;
        RECT 73.625 157.965 73.915 158.195 ;
        RECT 74.070 157.950 74.390 158.210 ;
        RECT 77.840 158.195 77.980 158.350 ;
        RECT 78.300 158.195 78.440 158.690 ;
        RECT 85.080 158.690 90.010 158.830 ;
        RECT 85.080 158.645 85.370 158.690 ;
        RECT 87.860 158.645 88.150 158.690 ;
        RECT 89.720 158.645 90.010 158.690 ;
        RECT 106.745 158.830 107.035 158.875 ;
        RECT 109.490 158.830 109.810 158.890 ;
        RECT 106.745 158.690 109.810 158.830 ;
        RECT 106.745 158.645 107.035 158.690 ;
        RECT 109.490 158.630 109.810 158.690 ;
        RECT 88.330 158.290 88.650 158.550 ;
        RECT 88.790 158.490 89.110 158.550 ;
        RECT 88.790 158.350 93.160 158.490 ;
        RECT 88.790 158.290 89.110 158.350 ;
        RECT 76.845 158.150 77.135 158.195 ;
        RECT 76.460 158.010 77.135 158.150 ;
        RECT 76.460 157.870 76.600 158.010 ;
        RECT 76.845 157.965 77.135 158.010 ;
        RECT 77.765 157.965 78.055 158.195 ;
        RECT 78.225 157.965 78.515 158.195 ;
        RECT 78.685 158.150 78.975 158.195 ;
        RECT 79.130 158.150 79.450 158.210 ;
        RECT 81.890 158.150 82.210 158.210 ;
        RECT 78.685 158.010 82.210 158.150 ;
        RECT 78.685 157.965 78.975 158.010 ;
        RECT 76.370 157.810 76.690 157.870 ;
        RECT 53.460 157.670 61.420 157.810 ;
        RECT 72.320 157.670 76.690 157.810 ;
        RECT 78.300 157.810 78.440 157.965 ;
        RECT 79.130 157.950 79.450 158.010 ;
        RECT 81.890 157.950 82.210 158.010 ;
        RECT 85.080 158.150 85.370 158.195 ;
        RECT 90.185 158.150 90.475 158.195 ;
        RECT 91.090 158.150 91.410 158.210 ;
        RECT 93.020 158.195 93.160 158.350 ;
        RECT 85.080 158.010 87.615 158.150 ;
        RECT 85.080 157.965 85.370 158.010 ;
        RECT 82.350 157.810 82.670 157.870 ;
        RECT 83.270 157.855 83.590 157.870 ;
        RECT 87.400 157.855 87.615 158.010 ;
        RECT 90.185 158.010 91.410 158.150 ;
        RECT 90.185 157.965 90.475 158.010 ;
        RECT 91.090 157.950 91.410 158.010 ;
        RECT 92.945 157.965 93.235 158.195 ;
        RECT 78.300 157.670 82.670 157.810 ;
        RECT 36.350 157.610 36.670 157.670 ;
        RECT 43.340 157.530 43.480 157.670 ;
        RECT 23.945 157.285 24.235 157.515 ;
        RECT 34.970 157.270 35.290 157.530 ;
        RECT 42.330 157.270 42.650 157.530 ;
        RECT 43.250 157.270 43.570 157.530 ;
        RECT 46.010 157.270 46.330 157.530 ;
        RECT 50.150 157.470 50.470 157.530 ;
        RECT 50.625 157.470 50.915 157.515 ;
        RECT 50.150 157.330 50.915 157.470 ;
        RECT 52.540 157.470 52.680 157.670 ;
        RECT 53.370 157.470 53.690 157.530 ;
        RECT 52.540 157.330 53.690 157.470 ;
        RECT 50.150 157.270 50.470 157.330 ;
        RECT 50.625 157.285 50.915 157.330 ;
        RECT 53.370 157.270 53.690 157.330 ;
        RECT 58.890 157.470 59.210 157.530 ;
        RECT 60.745 157.470 61.035 157.515 ;
        RECT 58.890 157.330 61.035 157.470 ;
        RECT 61.280 157.470 61.420 157.670 ;
        RECT 76.370 157.610 76.690 157.670 ;
        RECT 82.350 157.610 82.670 157.670 ;
        RECT 83.220 157.810 83.590 157.855 ;
        RECT 86.480 157.810 86.770 157.855 ;
        RECT 83.220 157.670 86.770 157.810 ;
        RECT 83.220 157.625 83.590 157.670 ;
        RECT 86.480 157.625 86.770 157.670 ;
        RECT 87.400 157.810 87.690 157.855 ;
        RECT 89.260 157.810 89.550 157.855 ;
        RECT 87.400 157.670 89.550 157.810 ;
        RECT 93.020 157.810 93.160 157.965 ;
        RECT 96.610 157.950 96.930 158.210 ;
        RECT 99.845 157.965 100.135 158.195 ;
        RECT 95.230 157.810 95.550 157.870 ;
        RECT 99.920 157.810 100.060 157.965 ;
        RECT 105.350 157.950 105.670 158.210 ;
        RECT 105.825 158.150 106.115 158.195 ;
        RECT 109.030 158.150 109.350 158.210 ;
        RECT 105.825 158.010 109.350 158.150 ;
        RECT 105.825 157.965 106.115 158.010 ;
        RECT 109.030 157.950 109.350 158.010 ;
        RECT 109.490 157.950 109.810 158.210 ;
        RECT 109.950 157.950 110.270 158.210 ;
        RECT 110.500 158.195 110.640 159.030 ;
        RECT 112.250 158.970 112.570 159.030 ;
        RECT 119.625 159.170 119.915 159.215 ;
        RECT 120.990 159.170 121.310 159.230 ;
        RECT 119.625 159.030 121.310 159.170 ;
        RECT 119.625 158.985 119.915 159.030 ;
        RECT 120.990 158.970 121.310 159.030 ;
        RECT 116.850 158.290 117.170 158.550 ;
        RECT 110.425 157.965 110.715 158.195 ;
        RECT 111.345 158.150 111.635 158.195 ;
        RECT 111.790 158.150 112.110 158.210 ;
        RECT 111.345 158.010 112.110 158.150 ;
        RECT 111.345 157.965 111.635 158.010 ;
        RECT 111.790 157.950 112.110 158.010 ;
        RECT 112.250 157.810 112.570 157.870 ;
        RECT 93.020 157.670 112.570 157.810 ;
        RECT 87.400 157.625 87.690 157.670 ;
        RECT 89.260 157.625 89.550 157.670 ;
        RECT 83.270 157.610 83.590 157.625 ;
        RECT 95.230 157.610 95.550 157.670 ;
        RECT 112.250 157.610 112.570 157.670 ;
        RECT 74.070 157.470 74.390 157.530 ;
        RECT 61.280 157.330 74.390 157.470 ;
        RECT 58.890 157.270 59.210 157.330 ;
        RECT 60.745 157.285 61.035 157.330 ;
        RECT 74.070 157.270 74.390 157.330 ;
        RECT 75.465 157.470 75.755 157.515 ;
        RECT 75.910 157.470 76.230 157.530 ;
        RECT 75.465 157.330 76.230 157.470 ;
        RECT 75.465 157.285 75.755 157.330 ;
        RECT 75.910 157.270 76.230 157.330 ;
        RECT 108.125 157.470 108.415 157.515 ;
        RECT 109.030 157.470 109.350 157.530 ;
        RECT 108.125 157.330 109.350 157.470 ;
        RECT 108.125 157.285 108.415 157.330 ;
        RECT 109.030 157.270 109.350 157.330 ;
        RECT 14.660 156.650 127.820 157.130 ;
        RECT 17.275 156.450 17.565 156.495 ;
        RECT 22.090 156.450 22.410 156.510 ;
        RECT 33.590 156.450 33.910 156.510 ;
        RECT 34.525 156.450 34.815 156.495 ;
        RECT 17.275 156.310 32.900 156.450 ;
        RECT 17.275 156.265 17.565 156.310 ;
        RECT 22.090 156.250 22.410 156.310 ;
        RECT 19.330 156.155 19.650 156.170 ;
        RECT 19.280 156.110 19.650 156.155 ;
        RECT 22.540 156.110 22.830 156.155 ;
        RECT 19.280 155.970 22.830 156.110 ;
        RECT 19.280 155.925 19.650 155.970 ;
        RECT 22.540 155.925 22.830 155.970 ;
        RECT 23.460 156.110 23.750 156.155 ;
        RECT 25.320 156.110 25.610 156.155 ;
        RECT 23.460 155.970 25.610 156.110 ;
        RECT 32.760 156.110 32.900 156.310 ;
        RECT 33.590 156.310 34.815 156.450 ;
        RECT 33.590 156.250 33.910 156.310 ;
        RECT 34.525 156.265 34.815 156.310 ;
        RECT 34.970 156.250 35.290 156.510 ;
        RECT 41.870 156.450 42.190 156.510 ;
        RECT 45.090 156.450 45.410 156.510 ;
        RECT 40.580 156.310 45.410 156.450 ;
        RECT 32.760 155.970 34.740 156.110 ;
        RECT 23.460 155.925 23.750 155.970 ;
        RECT 25.320 155.925 25.610 155.970 ;
        RECT 19.330 155.910 19.650 155.925 ;
        RECT 21.140 155.770 21.430 155.815 ;
        RECT 23.460 155.770 23.675 155.925 ;
        RECT 21.140 155.630 23.675 155.770 ;
        RECT 26.245 155.770 26.535 155.815 ;
        RECT 27.150 155.770 27.470 155.830 ;
        RECT 26.245 155.630 27.470 155.770 ;
        RECT 21.140 155.585 21.430 155.630 ;
        RECT 26.245 155.585 26.535 155.630 ;
        RECT 27.150 155.570 27.470 155.630 ;
        RECT 27.610 155.570 27.930 155.830 ;
        RECT 31.290 155.770 31.610 155.830 ;
        RECT 33.590 155.770 33.910 155.830 ;
        RECT 31.290 155.630 33.910 155.770 ;
        RECT 31.290 155.570 31.610 155.630 ;
        RECT 33.590 155.570 33.910 155.630 ;
        RECT 24.405 155.430 24.695 155.475 ;
        RECT 30.830 155.430 31.150 155.490 ;
        RECT 34.050 155.430 34.370 155.490 ;
        RECT 24.405 155.290 26.920 155.430 ;
        RECT 24.405 155.245 24.695 155.290 ;
        RECT 26.780 155.135 26.920 155.290 ;
        RECT 30.830 155.290 34.370 155.430 ;
        RECT 34.600 155.430 34.740 155.970 ;
        RECT 40.580 155.770 40.720 156.310 ;
        RECT 41.870 156.250 42.190 156.310 ;
        RECT 45.090 156.250 45.410 156.310 ;
        RECT 49.230 156.450 49.550 156.510 ;
        RECT 50.610 156.450 50.930 156.510 ;
        RECT 67.170 156.450 67.490 156.510 ;
        RECT 102.590 156.450 102.910 156.510 ;
        RECT 108.570 156.450 108.890 156.510 ;
        RECT 111.790 156.450 112.110 156.510 ;
        RECT 49.230 156.310 49.920 156.450 ;
        RECT 49.230 156.250 49.550 156.310 ;
        RECT 40.950 156.110 41.270 156.170 ;
        RECT 45.180 156.110 45.320 156.250 ;
        RECT 40.950 155.970 43.480 156.110 ;
        RECT 40.950 155.910 41.270 155.970 ;
        RECT 41.425 155.770 41.715 155.815 ;
        RECT 40.580 155.630 41.715 155.770 ;
        RECT 41.425 155.585 41.715 155.630 ;
        RECT 41.870 155.570 42.190 155.830 ;
        RECT 43.340 155.815 43.480 155.970 ;
        RECT 45.180 155.970 49.000 156.110 ;
        RECT 45.180 155.815 45.320 155.970 ;
        RECT 42.345 155.585 42.635 155.815 ;
        RECT 43.265 155.585 43.555 155.815 ;
        RECT 45.105 155.585 45.395 155.815 ;
        RECT 45.550 155.585 45.840 155.815 ;
        RECT 46.050 155.585 46.340 155.815 ;
        RECT 42.420 155.430 42.560 155.585 ;
        RECT 34.600 155.290 42.560 155.430 ;
        RECT 43.710 155.430 44.030 155.490 ;
        RECT 45.640 155.430 45.780 155.585 ;
        RECT 43.710 155.290 45.780 155.430 ;
        RECT 30.830 155.230 31.150 155.290 ;
        RECT 34.050 155.230 34.370 155.290 ;
        RECT 43.710 155.230 44.030 155.290 ;
        RECT 21.140 155.090 21.430 155.135 ;
        RECT 23.920 155.090 24.210 155.135 ;
        RECT 25.780 155.090 26.070 155.135 ;
        RECT 21.140 154.950 26.070 155.090 ;
        RECT 21.140 154.905 21.430 154.950 ;
        RECT 23.920 154.905 24.210 154.950 ;
        RECT 25.780 154.905 26.070 154.950 ;
        RECT 26.705 154.905 26.995 155.135 ;
        RECT 32.210 155.090 32.530 155.150 ;
        RECT 46.100 155.090 46.240 155.585 ;
        RECT 46.930 155.570 47.250 155.830 ;
        RECT 48.860 155.815 49.000 155.970 ;
        RECT 49.780 155.815 49.920 156.310 ;
        RECT 50.610 156.310 85.110 156.450 ;
        RECT 50.610 156.250 50.930 156.310 ;
        RECT 67.170 156.250 67.490 156.310 ;
        RECT 53.370 156.110 53.690 156.170 ;
        RECT 58.890 156.155 59.210 156.170 ;
        RECT 50.240 155.970 53.690 156.110 ;
        RECT 48.785 155.585 49.075 155.815 ;
        RECT 49.245 155.585 49.535 155.815 ;
        RECT 49.705 155.585 49.995 155.815 ;
        RECT 49.320 155.430 49.460 155.585 ;
        RECT 50.240 155.430 50.380 155.970 ;
        RECT 53.370 155.910 53.690 155.970 ;
        RECT 55.620 156.110 55.910 156.155 ;
        RECT 58.880 156.110 59.210 156.155 ;
        RECT 55.620 155.970 59.210 156.110 ;
        RECT 55.620 155.925 55.910 155.970 ;
        RECT 58.880 155.925 59.210 155.970 ;
        RECT 58.890 155.910 59.210 155.925 ;
        RECT 59.800 156.110 60.090 156.155 ;
        RECT 61.660 156.110 61.950 156.155 ;
        RECT 59.800 155.970 61.950 156.110 ;
        RECT 59.800 155.925 60.090 155.970 ;
        RECT 61.660 155.925 61.950 155.970 ;
        RECT 74.070 156.110 74.390 156.170 ;
        RECT 80.970 156.110 81.290 156.170 ;
        RECT 74.070 155.970 78.440 156.110 ;
        RECT 50.625 155.770 50.915 155.815 ;
        RECT 53.830 155.770 54.150 155.830 ;
        RECT 50.625 155.630 54.150 155.770 ;
        RECT 50.625 155.585 50.915 155.630 ;
        RECT 49.320 155.290 50.380 155.430 ;
        RECT 32.210 154.950 46.240 155.090 ;
        RECT 46.930 155.090 47.250 155.150 ;
        RECT 50.700 155.090 50.840 155.585 ;
        RECT 53.830 155.570 54.150 155.630 ;
        RECT 57.480 155.770 57.770 155.815 ;
        RECT 59.800 155.770 60.015 155.925 ;
        RECT 74.070 155.910 74.390 155.970 ;
        RECT 78.300 155.830 78.440 155.970 ;
        RECT 79.680 155.970 81.290 156.110 ;
        RECT 84.970 156.110 85.110 156.310 ;
        RECT 102.590 156.310 112.110 156.450 ;
        RECT 102.590 156.250 102.910 156.310 ;
        RECT 103.050 156.110 103.370 156.170 ;
        RECT 84.970 155.970 98.220 156.110 ;
        RECT 57.480 155.630 60.015 155.770 ;
        RECT 62.585 155.770 62.875 155.815 ;
        RECT 63.950 155.770 64.270 155.830 ;
        RECT 62.585 155.630 64.270 155.770 ;
        RECT 57.480 155.585 57.770 155.630 ;
        RECT 62.585 155.585 62.875 155.630 ;
        RECT 63.950 155.570 64.270 155.630 ;
        RECT 74.530 155.570 74.850 155.830 ;
        RECT 78.210 155.570 78.530 155.830 ;
        RECT 78.670 155.570 78.990 155.830 ;
        RECT 79.145 155.770 79.435 155.815 ;
        RECT 79.680 155.770 79.820 155.970 ;
        RECT 80.970 155.910 81.290 155.970 ;
        RECT 79.145 155.630 79.820 155.770 ;
        RECT 79.145 155.585 79.435 155.630 ;
        RECT 80.065 155.585 80.355 155.815 ;
        RECT 60.745 155.430 61.035 155.475 ;
        RECT 61.190 155.430 61.510 155.490 ;
        RECT 60.745 155.290 61.510 155.430 ;
        RECT 60.745 155.245 61.035 155.290 ;
        RECT 61.190 155.230 61.510 155.290 ;
        RECT 65.790 155.230 66.110 155.490 ;
        RECT 76.370 155.430 76.690 155.490 ;
        RECT 80.140 155.430 80.280 155.585 ;
        RECT 81.890 155.570 82.210 155.830 ;
        RECT 82.350 155.570 82.670 155.830 ;
        RECT 82.810 155.570 83.130 155.830 ;
        RECT 83.745 155.585 84.035 155.815 ;
        RECT 84.650 155.770 84.970 155.830 ;
        RECT 97.545 155.770 97.835 155.815 ;
        RECT 84.650 155.630 97.835 155.770 ;
        RECT 83.820 155.430 83.960 155.585 ;
        RECT 84.650 155.570 84.970 155.630 ;
        RECT 97.545 155.585 97.835 155.630 ;
        RECT 76.370 155.290 83.960 155.430 ;
        RECT 76.370 155.230 76.690 155.290 ;
        RECT 46.930 154.950 50.840 155.090 ;
        RECT 57.480 155.090 57.770 155.135 ;
        RECT 60.260 155.090 60.550 155.135 ;
        RECT 62.120 155.090 62.410 155.135 ;
        RECT 57.480 154.950 62.410 155.090 ;
        RECT 32.210 154.890 32.530 154.950 ;
        RECT 46.930 154.890 47.250 154.950 ;
        RECT 57.480 154.905 57.770 154.950 ;
        RECT 60.260 154.905 60.550 154.950 ;
        RECT 62.120 154.905 62.410 154.950 ;
        RECT 78.670 155.090 78.990 155.150 ;
        RECT 82.350 155.090 82.670 155.150 ;
        RECT 78.670 154.950 82.670 155.090 ;
        RECT 97.620 155.090 97.760 155.585 ;
        RECT 98.080 155.430 98.220 155.970 ;
        RECT 103.050 155.970 106.500 156.110 ;
        RECT 103.050 155.910 103.370 155.970 ;
        RECT 98.450 155.570 98.770 155.830 ;
        RECT 98.910 155.570 99.230 155.830 ;
        RECT 99.385 155.770 99.675 155.815 ;
        RECT 104.905 155.770 105.195 155.815 ;
        RECT 99.385 155.630 105.195 155.770 ;
        RECT 99.385 155.585 99.675 155.630 ;
        RECT 104.905 155.585 105.195 155.630 ;
        RECT 99.460 155.430 99.600 155.585 ;
        RECT 98.080 155.290 99.600 155.430 ;
        RECT 102.590 155.090 102.910 155.150 ;
        RECT 97.620 154.950 102.910 155.090 ;
        RECT 78.670 154.890 78.990 154.950 ;
        RECT 82.350 154.890 82.670 154.950 ;
        RECT 102.590 154.890 102.910 154.950 ;
        RECT 35.890 154.750 36.210 154.810 ;
        RECT 36.825 154.750 37.115 154.795 ;
        RECT 35.890 154.610 37.115 154.750 ;
        RECT 35.890 154.550 36.210 154.610 ;
        RECT 36.825 154.565 37.115 154.610 ;
        RECT 40.030 154.550 40.350 154.810 ;
        RECT 43.710 154.550 44.030 154.810 ;
        RECT 45.090 154.750 45.410 154.810 ;
        RECT 47.020 154.750 47.160 154.890 ;
        RECT 45.090 154.610 47.160 154.750 ;
        RECT 47.405 154.750 47.695 154.795 ;
        RECT 49.230 154.750 49.550 154.810 ;
        RECT 53.830 154.795 54.150 154.810 ;
        RECT 47.405 154.610 49.550 154.750 ;
        RECT 45.090 154.550 45.410 154.610 ;
        RECT 47.405 154.565 47.695 154.610 ;
        RECT 49.230 154.550 49.550 154.610 ;
        RECT 53.615 154.565 54.150 154.795 ;
        RECT 53.830 154.550 54.150 154.565 ;
        RECT 54.290 154.750 54.610 154.810 ;
        RECT 69.930 154.750 70.250 154.810 ;
        RECT 54.290 154.610 70.250 154.750 ;
        RECT 54.290 154.550 54.610 154.610 ;
        RECT 69.930 154.550 70.250 154.610 ;
        RECT 76.370 154.750 76.690 154.810 ;
        RECT 76.845 154.750 77.135 154.795 ;
        RECT 76.370 154.610 77.135 154.750 ;
        RECT 76.370 154.550 76.690 154.610 ;
        RECT 76.845 154.565 77.135 154.610 ;
        RECT 80.510 154.550 80.830 154.810 ;
        RECT 99.830 154.750 100.150 154.810 ;
        RECT 100.765 154.750 101.055 154.795 ;
        RECT 99.830 154.610 101.055 154.750 ;
        RECT 99.830 154.550 100.150 154.610 ;
        RECT 100.765 154.565 101.055 154.610 ;
        RECT 103.525 154.750 103.815 154.795 ;
        RECT 103.970 154.750 104.290 154.810 ;
        RECT 103.525 154.610 104.290 154.750 ;
        RECT 104.980 154.750 105.120 155.585 ;
        RECT 105.350 155.570 105.670 155.830 ;
        RECT 105.825 155.770 106.115 155.815 ;
        RECT 106.360 155.770 106.500 155.970 ;
        RECT 106.820 155.815 106.960 156.310 ;
        RECT 108.570 156.250 108.890 156.310 ;
        RECT 111.790 156.250 112.110 156.310 ;
        RECT 110.870 156.110 111.190 156.170 ;
        RECT 108.200 155.970 111.190 156.110 ;
        RECT 108.200 155.815 108.340 155.970 ;
        RECT 110.870 155.910 111.190 155.970 ;
        RECT 105.825 155.630 106.500 155.770 ;
        RECT 106.745 155.770 107.035 155.815 ;
        RECT 107.205 155.770 107.495 155.815 ;
        RECT 106.745 155.630 107.495 155.770 ;
        RECT 105.825 155.585 106.115 155.630 ;
        RECT 106.745 155.585 107.035 155.630 ;
        RECT 107.205 155.585 107.495 155.630 ;
        RECT 108.125 155.585 108.415 155.815 ;
        RECT 108.585 155.585 108.875 155.815 ;
        RECT 109.045 155.770 109.335 155.815 ;
        RECT 109.490 155.770 109.810 155.830 ;
        RECT 109.045 155.630 109.810 155.770 ;
        RECT 109.045 155.585 109.335 155.630 ;
        RECT 105.440 155.430 105.580 155.570 ;
        RECT 108.660 155.430 108.800 155.585 ;
        RECT 105.440 155.290 108.800 155.430 ;
        RECT 109.120 155.090 109.260 155.585 ;
        RECT 109.490 155.570 109.810 155.630 ;
        RECT 113.170 155.770 113.490 155.830 ;
        RECT 116.405 155.770 116.695 155.815 ;
        RECT 113.170 155.630 116.695 155.770 ;
        RECT 113.170 155.570 113.490 155.630 ;
        RECT 116.405 155.585 116.695 155.630 ;
        RECT 117.770 155.230 118.090 155.490 ;
        RECT 108.660 154.950 109.260 155.090 ;
        RECT 106.730 154.750 107.050 154.810 ;
        RECT 108.660 154.750 108.800 154.950 ;
        RECT 104.980 154.610 108.800 154.750 ;
        RECT 110.425 154.750 110.715 154.795 ;
        RECT 110.870 154.750 111.190 154.810 ;
        RECT 110.425 154.610 111.190 154.750 ;
        RECT 103.525 154.565 103.815 154.610 ;
        RECT 103.970 154.550 104.290 154.610 ;
        RECT 106.730 154.550 107.050 154.610 ;
        RECT 110.425 154.565 110.715 154.610 ;
        RECT 110.870 154.550 111.190 154.610 ;
        RECT 14.660 153.930 127.820 154.410 ;
        RECT 23.945 153.730 24.235 153.775 ;
        RECT 27.610 153.730 27.930 153.790 ;
        RECT 23.945 153.590 27.930 153.730 ;
        RECT 23.945 153.545 24.235 153.590 ;
        RECT 27.610 153.530 27.930 153.590 ;
        RECT 70.390 153.730 70.710 153.790 ;
        RECT 72.245 153.730 72.535 153.775 ;
        RECT 70.390 153.590 72.535 153.730 ;
        RECT 70.390 153.530 70.710 153.590 ;
        RECT 72.245 153.545 72.535 153.590 ;
        RECT 73.610 153.530 73.930 153.790 ;
        RECT 98.910 153.730 99.230 153.790 ;
        RECT 84.970 153.590 99.230 153.730 ;
        RECT 34.020 153.390 34.310 153.435 ;
        RECT 36.800 153.390 37.090 153.435 ;
        RECT 38.660 153.390 38.950 153.435 ;
        RECT 54.290 153.390 54.610 153.450 ;
        RECT 34.020 153.250 38.950 153.390 ;
        RECT 34.020 153.205 34.310 153.250 ;
        RECT 36.800 153.205 37.090 153.250 ;
        RECT 38.660 153.205 38.950 153.250 ;
        RECT 42.420 153.250 54.610 153.390 ;
        RECT 21.170 152.850 21.490 153.110 ;
        RECT 21.645 153.050 21.935 153.095 ;
        RECT 22.090 153.050 22.410 153.110 ;
        RECT 21.645 152.910 22.410 153.050 ;
        RECT 21.645 152.865 21.935 152.910 ;
        RECT 22.090 152.850 22.410 152.910 ;
        RECT 37.270 152.850 37.590 153.110 ;
        RECT 37.730 153.050 38.050 153.110 ;
        RECT 37.730 152.910 42.100 153.050 ;
        RECT 37.730 152.850 38.050 152.910 ;
        RECT 34.020 152.710 34.310 152.755 ;
        RECT 36.810 152.710 37.130 152.770 ;
        RECT 41.960 152.755 42.100 152.910 ;
        RECT 39.125 152.710 39.415 152.755 ;
        RECT 34.020 152.570 36.555 152.710 ;
        RECT 34.020 152.525 34.310 152.570 ;
        RECT 32.160 152.370 32.450 152.415 ;
        RECT 33.590 152.370 33.910 152.430 ;
        RECT 36.340 152.415 36.555 152.570 ;
        RECT 36.810 152.570 39.415 152.710 ;
        RECT 36.810 152.510 37.130 152.570 ;
        RECT 39.125 152.525 39.415 152.570 ;
        RECT 40.965 152.525 41.255 152.755 ;
        RECT 41.425 152.525 41.715 152.755 ;
        RECT 41.885 152.525 42.175 152.755 ;
        RECT 35.420 152.370 35.710 152.415 ;
        RECT 32.160 152.230 35.710 152.370 ;
        RECT 32.160 152.185 32.450 152.230 ;
        RECT 33.590 152.170 33.910 152.230 ;
        RECT 35.420 152.185 35.710 152.230 ;
        RECT 36.340 152.370 36.630 152.415 ;
        RECT 38.200 152.370 38.490 152.415 ;
        RECT 36.340 152.230 38.490 152.370 ;
        RECT 36.340 152.185 36.630 152.230 ;
        RECT 38.200 152.185 38.490 152.230 ;
        RECT 22.105 152.030 22.395 152.075 ;
        RECT 22.550 152.030 22.870 152.090 ;
        RECT 22.105 151.890 22.870 152.030 ;
        RECT 22.105 151.845 22.395 151.890 ;
        RECT 22.550 151.830 22.870 151.890 ;
        RECT 30.155 152.030 30.445 152.075 ;
        RECT 31.290 152.030 31.610 152.090 ;
        RECT 30.155 151.890 31.610 152.030 ;
        RECT 30.155 151.845 30.445 151.890 ;
        RECT 31.290 151.830 31.610 151.890 ;
        RECT 34.970 152.030 35.290 152.090 ;
        RECT 39.585 152.030 39.875 152.075 ;
        RECT 34.970 151.890 39.875 152.030 ;
        RECT 41.040 152.030 41.180 152.525 ;
        RECT 41.500 152.370 41.640 152.525 ;
        RECT 42.420 152.370 42.560 153.250 ;
        RECT 54.290 153.190 54.610 153.250 ;
        RECT 62.540 153.390 62.830 153.435 ;
        RECT 65.320 153.390 65.610 153.435 ;
        RECT 67.180 153.390 67.470 153.435 ;
        RECT 62.540 153.250 67.470 153.390 ;
        RECT 62.540 153.205 62.830 153.250 ;
        RECT 65.320 153.205 65.610 153.250 ;
        RECT 67.180 153.205 67.470 153.250 ;
        RECT 69.930 153.390 70.250 153.450 ;
        RECT 84.970 153.390 85.110 153.590 ;
        RECT 98.910 153.530 99.230 153.590 ;
        RECT 103.050 153.730 103.370 153.790 ;
        RECT 103.525 153.730 103.815 153.775 ;
        RECT 109.950 153.730 110.270 153.790 ;
        RECT 103.050 153.590 103.815 153.730 ;
        RECT 103.050 153.530 103.370 153.590 ;
        RECT 103.525 153.545 103.815 153.590 ;
        RECT 107.280 153.590 110.270 153.730 ;
        RECT 69.930 153.250 85.110 153.390 ;
        RECT 90.600 153.390 90.890 153.435 ;
        RECT 93.380 153.390 93.670 153.435 ;
        RECT 95.240 153.390 95.530 153.435 ;
        RECT 90.600 153.250 95.530 153.390 ;
        RECT 99.000 153.390 99.140 153.530 ;
        RECT 105.350 153.390 105.670 153.450 ;
        RECT 99.000 153.250 105.670 153.390 ;
        RECT 69.930 153.190 70.250 153.250 ;
        RECT 90.600 153.205 90.890 153.250 ;
        RECT 93.380 153.205 93.670 153.250 ;
        RECT 95.240 153.205 95.530 153.250 ;
        RECT 105.350 153.190 105.670 153.250 ;
        RECT 64.410 153.050 64.730 153.110 ;
        RECT 69.470 153.050 69.790 153.110 ;
        RECT 74.070 153.050 74.390 153.110 ;
        RECT 74.545 153.050 74.835 153.095 ;
        RECT 64.410 152.910 69.240 153.050 ;
        RECT 64.410 152.850 64.730 152.910 ;
        RECT 42.805 152.710 43.095 152.755 ;
        RECT 44.630 152.710 44.950 152.770 ;
        RECT 42.805 152.570 44.950 152.710 ;
        RECT 42.805 152.525 43.095 152.570 ;
        RECT 44.630 152.510 44.950 152.570 ;
        RECT 51.070 152.710 51.390 152.770 ;
        RECT 57.050 152.710 57.370 152.770 ;
        RECT 51.070 152.570 57.370 152.710 ;
        RECT 51.070 152.510 51.390 152.570 ;
        RECT 57.050 152.510 57.370 152.570 ;
        RECT 62.540 152.710 62.830 152.755 ;
        RECT 62.540 152.570 65.075 152.710 ;
        RECT 62.540 152.525 62.830 152.570 ;
        RECT 43.250 152.370 43.570 152.430 ;
        RECT 64.860 152.415 65.075 152.570 ;
        RECT 65.790 152.510 66.110 152.770 ;
        RECT 67.645 152.710 67.935 152.755 ;
        RECT 68.550 152.710 68.870 152.770 ;
        RECT 67.645 152.570 68.870 152.710 ;
        RECT 69.100 152.710 69.240 152.910 ;
        RECT 69.470 152.910 73.840 153.050 ;
        RECT 69.470 152.850 69.790 152.910 ;
        RECT 70.850 152.710 71.170 152.770 ;
        RECT 69.100 152.570 71.170 152.710 ;
        RECT 67.645 152.525 67.935 152.570 ;
        RECT 68.550 152.510 68.870 152.570 ;
        RECT 70.850 152.510 71.170 152.570 ;
        RECT 71.325 152.525 71.615 152.755 ;
        RECT 71.770 152.710 72.090 152.770 ;
        RECT 73.165 152.710 73.455 152.755 ;
        RECT 71.770 152.570 73.455 152.710 ;
        RECT 73.700 152.710 73.840 152.910 ;
        RECT 74.070 152.910 74.835 153.050 ;
        RECT 74.070 152.850 74.390 152.910 ;
        RECT 74.545 152.865 74.835 152.910 ;
        RECT 92.010 153.050 92.330 153.110 ;
        RECT 92.010 152.910 93.620 153.050 ;
        RECT 92.010 152.850 92.330 152.910 ;
        RECT 75.005 152.710 75.295 152.755 ;
        RECT 73.700 152.570 75.295 152.710 ;
        RECT 41.500 152.230 43.570 152.370 ;
        RECT 43.250 152.170 43.570 152.230 ;
        RECT 57.525 152.370 57.815 152.415 ;
        RECT 60.680 152.370 60.970 152.415 ;
        RECT 63.940 152.370 64.230 152.415 ;
        RECT 57.525 152.230 64.230 152.370 ;
        RECT 57.525 152.185 57.815 152.230 ;
        RECT 60.680 152.185 60.970 152.230 ;
        RECT 63.940 152.185 64.230 152.230 ;
        RECT 64.860 152.370 65.150 152.415 ;
        RECT 66.720 152.370 67.010 152.415 ;
        RECT 64.860 152.230 67.010 152.370 ;
        RECT 71.400 152.370 71.540 152.525 ;
        RECT 71.770 152.510 72.090 152.570 ;
        RECT 73.165 152.525 73.455 152.570 ;
        RECT 75.005 152.525 75.295 152.570 ;
        RECT 90.600 152.710 90.890 152.755 ;
        RECT 93.480 152.710 93.620 152.910 ;
        RECT 93.850 152.850 94.170 153.110 ;
        RECT 104.430 152.850 104.750 153.110 ;
        RECT 105.440 153.050 105.580 153.190 ;
        RECT 107.280 153.050 107.420 153.590 ;
        RECT 109.950 153.530 110.270 153.590 ;
        RECT 108.110 153.390 108.430 153.450 ;
        RECT 114.550 153.390 114.870 153.450 ;
        RECT 108.110 153.250 114.870 153.390 ;
        RECT 108.110 153.190 108.430 153.250 ;
        RECT 114.550 153.190 114.870 153.250 ;
        RECT 105.440 152.910 107.420 153.050 ;
        RECT 95.705 152.710 95.995 152.755 ;
        RECT 90.600 152.570 93.135 152.710 ;
        RECT 93.480 152.570 95.995 152.710 ;
        RECT 90.600 152.525 90.890 152.570 ;
        RECT 72.230 152.370 72.550 152.430 ;
        RECT 73.610 152.370 73.930 152.430 ;
        RECT 87.870 152.370 88.190 152.430 ;
        RECT 92.920 152.415 93.135 152.570 ;
        RECT 95.705 152.525 95.995 152.570 ;
        RECT 103.525 152.710 103.815 152.755 ;
        RECT 103.525 152.570 106.500 152.710 ;
        RECT 103.525 152.525 103.815 152.570 ;
        RECT 71.400 152.230 73.930 152.370 ;
        RECT 64.860 152.185 65.150 152.230 ;
        RECT 66.720 152.185 67.010 152.230 ;
        RECT 72.230 152.170 72.550 152.230 ;
        RECT 73.610 152.170 73.930 152.230 ;
        RECT 74.620 152.230 88.190 152.370 ;
        RECT 41.870 152.030 42.190 152.090 ;
        RECT 50.610 152.030 50.930 152.090 ;
        RECT 58.890 152.075 59.210 152.090 ;
        RECT 41.040 151.890 50.930 152.030 ;
        RECT 34.970 151.830 35.290 151.890 ;
        RECT 39.585 151.845 39.875 151.890 ;
        RECT 41.870 151.830 42.190 151.890 ;
        RECT 50.610 151.830 50.930 151.890 ;
        RECT 58.675 151.845 59.210 152.075 ;
        RECT 58.890 151.830 59.210 151.845 ;
        RECT 70.390 152.030 70.710 152.090 ;
        RECT 74.620 152.030 74.760 152.230 ;
        RECT 87.870 152.170 88.190 152.230 ;
        RECT 88.740 152.370 89.030 152.415 ;
        RECT 92.000 152.370 92.290 152.415 ;
        RECT 92.920 152.370 93.210 152.415 ;
        RECT 94.780 152.370 95.070 152.415 ;
        RECT 88.740 152.230 92.700 152.370 ;
        RECT 88.740 152.185 89.030 152.230 ;
        RECT 92.000 152.185 92.290 152.230 ;
        RECT 70.390 151.890 74.760 152.030 ;
        RECT 70.390 151.830 70.710 151.890 ;
        RECT 74.990 151.830 75.310 152.090 ;
        RECT 86.490 152.075 86.810 152.090 ;
        RECT 86.490 151.845 87.025 152.075 ;
        RECT 92.560 152.030 92.700 152.230 ;
        RECT 92.920 152.230 95.070 152.370 ;
        RECT 92.920 152.185 93.210 152.230 ;
        RECT 94.780 152.185 95.070 152.230 ;
        RECT 104.890 152.170 105.210 152.430 ;
        RECT 106.360 152.370 106.500 152.570 ;
        RECT 106.730 152.510 107.050 152.770 ;
        RECT 107.280 152.755 107.420 152.910 ;
        RECT 109.950 153.050 110.270 153.110 ;
        RECT 116.390 153.050 116.710 153.110 ;
        RECT 109.950 152.910 111.100 153.050 ;
        RECT 109.950 152.850 110.270 152.910 ;
        RECT 107.205 152.525 107.495 152.755 ;
        RECT 107.650 152.510 107.970 152.770 ;
        RECT 108.570 152.510 108.890 152.770 ;
        RECT 109.490 152.710 109.810 152.770 ;
        RECT 110.960 152.755 111.100 152.910 ;
        RECT 111.420 152.910 116.710 153.050 ;
        RECT 111.420 152.755 111.560 152.910 ;
        RECT 116.390 152.850 116.710 152.910 ;
        RECT 110.425 152.710 110.715 152.755 ;
        RECT 109.490 152.570 110.715 152.710 ;
        RECT 109.490 152.510 109.810 152.570 ;
        RECT 110.425 152.525 110.715 152.570 ;
        RECT 110.885 152.525 111.175 152.755 ;
        RECT 111.345 152.525 111.635 152.755 ;
        RECT 112.265 152.710 112.555 152.755 ;
        RECT 119.610 152.710 119.930 152.770 ;
        RECT 111.880 152.570 112.555 152.710 ;
        RECT 109.045 152.370 109.335 152.415 ;
        RECT 106.360 152.230 109.335 152.370 ;
        RECT 109.045 152.185 109.335 152.230 ;
        RECT 93.850 152.030 94.170 152.090 ;
        RECT 92.560 151.890 94.170 152.030 ;
        RECT 86.490 151.830 86.810 151.845 ;
        RECT 93.850 151.830 94.170 151.890 ;
        RECT 101.670 152.030 101.990 152.090 ;
        RECT 102.605 152.030 102.895 152.075 ;
        RECT 101.670 151.890 102.895 152.030 ;
        RECT 101.670 151.830 101.990 151.890 ;
        RECT 102.605 151.845 102.895 151.890 ;
        RECT 105.350 151.830 105.670 152.090 ;
        RECT 108.570 152.030 108.890 152.090 ;
        RECT 111.880 152.030 112.020 152.570 ;
        RECT 112.265 152.525 112.555 152.570 ;
        RECT 112.800 152.570 119.930 152.710 ;
        RECT 108.570 151.890 112.020 152.030 ;
        RECT 112.250 152.030 112.570 152.090 ;
        RECT 112.800 152.030 112.940 152.570 ;
        RECT 119.610 152.510 119.930 152.570 ;
        RECT 120.545 152.525 120.835 152.755 ;
        RECT 115.930 152.370 116.250 152.430 ;
        RECT 120.620 152.370 120.760 152.525 ;
        RECT 115.930 152.230 120.760 152.370 ;
        RECT 115.930 152.170 116.250 152.230 ;
        RECT 112.250 151.890 112.940 152.030 ;
        RECT 118.230 152.030 118.550 152.090 ;
        RECT 119.165 152.030 119.455 152.075 ;
        RECT 118.230 151.890 119.455 152.030 ;
        RECT 108.570 151.830 108.890 151.890 ;
        RECT 112.250 151.830 112.570 151.890 ;
        RECT 118.230 151.830 118.550 151.890 ;
        RECT 119.165 151.845 119.455 151.890 ;
        RECT 121.465 152.030 121.755 152.075 ;
        RECT 123.290 152.030 123.610 152.090 ;
        RECT 121.465 151.890 123.610 152.030 ;
        RECT 121.465 151.845 121.755 151.890 ;
        RECT 123.290 151.830 123.610 151.890 ;
        RECT 14.660 151.210 127.820 151.690 ;
        RECT 33.590 150.810 33.910 151.070 ;
        RECT 36.825 151.010 37.115 151.055 ;
        RECT 37.270 151.010 37.590 151.070 ;
        RECT 36.825 150.870 37.590 151.010 ;
        RECT 36.825 150.825 37.115 150.870 ;
        RECT 37.270 150.810 37.590 150.870 ;
        RECT 60.745 150.825 61.035 151.055 ;
        RECT 61.190 151.010 61.510 151.070 ;
        RECT 61.665 151.010 61.955 151.055 ;
        RECT 61.190 150.870 61.955 151.010 ;
        RECT 18.820 150.670 19.110 150.715 ;
        RECT 20.250 150.670 20.570 150.730 ;
        RECT 22.080 150.670 22.370 150.715 ;
        RECT 18.820 150.530 22.370 150.670 ;
        RECT 18.820 150.485 19.110 150.530 ;
        RECT 20.250 150.470 20.570 150.530 ;
        RECT 22.080 150.485 22.370 150.530 ;
        RECT 23.000 150.670 23.290 150.715 ;
        RECT 24.860 150.670 25.150 150.715 ;
        RECT 23.000 150.530 25.150 150.670 ;
        RECT 23.000 150.485 23.290 150.530 ;
        RECT 24.860 150.485 25.150 150.530 ;
        RECT 31.290 150.670 31.610 150.730 ;
        RECT 58.445 150.670 58.735 150.715 ;
        RECT 31.290 150.530 43.940 150.670 ;
        RECT 20.680 150.330 20.970 150.375 ;
        RECT 23.000 150.330 23.215 150.485 ;
        RECT 31.290 150.470 31.610 150.530 ;
        RECT 20.680 150.190 23.215 150.330 ;
        RECT 29.910 150.330 30.230 150.390 ;
        RECT 33.145 150.330 33.435 150.375 ;
        RECT 29.910 150.190 33.435 150.330 ;
        RECT 20.680 150.145 20.970 150.190 ;
        RECT 29.910 150.130 30.230 150.190 ;
        RECT 33.145 150.145 33.435 150.190 ;
        RECT 35.890 150.130 36.210 150.390 ;
        RECT 41.870 150.330 42.190 150.390 ;
        RECT 42.805 150.330 43.095 150.375 ;
        RECT 41.870 150.190 43.095 150.330 ;
        RECT 41.870 150.130 42.190 150.190 ;
        RECT 42.805 150.145 43.095 150.190 ;
        RECT 43.250 150.130 43.570 150.390 ;
        RECT 43.800 150.375 43.940 150.530 ;
        RECT 53.920 150.530 58.735 150.670 ;
        RECT 53.920 150.390 54.060 150.530 ;
        RECT 58.445 150.485 58.735 150.530 ;
        RECT 43.725 150.145 44.015 150.375 ;
        RECT 44.645 150.330 44.935 150.375 ;
        RECT 45.090 150.330 45.410 150.390 ;
        RECT 44.645 150.190 45.410 150.330 ;
        RECT 44.645 150.145 44.935 150.190 ;
        RECT 45.090 150.130 45.410 150.190 ;
        RECT 48.785 150.145 49.075 150.375 ;
        RECT 16.815 149.990 17.105 150.035 ;
        RECT 22.550 149.990 22.870 150.050 ;
        RECT 16.815 149.850 22.870 149.990 ;
        RECT 16.815 149.805 17.105 149.850 ;
        RECT 22.550 149.790 22.870 149.850 ;
        RECT 23.945 149.990 24.235 150.035 ;
        RECT 24.850 149.990 25.170 150.050 ;
        RECT 23.945 149.850 25.170 149.990 ;
        RECT 23.945 149.805 24.235 149.850 ;
        RECT 24.850 149.790 25.170 149.850 ;
        RECT 25.785 149.990 26.075 150.035 ;
        RECT 36.350 149.990 36.670 150.050 ;
        RECT 25.785 149.850 36.670 149.990 ;
        RECT 48.860 149.990 49.000 150.145 ;
        RECT 49.690 150.130 50.010 150.390 ;
        RECT 50.150 150.130 50.470 150.390 ;
        RECT 52.925 150.145 53.215 150.375 ;
        RECT 50.610 149.990 50.930 150.050 ;
        RECT 48.860 149.850 50.930 149.990 ;
        RECT 53.000 149.990 53.140 150.145 ;
        RECT 53.370 150.130 53.690 150.390 ;
        RECT 53.830 150.130 54.150 150.390 ;
        RECT 54.765 150.330 55.055 150.375 ;
        RECT 56.590 150.330 56.910 150.390 ;
        RECT 54.765 150.190 56.910 150.330 ;
        RECT 54.765 150.145 55.055 150.190 ;
        RECT 56.590 150.130 56.910 150.190 ;
        RECT 58.890 150.130 59.210 150.390 ;
        RECT 60.820 150.330 60.960 150.825 ;
        RECT 61.190 150.810 61.510 150.870 ;
        RECT 61.665 150.825 61.955 150.870 ;
        RECT 64.885 151.010 65.175 151.055 ;
        RECT 65.790 151.010 66.110 151.070 ;
        RECT 64.885 150.870 66.110 151.010 ;
        RECT 64.885 150.825 65.175 150.870 ;
        RECT 65.790 150.810 66.110 150.870 ;
        RECT 68.565 151.010 68.855 151.055 ;
        RECT 86.045 151.010 86.335 151.055 ;
        RECT 86.490 151.010 86.810 151.070 ;
        RECT 88.345 151.010 88.635 151.055 ;
        RECT 92.945 151.010 93.235 151.055 ;
        RECT 93.390 151.010 93.710 151.070 ;
        RECT 68.565 150.870 71.540 151.010 ;
        RECT 68.565 150.825 68.855 150.870 ;
        RECT 62.585 150.330 62.875 150.375 ;
        RECT 60.820 150.190 62.875 150.330 ;
        RECT 62.585 150.145 62.875 150.190 ;
        RECT 63.950 150.130 64.270 150.390 ;
        RECT 67.645 150.330 67.935 150.375 ;
        RECT 69.470 150.330 69.790 150.390 ;
        RECT 67.645 150.190 69.790 150.330 ;
        RECT 67.645 150.145 67.935 150.190 ;
        RECT 69.470 150.130 69.790 150.190 ;
        RECT 70.850 150.130 71.170 150.390 ;
        RECT 54.290 149.990 54.610 150.050 ;
        RECT 53.000 149.850 54.610 149.990 ;
        RECT 25.785 149.805 26.075 149.850 ;
        RECT 36.350 149.790 36.670 149.850 ;
        RECT 50.610 149.790 50.930 149.850 ;
        RECT 54.290 149.790 54.610 149.850 ;
        RECT 57.985 149.990 58.275 150.035 ;
        RECT 65.790 149.990 66.110 150.050 ;
        RECT 57.985 149.850 65.100 149.990 ;
        RECT 57.985 149.805 58.275 149.850 ;
        RECT 64.960 149.710 65.100 149.850 ;
        RECT 65.790 149.850 71.080 149.990 ;
        RECT 65.790 149.790 66.110 149.850 ;
        RECT 20.680 149.650 20.970 149.695 ;
        RECT 23.460 149.650 23.750 149.695 ;
        RECT 25.320 149.650 25.610 149.695 ;
        RECT 20.680 149.510 25.610 149.650 ;
        RECT 20.680 149.465 20.970 149.510 ;
        RECT 23.460 149.465 23.750 149.510 ;
        RECT 25.320 149.465 25.610 149.510 ;
        RECT 51.085 149.650 51.375 149.695 ;
        RECT 60.270 149.650 60.590 149.710 ;
        RECT 51.085 149.510 60.590 149.650 ;
        RECT 51.085 149.465 51.375 149.510 ;
        RECT 60.270 149.450 60.590 149.510 ;
        RECT 64.870 149.650 65.190 149.710 ;
        RECT 70.940 149.650 71.080 149.850 ;
        RECT 71.400 149.650 71.540 150.870 ;
        RECT 86.045 150.870 87.180 151.010 ;
        RECT 86.045 150.825 86.335 150.870 ;
        RECT 86.490 150.810 86.810 150.870 ;
        RECT 73.165 150.670 73.455 150.715 ;
        RECT 74.990 150.670 75.310 150.730 ;
        RECT 75.465 150.670 75.755 150.715 ;
        RECT 73.165 150.530 75.755 150.670 ;
        RECT 73.165 150.485 73.455 150.530 ;
        RECT 74.990 150.470 75.310 150.530 ;
        RECT 75.465 150.485 75.755 150.530 ;
        RECT 77.305 150.670 77.595 150.715 ;
        RECT 77.305 150.530 85.340 150.670 ;
        RECT 77.305 150.485 77.595 150.530 ;
        RECT 75.910 150.330 76.230 150.390 ;
        RECT 78.685 150.330 78.975 150.375 ;
        RECT 75.910 150.190 78.975 150.330 ;
        RECT 75.910 150.130 76.230 150.190 ;
        RECT 78.685 150.145 78.975 150.190 ;
        RECT 80.050 150.130 80.370 150.390 ;
        RECT 85.200 150.050 85.340 150.530 ;
        RECT 86.030 150.330 86.350 150.390 ;
        RECT 86.505 150.330 86.795 150.375 ;
        RECT 86.030 150.190 86.795 150.330 ;
        RECT 86.030 150.130 86.350 150.190 ;
        RECT 86.505 150.145 86.795 150.190 ;
        RECT 79.590 149.790 79.910 150.050 ;
        RECT 85.110 149.790 85.430 150.050 ;
        RECT 78.210 149.650 78.530 149.710 ;
        RECT 64.870 149.510 70.620 149.650 ;
        RECT 70.940 149.510 78.530 149.650 ;
        RECT 87.040 149.650 87.180 150.870 ;
        RECT 88.345 150.870 92.240 151.010 ;
        RECT 88.345 150.825 88.635 150.870 ;
        RECT 92.100 150.495 92.240 150.870 ;
        RECT 92.945 150.870 93.710 151.010 ;
        RECT 92.945 150.825 93.235 150.870 ;
        RECT 93.390 150.810 93.710 150.870 ;
        RECT 93.850 150.810 94.170 151.070 ;
        RECT 104.890 151.010 105.210 151.070 ;
        RECT 107.205 151.010 107.495 151.055 ;
        RECT 94.400 150.870 104.660 151.010 ;
        RECT 90.645 150.145 90.935 150.375 ;
        RECT 92.025 150.265 92.315 150.495 ;
        RECT 94.400 150.375 94.540 150.870 ;
        RECT 95.690 150.670 96.010 150.730 ;
        RECT 98.105 150.670 98.395 150.715 ;
        RECT 101.345 150.670 101.995 150.715 ;
        RECT 95.690 150.530 101.995 150.670 ;
        RECT 95.690 150.470 96.010 150.530 ;
        RECT 98.105 150.485 98.695 150.530 ;
        RECT 101.345 150.485 101.995 150.530 ;
        RECT 103.510 150.670 103.830 150.730 ;
        RECT 103.985 150.670 104.275 150.715 ;
        RECT 103.510 150.530 104.275 150.670 ;
        RECT 104.520 150.670 104.660 150.870 ;
        RECT 104.890 150.870 107.495 151.010 ;
        RECT 104.890 150.810 105.210 150.870 ;
        RECT 107.205 150.825 107.495 150.870 ;
        RECT 116.850 150.670 117.170 150.730 ;
        RECT 104.520 150.530 117.170 150.670 ;
        RECT 94.325 150.330 94.615 150.375 ;
        RECT 92.560 150.190 94.615 150.330 ;
        RECT 90.720 149.990 90.860 150.145 ;
        RECT 92.560 149.990 92.700 150.190 ;
        RECT 94.325 150.145 94.615 150.190 ;
        RECT 98.405 150.170 98.695 150.485 ;
        RECT 103.510 150.470 103.830 150.530 ;
        RECT 103.985 150.485 104.275 150.530 ;
        RECT 116.850 150.470 117.170 150.530 ;
        RECT 117.425 150.670 117.715 150.715 ;
        RECT 118.230 150.670 118.550 150.730 ;
        RECT 120.665 150.670 121.315 150.715 ;
        RECT 117.425 150.530 121.315 150.670 ;
        RECT 117.425 150.485 118.015 150.530 ;
        RECT 99.485 150.330 99.775 150.375 ;
        RECT 103.065 150.330 103.355 150.375 ;
        RECT 104.900 150.330 105.190 150.375 ;
        RECT 99.485 150.190 105.190 150.330 ;
        RECT 99.485 150.145 99.775 150.190 ;
        RECT 103.065 150.145 103.355 150.190 ;
        RECT 104.900 150.145 105.190 150.190 ;
        RECT 108.110 150.330 108.430 150.390 ;
        RECT 108.585 150.330 108.875 150.375 ;
        RECT 108.110 150.190 108.875 150.330 ;
        RECT 108.110 150.130 108.430 150.190 ;
        RECT 108.585 150.145 108.875 150.190 ;
        RECT 109.045 150.145 109.335 150.375 ;
        RECT 109.505 150.145 109.795 150.375 ;
        RECT 109.950 150.330 110.270 150.390 ;
        RECT 110.425 150.330 110.715 150.375 ;
        RECT 109.950 150.190 110.715 150.330 ;
        RECT 105.365 149.990 105.655 150.035 ;
        RECT 90.720 149.850 92.700 149.990 ;
        RECT 94.400 149.850 105.655 149.990 ;
        RECT 94.400 149.710 94.540 149.850 ;
        RECT 105.365 149.805 105.655 149.850 ;
        RECT 107.650 149.990 107.970 150.050 ;
        RECT 109.120 149.990 109.260 150.145 ;
        RECT 107.650 149.850 109.260 149.990 ;
        RECT 109.580 149.990 109.720 150.145 ;
        RECT 109.950 150.130 110.270 150.190 ;
        RECT 110.425 150.145 110.715 150.190 ;
        RECT 117.725 150.170 118.015 150.485 ;
        RECT 118.230 150.470 118.550 150.530 ;
        RECT 120.665 150.485 121.315 150.530 ;
        RECT 123.290 150.470 123.610 150.730 ;
        RECT 118.805 150.330 119.095 150.375 ;
        RECT 122.385 150.330 122.675 150.375 ;
        RECT 124.220 150.330 124.510 150.375 ;
        RECT 118.805 150.190 124.510 150.330 ;
        RECT 118.805 150.145 119.095 150.190 ;
        RECT 122.385 150.145 122.675 150.190 ;
        RECT 124.220 150.145 124.510 150.190 ;
        RECT 111.345 149.990 111.635 150.035 ;
        RECT 115.945 149.990 116.235 150.035 ;
        RECT 109.580 149.850 116.235 149.990 ;
        RECT 107.650 149.790 107.970 149.850 ;
        RECT 93.850 149.650 94.170 149.710 ;
        RECT 87.040 149.510 94.170 149.650 ;
        RECT 64.870 149.450 65.190 149.510 ;
        RECT 40.950 149.310 41.270 149.370 ;
        RECT 41.425 149.310 41.715 149.355 ;
        RECT 40.950 149.170 41.715 149.310 ;
        RECT 40.950 149.110 41.270 149.170 ;
        RECT 41.425 149.125 41.715 149.170 ;
        RECT 44.170 149.310 44.490 149.370 ;
        RECT 48.785 149.310 49.075 149.355 ;
        RECT 44.170 149.170 49.075 149.310 ;
        RECT 44.170 149.110 44.490 149.170 ;
        RECT 48.785 149.125 49.075 149.170 ;
        RECT 51.530 149.110 51.850 149.370 ;
        RECT 65.330 149.310 65.650 149.370 ;
        RECT 69.945 149.310 70.235 149.355 ;
        RECT 65.330 149.170 70.235 149.310 ;
        RECT 70.480 149.310 70.620 149.510 ;
        RECT 78.210 149.450 78.530 149.510 ;
        RECT 93.850 149.450 94.170 149.510 ;
        RECT 94.310 149.450 94.630 149.710 ;
        RECT 99.485 149.650 99.775 149.695 ;
        RECT 102.605 149.650 102.895 149.695 ;
        RECT 104.495 149.650 104.785 149.695 ;
        RECT 99.485 149.510 104.785 149.650 ;
        RECT 109.120 149.650 109.260 149.850 ;
        RECT 111.345 149.805 111.635 149.850 ;
        RECT 115.945 149.805 116.235 149.850 ;
        RECT 124.685 149.990 124.975 150.035 ;
        RECT 126.050 149.990 126.370 150.050 ;
        RECT 124.685 149.850 126.370 149.990 ;
        RECT 124.685 149.805 124.975 149.850 ;
        RECT 126.050 149.790 126.370 149.850 ;
        RECT 111.790 149.650 112.110 149.710 ;
        RECT 109.120 149.510 112.110 149.650 ;
        RECT 99.485 149.465 99.775 149.510 ;
        RECT 102.605 149.465 102.895 149.510 ;
        RECT 104.495 149.465 104.785 149.510 ;
        RECT 111.790 149.450 112.110 149.510 ;
        RECT 118.805 149.650 119.095 149.695 ;
        RECT 121.925 149.650 122.215 149.695 ;
        RECT 123.815 149.650 124.105 149.695 ;
        RECT 118.805 149.510 124.105 149.650 ;
        RECT 118.805 149.465 119.095 149.510 ;
        RECT 121.925 149.465 122.215 149.510 ;
        RECT 123.815 149.465 124.105 149.510 ;
        RECT 71.785 149.310 72.075 149.355 ;
        RECT 70.480 149.170 72.075 149.310 ;
        RECT 65.330 149.110 65.650 149.170 ;
        RECT 69.945 149.125 70.235 149.170 ;
        RECT 71.785 149.125 72.075 149.170 ;
        RECT 75.910 149.310 76.230 149.370 ;
        RECT 77.765 149.310 78.055 149.355 ;
        RECT 75.910 149.170 78.055 149.310 ;
        RECT 75.910 149.110 76.230 149.170 ;
        RECT 77.765 149.125 78.055 149.170 ;
        RECT 80.065 149.310 80.355 149.355 ;
        RECT 81.890 149.310 82.210 149.370 ;
        RECT 80.065 149.170 82.210 149.310 ;
        RECT 80.065 149.125 80.355 149.170 ;
        RECT 81.890 149.110 82.210 149.170 ;
        RECT 90.185 149.310 90.475 149.355 ;
        RECT 90.630 149.310 90.950 149.370 ;
        RECT 90.185 149.170 90.950 149.310 ;
        RECT 90.185 149.125 90.475 149.170 ;
        RECT 90.630 149.110 90.950 149.170 ;
        RECT 96.610 149.110 96.930 149.370 ;
        RECT 114.090 149.110 114.410 149.370 ;
        RECT 14.660 148.490 127.820 148.970 ;
        RECT 24.850 148.090 25.170 148.350 ;
        RECT 35.890 148.290 36.210 148.350 ;
        RECT 48.785 148.290 49.075 148.335 ;
        RECT 49.230 148.290 49.550 148.350 ;
        RECT 35.890 148.150 43.020 148.290 ;
        RECT 35.890 148.090 36.210 148.150 ;
        RECT 23.945 147.765 24.235 147.995 ;
        RECT 28.530 147.950 28.850 148.010 ;
        RECT 28.530 147.810 34.740 147.950 ;
        RECT 21.170 147.410 21.490 147.670 ;
        RECT 24.020 147.270 24.160 147.765 ;
        RECT 28.530 147.750 28.850 147.810 ;
        RECT 32.685 147.610 32.975 147.655 ;
        RECT 34.050 147.610 34.370 147.670 ;
        RECT 26.320 147.470 31.980 147.610 ;
        RECT 25.785 147.270 26.075 147.315 ;
        RECT 24.020 147.130 26.075 147.270 ;
        RECT 25.785 147.085 26.075 147.130 ;
        RECT 22.105 146.930 22.395 146.975 ;
        RECT 23.010 146.930 23.330 146.990 ;
        RECT 26.320 146.930 26.460 147.470 ;
        RECT 28.085 147.270 28.375 147.315 ;
        RECT 28.085 147.130 30.140 147.270 ;
        RECT 28.085 147.085 28.375 147.130 ;
        RECT 22.105 146.790 26.460 146.930 ;
        RECT 22.105 146.745 22.395 146.790 ;
        RECT 23.010 146.730 23.330 146.790 ;
        RECT 21.645 146.590 21.935 146.635 ;
        RECT 22.550 146.590 22.870 146.650 ;
        RECT 28.530 146.590 28.850 146.650 ;
        RECT 21.645 146.450 28.850 146.590 ;
        RECT 21.645 146.405 21.935 146.450 ;
        RECT 22.550 146.390 22.870 146.450 ;
        RECT 28.530 146.390 28.850 146.450 ;
        RECT 28.990 146.390 29.310 146.650 ;
        RECT 29.465 146.590 29.755 146.635 ;
        RECT 30.000 146.590 30.140 147.130 ;
        RECT 31.290 147.070 31.610 147.330 ;
        RECT 31.840 146.975 31.980 147.470 ;
        RECT 32.685 147.470 34.370 147.610 ;
        RECT 34.600 147.610 34.740 147.810 ;
        RECT 36.900 147.810 42.100 147.950 ;
        RECT 36.900 147.610 37.040 147.810 ;
        RECT 34.600 147.470 37.040 147.610 ;
        RECT 37.360 147.470 41.640 147.610 ;
        RECT 32.685 147.425 32.975 147.470 ;
        RECT 34.050 147.410 34.370 147.470 ;
        RECT 35.890 147.070 36.210 147.330 ;
        RECT 37.360 147.315 37.500 147.470 ;
        RECT 41.500 147.315 41.640 147.470 ;
        RECT 41.960 147.315 42.100 147.810 ;
        RECT 42.880 147.315 43.020 148.150 ;
        RECT 48.785 148.150 49.550 148.290 ;
        RECT 48.785 148.105 49.075 148.150 ;
        RECT 49.230 148.090 49.550 148.150 ;
        RECT 50.610 148.290 50.930 148.350 ;
        RECT 53.385 148.290 53.675 148.335 ;
        RECT 50.610 148.150 53.675 148.290 ;
        RECT 50.610 148.090 50.930 148.150 ;
        RECT 53.385 148.105 53.675 148.150 ;
        RECT 54.750 148.290 55.070 148.350 ;
        RECT 73.610 148.290 73.930 148.350 ;
        RECT 54.750 148.150 73.930 148.290 ;
        RECT 54.750 148.090 55.070 148.150 ;
        RECT 73.610 148.090 73.930 148.150 ;
        RECT 80.050 148.090 80.370 148.350 ;
        RECT 85.110 148.290 85.430 148.350 ;
        RECT 85.110 148.150 95.460 148.290 ;
        RECT 85.110 148.090 85.430 148.150 ;
        RECT 49.705 147.950 49.995 147.995 ;
        RECT 57.050 147.950 57.370 148.010 ;
        RECT 78.210 147.950 78.530 148.010 ;
        RECT 83.270 147.950 83.590 148.010 ;
        RECT 49.705 147.810 57.370 147.950 ;
        RECT 49.705 147.765 49.995 147.810 ;
        RECT 57.050 147.750 57.370 147.810 ;
        RECT 57.600 147.810 66.480 147.950 ;
        RECT 48.325 147.610 48.615 147.655 ;
        RECT 52.450 147.610 52.770 147.670 ;
        RECT 48.325 147.470 52.770 147.610 ;
        RECT 48.325 147.425 48.615 147.470 ;
        RECT 52.450 147.410 52.770 147.470 ;
        RECT 53.370 147.610 53.690 147.670 ;
        RECT 57.600 147.610 57.740 147.810 ;
        RECT 53.370 147.470 57.740 147.610 ;
        RECT 60.745 147.610 61.035 147.655 ;
        RECT 64.870 147.610 65.190 147.670 ;
        RECT 60.745 147.470 65.190 147.610 ;
        RECT 53.370 147.410 53.690 147.470 ;
        RECT 36.825 147.085 37.115 147.315 ;
        RECT 37.285 147.085 37.575 147.315 ;
        RECT 37.745 147.270 38.035 147.315 ;
        RECT 40.965 147.270 41.255 147.315 ;
        RECT 37.745 147.130 41.255 147.270 ;
        RECT 37.745 147.085 38.035 147.130 ;
        RECT 40.965 147.085 41.255 147.130 ;
        RECT 41.425 147.085 41.715 147.315 ;
        RECT 41.885 147.085 42.175 147.315 ;
        RECT 42.805 147.270 43.095 147.315 ;
        RECT 44.630 147.270 44.950 147.330 ;
        RECT 42.805 147.130 44.950 147.270 ;
        RECT 42.805 147.085 43.095 147.130 ;
        RECT 31.765 146.930 32.055 146.975 ;
        RECT 36.900 146.930 37.040 147.085 ;
        RECT 39.585 146.930 39.875 146.975 ;
        RECT 31.765 146.790 37.040 146.930 ;
        RECT 37.820 146.790 39.875 146.930 ;
        RECT 31.765 146.745 32.055 146.790 ;
        RECT 29.465 146.450 30.140 146.590 ;
        RECT 36.810 146.590 37.130 146.650 ;
        RECT 37.820 146.590 37.960 146.790 ;
        RECT 39.585 146.745 39.875 146.790 ;
        RECT 36.810 146.450 37.960 146.590 ;
        RECT 38.650 146.590 38.970 146.650 ;
        RECT 39.125 146.590 39.415 146.635 ;
        RECT 38.650 146.450 39.415 146.590 ;
        RECT 41.040 146.590 41.180 147.085 ;
        RECT 41.500 146.930 41.640 147.085 ;
        RECT 44.630 147.070 44.950 147.130 ;
        RECT 48.770 147.070 49.090 147.330 ;
        RECT 51.990 147.070 52.310 147.330 ;
        RECT 54.750 147.070 55.070 147.330 ;
        RECT 55.300 147.315 55.440 147.470 ;
        RECT 60.745 147.425 61.035 147.470 ;
        RECT 64.870 147.410 65.190 147.470 ;
        RECT 55.225 147.085 55.515 147.315 ;
        RECT 55.685 147.085 55.975 147.315 ;
        RECT 56.590 147.270 56.910 147.330 ;
        RECT 65.790 147.270 66.110 147.330 ;
        RECT 56.590 147.130 66.110 147.270 ;
        RECT 66.340 147.270 66.480 147.810 ;
        RECT 76.460 147.810 83.590 147.950 ;
        RECT 70.850 147.610 71.170 147.670 ;
        RECT 70.850 147.470 72.920 147.610 ;
        RECT 70.850 147.410 71.170 147.470 ;
        RECT 66.340 147.130 71.310 147.270 ;
        RECT 43.250 146.930 43.570 146.990 ;
        RECT 41.500 146.790 43.570 146.930 ;
        RECT 43.250 146.730 43.570 146.790 ;
        RECT 47.405 146.930 47.695 146.975 ;
        RECT 51.530 146.930 51.850 146.990 ;
        RECT 47.405 146.790 51.850 146.930 ;
        RECT 55.760 146.930 55.900 147.085 ;
        RECT 56.590 147.070 56.910 147.130 ;
        RECT 65.790 147.070 66.110 147.130 ;
        RECT 58.890 146.930 59.210 146.990 ;
        RECT 61.205 146.930 61.495 146.975 ;
        RECT 55.760 146.790 61.495 146.930 ;
        RECT 71.170 146.930 71.310 147.130 ;
        RECT 72.230 147.070 72.550 147.330 ;
        RECT 72.780 147.315 72.920 147.470 ;
        RECT 76.460 147.315 76.600 147.810 ;
        RECT 78.210 147.750 78.530 147.810 ;
        RECT 83.270 147.750 83.590 147.810 ;
        RECT 89.220 147.950 89.510 147.995 ;
        RECT 92.000 147.950 92.290 147.995 ;
        RECT 93.860 147.950 94.150 147.995 ;
        RECT 89.220 147.810 94.150 147.950 ;
        RECT 95.320 147.950 95.460 148.150 ;
        RECT 95.690 148.090 96.010 148.350 ;
        RECT 96.610 148.290 96.930 148.350 ;
        RECT 103.065 148.290 103.355 148.335 ;
        RECT 103.510 148.290 103.830 148.350 ;
        RECT 96.610 148.150 100.980 148.290 ;
        RECT 96.610 148.090 96.930 148.150 ;
        RECT 95.320 147.810 97.300 147.950 ;
        RECT 89.220 147.765 89.510 147.810 ;
        RECT 92.000 147.765 92.290 147.810 ;
        RECT 93.860 147.765 94.150 147.810 ;
        RECT 86.490 147.610 86.810 147.670 ;
        RECT 77.380 147.470 86.810 147.610 ;
        RECT 77.380 147.315 77.520 147.470 ;
        RECT 86.490 147.410 86.810 147.470 ;
        RECT 91.090 147.610 91.410 147.670 ;
        RECT 97.160 147.655 97.300 147.810 ;
        RECT 100.305 147.765 100.595 147.995 ;
        RECT 100.840 147.950 100.980 148.150 ;
        RECT 103.065 148.150 103.830 148.290 ;
        RECT 103.065 148.105 103.355 148.150 ;
        RECT 103.510 148.090 103.830 148.150 ;
        RECT 103.985 148.290 104.275 148.335 ;
        RECT 104.430 148.290 104.750 148.350 ;
        RECT 103.985 148.150 104.750 148.290 ;
        RECT 103.985 148.105 104.275 148.150 ;
        RECT 104.430 148.090 104.750 148.150 ;
        RECT 106.270 148.090 106.590 148.350 ;
        RECT 115.930 148.090 116.250 148.350 ;
        RECT 120.500 147.950 120.790 147.995 ;
        RECT 123.280 147.950 123.570 147.995 ;
        RECT 125.140 147.950 125.430 147.995 ;
        RECT 100.840 147.810 109.260 147.950 ;
        RECT 92.485 147.610 92.775 147.655 ;
        RECT 91.090 147.470 92.775 147.610 ;
        RECT 91.090 147.410 91.410 147.470 ;
        RECT 92.485 147.425 92.775 147.470 ;
        RECT 97.085 147.425 97.375 147.655 ;
        RECT 72.705 147.085 72.995 147.315 ;
        RECT 76.385 147.085 76.675 147.315 ;
        RECT 77.305 147.085 77.595 147.315 ;
        RECT 77.765 147.085 78.055 147.315 ;
        RECT 78.210 147.270 78.530 147.330 ;
        RECT 80.050 147.270 80.370 147.330 ;
        RECT 81.445 147.270 81.735 147.315 ;
        RECT 78.210 147.130 81.735 147.270 ;
        RECT 77.840 146.930 77.980 147.085 ;
        RECT 78.210 147.070 78.530 147.130 ;
        RECT 80.050 147.070 80.370 147.130 ;
        RECT 81.445 147.085 81.735 147.130 ;
        RECT 81.905 147.085 82.195 147.315 ;
        RECT 81.980 146.930 82.120 147.085 ;
        RECT 82.350 147.070 82.670 147.330 ;
        RECT 83.270 147.070 83.590 147.330 ;
        RECT 89.220 147.270 89.510 147.315 ;
        RECT 89.220 147.130 91.755 147.270 ;
        RECT 89.220 147.085 89.510 147.130 ;
        RECT 82.810 146.930 83.130 146.990 ;
        RECT 90.630 146.975 90.950 146.990 ;
        RECT 71.170 146.790 83.130 146.930 ;
        RECT 47.405 146.745 47.695 146.790 ;
        RECT 51.530 146.730 51.850 146.790 ;
        RECT 58.890 146.730 59.210 146.790 ;
        RECT 61.205 146.745 61.495 146.790 ;
        RECT 41.870 146.590 42.190 146.650 ;
        RECT 41.040 146.450 42.190 146.590 ;
        RECT 29.465 146.405 29.755 146.450 ;
        RECT 36.810 146.390 37.130 146.450 ;
        RECT 38.650 146.390 38.970 146.450 ;
        RECT 39.125 146.405 39.415 146.450 ;
        RECT 41.870 146.390 42.190 146.450 ;
        RECT 49.690 146.590 50.010 146.650 ;
        RECT 51.085 146.590 51.375 146.635 ;
        RECT 49.690 146.450 51.375 146.590 ;
        RECT 49.690 146.390 50.010 146.450 ;
        RECT 51.085 146.405 51.375 146.450 ;
        RECT 59.350 146.590 59.670 146.650 ;
        RECT 61.665 146.590 61.955 146.635 ;
        RECT 59.350 146.450 61.955 146.590 ;
        RECT 59.350 146.390 59.670 146.450 ;
        RECT 61.665 146.405 61.955 146.450 ;
        RECT 63.505 146.590 63.795 146.635 ;
        RECT 63.950 146.590 64.270 146.650 ;
        RECT 71.400 146.635 71.540 146.790 ;
        RECT 82.810 146.730 83.130 146.790 ;
        RECT 87.360 146.930 87.650 146.975 ;
        RECT 90.620 146.930 90.950 146.975 ;
        RECT 87.360 146.790 90.950 146.930 ;
        RECT 87.360 146.745 87.650 146.790 ;
        RECT 90.620 146.745 90.950 146.790 ;
        RECT 91.540 146.975 91.755 147.130 ;
        RECT 94.310 147.070 94.630 147.330 ;
        RECT 95.230 147.070 95.550 147.330 ;
        RECT 98.465 147.085 98.755 147.315 ;
        RECT 100.380 147.270 100.520 147.765 ;
        RECT 103.050 147.610 103.370 147.670 ;
        RECT 105.825 147.610 106.115 147.655 ;
        RECT 103.050 147.470 106.115 147.610 ;
        RECT 103.050 147.410 103.370 147.470 ;
        RECT 105.825 147.425 106.115 147.470 ;
        RECT 107.650 147.610 107.970 147.670 ;
        RECT 107.650 147.470 108.800 147.610 ;
        RECT 107.650 147.410 107.970 147.470 ;
        RECT 102.145 147.270 102.435 147.315 ;
        RECT 100.380 147.130 102.435 147.270 ;
        RECT 102.145 147.085 102.435 147.130 ;
        RECT 104.905 147.270 105.195 147.315 ;
        RECT 105.350 147.270 105.670 147.330 ;
        RECT 104.905 147.130 105.670 147.270 ;
        RECT 104.905 147.085 105.195 147.130 ;
        RECT 91.540 146.930 91.830 146.975 ;
        RECT 93.400 146.930 93.690 146.975 ;
        RECT 91.540 146.790 93.690 146.930 ;
        RECT 91.540 146.745 91.830 146.790 ;
        RECT 93.400 146.745 93.690 146.790 ;
        RECT 93.850 146.930 94.170 146.990 ;
        RECT 98.540 146.930 98.680 147.085 ;
        RECT 105.350 147.070 105.670 147.130 ;
        RECT 108.110 147.070 108.430 147.330 ;
        RECT 108.660 147.315 108.800 147.470 ;
        RECT 109.120 147.315 109.260 147.810 ;
        RECT 120.500 147.810 125.430 147.950 ;
        RECT 120.500 147.765 120.790 147.810 ;
        RECT 123.280 147.765 123.570 147.810 ;
        RECT 125.140 147.765 125.430 147.810 ;
        RECT 113.170 147.410 113.490 147.670 ;
        RECT 108.585 147.085 108.875 147.315 ;
        RECT 109.045 147.085 109.335 147.315 ;
        RECT 109.950 147.270 110.270 147.330 ;
        RECT 112.250 147.270 112.570 147.330 ;
        RECT 109.950 147.130 112.570 147.270 ;
        RECT 109.950 147.070 110.270 147.130 ;
        RECT 112.250 147.070 112.570 147.130 ;
        RECT 114.105 147.085 114.395 147.315 ;
        RECT 120.500 147.270 120.790 147.315 ;
        RECT 120.500 147.130 123.035 147.270 ;
        RECT 120.500 147.085 120.790 147.130 ;
        RECT 93.850 146.790 98.680 146.930 ;
        RECT 106.285 146.930 106.575 146.975 ;
        RECT 106.745 146.930 107.035 146.975 ;
        RECT 114.180 146.930 114.320 147.085 ;
        RECT 106.285 146.790 107.035 146.930 ;
        RECT 90.630 146.730 90.950 146.745 ;
        RECT 93.850 146.730 94.170 146.790 ;
        RECT 106.285 146.745 106.575 146.790 ;
        RECT 106.745 146.745 107.035 146.790 ;
        RECT 107.280 146.790 114.320 146.930 ;
        RECT 116.635 146.930 116.925 146.975 ;
        RECT 117.770 146.930 118.090 146.990 ;
        RECT 116.635 146.790 118.090 146.930 ;
        RECT 63.505 146.450 64.270 146.590 ;
        RECT 63.505 146.405 63.795 146.450 ;
        RECT 63.950 146.390 64.270 146.450 ;
        RECT 71.325 146.405 71.615 146.635 ;
        RECT 73.610 146.590 73.930 146.650 ;
        RECT 78.210 146.590 78.530 146.650 ;
        RECT 73.610 146.450 78.530 146.590 ;
        RECT 73.610 146.390 73.930 146.450 ;
        RECT 78.210 146.390 78.530 146.450 ;
        RECT 79.590 146.390 79.910 146.650 ;
        RECT 82.350 146.590 82.670 146.650 ;
        RECT 85.355 146.590 85.645 146.635 ;
        RECT 86.030 146.590 86.350 146.650 ;
        RECT 82.350 146.450 86.350 146.590 ;
        RECT 82.350 146.390 82.670 146.450 ;
        RECT 85.355 146.405 85.645 146.450 ;
        RECT 86.030 146.390 86.350 146.450 ;
        RECT 97.070 146.590 97.390 146.650 ;
        RECT 98.005 146.590 98.295 146.635 ;
        RECT 107.280 146.590 107.420 146.790 ;
        RECT 116.635 146.745 116.925 146.790 ;
        RECT 117.770 146.730 118.090 146.790 ;
        RECT 118.640 146.930 118.930 146.975 ;
        RECT 120.070 146.930 120.390 146.990 ;
        RECT 122.820 146.975 123.035 147.130 ;
        RECT 123.750 147.070 124.070 147.330 ;
        RECT 125.605 147.270 125.895 147.315 ;
        RECT 126.050 147.270 126.370 147.330 ;
        RECT 125.605 147.130 126.370 147.270 ;
        RECT 125.605 147.085 125.895 147.130 ;
        RECT 126.050 147.070 126.370 147.130 ;
        RECT 121.900 146.930 122.190 146.975 ;
        RECT 118.640 146.790 122.190 146.930 ;
        RECT 118.640 146.745 118.930 146.790 ;
        RECT 120.070 146.730 120.390 146.790 ;
        RECT 121.900 146.745 122.190 146.790 ;
        RECT 122.820 146.930 123.110 146.975 ;
        RECT 124.680 146.930 124.970 146.975 ;
        RECT 122.820 146.790 124.970 146.930 ;
        RECT 122.820 146.745 123.110 146.790 ;
        RECT 124.680 146.745 124.970 146.790 ;
        RECT 97.070 146.450 107.420 146.590 ;
        RECT 108.110 146.590 108.430 146.650 ;
        RECT 109.490 146.590 109.810 146.650 ;
        RECT 108.110 146.450 109.810 146.590 ;
        RECT 97.070 146.390 97.390 146.450 ;
        RECT 98.005 146.405 98.295 146.450 ;
        RECT 108.110 146.390 108.430 146.450 ;
        RECT 109.490 146.390 109.810 146.450 ;
        RECT 113.645 146.590 113.935 146.635 ;
        RECT 114.090 146.590 114.410 146.650 ;
        RECT 117.310 146.590 117.630 146.650 ;
        RECT 113.645 146.450 117.630 146.590 ;
        RECT 113.645 146.405 113.935 146.450 ;
        RECT 114.090 146.390 114.410 146.450 ;
        RECT 117.310 146.390 117.630 146.450 ;
        RECT 14.660 145.770 127.820 146.250 ;
        RECT 20.250 145.370 20.570 145.630 ;
        RECT 23.010 145.615 23.330 145.630 ;
        RECT 22.795 145.385 23.330 145.615 ;
        RECT 51.070 145.570 51.390 145.630 ;
        RECT 23.010 145.370 23.330 145.385 ;
        RECT 41.040 145.430 51.390 145.570 ;
        RECT 21.645 145.230 21.935 145.275 ;
        RECT 24.800 145.230 25.090 145.275 ;
        RECT 28.060 145.230 28.350 145.275 ;
        RECT 21.645 145.090 28.350 145.230 ;
        RECT 21.645 145.045 21.935 145.090 ;
        RECT 24.800 145.045 25.090 145.090 ;
        RECT 28.060 145.045 28.350 145.090 ;
        RECT 28.980 145.230 29.270 145.275 ;
        RECT 30.840 145.230 31.130 145.275 ;
        RECT 28.980 145.090 31.130 145.230 ;
        RECT 28.980 145.045 29.270 145.090 ;
        RECT 30.840 145.045 31.130 145.090 ;
        RECT 19.805 144.890 20.095 144.935 ;
        RECT 21.185 144.890 21.475 144.935 ;
        RECT 19.805 144.750 21.475 144.890 ;
        RECT 19.805 144.705 20.095 144.750 ;
        RECT 21.185 144.705 21.475 144.750 ;
        RECT 26.660 144.890 26.950 144.935 ;
        RECT 28.980 144.890 29.195 145.045 ;
        RECT 26.660 144.750 29.195 144.890 ;
        RECT 30.370 144.890 30.690 144.950 ;
        RECT 41.040 144.935 41.180 145.430 ;
        RECT 51.070 145.370 51.390 145.430 ;
        RECT 51.990 145.370 52.310 145.630 ;
        RECT 53.830 145.370 54.150 145.630 ;
        RECT 80.970 145.570 81.290 145.630 ;
        RECT 80.600 145.430 81.290 145.570 ;
        RECT 41.425 145.230 41.715 145.275 ;
        RECT 44.580 145.230 44.870 145.275 ;
        RECT 47.840 145.230 48.130 145.275 ;
        RECT 41.425 145.090 48.130 145.230 ;
        RECT 41.425 145.045 41.715 145.090 ;
        RECT 44.580 145.045 44.870 145.090 ;
        RECT 47.840 145.045 48.130 145.090 ;
        RECT 48.760 145.230 49.050 145.275 ;
        RECT 50.620 145.230 50.910 145.275 ;
        RECT 48.760 145.090 50.910 145.230 ;
        RECT 51.160 145.230 51.300 145.370 ;
        RECT 55.210 145.230 55.530 145.290 ;
        RECT 59.350 145.230 59.670 145.290 ;
        RECT 65.345 145.230 65.635 145.275 ;
        RECT 51.160 145.090 58.660 145.230 ;
        RECT 48.760 145.045 49.050 145.090 ;
        RECT 50.620 145.045 50.910 145.090 ;
        RECT 40.965 144.890 41.255 144.935 ;
        RECT 30.370 144.750 41.255 144.890 ;
        RECT 26.660 144.705 26.950 144.750 ;
        RECT 21.260 143.870 21.400 144.705 ;
        RECT 30.370 144.690 30.690 144.750 ;
        RECT 40.965 144.705 41.255 144.750 ;
        RECT 46.440 144.890 46.730 144.935 ;
        RECT 48.760 144.890 48.975 145.045 ;
        RECT 55.210 145.030 55.530 145.090 ;
        RECT 46.440 144.750 48.975 144.890 ;
        RECT 46.440 144.705 46.730 144.750 ;
        RECT 49.690 144.690 50.010 144.950 ;
        RECT 58.520 144.935 58.660 145.090 ;
        RECT 59.350 145.090 65.635 145.230 ;
        RECT 59.350 145.030 59.670 145.090 ;
        RECT 65.345 145.045 65.635 145.090 ;
        RECT 79.590 145.030 79.910 145.290 ;
        RECT 54.305 144.890 54.595 144.935 ;
        RECT 50.240 144.750 54.595 144.890 ;
        RECT 28.990 144.550 29.310 144.610 ;
        RECT 29.925 144.550 30.215 144.595 ;
        RECT 28.990 144.410 30.215 144.550 ;
        RECT 28.990 144.350 29.310 144.410 ;
        RECT 29.925 144.365 30.215 144.410 ;
        RECT 31.765 144.550 32.055 144.595 ;
        RECT 36.350 144.550 36.670 144.610 ;
        RECT 31.765 144.410 36.670 144.550 ;
        RECT 31.765 144.365 32.055 144.410 ;
        RECT 36.350 144.350 36.670 144.410 ;
        RECT 42.575 144.550 42.865 144.595 ;
        RECT 50.240 144.550 50.380 144.750 ;
        RECT 54.305 144.705 54.595 144.750 ;
        RECT 58.445 144.705 58.735 144.935 ;
        RECT 65.790 144.690 66.110 144.950 ;
        RECT 80.600 144.935 80.740 145.430 ;
        RECT 80.970 145.370 81.290 145.430 ;
        RECT 86.030 145.370 86.350 145.630 ;
        RECT 91.090 145.370 91.410 145.630 ;
        RECT 97.070 145.370 97.390 145.630 ;
        RECT 117.310 145.370 117.630 145.630 ;
        RECT 120.070 145.370 120.390 145.630 ;
        RECT 122.385 145.570 122.675 145.615 ;
        RECT 123.750 145.570 124.070 145.630 ;
        RECT 122.385 145.430 124.070 145.570 ;
        RECT 122.385 145.385 122.675 145.430 ;
        RECT 123.750 145.370 124.070 145.430 ;
        RECT 107.205 145.230 107.495 145.275 ;
        RECT 109.965 145.230 110.255 145.275 ;
        RECT 107.205 145.090 110.255 145.230 ;
        RECT 107.205 145.045 107.495 145.090 ;
        RECT 109.965 145.045 110.255 145.090 ;
        RECT 112.340 145.090 117.080 145.230 ;
        RECT 80.525 144.705 80.815 144.935 ;
        RECT 80.985 144.890 81.275 144.935 ;
        RECT 81.430 144.890 81.750 144.950 ;
        RECT 80.985 144.750 81.750 144.890 ;
        RECT 80.985 144.705 81.275 144.750 ;
        RECT 81.430 144.690 81.750 144.750 ;
        RECT 84.650 144.890 84.970 144.950 ;
        RECT 86.505 144.890 86.795 144.935 ;
        RECT 90.185 144.890 90.475 144.935 ;
        RECT 84.650 144.750 86.795 144.890 ;
        RECT 84.650 144.690 84.970 144.750 ;
        RECT 86.505 144.705 86.795 144.750 ;
        RECT 88.420 144.750 90.475 144.890 ;
        RECT 50.610 144.550 50.930 144.610 ;
        RECT 42.575 144.410 50.930 144.550 ;
        RECT 42.575 144.365 42.865 144.410 ;
        RECT 50.610 144.350 50.930 144.410 ;
        RECT 51.545 144.365 51.835 144.595 ;
        RECT 54.750 144.550 55.070 144.610 ;
        RECT 55.225 144.550 55.515 144.595 ;
        RECT 64.870 144.550 65.190 144.610 ;
        RECT 69.470 144.550 69.790 144.610 ;
        RECT 54.750 144.410 69.790 144.550 ;
        RECT 26.660 144.210 26.950 144.255 ;
        RECT 29.440 144.210 29.730 144.255 ;
        RECT 31.300 144.210 31.590 144.255 ;
        RECT 26.660 144.070 31.590 144.210 ;
        RECT 26.660 144.025 26.950 144.070 ;
        RECT 29.440 144.025 29.730 144.070 ;
        RECT 31.300 144.025 31.590 144.070 ;
        RECT 46.440 144.210 46.730 144.255 ;
        RECT 49.220 144.210 49.510 144.255 ;
        RECT 51.080 144.210 51.370 144.255 ;
        RECT 46.440 144.070 51.370 144.210 ;
        RECT 51.620 144.210 51.760 144.365 ;
        RECT 54.750 144.350 55.070 144.410 ;
        RECT 55.225 144.365 55.515 144.410 ;
        RECT 64.870 144.350 65.190 144.410 ;
        RECT 69.470 144.350 69.790 144.410 ;
        RECT 85.110 144.350 85.430 144.610 ;
        RECT 63.950 144.210 64.270 144.270 ;
        RECT 51.620 144.070 64.270 144.210 ;
        RECT 46.440 144.025 46.730 144.070 ;
        RECT 49.220 144.025 49.510 144.070 ;
        RECT 51.080 144.025 51.370 144.070 ;
        RECT 63.950 144.010 64.270 144.070 ;
        RECT 69.010 144.210 69.330 144.270 ;
        RECT 70.850 144.210 71.170 144.270 ;
        RECT 69.010 144.070 71.170 144.210 ;
        RECT 69.010 144.010 69.330 144.070 ;
        RECT 70.850 144.010 71.170 144.070 ;
        RECT 75.450 144.210 75.770 144.270 ;
        RECT 88.420 144.255 88.560 144.750 ;
        RECT 90.185 144.705 90.475 144.750 ;
        RECT 94.325 144.890 94.615 144.935 ;
        RECT 96.610 144.890 96.930 144.950 ;
        RECT 94.325 144.750 96.930 144.890 ;
        RECT 94.325 144.705 94.615 144.750 ;
        RECT 96.610 144.690 96.930 144.750 ;
        RECT 108.585 144.890 108.875 144.935 ;
        RECT 109.030 144.890 109.350 144.950 ;
        RECT 108.585 144.750 109.350 144.890 ;
        RECT 108.585 144.705 108.875 144.750 ;
        RECT 109.030 144.690 109.350 144.750 ;
        RECT 109.490 144.890 109.810 144.950 ;
        RECT 111.345 144.890 111.635 144.935 ;
        RECT 109.490 144.750 111.635 144.890 ;
        RECT 109.490 144.690 109.810 144.750 ;
        RECT 111.345 144.705 111.635 144.750 ;
        RECT 108.125 144.550 108.415 144.595 ;
        RECT 110.410 144.550 110.730 144.610 ;
        RECT 108.125 144.410 110.730 144.550 ;
        RECT 108.125 144.365 108.415 144.410 ;
        RECT 110.410 144.350 110.730 144.410 ;
        RECT 81.905 144.210 82.195 144.255 ;
        RECT 75.450 144.070 82.195 144.210 ;
        RECT 75.450 144.010 75.770 144.070 ;
        RECT 81.905 144.025 82.195 144.070 ;
        RECT 88.345 144.025 88.635 144.255 ;
        RECT 109.030 144.210 109.350 144.270 ;
        RECT 109.505 144.210 109.795 144.255 ;
        RECT 111.420 144.210 111.560 144.705 ;
        RECT 111.790 144.690 112.110 144.950 ;
        RECT 112.340 144.935 112.480 145.090 ;
        RECT 112.265 144.705 112.555 144.935 ;
        RECT 112.710 144.890 113.030 144.950 ;
        RECT 113.185 144.890 113.475 144.935 ;
        RECT 112.710 144.750 113.475 144.890 ;
        RECT 112.710 144.690 113.030 144.750 ;
        RECT 113.185 144.705 113.475 144.750 ;
        RECT 113.630 144.550 113.950 144.610 ;
        RECT 116.940 144.595 117.080 145.090 ;
        RECT 119.610 144.690 119.930 144.950 ;
        RECT 121.465 144.705 121.755 144.935 ;
        RECT 115.945 144.550 116.235 144.595 ;
        RECT 113.630 144.410 116.235 144.550 ;
        RECT 113.630 144.350 113.950 144.410 ;
        RECT 115.945 144.365 116.235 144.410 ;
        RECT 116.865 144.550 117.155 144.595 ;
        RECT 117.770 144.550 118.090 144.610 ;
        RECT 121.540 144.550 121.680 144.705 ;
        RECT 116.865 144.410 118.090 144.550 ;
        RECT 116.865 144.365 117.155 144.410 ;
        RECT 117.770 144.350 118.090 144.410 ;
        RECT 119.240 144.410 121.680 144.550 ;
        RECT 119.240 144.255 119.380 144.410 ;
        RECT 109.030 144.070 109.795 144.210 ;
        RECT 109.030 144.010 109.350 144.070 ;
        RECT 109.505 144.025 109.795 144.070 ;
        RECT 110.500 144.070 111.560 144.210 ;
        RECT 110.500 143.930 110.640 144.070 ;
        RECT 119.165 144.025 119.455 144.255 ;
        RECT 29.910 143.870 30.230 143.930 ;
        RECT 21.260 143.730 30.230 143.870 ;
        RECT 29.910 143.670 30.230 143.730 ;
        RECT 58.890 143.670 59.210 143.930 ;
        RECT 67.645 143.870 67.935 143.915 ;
        RECT 69.930 143.870 70.250 143.930 ;
        RECT 67.645 143.730 70.250 143.870 ;
        RECT 67.645 143.685 67.935 143.730 ;
        RECT 69.930 143.670 70.250 143.730 ;
        RECT 80.970 143.670 81.290 143.930 ;
        RECT 108.585 143.870 108.875 143.915 ;
        RECT 109.950 143.870 110.270 143.930 ;
        RECT 108.585 143.730 110.270 143.870 ;
        RECT 108.585 143.685 108.875 143.730 ;
        RECT 109.950 143.670 110.270 143.730 ;
        RECT 110.410 143.670 110.730 143.930 ;
        RECT 14.660 143.050 127.820 143.530 ;
        RECT 35.890 142.650 36.210 142.910 ;
        RECT 48.325 142.665 48.615 142.895 ;
        RECT 45.090 142.510 45.410 142.570 ;
        RECT 48.400 142.510 48.540 142.665 ;
        RECT 59.350 142.650 59.670 142.910 ;
        RECT 109.030 142.850 109.350 142.910 ;
        RECT 111.790 142.850 112.110 142.910 ;
        RECT 109.030 142.710 112.110 142.850 ;
        RECT 109.030 142.650 109.350 142.710 ;
        RECT 111.790 142.650 112.110 142.710 ;
        RECT 45.090 142.370 48.540 142.510 ;
        RECT 62.685 142.510 62.975 142.555 ;
        RECT 65.805 142.510 66.095 142.555 ;
        RECT 67.695 142.510 67.985 142.555 ;
        RECT 69.010 142.510 69.330 142.570 ;
        RECT 62.685 142.370 67.985 142.510 ;
        RECT 45.090 142.310 45.410 142.370 ;
        RECT 62.685 142.325 62.975 142.370 ;
        RECT 65.805 142.325 66.095 142.370 ;
        RECT 67.695 142.325 67.985 142.370 ;
        RECT 68.180 142.370 69.330 142.510 ;
        RECT 34.510 142.170 34.830 142.230 ;
        RECT 35.905 142.170 36.195 142.215 ;
        RECT 34.510 142.030 36.195 142.170 ;
        RECT 34.510 141.970 34.830 142.030 ;
        RECT 35.905 141.985 36.195 142.030 ;
        RECT 46.470 142.170 46.790 142.230 ;
        RECT 48.785 142.170 49.075 142.215 ;
        RECT 46.470 142.030 49.075 142.170 ;
        RECT 46.470 141.970 46.790 142.030 ;
        RECT 48.785 141.985 49.075 142.030 ;
        RECT 53.370 142.170 53.690 142.230 ;
        RECT 56.605 142.170 56.895 142.215 ;
        RECT 59.825 142.170 60.115 142.215 ;
        RECT 68.180 142.170 68.320 142.370 ;
        RECT 69.010 142.310 69.330 142.370 ;
        RECT 53.370 142.030 54.520 142.170 ;
        RECT 53.370 141.970 53.690 142.030 ;
        RECT 34.970 141.830 35.290 141.890 ;
        RECT 35.445 141.830 35.735 141.875 ;
        RECT 34.970 141.690 35.735 141.830 ;
        RECT 34.970 141.630 35.290 141.690 ;
        RECT 35.445 141.645 35.735 141.690 ;
        RECT 46.010 141.830 46.330 141.890 ;
        RECT 48.325 141.830 48.615 141.875 ;
        RECT 46.010 141.690 48.615 141.830 ;
        RECT 46.010 141.630 46.330 141.690 ;
        RECT 48.325 141.645 48.615 141.690 ;
        RECT 53.830 141.630 54.150 141.890 ;
        RECT 54.380 141.875 54.520 142.030 ;
        RECT 54.840 142.030 60.115 142.170 ;
        RECT 54.840 141.875 54.980 142.030 ;
        RECT 56.605 141.985 56.895 142.030 ;
        RECT 59.825 141.985 60.115 142.030 ;
        RECT 60.360 142.030 68.320 142.170 ;
        RECT 54.305 141.645 54.595 141.875 ;
        RECT 54.765 141.645 55.055 141.875 ;
        RECT 55.685 141.830 55.975 141.875 ;
        RECT 56.130 141.830 56.450 141.890 ;
        RECT 60.360 141.830 60.500 142.030 ;
        RECT 68.550 141.970 68.870 142.230 ;
        RECT 113.170 142.170 113.490 142.230 ;
        RECT 116.405 142.170 116.695 142.215 ;
        RECT 113.170 142.030 116.695 142.170 ;
        RECT 113.170 141.970 113.490 142.030 ;
        RECT 116.405 141.985 116.695 142.030 ;
        RECT 55.685 141.690 56.450 141.830 ;
        RECT 55.685 141.645 55.975 141.690 ;
        RECT 56.130 141.630 56.450 141.690 ;
        RECT 58.060 141.690 60.500 141.830 ;
        RECT 36.825 141.490 37.115 141.535 ;
        RECT 39.570 141.490 39.890 141.550 ;
        RECT 36.825 141.350 39.890 141.490 ;
        RECT 36.825 141.305 37.115 141.350 ;
        RECT 39.570 141.290 39.890 141.350 ;
        RECT 49.705 141.490 49.995 141.535 ;
        RECT 52.465 141.490 52.755 141.535 ;
        RECT 49.705 141.350 52.755 141.490 ;
        RECT 49.705 141.305 49.995 141.350 ;
        RECT 52.465 141.305 52.755 141.350 ;
        RECT 29.450 141.150 29.770 141.210 ;
        RECT 34.525 141.150 34.815 141.195 ;
        RECT 29.450 141.010 34.815 141.150 ;
        RECT 29.450 140.950 29.770 141.010 ;
        RECT 34.525 140.965 34.815 141.010 ;
        RECT 47.405 141.150 47.695 141.195 ;
        RECT 58.060 141.150 58.200 141.690 ;
        RECT 58.890 141.490 59.210 141.550 ;
        RECT 61.605 141.535 61.895 141.850 ;
        RECT 62.685 141.830 62.975 141.875 ;
        RECT 66.265 141.830 66.555 141.875 ;
        RECT 68.100 141.830 68.390 141.875 ;
        RECT 62.685 141.690 68.390 141.830 ;
        RECT 62.685 141.645 62.975 141.690 ;
        RECT 66.265 141.645 66.555 141.690 ;
        RECT 68.100 141.645 68.390 141.690 ;
        RECT 69.930 141.630 70.250 141.890 ;
        RECT 70.850 141.830 71.170 141.890 ;
        RECT 72.705 141.830 72.995 141.875 ;
        RECT 70.850 141.690 72.995 141.830 ;
        RECT 70.850 141.630 71.170 141.690 ;
        RECT 72.705 141.645 72.995 141.690 ;
        RECT 117.770 141.630 118.090 141.890 ;
        RECT 119.610 141.830 119.930 141.890 ;
        RECT 120.085 141.830 120.375 141.875 ;
        RECT 119.610 141.690 120.375 141.830 ;
        RECT 119.610 141.630 119.930 141.690 ;
        RECT 120.085 141.645 120.375 141.690 ;
        RECT 61.305 141.490 61.895 141.535 ;
        RECT 64.545 141.490 65.195 141.535 ;
        RECT 58.890 141.350 65.195 141.490 ;
        RECT 58.890 141.290 59.210 141.350 ;
        RECT 61.305 141.305 61.595 141.350 ;
        RECT 64.545 141.305 65.195 141.350 ;
        RECT 67.185 141.490 67.475 141.535 ;
        RECT 67.185 141.350 69.240 141.490 ;
        RECT 67.185 141.305 67.475 141.350 ;
        RECT 47.405 141.010 58.200 141.150 ;
        RECT 63.950 141.150 64.270 141.210 ;
        RECT 68.550 141.150 68.870 141.210 ;
        RECT 69.100 141.195 69.240 141.350 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 63.950 141.010 68.870 141.150 ;
        RECT 47.405 140.965 47.695 141.010 ;
        RECT 63.950 140.950 64.270 141.010 ;
        RECT 68.550 140.950 68.870 141.010 ;
        RECT 69.025 140.965 69.315 141.195 ;
        RECT 72.230 140.950 72.550 141.210 ;
        RECT 117.310 140.950 117.630 141.210 ;
        RECT 119.610 140.950 119.930 141.210 ;
        RECT 120.530 140.950 120.850 141.210 ;
        RECT 14.660 140.330 127.820 140.810 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 35.890 139.930 36.210 140.190 ;
        RECT 38.665 139.945 38.955 140.175 ;
        RECT 39.570 140.130 39.890 140.190 ;
        RECT 59.365 140.130 59.655 140.175 ;
        RECT 61.190 140.130 61.510 140.190 ;
        RECT 63.965 140.130 64.255 140.175 ;
        RECT 39.570 139.990 59.655 140.130 ;
        RECT 18.360 139.790 18.650 139.835 ;
        RECT 19.330 139.790 19.650 139.850 ;
        RECT 21.620 139.790 21.910 139.835 ;
        RECT 18.360 139.650 21.910 139.790 ;
        RECT 18.360 139.605 18.650 139.650 ;
        RECT 19.330 139.590 19.650 139.650 ;
        RECT 21.620 139.605 21.910 139.650 ;
        RECT 22.540 139.790 22.830 139.835 ;
        RECT 24.400 139.790 24.690 139.835 ;
        RECT 38.740 139.790 38.880 139.945 ;
        RECT 39.570 139.930 39.890 139.990 ;
        RECT 59.365 139.945 59.655 139.990 ;
        RECT 59.900 139.990 64.255 140.130 ;
        RECT 22.540 139.650 24.690 139.790 ;
        RECT 22.540 139.605 22.830 139.650 ;
        RECT 24.400 139.605 24.690 139.650 ;
        RECT 36.670 139.650 38.880 139.790 ;
        RECT 40.965 139.790 41.255 139.835 ;
        RECT 41.410 139.790 41.730 139.850 ;
        RECT 59.900 139.790 60.040 139.990 ;
        RECT 61.190 139.930 61.510 139.990 ;
        RECT 63.965 139.945 64.255 139.990 ;
        RECT 65.790 140.130 66.110 140.190 ;
        RECT 67.875 140.130 68.165 140.175 ;
        RECT 65.790 139.990 68.165 140.130 ;
        RECT 65.790 139.930 66.110 139.990 ;
        RECT 67.875 139.945 68.165 139.990 ;
        RECT 81.430 139.930 81.750 140.190 ;
        RECT 84.650 140.130 84.970 140.190 ;
        RECT 86.045 140.130 86.335 140.175 ;
        RECT 84.650 139.990 86.335 140.130 ;
        RECT 84.650 139.930 84.970 139.990 ;
        RECT 86.045 139.945 86.335 139.990 ;
        RECT 88.345 139.945 88.635 140.175 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 65.880 139.790 66.020 139.930 ;
        RECT 40.965 139.650 41.730 139.790 ;
        RECT 20.220 139.450 20.510 139.495 ;
        RECT 22.540 139.450 22.755 139.605 ;
        RECT 20.220 139.310 22.755 139.450 ;
        RECT 34.970 139.450 35.290 139.510 ;
        RECT 35.890 139.450 36.210 139.510 ;
        RECT 36.670 139.450 36.810 139.650 ;
        RECT 40.965 139.605 41.255 139.650 ;
        RECT 41.410 139.590 41.730 139.650 ;
        RECT 55.300 139.650 60.040 139.790 ;
        RECT 61.740 139.650 66.020 139.790 ;
        RECT 69.880 139.790 70.170 139.835 ;
        RECT 72.230 139.790 72.550 139.850 ;
        RECT 73.140 139.790 73.430 139.835 ;
        RECT 69.880 139.650 73.430 139.790 ;
        RECT 34.970 139.310 35.485 139.450 ;
        RECT 35.890 139.310 36.810 139.450 ;
        RECT 39.585 139.450 39.875 139.495 ;
        RECT 55.300 139.450 55.440 139.650 ;
        RECT 39.585 139.310 55.440 139.450 ;
        RECT 20.220 139.265 20.510 139.310 ;
        RECT 34.970 139.250 35.290 139.310 ;
        RECT 35.890 139.250 36.210 139.310 ;
        RECT 39.585 139.265 39.875 139.310 ;
        RECT 55.685 139.265 55.975 139.495 ;
        RECT 23.470 138.910 23.790 139.170 ;
        RECT 25.325 139.110 25.615 139.155 ;
        RECT 29.910 139.110 30.230 139.170 ;
        RECT 25.325 138.970 30.230 139.110 ;
        RECT 25.325 138.925 25.615 138.970 ;
        RECT 29.910 138.910 30.230 138.970 ;
        RECT 30.370 139.110 30.690 139.170 ;
        RECT 34.065 139.110 34.355 139.155 ;
        RECT 30.370 138.970 34.355 139.110 ;
        RECT 30.370 138.910 30.690 138.970 ;
        RECT 34.065 138.925 34.355 138.970 ;
        RECT 40.030 138.910 40.350 139.170 ;
        RECT 55.210 139.110 55.530 139.170 ;
        RECT 55.760 139.110 55.900 139.265 ;
        RECT 56.130 139.250 56.450 139.510 ;
        RECT 60.730 139.250 61.050 139.510 ;
        RECT 61.740 139.495 61.880 139.650 ;
        RECT 69.880 139.605 70.170 139.650 ;
        RECT 72.230 139.590 72.550 139.650 ;
        RECT 73.140 139.605 73.430 139.650 ;
        RECT 74.060 139.790 74.350 139.835 ;
        RECT 75.920 139.790 76.210 139.835 ;
        RECT 74.060 139.650 76.210 139.790 ;
        RECT 74.060 139.605 74.350 139.650 ;
        RECT 75.920 139.605 76.210 139.650 ;
        RECT 80.050 139.790 80.370 139.850 ;
        RECT 81.520 139.790 81.660 139.930 ;
        RECT 84.740 139.790 84.880 139.930 ;
        RECT 80.050 139.650 81.660 139.790 ;
        RECT 81.980 139.650 84.880 139.790 ;
        RECT 61.205 139.265 61.495 139.495 ;
        RECT 61.665 139.265 61.955 139.495 ;
        RECT 62.585 139.265 62.875 139.495 ;
        RECT 55.210 138.970 55.900 139.110 ;
        RECT 55.210 138.910 55.530 138.970 ;
        RECT 20.220 138.770 20.510 138.815 ;
        RECT 23.000 138.770 23.290 138.815 ;
        RECT 24.860 138.770 25.150 138.815 ;
        RECT 20.220 138.630 25.150 138.770 ;
        RECT 20.220 138.585 20.510 138.630 ;
        RECT 23.000 138.585 23.290 138.630 ;
        RECT 24.860 138.585 25.150 138.630 ;
        RECT 16.355 138.430 16.645 138.475 ;
        RECT 22.550 138.430 22.870 138.490 ;
        RECT 16.355 138.290 22.870 138.430 ;
        RECT 16.355 138.245 16.645 138.290 ;
        RECT 22.550 138.230 22.870 138.290 ;
        RECT 34.510 138.430 34.830 138.490 ;
        RECT 39.585 138.430 39.875 138.475 ;
        RECT 34.510 138.290 39.875 138.430 ;
        RECT 34.510 138.230 34.830 138.290 ;
        RECT 39.585 138.245 39.875 138.290 ;
        RECT 47.850 138.430 48.170 138.490 ;
        RECT 50.150 138.430 50.470 138.490 ;
        RECT 53.830 138.430 54.150 138.490 ;
        RECT 47.850 138.290 54.150 138.430 ;
        RECT 61.280 138.430 61.420 139.265 ;
        RECT 62.660 138.770 62.800 139.265 ;
        RECT 65.330 139.250 65.650 139.510 ;
        RECT 65.805 139.265 66.095 139.495 ;
        RECT 65.880 139.110 66.020 139.265 ;
        RECT 66.250 139.250 66.570 139.510 ;
        RECT 67.185 139.450 67.475 139.495 ;
        RECT 68.090 139.450 68.410 139.510 ;
        RECT 67.185 139.310 68.410 139.450 ;
        RECT 67.185 139.265 67.475 139.310 ;
        RECT 68.090 139.250 68.410 139.310 ;
        RECT 71.740 139.450 72.030 139.495 ;
        RECT 74.060 139.450 74.275 139.605 ;
        RECT 80.050 139.590 80.370 139.650 ;
        RECT 81.060 139.495 81.200 139.650 ;
        RECT 81.980 139.495 82.120 139.650 ;
        RECT 71.740 139.310 74.275 139.450 ;
        RECT 71.740 139.265 72.030 139.310 ;
        RECT 80.985 139.265 81.275 139.495 ;
        RECT 81.445 139.265 81.735 139.495 ;
        RECT 81.905 139.265 82.195 139.495 ;
        RECT 82.825 139.265 83.115 139.495 ;
        RECT 70.390 139.110 70.710 139.170 ;
        RECT 65.880 138.970 70.710 139.110 ;
        RECT 64.410 138.770 64.730 138.830 ;
        RECT 67.630 138.770 67.950 138.830 ;
        RECT 62.660 138.630 67.950 138.770 ;
        RECT 64.410 138.570 64.730 138.630 ;
        RECT 67.630 138.570 67.950 138.630 ;
        RECT 66.710 138.430 67.030 138.490 ;
        RECT 68.180 138.430 68.320 138.970 ;
        RECT 70.390 138.910 70.710 138.970 ;
        RECT 74.990 138.910 75.310 139.170 ;
        RECT 76.845 138.925 77.135 139.155 ;
        RECT 81.520 139.110 81.660 139.265 ;
        RECT 82.350 139.110 82.670 139.170 ;
        RECT 81.520 138.970 82.670 139.110 ;
        RECT 82.900 139.110 83.040 139.265 ;
        RECT 86.490 139.250 86.810 139.510 ;
        RECT 88.420 139.450 88.560 139.945 ;
        RECT 100.240 139.790 100.530 139.835 ;
        RECT 102.590 139.790 102.910 139.850 ;
        RECT 103.500 139.790 103.790 139.835 ;
        RECT 100.240 139.650 103.790 139.790 ;
        RECT 100.240 139.605 100.530 139.650 ;
        RECT 102.590 139.590 102.910 139.650 ;
        RECT 103.500 139.605 103.790 139.650 ;
        RECT 104.420 139.790 104.710 139.835 ;
        RECT 106.280 139.790 106.570 139.835 ;
        RECT 104.420 139.650 106.570 139.790 ;
        RECT 104.420 139.605 104.710 139.650 ;
        RECT 106.280 139.605 106.570 139.650 ;
        RECT 110.410 139.790 110.730 139.850 ;
        RECT 112.250 139.790 112.570 139.850 ;
        RECT 117.310 139.835 117.630 139.850 ;
        RECT 113.185 139.790 113.475 139.835 ;
        RECT 117.095 139.790 117.630 139.835 ;
        RECT 110.410 139.650 112.020 139.790 ;
        RECT 89.265 139.450 89.555 139.495 ;
        RECT 88.420 139.310 89.555 139.450 ;
        RECT 89.265 139.265 89.555 139.310 ;
        RECT 102.100 139.450 102.390 139.495 ;
        RECT 104.420 139.450 104.635 139.605 ;
        RECT 110.410 139.590 110.730 139.650 ;
        RECT 102.100 139.310 104.635 139.450 ;
        RECT 109.490 139.450 109.810 139.510 ;
        RECT 109.965 139.450 110.255 139.495 ;
        RECT 109.490 139.310 110.255 139.450 ;
        RECT 110.885 139.440 111.175 139.510 ;
        RECT 111.880 139.495 112.020 139.650 ;
        RECT 112.250 139.650 113.475 139.790 ;
        RECT 112.250 139.590 112.570 139.650 ;
        RECT 113.185 139.605 113.475 139.650 ;
        RECT 114.180 139.650 117.630 139.790 ;
        RECT 102.100 139.265 102.390 139.310 ;
        RECT 109.490 139.250 109.810 139.310 ;
        RECT 109.965 139.265 110.255 139.310 ;
        RECT 110.500 139.300 111.175 139.440 ;
        RECT 83.270 139.110 83.590 139.170 ;
        RECT 82.900 138.970 83.590 139.110 ;
        RECT 71.740 138.770 72.030 138.815 ;
        RECT 74.520 138.770 74.810 138.815 ;
        RECT 76.380 138.770 76.670 138.815 ;
        RECT 71.740 138.630 76.670 138.770 ;
        RECT 76.920 138.770 77.060 138.925 ;
        RECT 82.350 138.910 82.670 138.970 ;
        RECT 83.270 138.910 83.590 138.970 ;
        RECT 85.110 138.910 85.430 139.170 ;
        RECT 98.235 139.110 98.525 139.155 ;
        RECT 98.910 139.110 99.230 139.170 ;
        RECT 98.235 138.970 99.230 139.110 ;
        RECT 98.235 138.925 98.525 138.970 ;
        RECT 98.910 138.910 99.230 138.970 ;
        RECT 105.350 138.910 105.670 139.170 ;
        RECT 107.205 138.925 107.495 139.155 ;
        RECT 94.310 138.770 94.630 138.830 ;
        RECT 76.920 138.630 94.630 138.770 ;
        RECT 71.740 138.585 72.030 138.630 ;
        RECT 74.520 138.585 74.810 138.630 ;
        RECT 76.380 138.585 76.670 138.630 ;
        RECT 94.310 138.570 94.630 138.630 ;
        RECT 102.100 138.770 102.390 138.815 ;
        RECT 104.880 138.770 105.170 138.815 ;
        RECT 106.740 138.770 107.030 138.815 ;
        RECT 102.100 138.630 107.030 138.770 ;
        RECT 102.100 138.585 102.390 138.630 ;
        RECT 104.880 138.585 105.170 138.630 ;
        RECT 106.740 138.585 107.030 138.630 ;
        RECT 61.280 138.290 68.320 138.430 ;
        RECT 47.850 138.230 48.170 138.290 ;
        RECT 50.150 138.230 50.470 138.290 ;
        RECT 53.830 138.230 54.150 138.290 ;
        RECT 66.710 138.230 67.030 138.290 ;
        RECT 79.590 138.230 79.910 138.490 ;
        RECT 90.185 138.430 90.475 138.475 ;
        RECT 91.090 138.430 91.410 138.490 ;
        RECT 90.185 138.290 91.410 138.430 ;
        RECT 90.185 138.245 90.475 138.290 ;
        RECT 91.090 138.230 91.410 138.290 ;
        RECT 98.450 138.430 98.770 138.490 ;
        RECT 107.280 138.430 107.420 138.925 ;
        RECT 110.500 138.770 110.640 139.300 ;
        RECT 110.885 139.280 111.175 139.300 ;
        RECT 111.345 139.265 111.635 139.495 ;
        RECT 111.805 139.265 112.095 139.495 ;
        RECT 111.420 139.110 111.560 139.265 ;
        RECT 112.710 139.250 113.030 139.510 ;
        RECT 112.800 139.110 112.940 139.250 ;
        RECT 111.420 138.970 112.940 139.110 ;
        RECT 112.710 138.770 113.030 138.830 ;
        RECT 114.180 138.770 114.320 139.650 ;
        RECT 117.095 139.605 117.630 139.650 ;
        RECT 119.100 139.790 119.390 139.835 ;
        RECT 120.530 139.790 120.850 139.850 ;
        RECT 122.360 139.790 122.650 139.835 ;
        RECT 119.100 139.650 122.650 139.790 ;
        RECT 119.100 139.605 119.390 139.650 ;
        RECT 117.310 139.590 117.630 139.605 ;
        RECT 120.530 139.590 120.850 139.650 ;
        RECT 122.360 139.605 122.650 139.650 ;
        RECT 123.280 139.790 123.570 139.835 ;
        RECT 125.140 139.790 125.430 139.835 ;
        RECT 123.280 139.650 125.430 139.790 ;
        RECT 123.280 139.605 123.570 139.650 ;
        RECT 125.140 139.605 125.430 139.650 ;
        RECT 115.485 139.265 115.775 139.495 ;
        RECT 110.500 138.630 114.320 138.770 ;
        RECT 115.560 138.770 115.700 139.265 ;
        RECT 115.930 139.250 116.250 139.510 ;
        RECT 120.960 139.450 121.250 139.495 ;
        RECT 123.280 139.450 123.495 139.605 ;
        RECT 120.960 139.310 123.495 139.450 ;
        RECT 120.960 139.265 121.250 139.310 ;
        RECT 124.210 139.250 124.530 139.510 ;
        RECT 129.090 139.190 134.150 139.405 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 126.050 138.910 126.370 139.170 ;
        RECT 120.070 138.770 120.390 138.830 ;
        RECT 115.560 138.630 120.390 138.770 ;
        RECT 112.710 138.570 113.030 138.630 ;
        RECT 120.070 138.570 120.390 138.630 ;
        RECT 120.960 138.770 121.250 138.815 ;
        RECT 123.740 138.770 124.030 138.815 ;
        RECT 125.600 138.770 125.890 138.815 ;
        RECT 120.960 138.630 125.890 138.770 ;
        RECT 120.960 138.585 121.250 138.630 ;
        RECT 123.740 138.585 124.030 138.630 ;
        RECT 125.600 138.585 125.890 138.630 ;
        RECT 121.450 138.430 121.770 138.490 ;
        RECT 124.670 138.430 124.990 138.490 ;
        RECT 126.140 138.430 126.280 138.910 ;
        RECT 98.450 138.290 126.280 138.430 ;
        RECT 129.090 138.530 144.510 139.190 ;
        RECT 98.450 138.230 98.770 138.290 ;
        RECT 121.450 138.230 121.770 138.290 ;
        RECT 124.670 138.230 124.990 138.290 ;
        RECT 129.090 138.225 134.150 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 14.660 137.610 127.820 138.090 ;
        RECT 34.510 137.210 34.830 137.470 ;
        RECT 35.905 137.225 36.195 137.455 ;
        RECT 38.190 137.410 38.510 137.470 ;
        RECT 38.665 137.410 38.955 137.455 ;
        RECT 38.190 137.270 38.955 137.410 ;
        RECT 34.050 137.070 34.370 137.130 ;
        RECT 35.980 137.070 36.120 137.225 ;
        RECT 38.190 137.210 38.510 137.270 ;
        RECT 38.665 137.225 38.955 137.270 ;
        RECT 44.630 137.210 44.950 137.470 ;
        RECT 48.310 137.410 48.630 137.470 ;
        RECT 51.070 137.410 51.390 137.470 ;
        RECT 53.370 137.410 53.690 137.470 ;
        RECT 48.310 137.270 53.690 137.410 ;
        RECT 48.310 137.210 48.630 137.270 ;
        RECT 51.070 137.210 51.390 137.270 ;
        RECT 53.370 137.210 53.690 137.270 ;
        RECT 60.730 137.410 61.050 137.470 ;
        RECT 60.730 137.270 62.800 137.410 ;
        RECT 60.730 137.210 61.050 137.270 ;
        RECT 61.205 137.070 61.495 137.115 ;
        RECT 34.050 136.930 36.120 137.070 ;
        RECT 40.120 136.930 61.495 137.070 ;
        RECT 34.050 136.870 34.370 136.930 ;
        RECT 21.630 136.730 21.950 136.790 ;
        RECT 23.025 136.730 23.315 136.775 ;
        RECT 21.630 136.590 23.315 136.730 ;
        RECT 21.630 136.530 21.950 136.590 ;
        RECT 23.025 136.545 23.315 136.590 ;
        RECT 31.290 136.530 31.610 136.790 ;
        RECT 35.430 136.730 35.750 136.790 ;
        RECT 36.365 136.730 36.655 136.775 ;
        RECT 35.430 136.590 36.655 136.730 ;
        RECT 35.430 136.530 35.750 136.590 ;
        RECT 36.365 136.545 36.655 136.590 ;
        RECT 39.110 136.530 39.430 136.790 ;
        RECT 22.105 136.390 22.395 136.435 ;
        RECT 22.550 136.390 22.870 136.450 ;
        RECT 22.105 136.250 22.870 136.390 ;
        RECT 22.105 136.205 22.395 136.250 ;
        RECT 22.550 136.190 22.870 136.250 ;
        RECT 32.685 136.205 32.975 136.435 ;
        RECT 33.590 136.390 33.910 136.450 ;
        RECT 34.970 136.390 35.290 136.450 ;
        RECT 33.590 136.250 35.290 136.390 ;
        RECT 30.370 136.050 30.690 136.110 ;
        RECT 22.640 135.910 30.690 136.050 ;
        RECT 18.870 135.710 19.190 135.770 ;
        RECT 20.265 135.710 20.555 135.755 ;
        RECT 18.870 135.570 20.555 135.710 ;
        RECT 18.870 135.510 19.190 135.570 ;
        RECT 20.265 135.525 20.555 135.570 ;
        RECT 22.090 135.710 22.410 135.770 ;
        RECT 22.640 135.755 22.780 135.910 ;
        RECT 30.370 135.850 30.690 135.910 ;
        RECT 32.760 135.770 32.900 136.205 ;
        RECT 33.590 136.190 33.910 136.250 ;
        RECT 34.970 136.190 35.290 136.250 ;
        RECT 35.905 136.390 36.195 136.435 ;
        RECT 36.810 136.390 37.130 136.450 ;
        RECT 35.905 136.250 37.130 136.390 ;
        RECT 35.905 136.205 36.195 136.250 ;
        RECT 36.810 136.190 37.130 136.250 ;
        RECT 38.650 136.190 38.970 136.450 ;
        RECT 40.120 136.435 40.260 136.930 ;
        RECT 61.205 136.885 61.495 136.930 ;
        RECT 62.660 137.070 62.800 137.270 ;
        RECT 65.330 137.210 65.650 137.470 ;
        RECT 71.325 137.410 71.615 137.455 ;
        RECT 74.990 137.410 75.310 137.470 ;
        RECT 71.325 137.270 75.310 137.410 ;
        RECT 71.325 137.225 71.615 137.270 ;
        RECT 74.990 137.210 75.310 137.270 ;
        RECT 79.605 137.410 79.895 137.455 ;
        RECT 80.050 137.410 80.370 137.470 ;
        RECT 83.975 137.410 84.265 137.455 ;
        RECT 84.650 137.410 84.970 137.470 ;
        RECT 79.605 137.270 80.370 137.410 ;
        RECT 79.605 137.225 79.895 137.270 ;
        RECT 80.050 137.210 80.370 137.270 ;
        RECT 81.520 137.270 83.040 137.410 ;
        RECT 65.420 137.070 65.560 137.210 ;
        RECT 74.530 137.070 74.850 137.130 ;
        RECT 62.660 136.930 74.850 137.070 ;
        RECT 45.550 136.530 45.870 136.790 ;
        RECT 50.610 136.730 50.930 136.790 ;
        RECT 48.860 136.590 50.930 136.730 ;
        RECT 40.045 136.205 40.335 136.435 ;
        RECT 42.330 136.390 42.650 136.450 ;
        RECT 44.645 136.390 44.935 136.435 ;
        RECT 42.330 136.250 44.935 136.390 ;
        RECT 42.330 136.190 42.650 136.250 ;
        RECT 44.645 136.205 44.935 136.250 ;
        RECT 45.640 136.250 47.620 136.390 ;
        RECT 37.285 136.050 37.575 136.095 ;
        RECT 45.640 136.050 45.780 136.250 ;
        RECT 37.285 135.910 45.780 136.050 ;
        RECT 46.025 136.050 46.315 136.095 ;
        RECT 46.485 136.050 46.775 136.095 ;
        RECT 46.025 135.910 46.775 136.050 ;
        RECT 47.480 136.050 47.620 136.250 ;
        RECT 47.850 136.190 48.170 136.450 ;
        RECT 48.310 136.190 48.630 136.450 ;
        RECT 48.860 136.435 49.000 136.590 ;
        RECT 50.610 136.530 50.930 136.590 ;
        RECT 54.305 136.730 54.595 136.775 ;
        RECT 54.750 136.730 55.070 136.790 ;
        RECT 54.305 136.590 55.070 136.730 ;
        RECT 54.305 136.545 54.595 136.590 ;
        RECT 54.750 136.530 55.070 136.590 ;
        RECT 48.785 136.205 49.075 136.435 ;
        RECT 49.705 136.205 49.995 136.435 ;
        RECT 50.700 136.390 50.840 136.530 ;
        RECT 62.660 136.435 62.800 136.930 ;
        RECT 74.530 136.870 74.850 136.930 ;
        RECT 77.305 137.070 77.595 137.115 ;
        RECT 81.520 137.070 81.660 137.270 ;
        RECT 82.350 137.070 82.670 137.130 ;
        RECT 77.305 136.930 81.660 137.070 ;
        RECT 81.980 136.930 82.670 137.070 ;
        RECT 82.900 137.070 83.040 137.270 ;
        RECT 83.975 137.270 84.970 137.410 ;
        RECT 83.975 137.225 84.265 137.270 ;
        RECT 84.650 137.210 84.970 137.270 ;
        RECT 85.110 137.410 85.430 137.470 ;
        RECT 105.350 137.410 105.670 137.470 ;
        RECT 107.205 137.410 107.495 137.455 ;
        RECT 85.110 137.270 95.920 137.410 ;
        RECT 85.110 137.210 85.430 137.270 ;
        RECT 86.950 137.070 87.270 137.130 ;
        RECT 82.900 136.930 87.270 137.070 ;
        RECT 77.305 136.885 77.595 136.930 ;
        RECT 65.345 136.730 65.635 136.775 ;
        RECT 65.790 136.730 66.110 136.790 ;
        RECT 74.070 136.730 74.390 136.790 ;
        RECT 63.120 136.590 64.180 136.730 ;
        RECT 63.120 136.435 63.260 136.590 ;
        RECT 55.225 136.390 55.515 136.435 ;
        RECT 57.985 136.390 58.275 136.435 ;
        RECT 50.700 136.250 55.515 136.390 ;
        RECT 55.225 136.205 55.515 136.250 ;
        RECT 57.140 136.250 58.275 136.390 ;
        RECT 49.230 136.050 49.550 136.110 ;
        RECT 47.480 135.910 49.550 136.050 ;
        RECT 49.780 136.050 49.920 136.205 ;
        RECT 50.610 136.050 50.930 136.110 ;
        RECT 52.450 136.050 52.770 136.110 ;
        RECT 55.670 136.050 55.990 136.110 ;
        RECT 49.780 135.910 55.990 136.050 ;
        RECT 37.285 135.865 37.575 135.910 ;
        RECT 46.025 135.865 46.315 135.910 ;
        RECT 46.485 135.865 46.775 135.910 ;
        RECT 49.230 135.850 49.550 135.910 ;
        RECT 50.610 135.850 50.930 135.910 ;
        RECT 52.450 135.850 52.770 135.910 ;
        RECT 55.670 135.850 55.990 135.910 ;
        RECT 22.565 135.710 22.855 135.755 ;
        RECT 22.090 135.570 22.855 135.710 ;
        RECT 22.090 135.510 22.410 135.570 ;
        RECT 22.565 135.525 22.855 135.570 ;
        RECT 28.530 135.510 28.850 135.770 ;
        RECT 30.830 135.710 31.150 135.770 ;
        RECT 32.670 135.710 32.990 135.770 ;
        RECT 30.830 135.570 32.990 135.710 ;
        RECT 30.830 135.510 31.150 135.570 ;
        RECT 32.670 135.510 32.990 135.570 ;
        RECT 34.510 135.710 34.830 135.770 ;
        RECT 34.985 135.710 35.275 135.755 ;
        RECT 34.510 135.570 35.275 135.710 ;
        RECT 34.510 135.510 34.830 135.570 ;
        RECT 34.985 135.525 35.275 135.570 ;
        RECT 37.745 135.710 38.035 135.755 ;
        RECT 38.650 135.710 38.970 135.770 ;
        RECT 37.745 135.570 38.970 135.710 ;
        RECT 37.745 135.525 38.035 135.570 ;
        RECT 38.650 135.510 38.970 135.570 ;
        RECT 43.725 135.710 44.015 135.755 ;
        RECT 51.990 135.710 52.310 135.770 ;
        RECT 43.725 135.570 52.310 135.710 ;
        RECT 43.725 135.525 44.015 135.570 ;
        RECT 51.990 135.510 52.310 135.570 ;
        RECT 54.765 135.710 55.055 135.755 ;
        RECT 56.590 135.710 56.910 135.770 ;
        RECT 57.140 135.755 57.280 136.250 ;
        RECT 57.985 136.205 58.275 136.250 ;
        RECT 62.585 136.205 62.875 136.435 ;
        RECT 63.045 136.205 63.335 136.435 ;
        RECT 63.505 136.205 63.795 136.435 ;
        RECT 60.730 136.050 61.050 136.110 ;
        RECT 63.580 136.050 63.720 136.205 ;
        RECT 60.730 135.910 63.720 136.050 ;
        RECT 64.040 136.050 64.180 136.590 ;
        RECT 65.345 136.590 66.110 136.730 ;
        RECT 65.345 136.545 65.635 136.590 ;
        RECT 65.790 136.530 66.110 136.590 ;
        RECT 70.020 136.590 74.390 136.730 ;
        RECT 64.410 136.190 64.730 136.450 ;
        RECT 68.105 136.390 68.395 136.435 ;
        RECT 68.565 136.390 68.855 136.435 ;
        RECT 68.105 136.250 68.855 136.390 ;
        RECT 68.105 136.205 68.395 136.250 ;
        RECT 68.565 136.205 68.855 136.250 ;
        RECT 69.470 136.190 69.790 136.450 ;
        RECT 70.020 136.435 70.160 136.590 ;
        RECT 74.070 136.530 74.390 136.590 ;
        RECT 69.945 136.205 70.235 136.435 ;
        RECT 70.405 136.205 70.695 136.435 ;
        RECT 76.370 136.390 76.690 136.450 ;
        RECT 78.225 136.390 78.515 136.435 ;
        RECT 76.370 136.250 78.515 136.390 ;
        RECT 65.330 136.050 65.650 136.110 ;
        RECT 66.710 136.050 67.030 136.110 ;
        RECT 70.480 136.050 70.620 136.205 ;
        RECT 76.370 136.190 76.690 136.250 ;
        RECT 78.225 136.205 78.515 136.250 ;
        RECT 78.685 136.205 78.975 136.435 ;
        RECT 64.040 135.910 67.030 136.050 ;
        RECT 60.730 135.850 61.050 135.910 ;
        RECT 65.330 135.850 65.650 135.910 ;
        RECT 66.710 135.850 67.030 135.910 ;
        RECT 70.020 135.910 70.620 136.050 ;
        RECT 78.760 136.050 78.900 136.205 ;
        RECT 79.590 136.190 79.910 136.450 ;
        RECT 81.430 136.190 81.750 136.450 ;
        RECT 81.980 136.435 82.120 136.930 ;
        RECT 82.350 136.870 82.670 136.930 ;
        RECT 86.950 136.870 87.270 136.930 ;
        RECT 87.840 137.070 88.130 137.115 ;
        RECT 90.620 137.070 90.910 137.115 ;
        RECT 92.480 137.070 92.770 137.115 ;
        RECT 87.840 136.930 92.770 137.070 ;
        RECT 95.780 137.070 95.920 137.270 ;
        RECT 105.350 137.270 107.495 137.410 ;
        RECT 105.350 137.210 105.670 137.270 ;
        RECT 107.205 137.225 107.495 137.270 ;
        RECT 119.610 137.410 119.930 137.470 ;
        RECT 119.610 137.270 123.520 137.410 ;
        RECT 119.610 137.210 119.930 137.270 ;
        RECT 113.170 137.070 113.490 137.130 ;
        RECT 95.780 136.930 96.380 137.070 ;
        RECT 87.840 136.885 88.130 136.930 ;
        RECT 90.620 136.885 90.910 136.930 ;
        RECT 92.480 136.885 92.770 136.930 ;
        RECT 86.490 136.730 86.810 136.790 ;
        RECT 82.440 136.590 86.810 136.730 ;
        RECT 82.440 136.435 82.580 136.590 ;
        RECT 86.490 136.530 86.810 136.590 ;
        RECT 91.090 136.530 91.410 136.790 ;
        RECT 91.550 136.730 91.870 136.790 ;
        RECT 96.240 136.775 96.380 136.930 ;
        RECT 103.600 136.930 113.490 137.070 ;
        RECT 103.600 136.775 103.740 136.930 ;
        RECT 110.040 136.775 110.180 136.930 ;
        RECT 113.170 136.870 113.490 136.930 ;
        RECT 117.740 137.070 118.030 137.115 ;
        RECT 120.520 137.070 120.810 137.115 ;
        RECT 122.380 137.070 122.670 137.115 ;
        RECT 117.740 136.930 122.670 137.070 ;
        RECT 117.740 136.885 118.030 136.930 ;
        RECT 120.520 136.885 120.810 136.930 ;
        RECT 122.380 136.885 122.670 136.930 ;
        RECT 95.705 136.730 95.995 136.775 ;
        RECT 91.550 136.590 95.995 136.730 ;
        RECT 91.550 136.530 91.870 136.590 ;
        RECT 95.705 136.545 95.995 136.590 ;
        RECT 96.165 136.730 96.455 136.775 ;
        RECT 103.525 136.730 103.815 136.775 ;
        RECT 96.165 136.590 103.815 136.730 ;
        RECT 96.165 136.545 96.455 136.590 ;
        RECT 103.525 136.545 103.815 136.590 ;
        RECT 104.980 136.590 109.260 136.730 ;
        RECT 81.905 136.205 82.195 136.435 ;
        RECT 82.365 136.205 82.655 136.435 ;
        RECT 83.270 136.190 83.590 136.450 ;
        RECT 87.840 136.390 88.130 136.435 ;
        RECT 87.840 136.250 90.375 136.390 ;
        RECT 87.840 136.205 88.130 136.250 ;
        RECT 84.190 136.050 84.510 136.110 ;
        RECT 78.760 135.910 84.510 136.050 ;
        RECT 54.765 135.570 56.910 135.710 ;
        RECT 54.765 135.525 55.055 135.570 ;
        RECT 56.590 135.510 56.910 135.570 ;
        RECT 57.065 135.525 57.355 135.755 ;
        RECT 58.905 135.710 59.195 135.755 ;
        RECT 59.810 135.710 60.130 135.770 ;
        RECT 58.905 135.570 60.130 135.710 ;
        RECT 58.905 135.525 59.195 135.570 ;
        RECT 59.810 135.510 60.130 135.570 ;
        RECT 61.190 135.710 61.510 135.770 ;
        RECT 70.020 135.710 70.160 135.910 ;
        RECT 84.190 135.850 84.510 135.910 ;
        RECT 85.980 136.050 86.270 136.095 ;
        RECT 88.330 136.050 88.650 136.110 ;
        RECT 90.160 136.095 90.375 136.250 ;
        RECT 92.945 136.205 93.235 136.435 ;
        RECT 93.390 136.390 93.710 136.450 ;
        RECT 97.990 136.390 98.310 136.450 ;
        RECT 93.390 136.250 98.310 136.390 ;
        RECT 89.240 136.050 89.530 136.095 ;
        RECT 85.980 135.910 89.530 136.050 ;
        RECT 85.980 135.865 86.270 135.910 ;
        RECT 88.330 135.850 88.650 135.910 ;
        RECT 89.240 135.865 89.530 135.910 ;
        RECT 90.160 136.050 90.450 136.095 ;
        RECT 92.020 136.050 92.310 136.095 ;
        RECT 90.160 135.910 92.310 136.050 ;
        RECT 93.020 136.050 93.160 136.205 ;
        RECT 93.390 136.190 93.710 136.250 ;
        RECT 97.990 136.190 98.310 136.250 ;
        RECT 98.910 136.190 99.230 136.450 ;
        RECT 99.370 136.190 99.690 136.450 ;
        RECT 99.845 136.390 100.135 136.435 ;
        RECT 100.290 136.390 100.610 136.450 ;
        RECT 104.980 136.435 105.120 136.590 ;
        RECT 104.445 136.390 104.735 136.435 ;
        RECT 99.845 136.250 100.610 136.390 ;
        RECT 99.845 136.205 100.135 136.250 ;
        RECT 100.290 136.190 100.610 136.250 ;
        RECT 100.840 136.250 104.735 136.390 ;
        RECT 94.310 136.050 94.630 136.110 ;
        RECT 98.450 136.050 98.770 136.110 ;
        RECT 93.020 135.910 98.770 136.050 ;
        RECT 90.160 135.865 90.450 135.910 ;
        RECT 92.020 135.865 92.310 135.910 ;
        RECT 94.310 135.850 94.630 135.910 ;
        RECT 98.450 135.850 98.770 135.910 ;
        RECT 99.000 136.050 99.140 136.190 ;
        RECT 100.840 136.050 100.980 136.250 ;
        RECT 104.445 136.205 104.735 136.250 ;
        RECT 104.905 136.205 105.195 136.435 ;
        RECT 108.125 136.390 108.415 136.435 ;
        RECT 106.820 136.250 108.415 136.390 ;
        RECT 99.000 135.910 100.980 136.050 ;
        RECT 61.190 135.570 70.160 135.710 ;
        RECT 79.130 135.710 79.450 135.770 ;
        RECT 80.065 135.710 80.355 135.755 ;
        RECT 79.130 135.570 80.355 135.710 ;
        RECT 61.190 135.510 61.510 135.570 ;
        RECT 79.130 135.510 79.450 135.570 ;
        RECT 80.065 135.525 80.355 135.570 ;
        RECT 85.110 135.710 85.430 135.770 ;
        RECT 92.930 135.710 93.250 135.770 ;
        RECT 85.110 135.570 93.250 135.710 ;
        RECT 85.110 135.510 85.430 135.570 ;
        RECT 92.930 135.510 93.250 135.570 ;
        RECT 93.405 135.710 93.695 135.755 ;
        RECT 93.850 135.710 94.170 135.770 ;
        RECT 93.405 135.570 94.170 135.710 ;
        RECT 93.405 135.525 93.695 135.570 ;
        RECT 93.850 135.510 94.170 135.570 ;
        RECT 95.245 135.710 95.535 135.755 ;
        RECT 99.000 135.710 99.140 135.910 ;
        RECT 95.245 135.570 99.140 135.710 ;
        RECT 95.245 135.525 95.535 135.570 ;
        RECT 101.210 135.510 101.530 135.770 ;
        RECT 106.820 135.755 106.960 136.250 ;
        RECT 108.125 136.205 108.415 136.250 ;
        RECT 109.120 136.110 109.260 136.590 ;
        RECT 109.965 136.545 110.255 136.775 ;
        RECT 121.450 136.730 121.770 136.790 ;
        RECT 122.845 136.730 123.135 136.775 ;
        RECT 121.450 136.590 123.135 136.730 ;
        RECT 121.450 136.530 121.770 136.590 ;
        RECT 122.845 136.545 123.135 136.590 ;
        RECT 111.345 136.390 111.635 136.435 ;
        RECT 112.710 136.390 113.030 136.450 ;
        RECT 111.345 136.250 113.030 136.390 ;
        RECT 111.345 136.205 111.635 136.250 ;
        RECT 112.710 136.190 113.030 136.250 ;
        RECT 117.740 136.390 118.030 136.435 ;
        RECT 117.740 136.250 120.275 136.390 ;
        RECT 117.740 136.205 118.030 136.250 ;
        RECT 109.030 136.050 109.350 136.110 ;
        RECT 115.930 136.095 116.250 136.110 ;
        RECT 120.060 136.095 120.275 136.250 ;
        RECT 120.990 136.190 121.310 136.450 ;
        RECT 123.380 136.435 123.520 137.270 ;
        RECT 124.210 137.210 124.530 137.470 ;
        RECT 123.305 136.205 123.595 136.435 ;
        RECT 110.885 136.050 111.175 136.095 ;
        RECT 113.875 136.050 114.165 136.095 ;
        RECT 109.030 135.910 114.165 136.050 ;
        RECT 109.030 135.850 109.350 135.910 ;
        RECT 110.885 135.865 111.175 135.910 ;
        RECT 113.875 135.865 114.165 135.910 ;
        RECT 115.880 136.050 116.250 136.095 ;
        RECT 119.140 136.050 119.430 136.095 ;
        RECT 115.880 135.910 119.430 136.050 ;
        RECT 115.880 135.865 116.250 135.910 ;
        RECT 119.140 135.865 119.430 135.910 ;
        RECT 120.060 136.050 120.350 136.095 ;
        RECT 121.920 136.050 122.210 136.095 ;
        RECT 120.060 135.910 122.210 136.050 ;
        RECT 120.060 135.865 120.350 135.910 ;
        RECT 121.920 135.865 122.210 135.910 ;
        RECT 115.930 135.850 116.250 135.865 ;
        RECT 106.745 135.525 107.035 135.755 ;
        RECT 113.170 135.510 113.490 135.770 ;
        RECT 14.660 134.890 127.820 135.370 ;
        RECT 19.330 134.490 19.650 134.750 ;
        RECT 20.955 134.690 21.245 134.735 ;
        RECT 22.090 134.690 22.410 134.750 ;
        RECT 20.955 134.550 22.410 134.690 ;
        RECT 20.955 134.505 21.245 134.550 ;
        RECT 22.090 134.490 22.410 134.550 ;
        RECT 32.685 134.690 32.975 134.735 ;
        RECT 34.050 134.690 34.370 134.750 ;
        RECT 32.685 134.550 34.370 134.690 ;
        RECT 32.685 134.505 32.975 134.550 ;
        RECT 34.050 134.490 34.370 134.550 ;
        RECT 50.610 134.490 50.930 134.750 ;
        RECT 52.695 134.690 52.985 134.735 ;
        RECT 56.590 134.690 56.910 134.750 ;
        RECT 51.160 134.550 56.910 134.690 ;
        RECT 17.045 134.350 17.335 134.395 ;
        RECT 19.420 134.350 19.560 134.490 ;
        RECT 17.045 134.210 19.560 134.350 ;
        RECT 19.805 134.350 20.095 134.395 ;
        RECT 22.960 134.350 23.250 134.395 ;
        RECT 26.220 134.350 26.510 134.395 ;
        RECT 19.805 134.210 26.510 134.350 ;
        RECT 17.045 134.165 17.335 134.210 ;
        RECT 19.805 134.165 20.095 134.210 ;
        RECT 22.960 134.165 23.250 134.210 ;
        RECT 26.220 134.165 26.510 134.210 ;
        RECT 27.140 134.350 27.430 134.395 ;
        RECT 29.000 134.350 29.290 134.395 ;
        RECT 36.350 134.350 36.670 134.410 ;
        RECT 27.140 134.210 29.290 134.350 ;
        RECT 27.140 134.165 27.430 134.210 ;
        RECT 29.000 134.165 29.290 134.210 ;
        RECT 30.000 134.210 36.670 134.350 ;
        RECT 17.505 133.825 17.795 134.055 ;
        RECT 17.965 134.010 18.255 134.055 ;
        RECT 18.870 134.010 19.190 134.070 ;
        RECT 17.965 133.870 19.190 134.010 ;
        RECT 17.965 133.825 18.255 133.870 ;
        RECT 17.580 133.670 17.720 133.825 ;
        RECT 18.870 133.810 19.190 133.870 ;
        RECT 19.345 134.010 19.635 134.055 ;
        RECT 24.820 134.010 25.110 134.055 ;
        RECT 27.140 134.010 27.355 134.165 ;
        RECT 30.000 134.070 30.140 134.210 ;
        RECT 36.350 134.150 36.670 134.210 ;
        RECT 42.345 134.350 42.635 134.395 ;
        RECT 48.785 134.350 49.075 134.395 ;
        RECT 50.700 134.350 50.840 134.490 ;
        RECT 42.345 134.210 49.075 134.350 ;
        RECT 42.345 134.165 42.635 134.210 ;
        RECT 48.785 134.165 49.075 134.210 ;
        RECT 49.780 134.210 50.840 134.350 ;
        RECT 19.345 133.870 20.020 134.010 ;
        RECT 19.345 133.825 19.635 133.870 ;
        RECT 19.880 133.730 20.020 133.870 ;
        RECT 24.820 133.870 27.355 134.010 ;
        RECT 27.700 133.870 29.680 134.010 ;
        RECT 24.820 133.825 25.110 133.870 ;
        RECT 19.790 133.670 20.110 133.730 ;
        RECT 17.580 133.530 20.110 133.670 ;
        RECT 19.790 133.470 20.110 133.530 ;
        RECT 22.090 133.670 22.410 133.730 ;
        RECT 27.700 133.670 27.840 133.870 ;
        RECT 22.090 133.530 27.840 133.670 ;
        RECT 28.085 133.670 28.375 133.715 ;
        RECT 28.990 133.670 29.310 133.730 ;
        RECT 28.085 133.530 29.310 133.670 ;
        RECT 29.540 133.670 29.680 133.870 ;
        RECT 29.910 133.810 30.230 134.070 ;
        RECT 31.290 134.010 31.610 134.070 ;
        RECT 30.460 133.870 31.610 134.010 ;
        RECT 30.460 133.670 30.600 133.870 ;
        RECT 31.290 133.810 31.610 133.870 ;
        RECT 31.765 134.010 32.055 134.055 ;
        RECT 32.210 134.010 32.530 134.070 ;
        RECT 31.765 133.870 32.530 134.010 ;
        RECT 31.765 133.825 32.055 133.870 ;
        RECT 32.210 133.810 32.530 133.870 ;
        RECT 32.670 134.010 32.990 134.070 ;
        RECT 34.985 134.010 35.275 134.055 ;
        RECT 32.670 133.870 35.275 134.010 ;
        RECT 32.670 133.810 32.990 133.870 ;
        RECT 34.985 133.825 35.275 133.870 ;
        RECT 39.585 133.825 39.875 134.055 ;
        RECT 29.540 133.530 30.600 133.670 ;
        RECT 22.090 133.470 22.410 133.530 ;
        RECT 28.085 133.485 28.375 133.530 ;
        RECT 28.990 133.470 29.310 133.530 ;
        RECT 30.845 133.485 31.135 133.715 ;
        RECT 31.380 133.670 31.520 133.810 ;
        RECT 33.605 133.670 33.895 133.715 ;
        RECT 31.380 133.530 33.895 133.670 ;
        RECT 33.605 133.485 33.895 133.530 ;
        RECT 34.525 133.485 34.815 133.715 ;
        RECT 39.660 133.670 39.800 133.825 ;
        RECT 40.490 133.810 40.810 134.070 ;
        RECT 40.950 133.810 41.270 134.070 ;
        RECT 42.790 134.010 43.110 134.070 ;
        RECT 43.265 134.010 43.555 134.055 ;
        RECT 42.790 133.870 43.555 134.010 ;
        RECT 42.790 133.810 43.110 133.870 ;
        RECT 43.265 133.825 43.555 133.870 ;
        RECT 43.710 133.810 44.030 134.070 ;
        RECT 46.470 133.810 46.790 134.070 ;
        RECT 46.945 133.825 47.235 134.055 ;
        RECT 47.405 133.825 47.695 134.055 ;
        RECT 48.325 134.010 48.615 134.055 ;
        RECT 49.780 134.010 49.920 134.210 ;
        RECT 48.325 133.870 49.920 134.010 ;
        RECT 48.325 133.825 48.615 133.870 ;
        RECT 45.105 133.670 45.395 133.715 ;
        RECT 39.660 133.530 45.395 133.670 ;
        RECT 45.105 133.485 45.395 133.530 ;
        RECT 18.885 133.330 19.175 133.375 ;
        RECT 23.470 133.330 23.790 133.390 ;
        RECT 18.885 133.190 23.790 133.330 ;
        RECT 18.885 133.145 19.175 133.190 ;
        RECT 23.470 133.130 23.790 133.190 ;
        RECT 24.820 133.330 25.110 133.375 ;
        RECT 27.600 133.330 27.890 133.375 ;
        RECT 29.460 133.330 29.750 133.375 ;
        RECT 24.820 133.190 29.750 133.330 ;
        RECT 30.920 133.330 31.060 133.485 ;
        RECT 34.600 133.330 34.740 133.485 ;
        RECT 34.970 133.330 35.290 133.390 ;
        RECT 30.920 133.190 35.290 133.330 ;
        RECT 24.820 133.145 25.110 133.190 ;
        RECT 27.600 133.145 27.890 133.190 ;
        RECT 29.460 133.145 29.750 133.190 ;
        RECT 34.970 133.130 35.290 133.190 ;
        RECT 31.290 132.990 31.610 133.050 ;
        RECT 35.890 132.990 36.210 133.050 ;
        RECT 31.290 132.850 36.210 132.990 ;
        RECT 31.290 132.790 31.610 132.850 ;
        RECT 35.890 132.790 36.210 132.850 ;
        RECT 36.825 132.990 37.115 133.035 ;
        RECT 39.570 132.990 39.890 133.050 ;
        RECT 36.825 132.850 39.890 132.990 ;
        RECT 36.825 132.805 37.115 132.850 ;
        RECT 39.570 132.790 39.890 132.850 ;
        RECT 40.490 132.790 40.810 133.050 ;
        RECT 41.410 132.990 41.730 133.050 ;
        RECT 41.885 132.990 42.175 133.035 ;
        RECT 41.410 132.850 42.175 132.990 ;
        RECT 41.410 132.790 41.730 132.850 ;
        RECT 41.885 132.805 42.175 132.850 ;
        RECT 43.250 132.790 43.570 133.050 ;
        RECT 44.170 132.990 44.490 133.050 ;
        RECT 44.645 132.990 44.935 133.035 ;
        RECT 44.170 132.850 44.935 132.990 ;
        RECT 47.020 132.990 47.160 133.825 ;
        RECT 47.480 133.330 47.620 133.825 ;
        RECT 50.150 133.810 50.470 134.070 ;
        RECT 50.610 133.810 50.930 134.070 ;
        RECT 51.160 134.055 51.300 134.550 ;
        RECT 52.695 134.505 52.985 134.550 ;
        RECT 56.590 134.490 56.910 134.550 ;
        RECT 74.530 134.690 74.850 134.750 ;
        RECT 87.885 134.690 88.175 134.735 ;
        RECT 88.330 134.690 88.650 134.750 ;
        RECT 100.290 134.690 100.610 134.750 ;
        RECT 102.145 134.690 102.435 134.735 ;
        RECT 102.590 134.690 102.910 134.750 ;
        RECT 74.530 134.550 87.640 134.690 ;
        RECT 74.530 134.490 74.850 134.550 ;
        RECT 54.700 134.350 54.990 134.395 ;
        RECT 56.130 134.350 56.450 134.410 ;
        RECT 57.960 134.350 58.250 134.395 ;
        RECT 54.700 134.210 58.250 134.350 ;
        RECT 54.700 134.165 54.990 134.210 ;
        RECT 56.130 134.150 56.450 134.210 ;
        RECT 57.960 134.165 58.250 134.210 ;
        RECT 58.880 134.350 59.170 134.395 ;
        RECT 60.740 134.350 61.030 134.395 ;
        RECT 58.880 134.210 61.030 134.350 ;
        RECT 58.880 134.165 59.170 134.210 ;
        RECT 60.740 134.165 61.030 134.210 ;
        RECT 64.410 134.350 64.730 134.410 ;
        RECT 64.410 134.210 66.940 134.350 ;
        RECT 51.085 133.825 51.375 134.055 ;
        RECT 52.005 134.010 52.295 134.055 ;
        RECT 52.450 134.010 52.770 134.070 ;
        RECT 52.005 133.870 52.770 134.010 ;
        RECT 52.005 133.825 52.295 133.870 ;
        RECT 52.450 133.810 52.770 133.870 ;
        RECT 56.560 134.010 56.850 134.055 ;
        RECT 58.880 134.010 59.095 134.165 ;
        RECT 64.410 134.150 64.730 134.210 ;
        RECT 56.560 133.870 59.095 134.010 ;
        RECT 56.560 133.825 56.850 133.870 ;
        RECT 59.810 133.810 60.130 134.070 ;
        RECT 61.665 134.010 61.955 134.055 ;
        RECT 63.950 134.010 64.270 134.070 ;
        RECT 61.665 133.870 64.270 134.010 ;
        RECT 61.665 133.825 61.955 133.870 ;
        RECT 63.950 133.810 64.270 133.870 ;
        RECT 64.870 133.810 65.190 134.070 ;
        RECT 65.330 133.810 65.650 134.070 ;
        RECT 65.790 133.810 66.110 134.070 ;
        RECT 66.800 134.055 66.940 134.210 ;
        RECT 79.130 134.150 79.450 134.410 ;
        RECT 85.110 134.350 85.430 134.410 ;
        RECT 80.140 134.210 85.430 134.350 ;
        RECT 87.500 134.350 87.640 134.550 ;
        RECT 87.885 134.550 88.650 134.690 ;
        RECT 87.885 134.505 88.175 134.550 ;
        RECT 88.330 134.490 88.650 134.550 ;
        RECT 90.260 134.550 101.900 134.690 ;
        RECT 90.260 134.350 90.400 134.550 ;
        RECT 100.290 134.490 100.610 134.550 ;
        RECT 87.500 134.210 90.400 134.350 ;
        RECT 90.630 134.350 90.950 134.410 ;
        RECT 91.500 134.350 91.790 134.395 ;
        RECT 94.760 134.350 95.050 134.395 ;
        RECT 90.630 134.210 95.050 134.350 ;
        RECT 66.725 134.010 67.015 134.055 ;
        RECT 80.140 134.010 80.280 134.210 ;
        RECT 85.110 134.150 85.430 134.210 ;
        RECT 90.630 134.150 90.950 134.210 ;
        RECT 91.500 134.165 91.790 134.210 ;
        RECT 94.760 134.165 95.050 134.210 ;
        RECT 95.680 134.350 95.970 134.395 ;
        RECT 97.540 134.350 97.830 134.395 ;
        RECT 95.680 134.210 97.830 134.350 ;
        RECT 95.680 134.165 95.970 134.210 ;
        RECT 97.540 134.165 97.830 134.210 ;
        RECT 66.725 133.870 80.280 134.010 ;
        RECT 66.725 133.825 67.015 133.870 ;
        RECT 80.510 133.810 80.830 134.070 ;
        RECT 88.330 133.810 88.650 134.070 ;
        RECT 93.360 134.010 93.650 134.055 ;
        RECT 95.680 134.010 95.895 134.165 ;
        RECT 101.210 134.150 101.530 134.410 ;
        RECT 101.760 134.350 101.900 134.550 ;
        RECT 102.145 134.550 102.910 134.690 ;
        RECT 102.145 134.505 102.435 134.550 ;
        RECT 102.590 134.490 102.910 134.550 ;
        RECT 120.085 134.690 120.375 134.735 ;
        RECT 120.990 134.690 121.310 134.750 ;
        RECT 120.085 134.550 121.310 134.690 ;
        RECT 120.085 134.505 120.375 134.550 ;
        RECT 120.990 134.490 121.310 134.550 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 105.825 134.350 106.115 134.395 ;
        RECT 106.285 134.350 106.575 134.395 ;
        RECT 110.410 134.350 110.730 134.410 ;
        RECT 101.760 134.210 105.020 134.350 ;
        RECT 93.360 133.870 95.895 134.010 ;
        RECT 93.360 133.825 93.650 133.870 ;
        RECT 97.990 133.810 98.310 134.070 ;
        RECT 98.450 133.810 98.770 134.070 ;
        RECT 99.830 133.810 100.150 134.070 ;
        RECT 102.590 133.810 102.910 134.070 ;
        RECT 103.970 134.010 104.290 134.070 ;
        RECT 104.445 134.010 104.735 134.055 ;
        RECT 103.970 133.870 104.735 134.010 ;
        RECT 104.880 134.010 105.020 134.210 ;
        RECT 105.825 134.210 106.575 134.350 ;
        RECT 105.825 134.165 106.115 134.210 ;
        RECT 106.285 134.165 106.575 134.210 ;
        RECT 107.740 134.210 110.730 134.350 ;
        RECT 107.740 134.055 107.880 134.210 ;
        RECT 110.410 134.150 110.730 134.210 ;
        RECT 112.250 134.150 112.570 134.410 ;
        RECT 107.665 134.010 107.955 134.055 ;
        RECT 104.880 133.870 107.955 134.010 ;
        RECT 103.970 133.810 104.290 133.870 ;
        RECT 104.445 133.825 104.735 133.870 ;
        RECT 107.665 133.825 107.955 133.870 ;
        RECT 108.110 133.810 108.430 134.070 ;
        RECT 108.585 134.010 108.875 134.055 ;
        RECT 109.030 134.010 109.350 134.070 ;
        RECT 108.585 133.870 109.350 134.010 ;
        RECT 108.585 133.825 108.875 133.870 ;
        RECT 109.030 133.810 109.350 133.870 ;
        RECT 109.490 133.810 109.810 134.070 ;
        RECT 110.870 133.810 111.190 134.070 ;
        RECT 111.330 133.810 111.650 134.070 ;
        RECT 113.170 134.010 113.490 134.070 ;
        RECT 119.165 134.010 119.455 134.055 ;
        RECT 113.170 133.870 119.455 134.010 ;
        RECT 113.170 133.810 113.490 133.870 ;
        RECT 119.165 133.825 119.455 133.870 ;
        RECT 49.230 133.670 49.550 133.730 ;
        RECT 63.505 133.670 63.795 133.715 ;
        RECT 49.230 133.530 63.795 133.670 ;
        RECT 49.230 133.470 49.550 133.530 ;
        RECT 63.505 133.485 63.795 133.530 ;
        RECT 80.065 133.670 80.355 133.715 ;
        RECT 83.730 133.670 84.050 133.730 ;
        RECT 80.065 133.530 84.050 133.670 ;
        RECT 80.065 133.485 80.355 133.530 ;
        RECT 83.730 133.470 84.050 133.530 ;
        RECT 86.490 133.670 86.810 133.730 ;
        RECT 89.495 133.670 89.785 133.715 ;
        RECT 91.550 133.670 91.870 133.730 ;
        RECT 86.490 133.530 91.870 133.670 ;
        RECT 86.490 133.470 86.810 133.530 ;
        RECT 89.495 133.485 89.785 133.530 ;
        RECT 91.550 133.470 91.870 133.530 ;
        RECT 95.230 133.670 95.550 133.730 ;
        RECT 96.625 133.670 96.915 133.715 ;
        RECT 95.230 133.530 96.915 133.670 ;
        RECT 98.080 133.670 98.220 133.810 ;
        RECT 98.080 133.530 100.520 133.670 ;
        RECT 95.230 133.470 95.550 133.530 ;
        RECT 96.625 133.485 96.915 133.530 ;
        RECT 55.670 133.330 55.990 133.390 ;
        RECT 47.480 133.190 55.990 133.330 ;
        RECT 55.670 133.130 55.990 133.190 ;
        RECT 56.560 133.330 56.850 133.375 ;
        RECT 59.340 133.330 59.630 133.375 ;
        RECT 61.200 133.330 61.490 133.375 ;
        RECT 56.560 133.190 61.490 133.330 ;
        RECT 56.560 133.145 56.850 133.190 ;
        RECT 59.340 133.145 59.630 133.190 ;
        RECT 61.200 133.145 61.490 133.190 ;
        RECT 81.445 133.330 81.735 133.375 ;
        RECT 93.360 133.330 93.650 133.375 ;
        RECT 96.140 133.330 96.430 133.375 ;
        RECT 98.000 133.330 98.290 133.375 ;
        RECT 81.445 133.190 88.100 133.330 ;
        RECT 81.445 133.145 81.735 133.190 ;
        RECT 50.610 132.990 50.930 133.050 ;
        RECT 47.020 132.850 50.930 132.990 ;
        RECT 44.170 132.790 44.490 132.850 ;
        RECT 44.645 132.805 44.935 132.850 ;
        RECT 50.610 132.790 50.930 132.850 ;
        RECT 80.525 132.990 80.815 133.035 ;
        RECT 83.270 132.990 83.590 133.050 ;
        RECT 80.525 132.850 83.590 132.990 ;
        RECT 87.960 132.990 88.100 133.190 ;
        RECT 93.360 133.190 98.290 133.330 ;
        RECT 100.380 133.330 100.520 133.530 ;
        RECT 100.750 133.470 101.070 133.730 ;
        RECT 102.130 133.670 102.450 133.730 ;
        RECT 104.905 133.670 105.195 133.715 ;
        RECT 102.130 133.530 105.195 133.670 ;
        RECT 102.130 133.470 102.450 133.530 ;
        RECT 104.905 133.485 105.195 133.530 ;
        RECT 109.580 133.330 109.720 133.810 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 100.380 133.190 109.720 133.330 ;
        RECT 93.360 133.145 93.650 133.190 ;
        RECT 96.140 133.145 96.430 133.190 ;
        RECT 98.000 133.145 98.290 133.190 ;
        RECT 94.770 132.990 95.090 133.050 ;
        RECT 87.960 132.850 95.090 132.990 ;
        RECT 80.525 132.805 80.815 132.850 ;
        RECT 83.270 132.790 83.590 132.850 ;
        RECT 94.770 132.790 95.090 132.850 ;
        RECT 98.925 132.990 99.215 133.035 ;
        RECT 99.830 132.990 100.150 133.050 ;
        RECT 98.925 132.850 100.150 132.990 ;
        RECT 98.925 132.805 99.215 132.850 ;
        RECT 99.830 132.790 100.150 132.850 ;
        RECT 101.210 132.790 101.530 133.050 ;
        RECT 103.510 132.790 103.830 133.050 ;
        RECT 104.890 132.790 105.210 133.050 ;
        RECT 109.965 132.990 110.255 133.035 ;
        RECT 110.410 132.990 110.730 133.050 ;
        RECT 109.965 132.850 110.730 132.990 ;
        RECT 109.965 132.805 110.255 132.850 ;
        RECT 110.410 132.790 110.730 132.850 ;
        RECT 111.330 132.790 111.650 133.050 ;
        RECT 14.660 132.170 127.820 132.650 ;
        RECT 28.990 131.770 29.310 132.030 ;
        RECT 30.830 132.015 31.150 132.030 ;
        RECT 30.615 131.785 31.150 132.015 ;
        RECT 30.830 131.770 31.150 131.785 ;
        RECT 34.050 131.970 34.370 132.030 ;
        RECT 78.685 131.970 78.975 132.015 ;
        RECT 80.050 131.970 80.370 132.030 ;
        RECT 34.050 131.830 40.260 131.970 ;
        RECT 34.050 131.770 34.370 131.830 ;
        RECT 40.120 131.690 40.260 131.830 ;
        RECT 78.685 131.830 80.370 131.970 ;
        RECT 78.685 131.785 78.975 131.830 ;
        RECT 80.050 131.770 80.370 131.830 ;
        RECT 89.725 131.970 90.015 132.015 ;
        RECT 90.630 131.970 90.950 132.030 ;
        RECT 89.725 131.830 90.950 131.970 ;
        RECT 89.725 131.785 90.015 131.830 ;
        RECT 90.630 131.770 90.950 131.830 ;
        RECT 109.950 131.770 110.270 132.030 ;
        RECT 34.480 131.630 34.770 131.675 ;
        RECT 37.260 131.630 37.550 131.675 ;
        RECT 39.120 131.630 39.410 131.675 ;
        RECT 34.480 131.490 39.410 131.630 ;
        RECT 34.480 131.445 34.770 131.490 ;
        RECT 37.260 131.445 37.550 131.490 ;
        RECT 39.120 131.445 39.410 131.490 ;
        RECT 40.030 131.630 40.350 131.690 ;
        RECT 69.945 131.630 70.235 131.675 ;
        RECT 100.290 131.630 100.610 131.690 ;
        RECT 40.030 131.490 100.610 131.630 ;
        RECT 40.030 131.430 40.350 131.490 ;
        RECT 69.945 131.445 70.235 131.490 ;
        RECT 100.290 131.430 100.610 131.490 ;
        RECT 102.590 131.630 102.910 131.690 ;
        RECT 118.230 131.630 118.550 131.690 ;
        RECT 102.590 131.490 118.550 131.630 ;
        RECT 102.590 131.430 102.910 131.490 ;
        RECT 118.230 131.430 118.550 131.490 ;
        RECT 21.185 131.290 21.475 131.335 ;
        RECT 22.090 131.290 22.410 131.350 ;
        RECT 21.185 131.150 22.410 131.290 ;
        RECT 21.185 131.105 21.475 131.150 ;
        RECT 22.090 131.090 22.410 131.150 ;
        RECT 36.350 131.290 36.670 131.350 ;
        RECT 36.350 131.150 37.500 131.290 ;
        RECT 36.350 131.090 36.670 131.150 ;
        RECT 28.530 130.950 28.850 131.010 ;
        RECT 29.925 130.950 30.215 130.995 ;
        RECT 28.530 130.810 30.215 130.950 ;
        RECT 28.530 130.750 28.850 130.810 ;
        RECT 29.925 130.765 30.215 130.810 ;
        RECT 34.480 130.950 34.770 130.995 ;
        RECT 37.360 130.950 37.500 131.150 ;
        RECT 37.730 131.090 38.050 131.350 ;
        RECT 64.870 131.290 65.190 131.350 ;
        RECT 66.725 131.290 67.015 131.335 ;
        RECT 69.470 131.290 69.790 131.350 ;
        RECT 64.870 131.150 69.790 131.290 ;
        RECT 64.870 131.090 65.190 131.150 ;
        RECT 66.725 131.105 67.015 131.150 ;
        RECT 69.470 131.090 69.790 131.150 ;
        RECT 73.625 131.290 73.915 131.335 ;
        RECT 74.070 131.290 74.390 131.350 ;
        RECT 73.625 131.150 74.390 131.290 ;
        RECT 73.625 131.105 73.915 131.150 ;
        RECT 74.070 131.090 74.390 131.150 ;
        RECT 39.585 130.950 39.875 130.995 ;
        RECT 70.865 130.950 71.155 130.995 ;
        RECT 72.690 130.950 73.010 131.010 ;
        RECT 74.545 130.950 74.835 130.995 ;
        RECT 79.605 130.950 79.895 130.995 ;
        RECT 34.480 130.810 37.015 130.950 ;
        RECT 37.360 130.810 42.560 130.950 ;
        RECT 34.480 130.765 34.770 130.810 ;
        RECT 22.105 130.610 22.395 130.655 ;
        RECT 23.470 130.610 23.790 130.670 ;
        RECT 22.105 130.470 23.790 130.610 ;
        RECT 22.105 130.425 22.395 130.470 ;
        RECT 23.470 130.410 23.790 130.470 ;
        RECT 32.620 130.610 32.910 130.655 ;
        RECT 34.050 130.610 34.370 130.670 ;
        RECT 36.800 130.655 37.015 130.810 ;
        RECT 39.585 130.765 39.875 130.810 ;
        RECT 35.880 130.610 36.170 130.655 ;
        RECT 32.620 130.470 36.170 130.610 ;
        RECT 32.620 130.425 32.910 130.470 ;
        RECT 34.050 130.410 34.370 130.470 ;
        RECT 35.880 130.425 36.170 130.470 ;
        RECT 36.800 130.610 37.090 130.655 ;
        RECT 38.660 130.610 38.950 130.655 ;
        RECT 36.800 130.470 38.950 130.610 ;
        RECT 36.800 130.425 37.090 130.470 ;
        RECT 38.660 130.425 38.950 130.470 ;
        RECT 21.645 130.270 21.935 130.315 ;
        RECT 22.550 130.270 22.870 130.330 ;
        RECT 21.645 130.130 22.870 130.270 ;
        RECT 21.645 130.085 21.935 130.130 ;
        RECT 22.550 130.070 22.870 130.130 ;
        RECT 23.010 130.270 23.330 130.330 ;
        RECT 42.420 130.315 42.560 130.810 ;
        RECT 70.865 130.810 74.835 130.950 ;
        RECT 70.865 130.765 71.155 130.810 ;
        RECT 72.690 130.750 73.010 130.810 ;
        RECT 74.545 130.765 74.835 130.810 ;
        RECT 75.080 130.810 79.895 130.950 ;
        RECT 48.785 130.610 49.075 130.655 ;
        RECT 49.230 130.610 49.550 130.670 ;
        RECT 48.785 130.470 49.550 130.610 ;
        RECT 48.785 130.425 49.075 130.470 ;
        RECT 49.230 130.410 49.550 130.470 ;
        RECT 64.410 130.610 64.730 130.670 ;
        RECT 65.790 130.610 66.110 130.670 ;
        RECT 67.645 130.610 67.935 130.655 ;
        RECT 64.410 130.470 67.935 130.610 ;
        RECT 64.410 130.410 64.730 130.470 ;
        RECT 65.790 130.410 66.110 130.470 ;
        RECT 67.645 130.425 67.935 130.470 ;
        RECT 68.090 130.610 68.410 130.670 ;
        RECT 75.080 130.610 75.220 130.810 ;
        RECT 79.605 130.765 79.895 130.810 ;
        RECT 80.050 130.750 80.370 131.010 ;
        RECT 88.330 130.950 88.650 131.010 ;
        RECT 89.265 130.950 89.555 130.995 ;
        RECT 91.090 130.950 91.410 131.010 ;
        RECT 88.330 130.810 91.410 130.950 ;
        RECT 88.330 130.750 88.650 130.810 ;
        RECT 89.265 130.765 89.555 130.810 ;
        RECT 91.090 130.750 91.410 130.810 ;
        RECT 98.450 130.950 98.770 131.010 ;
        RECT 100.305 130.950 100.595 130.995 ;
        RECT 98.450 130.810 100.595 130.950 ;
        RECT 98.450 130.750 98.770 130.810 ;
        RECT 100.305 130.765 100.595 130.810 ;
        RECT 110.870 130.750 111.190 131.010 ;
        RECT 111.805 130.950 112.095 130.995 ;
        RECT 112.250 130.950 112.570 131.010 ;
        RECT 111.805 130.810 112.570 130.950 ;
        RECT 111.805 130.765 112.095 130.810 ;
        RECT 112.250 130.750 112.570 130.810 ;
        RECT 68.090 130.470 75.220 130.610 ;
        RECT 68.090 130.410 68.410 130.470 ;
        RECT 75.080 130.330 75.220 130.470 ;
        RECT 23.945 130.270 24.235 130.315 ;
        RECT 23.010 130.130 24.235 130.270 ;
        RECT 23.010 130.070 23.330 130.130 ;
        RECT 23.945 130.085 24.235 130.130 ;
        RECT 42.345 130.270 42.635 130.315 ;
        RECT 42.790 130.270 43.110 130.330 ;
        RECT 42.345 130.130 43.110 130.270 ;
        RECT 42.345 130.085 42.635 130.130 ;
        RECT 42.790 130.070 43.110 130.130 ;
        RECT 66.250 130.270 66.570 130.330 ;
        RECT 67.185 130.270 67.475 130.315 ;
        RECT 66.250 130.130 67.475 130.270 ;
        RECT 66.250 130.070 66.570 130.130 ;
        RECT 67.185 130.085 67.475 130.130 ;
        RECT 69.485 130.270 69.775 130.315 ;
        RECT 70.390 130.270 70.710 130.330 ;
        RECT 69.485 130.130 70.710 130.270 ;
        RECT 69.485 130.085 69.775 130.130 ;
        RECT 70.390 130.070 70.710 130.130 ;
        RECT 71.770 130.070 72.090 130.330 ;
        RECT 74.990 130.070 75.310 130.330 ;
        RECT 14.660 129.450 127.820 129.930 ;
        RECT 17.735 129.250 18.025 129.295 ;
        RECT 23.470 129.250 23.790 129.310 ;
        RECT 17.735 129.110 27.840 129.250 ;
        RECT 17.735 129.065 18.025 129.110 ;
        RECT 23.470 129.050 23.790 129.110 ;
        RECT 19.740 128.910 20.030 128.955 ;
        RECT 21.170 128.910 21.490 128.970 ;
        RECT 23.000 128.910 23.290 128.955 ;
        RECT 19.740 128.770 23.290 128.910 ;
        RECT 19.740 128.725 20.030 128.770 ;
        RECT 21.170 128.710 21.490 128.770 ;
        RECT 23.000 128.725 23.290 128.770 ;
        RECT 23.920 128.910 24.210 128.955 ;
        RECT 25.780 128.910 26.070 128.955 ;
        RECT 23.920 128.770 26.070 128.910 ;
        RECT 27.700 128.910 27.840 129.110 ;
        RECT 34.050 129.050 34.370 129.310 ;
        RECT 37.730 129.250 38.050 129.310 ;
        RECT 38.665 129.250 38.955 129.295 ;
        RECT 37.730 129.110 38.955 129.250 ;
        RECT 37.730 129.050 38.050 129.110 ;
        RECT 38.665 129.065 38.955 129.110 ;
        RECT 41.885 129.250 42.175 129.295 ;
        RECT 43.710 129.250 44.030 129.310 ;
        RECT 41.885 129.110 44.030 129.250 ;
        RECT 41.885 129.065 42.175 129.110 ;
        RECT 43.710 129.050 44.030 129.110 ;
        RECT 44.185 129.250 44.475 129.295 ;
        RECT 45.090 129.250 45.410 129.310 ;
        RECT 44.185 129.110 45.410 129.250 ;
        RECT 44.185 129.065 44.475 129.110 ;
        RECT 45.090 129.050 45.410 129.110 ;
        RECT 49.245 129.250 49.535 129.295 ;
        RECT 49.690 129.250 50.010 129.310 ;
        RECT 49.245 129.110 50.010 129.250 ;
        RECT 49.245 129.065 49.535 129.110 ;
        RECT 49.690 129.050 50.010 129.110 ;
        RECT 55.670 129.250 55.990 129.310 ;
        RECT 56.145 129.250 56.435 129.295 ;
        RECT 55.670 129.110 56.435 129.250 ;
        RECT 55.670 129.050 55.990 129.110 ;
        RECT 56.145 129.065 56.435 129.110 ;
        RECT 56.590 129.050 56.910 129.310 ;
        RECT 65.115 129.250 65.405 129.295 ;
        RECT 66.250 129.250 66.570 129.310 ;
        RECT 65.115 129.110 66.570 129.250 ;
        RECT 65.115 129.065 65.405 129.110 ;
        RECT 66.250 129.050 66.570 129.110 ;
        RECT 77.840 129.110 81.660 129.250 ;
        RECT 42.790 128.910 43.110 128.970 ;
        RECT 46.945 128.910 47.235 128.955 ;
        RECT 63.950 128.910 64.270 128.970 ;
        RECT 27.700 128.770 40.260 128.910 ;
        RECT 23.920 128.725 24.210 128.770 ;
        RECT 25.780 128.725 26.070 128.770 ;
        RECT 21.600 128.570 21.890 128.615 ;
        RECT 23.920 128.570 24.135 128.725 ;
        RECT 21.600 128.430 24.135 128.570 ;
        RECT 26.705 128.570 26.995 128.615 ;
        RECT 29.910 128.570 30.230 128.630 ;
        RECT 26.705 128.430 30.230 128.570 ;
        RECT 21.600 128.385 21.890 128.430 ;
        RECT 26.705 128.385 26.995 128.430 ;
        RECT 29.910 128.370 30.230 128.430 ;
        RECT 30.370 128.570 30.690 128.630 ;
        RECT 33.605 128.570 33.895 128.615 ;
        RECT 30.370 128.430 33.895 128.570 ;
        RECT 30.370 128.370 30.690 128.430 ;
        RECT 33.605 128.385 33.895 128.430 ;
        RECT 39.570 128.370 39.890 128.630 ;
        RECT 40.120 128.615 40.260 128.770 ;
        RECT 42.790 128.770 64.270 128.910 ;
        RECT 42.790 128.710 43.110 128.770 ;
        RECT 46.945 128.725 47.235 128.770 ;
        RECT 63.950 128.710 64.270 128.770 ;
        RECT 67.120 128.910 67.410 128.955 ;
        RECT 68.550 128.910 68.870 128.970 ;
        RECT 70.380 128.910 70.670 128.955 ;
        RECT 67.120 128.770 70.670 128.910 ;
        RECT 67.120 128.725 67.410 128.770 ;
        RECT 68.550 128.710 68.870 128.770 ;
        RECT 70.380 128.725 70.670 128.770 ;
        RECT 71.300 128.910 71.590 128.955 ;
        RECT 73.160 128.910 73.450 128.955 ;
        RECT 71.300 128.770 73.450 128.910 ;
        RECT 71.300 128.725 71.590 128.770 ;
        RECT 73.160 128.725 73.450 128.770 ;
        RECT 40.045 128.385 40.335 128.615 ;
        RECT 40.965 128.570 41.255 128.615 ;
        RECT 43.265 128.570 43.555 128.615 ;
        RECT 46.010 128.570 46.330 128.630 ;
        RECT 48.325 128.570 48.615 128.615 ;
        RECT 68.090 128.570 68.410 128.630 ;
        RECT 40.965 128.430 68.410 128.570 ;
        RECT 40.965 128.385 41.255 128.430 ;
        RECT 43.265 128.385 43.555 128.430 ;
        RECT 46.010 128.370 46.330 128.430 ;
        RECT 48.325 128.385 48.615 128.430 ;
        RECT 68.090 128.370 68.410 128.430 ;
        RECT 68.980 128.570 69.270 128.615 ;
        RECT 71.300 128.570 71.515 128.725 ;
        RECT 68.980 128.430 71.515 128.570 ;
        RECT 68.980 128.385 69.270 128.430 ;
        RECT 72.230 128.370 72.550 128.630 ;
        RECT 74.990 128.570 75.310 128.630 ;
        RECT 77.840 128.615 77.980 129.110 ;
        RECT 78.685 128.910 78.975 128.955 ;
        RECT 80.510 128.910 80.830 128.970 ;
        RECT 78.685 128.770 80.830 128.910 ;
        RECT 81.520 128.910 81.660 129.110 ;
        RECT 83.270 129.050 83.590 129.310 ;
        RECT 88.330 129.050 88.650 129.310 ;
        RECT 89.725 129.065 90.015 129.295 ;
        RECT 81.520 128.770 84.420 128.910 ;
        RECT 78.685 128.725 78.975 128.770 ;
        RECT 80.510 128.710 80.830 128.770 ;
        RECT 84.280 128.615 84.420 128.770 ;
        RECT 84.740 128.770 85.800 128.910 ;
        RECT 75.465 128.570 75.755 128.615 ;
        RECT 77.765 128.570 78.055 128.615 ;
        RECT 80.985 128.570 81.275 128.615 ;
        RECT 74.990 128.430 78.055 128.570 ;
        RECT 74.990 128.370 75.310 128.430 ;
        RECT 75.465 128.385 75.755 128.430 ;
        RECT 77.765 128.385 78.055 128.430 ;
        RECT 79.220 128.430 81.275 128.570 ;
        RECT 23.930 128.230 24.250 128.290 ;
        RECT 24.865 128.230 25.155 128.275 ;
        RECT 23.930 128.090 25.155 128.230 ;
        RECT 23.930 128.030 24.250 128.090 ;
        RECT 24.865 128.045 25.155 128.090 ;
        RECT 42.345 128.045 42.635 128.275 ;
        RECT 42.790 128.230 43.110 128.290 ;
        RECT 47.405 128.230 47.695 128.275 ;
        RECT 42.790 128.090 47.695 128.230 ;
        RECT 21.600 127.890 21.890 127.935 ;
        RECT 24.380 127.890 24.670 127.935 ;
        RECT 26.240 127.890 26.530 127.935 ;
        RECT 21.600 127.750 26.530 127.890 ;
        RECT 21.600 127.705 21.890 127.750 ;
        RECT 24.380 127.705 24.670 127.750 ;
        RECT 26.240 127.705 26.530 127.750 ;
        RECT 22.550 127.550 22.870 127.610 ;
        RECT 42.420 127.550 42.560 128.045 ;
        RECT 42.790 128.030 43.110 128.090 ;
        RECT 47.405 128.045 47.695 128.090 ;
        RECT 54.750 128.230 55.070 128.290 ;
        RECT 55.225 128.230 55.515 128.275 ;
        RECT 54.750 128.090 55.515 128.230 ;
        RECT 54.750 128.030 55.070 128.090 ;
        RECT 55.225 128.045 55.515 128.090 ;
        RECT 63.950 128.230 64.270 128.290 ;
        RECT 74.085 128.230 74.375 128.275 ;
        RECT 63.950 128.090 74.375 128.230 ;
        RECT 63.950 128.030 64.270 128.090 ;
        RECT 74.085 128.045 74.375 128.090 ;
        RECT 74.545 128.045 74.835 128.275 ;
        RECT 76.845 128.230 77.135 128.275 ;
        RECT 78.670 128.230 78.990 128.290 ;
        RECT 79.220 128.230 79.360 128.430 ;
        RECT 80.985 128.385 81.275 128.430 ;
        RECT 84.205 128.385 84.495 128.615 ;
        RECT 76.845 128.090 79.360 128.230 ;
        RECT 76.845 128.045 77.135 128.090 ;
        RECT 68.980 127.890 69.270 127.935 ;
        RECT 71.760 127.890 72.050 127.935 ;
        RECT 73.620 127.890 73.910 127.935 ;
        RECT 68.980 127.750 73.910 127.890 ;
        RECT 74.620 127.890 74.760 128.045 ;
        RECT 78.670 128.030 78.990 128.090 ;
        RECT 80.065 128.045 80.355 128.275 ;
        RECT 79.130 127.890 79.450 127.950 ;
        RECT 74.620 127.750 79.450 127.890 ;
        RECT 80.140 127.890 80.280 128.045 ;
        RECT 80.510 128.030 80.830 128.290 ;
        RECT 81.060 128.230 81.200 128.385 ;
        RECT 84.740 128.230 84.880 128.770 ;
        RECT 85.125 128.385 85.415 128.615 ;
        RECT 81.060 128.090 84.880 128.230 ;
        RECT 85.200 127.890 85.340 128.385 ;
        RECT 85.660 128.230 85.800 128.770 ;
        RECT 87.425 128.570 87.715 128.615 ;
        RECT 89.800 128.570 89.940 129.065 ;
        RECT 95.230 129.050 95.550 129.310 ;
        RECT 98.450 129.250 98.770 129.310 ;
        RECT 102.145 129.250 102.435 129.295 ;
        RECT 98.450 129.110 102.435 129.250 ;
        RECT 98.450 129.050 98.770 129.110 ;
        RECT 102.145 129.065 102.435 129.110 ;
        RECT 104.890 129.050 105.210 129.310 ;
        RECT 106.270 129.250 106.590 129.310 ;
        RECT 107.205 129.250 107.495 129.295 ;
        RECT 106.270 129.110 107.495 129.250 ;
        RECT 106.270 129.050 106.590 129.110 ;
        RECT 107.205 129.065 107.495 129.110 ;
        RECT 111.330 129.050 111.650 129.310 ;
        RECT 95.690 128.710 96.010 128.970 ;
        RECT 105.900 128.770 108.340 128.910 ;
        RECT 87.425 128.430 89.940 128.570 ;
        RECT 91.565 128.570 91.855 128.615 ;
        RECT 93.850 128.570 94.170 128.630 ;
        RECT 94.325 128.570 94.615 128.615 ;
        RECT 91.565 128.430 93.620 128.570 ;
        RECT 87.425 128.385 87.715 128.430 ;
        RECT 91.565 128.385 91.855 128.430 ;
        RECT 92.025 128.230 92.315 128.275 ;
        RECT 85.660 128.090 92.315 128.230 ;
        RECT 92.025 128.045 92.315 128.090 ;
        RECT 92.485 128.045 92.775 128.275 ;
        RECT 93.480 128.230 93.620 128.430 ;
        RECT 93.850 128.430 94.615 128.570 ;
        RECT 93.850 128.370 94.170 128.430 ;
        RECT 94.325 128.385 94.615 128.430 ;
        RECT 100.290 128.570 100.610 128.630 ;
        RECT 105.900 128.615 106.040 128.770 ;
        RECT 105.825 128.570 106.115 128.615 ;
        RECT 100.290 128.430 106.115 128.570 ;
        RECT 100.290 128.370 100.610 128.430 ;
        RECT 105.825 128.385 106.115 128.430 ;
        RECT 106.270 128.370 106.590 128.630 ;
        RECT 108.200 128.615 108.340 128.770 ;
        RECT 108.125 128.570 108.415 128.615 ;
        RECT 110.425 128.570 110.715 128.615 ;
        RECT 110.870 128.570 111.190 128.630 ;
        RECT 112.725 128.570 113.015 128.615 ;
        RECT 108.125 128.430 113.015 128.570 ;
        RECT 108.125 128.385 108.415 128.430 ;
        RECT 110.425 128.385 110.715 128.430 ;
        RECT 110.870 128.370 111.190 128.430 ;
        RECT 112.725 128.385 113.015 128.430 ;
        RECT 113.170 128.370 113.490 128.630 ;
        RECT 118.230 128.370 118.550 128.630 ;
        RECT 119.625 128.385 119.915 128.615 ;
        RECT 98.910 128.230 99.230 128.290 ;
        RECT 105.350 128.230 105.670 128.290 ;
        RECT 109.045 128.230 109.335 128.275 ;
        RECT 93.480 128.090 109.335 128.230 ;
        RECT 91.550 127.890 91.870 127.950 ;
        RECT 80.140 127.750 84.880 127.890 ;
        RECT 85.200 127.750 91.870 127.890 ;
        RECT 68.980 127.705 69.270 127.750 ;
        RECT 71.760 127.705 72.050 127.750 ;
        RECT 73.620 127.705 73.910 127.750 ;
        RECT 79.130 127.690 79.450 127.750 ;
        RECT 84.740 127.610 84.880 127.750 ;
        RECT 91.550 127.690 91.870 127.750 ;
        RECT 22.550 127.410 42.560 127.550 ;
        RECT 57.970 127.550 58.290 127.610 ;
        RECT 58.445 127.550 58.735 127.595 ;
        RECT 57.970 127.410 58.735 127.550 ;
        RECT 22.550 127.350 22.870 127.410 ;
        RECT 57.970 127.350 58.290 127.410 ;
        RECT 58.445 127.365 58.735 127.410 ;
        RECT 76.385 127.550 76.675 127.595 ;
        RECT 81.890 127.550 82.210 127.610 ;
        RECT 76.385 127.410 82.210 127.550 ;
        RECT 76.385 127.365 76.675 127.410 ;
        RECT 81.890 127.350 82.210 127.410 ;
        RECT 82.825 127.550 83.115 127.595 ;
        RECT 83.730 127.550 84.050 127.610 ;
        RECT 82.825 127.410 84.050 127.550 ;
        RECT 82.825 127.365 83.115 127.410 ;
        RECT 83.730 127.350 84.050 127.410 ;
        RECT 84.650 127.550 84.970 127.610 ;
        RECT 92.560 127.550 92.700 128.045 ;
        RECT 98.910 128.030 99.230 128.090 ;
        RECT 105.350 128.030 105.670 128.090 ;
        RECT 109.045 128.045 109.335 128.090 ;
        RECT 109.490 128.030 109.810 128.290 ;
        RECT 115.010 128.230 115.330 128.290 ;
        RECT 119.700 128.230 119.840 128.385 ;
        RECT 115.010 128.090 119.840 128.230 ;
        RECT 115.010 128.030 115.330 128.090 ;
        RECT 103.050 127.890 103.370 127.950 ;
        RECT 111.805 127.890 112.095 127.935 ;
        RECT 103.050 127.750 112.095 127.890 ;
        RECT 103.050 127.690 103.370 127.750 ;
        RECT 111.805 127.705 112.095 127.750 ;
        RECT 84.650 127.410 92.700 127.550 ;
        RECT 84.650 127.350 84.970 127.410 ;
        RECT 118.690 127.350 119.010 127.610 ;
        RECT 120.530 127.350 120.850 127.610 ;
        RECT 14.660 126.730 127.820 127.210 ;
        RECT 23.930 126.330 24.250 126.590 ;
        RECT 71.325 126.530 71.615 126.575 ;
        RECT 72.230 126.530 72.550 126.590 ;
        RECT 78.670 126.575 78.990 126.590 ;
        RECT 71.325 126.390 72.550 126.530 ;
        RECT 71.325 126.345 71.615 126.390 ;
        RECT 72.230 126.330 72.550 126.390 ;
        RECT 78.455 126.345 78.990 126.575 ;
        RECT 78.670 126.330 78.990 126.345 ;
        RECT 79.130 126.530 79.450 126.590 ;
        RECT 80.510 126.530 80.830 126.590 ;
        RECT 98.910 126.575 99.230 126.590 ;
        RECT 79.130 126.390 80.830 126.530 ;
        RECT 79.130 126.330 79.450 126.390 ;
        RECT 80.510 126.330 80.830 126.390 ;
        RECT 98.695 126.345 99.230 126.575 ;
        RECT 98.910 126.330 99.230 126.345 ;
        RECT 115.010 126.330 115.330 126.590 ;
        RECT 55.670 126.190 55.990 126.250 ;
        RECT 82.320 126.190 82.610 126.235 ;
        RECT 85.100 126.190 85.390 126.235 ;
        RECT 86.960 126.190 87.250 126.235 ;
        RECT 55.670 126.050 60.960 126.190 ;
        RECT 55.670 125.990 55.990 126.050 ;
        RECT 19.790 125.850 20.110 125.910 ;
        RECT 30.370 125.850 30.690 125.910 ;
        RECT 19.790 125.710 30.690 125.850 ;
        RECT 19.790 125.650 20.110 125.710 ;
        RECT 21.170 125.510 21.490 125.570 ;
        RECT 22.180 125.555 22.320 125.710 ;
        RECT 30.370 125.650 30.690 125.710 ;
        RECT 35.890 125.850 36.210 125.910 ;
        RECT 42.805 125.850 43.095 125.895 ;
        RECT 54.750 125.850 55.070 125.910 ;
        RECT 59.825 125.850 60.115 125.895 ;
        RECT 35.890 125.710 43.095 125.850 ;
        RECT 35.890 125.650 36.210 125.710 ;
        RECT 42.805 125.665 43.095 125.710 ;
        RECT 43.800 125.710 46.240 125.850 ;
        RECT 21.645 125.510 21.935 125.555 ;
        RECT 21.170 125.370 21.935 125.510 ;
        RECT 21.170 125.310 21.490 125.370 ;
        RECT 21.645 125.325 21.935 125.370 ;
        RECT 22.105 125.325 22.395 125.555 ;
        RECT 23.010 125.310 23.330 125.570 ;
        RECT 36.810 125.310 37.130 125.570 ;
        RECT 37.745 125.325 38.035 125.555 ;
        RECT 38.190 125.510 38.510 125.570 ;
        RECT 38.665 125.510 38.955 125.555 ;
        RECT 38.190 125.370 38.955 125.510 ;
        RECT 37.820 125.170 37.960 125.325 ;
        RECT 38.190 125.310 38.510 125.370 ;
        RECT 38.665 125.325 38.955 125.370 ;
        RECT 40.490 125.310 40.810 125.570 ;
        RECT 41.425 125.325 41.715 125.555 ;
        RECT 40.030 125.170 40.350 125.230 ;
        RECT 37.820 125.030 40.350 125.170 ;
        RECT 41.500 125.170 41.640 125.325 ;
        RECT 42.330 125.310 42.650 125.570 ;
        RECT 43.800 125.555 43.940 125.710 ;
        RECT 46.100 125.570 46.240 125.710 ;
        RECT 54.750 125.710 60.115 125.850 ;
        RECT 60.820 125.850 60.960 126.050 ;
        RECT 82.320 126.050 87.250 126.190 ;
        RECT 82.320 126.005 82.610 126.050 ;
        RECT 85.100 126.005 85.390 126.050 ;
        RECT 86.960 126.005 87.250 126.050 ;
        RECT 90.190 126.190 90.480 126.235 ;
        RECT 92.050 126.190 92.340 126.235 ;
        RECT 94.830 126.190 95.120 126.235 ;
        RECT 90.190 126.050 95.120 126.190 ;
        RECT 90.190 126.005 90.480 126.050 ;
        RECT 92.050 126.005 92.340 126.050 ;
        RECT 94.830 126.005 95.120 126.050 ;
        RECT 119.580 126.190 119.870 126.235 ;
        RECT 122.360 126.190 122.650 126.235 ;
        RECT 124.220 126.190 124.510 126.235 ;
        RECT 119.580 126.050 124.510 126.190 ;
        RECT 119.580 126.005 119.870 126.050 ;
        RECT 122.360 126.005 122.650 126.050 ;
        RECT 124.220 126.005 124.510 126.050 ;
        RECT 74.545 125.850 74.835 125.895 ;
        RECT 79.590 125.850 79.910 125.910 ;
        RECT 84.650 125.850 84.970 125.910 ;
        RECT 60.820 125.710 61.420 125.850 ;
        RECT 54.750 125.650 55.070 125.710 ;
        RECT 59.825 125.665 60.115 125.710 ;
        RECT 43.725 125.510 44.015 125.555 ;
        RECT 42.880 125.370 44.015 125.510 ;
        RECT 42.880 125.170 43.020 125.370 ;
        RECT 43.725 125.325 44.015 125.370 ;
        RECT 44.630 125.310 44.950 125.570 ;
        RECT 46.010 125.310 46.330 125.570 ;
        RECT 46.470 125.310 46.790 125.570 ;
        RECT 57.970 125.310 58.290 125.570 ;
        RECT 60.730 125.310 61.050 125.570 ;
        RECT 61.280 125.555 61.420 125.710 ;
        RECT 74.545 125.710 84.970 125.850 ;
        RECT 74.545 125.665 74.835 125.710 ;
        RECT 79.590 125.650 79.910 125.710 ;
        RECT 84.650 125.650 84.970 125.710 ;
        RECT 88.330 125.850 88.650 125.910 ;
        RECT 91.565 125.850 91.855 125.895 ;
        RECT 98.450 125.850 98.770 125.910 ;
        RECT 88.330 125.710 91.855 125.850 ;
        RECT 88.330 125.650 88.650 125.710 ;
        RECT 91.565 125.665 91.855 125.710 ;
        RECT 92.100 125.710 98.770 125.850 ;
        RECT 61.205 125.325 61.495 125.555 ;
        RECT 68.550 125.510 68.870 125.570 ;
        RECT 69.025 125.510 69.315 125.555 ;
        RECT 68.550 125.370 69.315 125.510 ;
        RECT 68.550 125.310 68.870 125.370 ;
        RECT 69.025 125.325 69.315 125.370 ;
        RECT 69.485 125.510 69.775 125.555 ;
        RECT 69.930 125.510 70.250 125.570 ;
        RECT 69.485 125.370 70.250 125.510 ;
        RECT 69.485 125.325 69.775 125.370 ;
        RECT 69.930 125.310 70.250 125.370 ;
        RECT 70.390 125.310 70.710 125.570 ;
        RECT 71.770 125.510 72.090 125.570 ;
        RECT 73.165 125.510 73.455 125.555 ;
        RECT 71.170 125.370 73.455 125.510 ;
        RECT 41.500 125.030 43.020 125.170 ;
        RECT 43.250 125.170 43.570 125.230 ;
        RECT 45.105 125.170 45.395 125.215 ;
        RECT 43.250 125.030 45.395 125.170 ;
        RECT 40.030 124.970 40.350 125.030 ;
        RECT 43.250 124.970 43.570 125.030 ;
        RECT 45.105 124.985 45.395 125.030 ;
        RECT 49.245 125.170 49.535 125.215 ;
        RECT 71.170 125.170 71.310 125.370 ;
        RECT 71.770 125.310 72.090 125.370 ;
        RECT 73.165 125.325 73.455 125.370 ;
        RECT 82.320 125.510 82.610 125.555 ;
        RECT 82.320 125.370 84.855 125.510 ;
        RECT 82.320 125.325 82.610 125.370 ;
        RECT 49.245 125.030 71.310 125.170 ;
        RECT 80.460 125.170 80.750 125.215 ;
        RECT 82.810 125.170 83.130 125.230 ;
        RECT 84.640 125.215 84.855 125.370 ;
        RECT 85.570 125.310 85.890 125.570 ;
        RECT 87.425 125.510 87.715 125.555 ;
        RECT 89.725 125.510 90.015 125.555 ;
        RECT 92.100 125.510 92.240 125.710 ;
        RECT 98.450 125.650 98.770 125.710 ;
        RECT 112.265 125.850 112.555 125.895 ;
        RECT 113.630 125.850 113.950 125.910 ;
        RECT 112.265 125.710 113.950 125.850 ;
        RECT 112.265 125.665 112.555 125.710 ;
        RECT 113.630 125.650 113.950 125.710 ;
        RECT 120.530 125.850 120.850 125.910 ;
        RECT 122.845 125.850 123.135 125.895 ;
        RECT 120.530 125.710 123.135 125.850 ;
        RECT 120.530 125.650 120.850 125.710 ;
        RECT 122.845 125.665 123.135 125.710 ;
        RECT 94.830 125.510 95.120 125.555 ;
        RECT 87.425 125.370 92.240 125.510 ;
        RECT 92.585 125.370 95.120 125.510 ;
        RECT 87.425 125.325 87.715 125.370 ;
        RECT 89.725 125.325 90.015 125.370 ;
        RECT 92.585 125.215 92.800 125.370 ;
        RECT 94.830 125.325 95.120 125.370 ;
        RECT 99.370 125.310 99.690 125.570 ;
        RECT 100.290 125.310 100.610 125.570 ;
        RECT 101.210 125.310 101.530 125.570 ;
        RECT 105.350 125.510 105.670 125.570 ;
        RECT 112.725 125.510 113.015 125.555 ;
        RECT 105.350 125.370 113.015 125.510 ;
        RECT 105.350 125.310 105.670 125.370 ;
        RECT 112.725 125.325 113.015 125.370 ;
        RECT 119.580 125.510 119.870 125.555 ;
        RECT 119.580 125.370 122.115 125.510 ;
        RECT 119.580 125.325 119.870 125.370 ;
        RECT 83.720 125.170 84.010 125.215 ;
        RECT 80.460 125.030 84.010 125.170 ;
        RECT 49.245 124.985 49.535 125.030 ;
        RECT 80.460 124.985 80.750 125.030 ;
        RECT 82.810 124.970 83.130 125.030 ;
        RECT 83.720 124.985 84.010 125.030 ;
        RECT 84.640 125.170 84.930 125.215 ;
        RECT 86.500 125.170 86.790 125.215 ;
        RECT 84.640 125.030 86.790 125.170 ;
        RECT 84.640 124.985 84.930 125.030 ;
        RECT 86.500 124.985 86.790 125.030 ;
        RECT 90.650 125.170 90.940 125.215 ;
        RECT 92.510 125.170 92.800 125.215 ;
        RECT 90.650 125.030 92.800 125.170 ;
        RECT 90.650 124.985 90.940 125.030 ;
        RECT 92.510 124.985 92.800 125.030 ;
        RECT 93.390 125.215 93.710 125.230 ;
        RECT 93.390 125.170 93.720 125.215 ;
        RECT 96.690 125.170 96.980 125.215 ;
        RECT 93.390 125.030 96.980 125.170 ;
        RECT 93.390 124.985 93.720 125.030 ;
        RECT 96.690 124.985 96.980 125.030 ;
        RECT 117.720 125.170 118.010 125.215 ;
        RECT 118.690 125.170 119.010 125.230 ;
        RECT 121.900 125.215 122.115 125.370 ;
        RECT 124.670 125.310 124.990 125.570 ;
        RECT 120.980 125.170 121.270 125.215 ;
        RECT 117.720 125.030 121.270 125.170 ;
        RECT 117.720 124.985 118.010 125.030 ;
        RECT 93.390 124.970 93.710 124.985 ;
        RECT 118.690 124.970 119.010 125.030 ;
        RECT 120.980 124.985 121.270 125.030 ;
        RECT 121.900 125.170 122.190 125.215 ;
        RECT 123.760 125.170 124.050 125.215 ;
        RECT 121.900 125.030 124.050 125.170 ;
        RECT 121.900 124.985 122.190 125.030 ;
        RECT 123.760 124.985 124.050 125.030 ;
        RECT 46.010 124.830 46.330 124.890 ;
        RECT 47.865 124.830 48.155 124.875 ;
        RECT 46.010 124.690 48.155 124.830 ;
        RECT 46.010 124.630 46.330 124.690 ;
        RECT 47.865 124.645 48.155 124.690 ;
        RECT 58.905 124.830 59.195 124.875 ;
        RECT 60.270 124.830 60.590 124.890 ;
        RECT 58.905 124.690 60.590 124.830 ;
        RECT 58.905 124.645 59.195 124.690 ;
        RECT 60.270 124.630 60.590 124.690 ;
        RECT 63.045 124.830 63.335 124.875 ;
        RECT 69.930 124.830 70.250 124.890 ;
        RECT 63.045 124.690 70.250 124.830 ;
        RECT 63.045 124.645 63.335 124.690 ;
        RECT 69.930 124.630 70.250 124.690 ;
        RECT 113.170 124.830 113.490 124.890 ;
        RECT 115.715 124.830 116.005 124.875 ;
        RECT 113.170 124.690 116.005 124.830 ;
        RECT 113.170 124.630 113.490 124.690 ;
        RECT 115.715 124.645 116.005 124.690 ;
        RECT 14.660 124.010 127.820 124.490 ;
        RECT 22.550 123.810 22.870 123.870 ;
        RECT 23.470 123.810 23.790 123.870 ;
        RECT 24.405 123.810 24.695 123.855 ;
        RECT 22.550 123.610 23.010 123.810 ;
        RECT 23.470 123.670 24.695 123.810 ;
        RECT 23.470 123.610 23.790 123.670 ;
        RECT 24.405 123.625 24.695 123.670 ;
        RECT 24.865 123.810 25.155 123.855 ;
        RECT 42.790 123.810 43.110 123.870 ;
        RECT 24.865 123.670 43.110 123.810 ;
        RECT 24.865 123.625 25.155 123.670 ;
        RECT 22.870 123.470 23.010 123.610 ;
        RECT 24.940 123.470 25.080 123.625 ;
        RECT 42.790 123.610 43.110 123.670 ;
        RECT 53.155 123.810 53.445 123.855 ;
        RECT 55.670 123.810 55.990 123.870 ;
        RECT 53.155 123.670 55.990 123.810 ;
        RECT 53.155 123.625 53.445 123.670 ;
        RECT 55.670 123.610 55.990 123.670 ;
        RECT 60.730 123.810 61.050 123.870 ;
        RECT 65.805 123.810 66.095 123.855 ;
        RECT 60.730 123.670 66.095 123.810 ;
        RECT 60.730 123.610 61.050 123.670 ;
        RECT 65.805 123.625 66.095 123.670 ;
        RECT 82.365 123.810 82.655 123.855 ;
        RECT 82.810 123.810 83.130 123.870 ;
        RECT 82.365 123.670 83.130 123.810 ;
        RECT 82.365 123.625 82.655 123.670 ;
        RECT 82.810 123.610 83.130 123.670 ;
        RECT 84.665 123.810 84.955 123.855 ;
        RECT 85.570 123.810 85.890 123.870 ;
        RECT 84.665 123.670 85.890 123.810 ;
        RECT 84.665 123.625 84.955 123.670 ;
        RECT 85.570 123.610 85.890 123.670 ;
        RECT 93.390 123.610 93.710 123.870 ;
        RECT 22.870 123.330 25.080 123.470 ;
        RECT 55.160 123.470 55.450 123.515 ;
        RECT 57.510 123.470 57.830 123.530 ;
        RECT 58.420 123.470 58.710 123.515 ;
        RECT 55.160 123.330 58.710 123.470 ;
        RECT 55.160 123.285 55.450 123.330 ;
        RECT 57.510 123.270 57.830 123.330 ;
        RECT 58.420 123.285 58.710 123.330 ;
        RECT 59.340 123.470 59.630 123.515 ;
        RECT 61.200 123.470 61.490 123.515 ;
        RECT 59.340 123.330 61.490 123.470 ;
        RECT 59.340 123.285 59.630 123.330 ;
        RECT 61.200 123.285 61.490 123.330 ;
        RECT 111.805 123.470 112.095 123.515 ;
        RECT 113.170 123.470 113.490 123.530 ;
        RECT 111.805 123.330 113.490 123.470 ;
        RECT 111.805 123.285 112.095 123.330 ;
        RECT 34.970 122.930 35.290 123.190 ;
        RECT 57.020 123.130 57.310 123.175 ;
        RECT 59.340 123.130 59.555 123.285 ;
        RECT 113.170 123.270 113.490 123.330 ;
        RECT 117.720 123.470 118.010 123.515 ;
        RECT 119.150 123.470 119.470 123.530 ;
        RECT 120.980 123.470 121.270 123.515 ;
        RECT 117.720 123.330 121.270 123.470 ;
        RECT 117.720 123.285 118.010 123.330 ;
        RECT 119.150 123.270 119.470 123.330 ;
        RECT 120.980 123.285 121.270 123.330 ;
        RECT 121.900 123.470 122.190 123.515 ;
        RECT 123.760 123.470 124.050 123.515 ;
        RECT 121.900 123.330 124.050 123.470 ;
        RECT 121.900 123.285 122.190 123.330 ;
        RECT 123.760 123.285 124.050 123.330 ;
        RECT 57.020 122.990 59.555 123.130 ;
        RECT 57.020 122.945 57.310 122.990 ;
        RECT 60.270 122.930 60.590 123.190 ;
        RECT 62.125 123.130 62.415 123.175 ;
        RECT 63.950 123.130 64.270 123.190 ;
        RECT 62.125 122.990 64.270 123.130 ;
        RECT 62.125 122.945 62.415 122.990 ;
        RECT 63.950 122.930 64.270 122.990 ;
        RECT 64.410 123.130 64.730 123.190 ;
        RECT 65.345 123.130 65.635 123.175 ;
        RECT 64.410 122.990 65.635 123.130 ;
        RECT 64.410 122.930 64.730 122.990 ;
        RECT 65.345 122.945 65.635 122.990 ;
        RECT 73.150 123.130 73.470 123.190 ;
        RECT 82.825 123.130 83.115 123.175 ;
        RECT 83.270 123.130 83.590 123.190 ;
        RECT 73.150 122.990 83.590 123.130 ;
        RECT 73.150 122.930 73.470 122.990 ;
        RECT 82.825 122.945 83.115 122.990 ;
        RECT 83.270 122.930 83.590 122.990 ;
        RECT 83.730 122.930 84.050 123.190 ;
        RECT 91.090 123.130 91.410 123.190 ;
        RECT 92.945 123.130 93.235 123.175 ;
        RECT 100.290 123.130 100.610 123.190 ;
        RECT 91.090 122.990 100.610 123.130 ;
        RECT 91.090 122.930 91.410 122.990 ;
        RECT 92.945 122.945 93.235 122.990 ;
        RECT 100.290 122.930 100.610 122.990 ;
        RECT 112.265 123.130 112.555 123.175 ;
        RECT 112.710 123.130 113.030 123.190 ;
        RECT 115.715 123.130 116.005 123.175 ;
        RECT 112.265 122.990 116.005 123.130 ;
        RECT 112.265 122.945 112.555 122.990 ;
        RECT 112.710 122.930 113.030 122.990 ;
        RECT 115.715 122.945 116.005 122.990 ;
        RECT 119.580 123.130 119.870 123.175 ;
        RECT 121.900 123.130 122.115 123.285 ;
        RECT 119.580 122.990 122.115 123.130 ;
        RECT 119.580 122.945 119.870 122.990 ;
        RECT 124.670 122.930 124.990 123.190 ;
        RECT 22.090 122.790 22.410 122.850 ;
        RECT 23.485 122.790 23.775 122.835 ;
        RECT 33.605 122.790 33.895 122.835 ;
        RECT 22.090 122.650 33.895 122.790 ;
        RECT 22.090 122.590 22.410 122.650 ;
        RECT 23.485 122.605 23.775 122.650 ;
        RECT 33.605 122.605 33.895 122.650 ;
        RECT 34.525 122.790 34.815 122.835 ;
        RECT 36.810 122.790 37.130 122.850 ;
        RECT 41.870 122.790 42.190 122.850 ;
        RECT 34.525 122.650 42.190 122.790 ;
        RECT 34.525 122.605 34.815 122.650 ;
        RECT 33.680 122.450 33.820 122.605 ;
        RECT 36.810 122.590 37.130 122.650 ;
        RECT 41.870 122.590 42.190 122.650 ;
        RECT 64.870 122.590 65.190 122.850 ;
        RECT 105.350 122.790 105.670 122.850 ;
        RECT 110.885 122.790 111.175 122.835 ;
        RECT 113.630 122.790 113.950 122.850 ;
        RECT 105.350 122.650 113.950 122.790 ;
        RECT 105.350 122.590 105.670 122.650 ;
        RECT 110.885 122.605 111.175 122.650 ;
        RECT 113.630 122.590 113.950 122.650 ;
        RECT 121.450 122.790 121.770 122.850 ;
        RECT 122.845 122.790 123.135 122.835 ;
        RECT 121.450 122.650 123.135 122.790 ;
        RECT 121.450 122.590 121.770 122.650 ;
        RECT 122.845 122.605 123.135 122.650 ;
        RECT 43.710 122.450 44.030 122.510 ;
        RECT 46.010 122.450 46.330 122.510 ;
        RECT 46.930 122.450 47.250 122.510 ;
        RECT 33.680 122.310 47.250 122.450 ;
        RECT 43.710 122.250 44.030 122.310 ;
        RECT 46.010 122.250 46.330 122.310 ;
        RECT 46.930 122.250 47.250 122.310 ;
        RECT 57.020 122.450 57.310 122.495 ;
        RECT 59.800 122.450 60.090 122.495 ;
        RECT 61.660 122.450 61.950 122.495 ;
        RECT 57.020 122.310 61.950 122.450 ;
        RECT 57.020 122.265 57.310 122.310 ;
        RECT 59.800 122.265 60.090 122.310 ;
        RECT 61.660 122.265 61.950 122.310 ;
        RECT 119.580 122.450 119.870 122.495 ;
        RECT 122.360 122.450 122.650 122.495 ;
        RECT 124.220 122.450 124.510 122.495 ;
        RECT 119.580 122.310 124.510 122.450 ;
        RECT 119.580 122.265 119.870 122.310 ;
        RECT 122.360 122.265 122.650 122.310 ;
        RECT 124.220 122.265 124.510 122.310 ;
        RECT 26.690 121.910 27.010 122.170 ;
        RECT 36.810 121.910 37.130 122.170 ;
        RECT 67.645 122.110 67.935 122.155 ;
        RECT 68.090 122.110 68.410 122.170 ;
        RECT 67.645 121.970 68.410 122.110 ;
        RECT 67.645 121.925 67.935 121.970 ;
        RECT 68.090 121.910 68.410 121.970 ;
        RECT 114.105 122.110 114.395 122.155 ;
        RECT 120.530 122.110 120.850 122.170 ;
        RECT 114.105 121.970 120.850 122.110 ;
        RECT 114.105 121.925 114.395 121.970 ;
        RECT 120.530 121.910 120.850 121.970 ;
        RECT 14.660 121.290 127.820 121.770 ;
        RECT 30.615 121.090 30.905 121.135 ;
        RECT 34.970 121.090 35.290 121.150 ;
        RECT 30.615 120.950 35.290 121.090 ;
        RECT 30.615 120.905 30.905 120.950 ;
        RECT 34.970 120.890 35.290 120.950 ;
        RECT 57.510 120.890 57.830 121.150 ;
        RECT 59.595 121.090 59.885 121.135 ;
        RECT 60.730 121.090 61.050 121.150 ;
        RECT 59.595 120.950 61.050 121.090 ;
        RECT 59.595 120.905 59.885 120.950 ;
        RECT 60.730 120.890 61.050 120.950 ;
        RECT 119.150 120.890 119.470 121.150 ;
        RECT 121.450 120.890 121.770 121.150 ;
        RECT 22.090 120.750 22.410 120.810 ;
        RECT 34.480 120.750 34.770 120.795 ;
        RECT 37.260 120.750 37.550 120.795 ;
        RECT 39.120 120.750 39.410 120.795 ;
        RECT 63.460 120.750 63.750 120.795 ;
        RECT 66.240 120.750 66.530 120.795 ;
        RECT 68.100 120.750 68.390 120.795 ;
        RECT 22.090 120.610 23.240 120.750 ;
        RECT 22.090 120.550 22.410 120.610 ;
        RECT 22.550 120.210 22.870 120.470 ;
        RECT 23.100 120.455 23.240 120.610 ;
        RECT 34.480 120.610 39.410 120.750 ;
        RECT 34.480 120.565 34.770 120.610 ;
        RECT 37.260 120.565 37.550 120.610 ;
        RECT 39.120 120.565 39.410 120.610 ;
        RECT 42.880 120.610 47.620 120.750 ;
        RECT 23.025 120.225 23.315 120.455 ;
        RECT 35.890 120.410 36.210 120.470 ;
        RECT 42.880 120.410 43.020 120.610 ;
        RECT 30.920 120.270 43.020 120.410 ;
        RECT 43.265 120.410 43.555 120.455 ;
        RECT 43.710 120.410 44.030 120.470 ;
        RECT 43.265 120.270 44.030 120.410 ;
        RECT 26.690 120.070 27.010 120.130 ;
        RECT 27.165 120.070 27.455 120.115 ;
        RECT 26.690 119.930 27.455 120.070 ;
        RECT 26.690 119.870 27.010 119.930 ;
        RECT 27.165 119.885 27.455 119.930 ;
        RECT 30.920 119.790 31.060 120.270 ;
        RECT 35.890 120.210 36.210 120.270 ;
        RECT 43.265 120.225 43.555 120.270 ;
        RECT 43.710 120.210 44.030 120.270 ;
        RECT 46.470 120.210 46.790 120.470 ;
        RECT 46.930 120.210 47.250 120.470 ;
        RECT 47.480 120.455 47.620 120.610 ;
        RECT 63.460 120.610 68.390 120.750 ;
        RECT 63.460 120.565 63.750 120.610 ;
        RECT 66.240 120.565 66.530 120.610 ;
        RECT 68.100 120.565 68.390 120.610 ;
        RECT 69.025 120.565 69.315 120.795 ;
        RECT 113.140 120.750 113.430 120.795 ;
        RECT 115.920 120.750 116.210 120.795 ;
        RECT 117.780 120.750 118.070 120.795 ;
        RECT 113.140 120.610 118.070 120.750 ;
        RECT 113.140 120.565 113.430 120.610 ;
        RECT 115.920 120.565 116.210 120.610 ;
        RECT 117.780 120.565 118.070 120.610 ;
        RECT 47.405 120.225 47.695 120.455 ;
        RECT 66.725 120.410 67.015 120.455 ;
        RECT 69.100 120.410 69.240 120.565 ;
        RECT 66.725 120.270 69.240 120.410 ;
        RECT 77.765 120.410 78.055 120.455 ;
        RECT 79.590 120.410 79.910 120.470 ;
        RECT 83.730 120.410 84.050 120.470 ;
        RECT 93.865 120.410 94.155 120.455 ;
        RECT 98.005 120.410 98.295 120.455 ;
        RECT 105.350 120.410 105.670 120.470 ;
        RECT 109.490 120.455 109.810 120.470 ;
        RECT 77.765 120.270 105.670 120.410 ;
        RECT 66.725 120.225 67.015 120.270 ;
        RECT 77.765 120.225 78.055 120.270 ;
        RECT 79.590 120.210 79.910 120.270 ;
        RECT 83.730 120.210 84.050 120.270 ;
        RECT 93.865 120.225 94.155 120.270 ;
        RECT 98.005 120.225 98.295 120.270 ;
        RECT 105.350 120.210 105.670 120.270 ;
        RECT 106.285 120.410 106.575 120.455 ;
        RECT 109.275 120.410 109.810 120.455 ;
        RECT 106.285 120.270 109.810 120.410 ;
        RECT 106.285 120.225 106.575 120.270 ;
        RECT 109.275 120.225 109.810 120.270 ;
        RECT 109.490 120.210 109.810 120.225 ;
        RECT 110.040 120.270 118.920 120.410 ;
        RECT 34.480 120.070 34.770 120.115 ;
        RECT 34.480 119.930 37.015 120.070 ;
        RECT 34.480 119.885 34.770 119.930 ;
        RECT 22.105 119.730 22.395 119.775 ;
        RECT 30.830 119.730 31.150 119.790 ;
        RECT 22.105 119.590 31.150 119.730 ;
        RECT 22.105 119.545 22.395 119.590 ;
        RECT 30.830 119.530 31.150 119.590 ;
        RECT 32.620 119.730 32.910 119.775 ;
        RECT 34.970 119.730 35.290 119.790 ;
        RECT 36.800 119.775 37.015 119.930 ;
        RECT 37.730 119.870 38.050 120.130 ;
        RECT 39.585 119.885 39.875 120.115 ;
        RECT 35.880 119.730 36.170 119.775 ;
        RECT 32.620 119.590 36.170 119.730 ;
        RECT 32.620 119.545 32.910 119.590 ;
        RECT 34.970 119.530 35.290 119.590 ;
        RECT 35.880 119.545 36.170 119.590 ;
        RECT 36.800 119.730 37.090 119.775 ;
        RECT 38.660 119.730 38.950 119.775 ;
        RECT 36.800 119.590 38.950 119.730 ;
        RECT 39.660 119.730 39.800 119.885 ;
        RECT 41.870 119.870 42.190 120.130 ;
        RECT 45.550 119.870 45.870 120.130 ;
        RECT 46.560 120.070 46.700 120.210 ;
        RECT 47.865 120.070 48.155 120.115 ;
        RECT 46.560 119.930 48.155 120.070 ;
        RECT 47.865 119.885 48.155 119.930 ;
        RECT 50.150 120.070 50.470 120.130 ;
        RECT 50.625 120.070 50.915 120.115 ;
        RECT 54.305 120.070 54.595 120.115 ;
        RECT 50.150 119.930 54.595 120.070 ;
        RECT 50.150 119.870 50.470 119.930 ;
        RECT 50.625 119.885 50.915 119.930 ;
        RECT 54.305 119.885 54.595 119.930 ;
        RECT 55.685 120.070 55.975 120.115 ;
        RECT 57.970 120.070 58.290 120.130 ;
        RECT 55.685 119.930 58.290 120.070 ;
        RECT 55.685 119.885 55.975 119.930 ;
        RECT 57.970 119.870 58.290 119.930 ;
        RECT 63.460 120.070 63.750 120.115 ;
        RECT 63.460 119.930 65.995 120.070 ;
        RECT 63.460 119.885 63.750 119.930 ;
        RECT 46.470 119.730 46.790 119.790 ;
        RECT 39.660 119.590 46.790 119.730 ;
        RECT 36.800 119.545 37.090 119.590 ;
        RECT 38.660 119.545 38.950 119.590 ;
        RECT 46.470 119.530 46.790 119.590 ;
        RECT 61.600 119.730 61.890 119.775 ;
        RECT 62.110 119.730 62.430 119.790 ;
        RECT 65.780 119.775 65.995 119.930 ;
        RECT 68.565 119.885 68.855 120.115 ;
        RECT 64.860 119.730 65.150 119.775 ;
        RECT 61.600 119.590 65.150 119.730 ;
        RECT 61.600 119.545 61.890 119.590 ;
        RECT 62.110 119.530 62.430 119.590 ;
        RECT 64.860 119.545 65.150 119.590 ;
        RECT 65.780 119.730 66.070 119.775 ;
        RECT 67.640 119.730 67.930 119.775 ;
        RECT 65.780 119.590 67.930 119.730 ;
        RECT 68.640 119.730 68.780 119.885 ;
        RECT 69.930 119.870 70.250 120.130 ;
        RECT 73.150 120.070 73.470 120.130 ;
        RECT 74.545 120.070 74.835 120.115 ;
        RECT 81.905 120.070 82.195 120.115 ;
        RECT 73.150 119.930 74.835 120.070 ;
        RECT 73.150 119.870 73.470 119.930 ;
        RECT 74.545 119.885 74.835 119.930 ;
        RECT 80.600 119.930 82.195 120.070 ;
        RECT 70.850 119.730 71.170 119.790 ;
        RECT 68.640 119.590 71.170 119.730 ;
        RECT 65.780 119.545 66.070 119.590 ;
        RECT 67.640 119.545 67.930 119.590 ;
        RECT 70.850 119.530 71.170 119.590 ;
        RECT 78.225 119.730 78.515 119.775 ;
        RECT 79.590 119.730 79.910 119.790 ;
        RECT 78.225 119.590 79.910 119.730 ;
        RECT 78.225 119.545 78.515 119.590 ;
        RECT 79.590 119.530 79.910 119.590 ;
        RECT 20.265 119.390 20.555 119.435 ;
        RECT 21.170 119.390 21.490 119.450 ;
        RECT 20.265 119.250 21.490 119.390 ;
        RECT 20.265 119.205 20.555 119.250 ;
        RECT 21.170 119.190 21.490 119.250 ;
        RECT 25.310 119.390 25.630 119.450 ;
        RECT 26.245 119.390 26.535 119.435 ;
        RECT 25.310 119.250 26.535 119.390 ;
        RECT 25.310 119.190 25.630 119.250 ;
        RECT 26.245 119.205 26.535 119.250 ;
        RECT 40.030 119.190 40.350 119.450 ;
        RECT 42.330 119.190 42.650 119.450 ;
        RECT 44.645 119.390 44.935 119.435 ;
        RECT 45.090 119.390 45.410 119.450 ;
        RECT 44.645 119.250 45.410 119.390 ;
        RECT 44.645 119.205 44.935 119.250 ;
        RECT 45.090 119.190 45.410 119.250 ;
        RECT 49.690 119.190 50.010 119.450 ;
        RECT 51.070 119.190 51.390 119.450 ;
        RECT 75.005 119.390 75.295 119.435 ;
        RECT 75.450 119.390 75.770 119.450 ;
        RECT 75.005 119.250 75.770 119.390 ;
        RECT 75.005 119.205 75.295 119.250 ;
        RECT 75.450 119.190 75.770 119.250 ;
        RECT 78.685 119.390 78.975 119.435 ;
        RECT 79.130 119.390 79.450 119.450 ;
        RECT 80.600 119.435 80.740 119.930 ;
        RECT 81.905 119.885 82.195 119.930 ;
        RECT 83.270 119.870 83.590 120.130 ;
        RECT 84.190 119.870 84.510 120.130 ;
        RECT 93.390 120.070 93.710 120.130 ;
        RECT 99.370 120.070 99.690 120.130 ;
        RECT 93.390 119.930 99.690 120.070 ;
        RECT 93.390 119.870 93.710 119.930 ;
        RECT 99.370 119.870 99.690 119.930 ;
        RECT 100.290 120.070 100.610 120.130 ;
        RECT 103.525 120.070 103.815 120.115 ;
        RECT 110.040 120.070 110.180 120.270 ;
        RECT 118.780 120.130 118.920 120.270 ;
        RECT 100.290 119.930 110.180 120.070 ;
        RECT 113.140 120.070 113.430 120.115 ;
        RECT 113.140 119.930 115.675 120.070 ;
        RECT 100.290 119.870 100.610 119.930 ;
        RECT 103.525 119.885 103.815 119.930 ;
        RECT 113.140 119.885 113.430 119.930 ;
        RECT 98.925 119.730 99.215 119.775 ;
        RECT 102.590 119.730 102.910 119.790 ;
        RECT 106.270 119.730 106.590 119.790 ;
        RECT 106.745 119.730 107.035 119.775 ;
        RECT 98.925 119.590 107.035 119.730 ;
        RECT 98.925 119.545 99.215 119.590 ;
        RECT 102.590 119.530 102.910 119.590 ;
        RECT 106.270 119.530 106.590 119.590 ;
        RECT 106.745 119.545 107.035 119.590 ;
        RECT 111.280 119.730 111.570 119.775 ;
        RECT 113.630 119.730 113.950 119.790 ;
        RECT 115.460 119.775 115.675 119.930 ;
        RECT 116.390 119.870 116.710 120.130 ;
        RECT 118.245 119.885 118.535 120.115 ;
        RECT 114.540 119.730 114.830 119.775 ;
        RECT 111.280 119.590 114.830 119.730 ;
        RECT 111.280 119.545 111.570 119.590 ;
        RECT 113.630 119.530 113.950 119.590 ;
        RECT 114.540 119.545 114.830 119.590 ;
        RECT 115.460 119.730 115.750 119.775 ;
        RECT 117.320 119.730 117.610 119.775 ;
        RECT 115.460 119.590 117.610 119.730 ;
        RECT 115.460 119.545 115.750 119.590 ;
        RECT 117.320 119.545 117.610 119.590 ;
        RECT 78.685 119.250 79.450 119.390 ;
        RECT 78.685 119.205 78.975 119.250 ;
        RECT 79.130 119.190 79.450 119.250 ;
        RECT 80.525 119.205 80.815 119.435 ;
        RECT 80.970 119.190 81.290 119.450 ;
        RECT 82.810 119.190 83.130 119.450 ;
        RECT 84.650 119.390 84.970 119.450 ;
        RECT 85.125 119.390 85.415 119.435 ;
        RECT 84.650 119.250 85.415 119.390 ;
        RECT 84.650 119.190 84.970 119.250 ;
        RECT 85.125 119.205 85.415 119.250 ;
        RECT 87.410 119.390 87.730 119.450 ;
        RECT 91.105 119.390 91.395 119.435 ;
        RECT 87.410 119.250 91.395 119.390 ;
        RECT 87.410 119.190 87.730 119.250 ;
        RECT 91.105 119.205 91.395 119.250 ;
        RECT 92.945 119.390 93.235 119.435 ;
        RECT 93.850 119.390 94.170 119.450 ;
        RECT 92.945 119.250 94.170 119.390 ;
        RECT 92.945 119.205 93.235 119.250 ;
        RECT 93.850 119.190 94.170 119.250 ;
        RECT 101.210 119.190 101.530 119.450 ;
        RECT 103.985 119.390 104.275 119.435 ;
        RECT 105.810 119.390 106.130 119.450 ;
        RECT 103.985 119.250 106.130 119.390 ;
        RECT 103.985 119.205 104.275 119.250 ;
        RECT 105.810 119.190 106.130 119.250 ;
        RECT 108.585 119.390 108.875 119.435 ;
        RECT 109.030 119.390 109.350 119.450 ;
        RECT 108.585 119.250 109.350 119.390 ;
        RECT 108.585 119.205 108.875 119.250 ;
        RECT 109.030 119.190 109.350 119.250 ;
        RECT 111.790 119.390 112.110 119.450 ;
        RECT 118.320 119.390 118.460 119.885 ;
        RECT 118.690 119.870 119.010 120.130 ;
        RECT 120.530 119.870 120.850 120.130 ;
        RECT 111.790 119.250 118.460 119.390 ;
        RECT 111.790 119.190 112.110 119.250 ;
        RECT 14.660 118.570 127.820 119.050 ;
        RECT 18.195 118.370 18.485 118.415 ;
        RECT 22.550 118.370 22.870 118.430 ;
        RECT 18.195 118.230 22.870 118.370 ;
        RECT 18.195 118.185 18.485 118.230 ;
        RECT 22.550 118.170 22.870 118.230 ;
        RECT 36.350 118.415 36.670 118.430 ;
        RECT 36.350 118.185 36.885 118.415 ;
        RECT 37.975 118.370 38.265 118.415 ;
        RECT 42.330 118.370 42.650 118.430 ;
        RECT 37.975 118.230 42.650 118.370 ;
        RECT 37.975 118.185 38.265 118.230 ;
        RECT 36.350 118.170 36.670 118.185 ;
        RECT 42.330 118.170 42.650 118.230 ;
        RECT 62.110 118.170 62.430 118.430 ;
        RECT 63.735 118.370 64.025 118.415 ;
        RECT 64.410 118.370 64.730 118.430 ;
        RECT 63.735 118.230 64.730 118.370 ;
        RECT 63.735 118.185 64.025 118.230 ;
        RECT 64.410 118.170 64.730 118.230 ;
        RECT 73.395 118.370 73.685 118.415 ;
        RECT 79.130 118.370 79.450 118.430 ;
        RECT 73.395 118.230 79.450 118.370 ;
        RECT 73.395 118.185 73.685 118.230 ;
        RECT 79.130 118.170 79.450 118.230 ;
        RECT 82.825 118.370 83.115 118.415 ;
        RECT 84.190 118.370 84.510 118.430 ;
        RECT 93.390 118.415 93.710 118.430 ;
        RECT 82.825 118.230 84.510 118.370 ;
        RECT 82.825 118.185 83.115 118.230 ;
        RECT 84.190 118.170 84.510 118.230 ;
        RECT 93.175 118.185 93.710 118.415 ;
        RECT 93.390 118.170 93.710 118.185 ;
        RECT 102.590 118.415 102.910 118.430 ;
        RECT 102.590 118.185 103.125 118.415 ;
        RECT 102.590 118.170 102.910 118.185 ;
        RECT 113.630 118.170 113.950 118.430 ;
        RECT 116.390 118.170 116.710 118.430 ;
        RECT 23.470 118.075 23.790 118.090 ;
        RECT 20.200 118.030 20.490 118.075 ;
        RECT 23.460 118.030 23.790 118.075 ;
        RECT 20.200 117.890 23.790 118.030 ;
        RECT 20.200 117.845 20.490 117.890 ;
        RECT 23.460 117.845 23.790 117.890 ;
        RECT 23.470 117.830 23.790 117.845 ;
        RECT 24.380 118.030 24.670 118.075 ;
        RECT 26.240 118.030 26.530 118.075 ;
        RECT 24.380 117.890 26.530 118.030 ;
        RECT 24.380 117.845 24.670 117.890 ;
        RECT 26.240 117.845 26.530 117.890 ;
        RECT 28.550 118.030 28.840 118.075 ;
        RECT 30.410 118.030 30.700 118.075 ;
        RECT 28.550 117.890 30.700 118.030 ;
        RECT 28.550 117.845 28.840 117.890 ;
        RECT 30.410 117.845 30.700 117.890 ;
        RECT 31.330 118.030 31.620 118.075 ;
        RECT 34.590 118.030 34.880 118.075 ;
        RECT 35.430 118.030 35.750 118.090 ;
        RECT 43.250 118.075 43.570 118.090 ;
        RECT 31.330 117.890 35.750 118.030 ;
        RECT 31.330 117.845 31.620 117.890 ;
        RECT 34.590 117.845 34.880 117.890 ;
        RECT 17.505 117.690 17.795 117.735 ;
        RECT 19.330 117.690 19.650 117.750 ;
        RECT 17.505 117.550 19.650 117.690 ;
        RECT 17.505 117.505 17.795 117.550 ;
        RECT 19.330 117.490 19.650 117.550 ;
        RECT 22.060 117.690 22.350 117.735 ;
        RECT 24.380 117.690 24.595 117.845 ;
        RECT 22.060 117.550 24.595 117.690 ;
        RECT 22.060 117.505 22.350 117.550 ;
        RECT 25.310 117.490 25.630 117.750 ;
        RECT 30.485 117.690 30.700 117.845 ;
        RECT 35.430 117.830 35.750 117.890 ;
        RECT 39.980 118.030 40.270 118.075 ;
        RECT 43.240 118.030 43.570 118.075 ;
        RECT 39.980 117.890 43.570 118.030 ;
        RECT 39.980 117.845 40.270 117.890 ;
        RECT 43.240 117.845 43.570 117.890 ;
        RECT 43.250 117.830 43.570 117.845 ;
        RECT 44.160 118.030 44.450 118.075 ;
        RECT 46.020 118.030 46.310 118.075 ;
        RECT 44.160 117.890 46.310 118.030 ;
        RECT 44.160 117.845 44.450 117.890 ;
        RECT 46.020 117.845 46.310 117.890 ;
        RECT 49.640 118.030 49.930 118.075 ;
        RECT 51.070 118.030 51.390 118.090 ;
        RECT 52.900 118.030 53.190 118.075 ;
        RECT 49.640 117.890 53.190 118.030 ;
        RECT 49.640 117.845 49.930 117.890 ;
        RECT 32.730 117.690 33.020 117.735 ;
        RECT 30.485 117.550 33.020 117.690 ;
        RECT 32.730 117.505 33.020 117.550 ;
        RECT 41.840 117.690 42.130 117.735 ;
        RECT 44.160 117.690 44.375 117.845 ;
        RECT 51.070 117.830 51.390 117.890 ;
        RECT 52.900 117.845 53.190 117.890 ;
        RECT 53.820 118.030 54.110 118.075 ;
        RECT 55.680 118.030 55.970 118.075 ;
        RECT 53.820 117.890 55.970 118.030 ;
        RECT 53.820 117.845 54.110 117.890 ;
        RECT 55.680 117.845 55.970 117.890 ;
        RECT 65.740 118.030 66.030 118.075 ;
        RECT 66.710 118.030 67.030 118.090 ;
        RECT 75.450 118.075 75.770 118.090 ;
        RECT 69.000 118.030 69.290 118.075 ;
        RECT 65.740 117.890 69.290 118.030 ;
        RECT 65.740 117.845 66.030 117.890 ;
        RECT 41.840 117.550 44.375 117.690 ;
        RECT 41.840 117.505 42.130 117.550 ;
        RECT 45.090 117.490 45.410 117.750 ;
        RECT 46.470 117.690 46.790 117.750 ;
        RECT 46.945 117.690 47.235 117.735 ;
        RECT 46.470 117.550 47.235 117.690 ;
        RECT 46.470 117.490 46.790 117.550 ;
        RECT 46.945 117.505 47.235 117.550 ;
        RECT 51.500 117.690 51.790 117.735 ;
        RECT 53.820 117.690 54.035 117.845 ;
        RECT 66.710 117.830 67.030 117.890 ;
        RECT 69.000 117.845 69.290 117.890 ;
        RECT 69.920 118.030 70.210 118.075 ;
        RECT 71.780 118.030 72.070 118.075 ;
        RECT 69.920 117.890 72.070 118.030 ;
        RECT 69.920 117.845 70.210 117.890 ;
        RECT 71.780 117.845 72.070 117.890 ;
        RECT 75.400 118.030 75.770 118.075 ;
        RECT 78.660 118.030 78.950 118.075 ;
        RECT 75.400 117.890 78.950 118.030 ;
        RECT 75.400 117.845 75.770 117.890 ;
        RECT 78.660 117.845 78.950 117.890 ;
        RECT 79.580 118.030 79.870 118.075 ;
        RECT 81.440 118.030 81.730 118.075 ;
        RECT 79.580 117.890 81.730 118.030 ;
        RECT 79.580 117.845 79.870 117.890 ;
        RECT 81.440 117.845 81.730 117.890 ;
        RECT 83.270 118.030 83.590 118.090 ;
        RECT 89.725 118.030 90.015 118.075 ;
        RECT 95.180 118.030 95.470 118.075 ;
        RECT 98.440 118.030 98.730 118.075 ;
        RECT 83.270 117.890 89.480 118.030 ;
        RECT 51.500 117.550 54.035 117.690 ;
        RECT 51.500 117.505 51.790 117.550 ;
        RECT 25.770 117.350 26.090 117.410 ;
        RECT 27.165 117.350 27.455 117.395 ;
        RECT 27.625 117.350 27.915 117.395 ;
        RECT 25.770 117.210 27.915 117.350 ;
        RECT 25.770 117.150 26.090 117.210 ;
        RECT 27.165 117.165 27.455 117.210 ;
        RECT 27.625 117.165 27.915 117.210 ;
        RECT 29.465 117.350 29.755 117.395 ;
        RECT 39.110 117.350 39.430 117.410 ;
        RECT 29.465 117.210 39.430 117.350 ;
        RECT 47.020 117.350 47.160 117.505 ;
        RECT 54.750 117.490 55.070 117.750 ;
        RECT 57.970 117.690 58.290 117.750 ;
        RECT 59.810 117.690 60.130 117.750 ;
        RECT 61.665 117.690 61.955 117.735 ;
        RECT 57.970 117.550 61.955 117.690 ;
        RECT 57.970 117.490 58.290 117.550 ;
        RECT 59.810 117.490 60.130 117.550 ;
        RECT 61.665 117.505 61.955 117.550 ;
        RECT 67.600 117.690 67.890 117.735 ;
        RECT 69.920 117.690 70.135 117.845 ;
        RECT 75.450 117.830 75.770 117.845 ;
        RECT 67.600 117.550 70.135 117.690 ;
        RECT 77.260 117.690 77.550 117.735 ;
        RECT 79.580 117.690 79.795 117.845 ;
        RECT 83.270 117.830 83.590 117.890 ;
        RECT 77.260 117.550 79.795 117.690 ;
        RECT 80.525 117.690 80.815 117.735 ;
        RECT 80.970 117.690 81.290 117.750 ;
        RECT 84.665 117.690 84.955 117.735 ;
        RECT 80.525 117.550 81.290 117.690 ;
        RECT 67.600 117.505 67.890 117.550 ;
        RECT 77.260 117.505 77.550 117.550 ;
        RECT 80.525 117.505 80.815 117.550 ;
        RECT 56.590 117.350 56.910 117.410 ;
        RECT 47.020 117.210 56.910 117.350 ;
        RECT 61.740 117.350 61.880 117.505 ;
        RECT 80.970 117.490 81.290 117.550 ;
        RECT 81.520 117.550 84.955 117.690 ;
        RECT 69.470 117.350 69.790 117.410 ;
        RECT 61.740 117.210 69.790 117.350 ;
        RECT 29.465 117.165 29.755 117.210 ;
        RECT 39.110 117.150 39.430 117.210 ;
        RECT 56.590 117.150 56.910 117.210 ;
        RECT 69.470 117.150 69.790 117.210 ;
        RECT 70.850 117.150 71.170 117.410 ;
        RECT 71.310 117.350 71.630 117.410 ;
        RECT 72.705 117.350 72.995 117.395 ;
        RECT 71.310 117.210 72.995 117.350 ;
        RECT 71.310 117.150 71.630 117.210 ;
        RECT 72.705 117.165 72.995 117.210 ;
        RECT 79.590 117.350 79.910 117.410 ;
        RECT 81.520 117.350 81.660 117.550 ;
        RECT 84.665 117.505 84.955 117.550 ;
        RECT 85.125 117.690 85.415 117.735 ;
        RECT 85.125 117.550 87.180 117.690 ;
        RECT 85.125 117.505 85.415 117.550 ;
        RECT 79.590 117.210 81.660 117.350 ;
        RECT 82.365 117.350 82.655 117.395 ;
        RECT 85.570 117.350 85.890 117.410 ;
        RECT 82.365 117.210 85.890 117.350 ;
        RECT 79.590 117.150 79.910 117.210 ;
        RECT 82.365 117.165 82.655 117.210 ;
        RECT 85.570 117.150 85.890 117.210 ;
        RECT 86.045 117.165 86.335 117.395 ;
        RECT 87.040 117.350 87.180 117.550 ;
        RECT 87.410 117.490 87.730 117.750 ;
        RECT 89.340 117.735 89.480 117.890 ;
        RECT 89.725 117.890 98.730 118.030 ;
        RECT 89.725 117.845 90.015 117.890 ;
        RECT 95.180 117.845 95.470 117.890 ;
        RECT 98.440 117.845 98.730 117.890 ;
        RECT 99.360 118.030 99.650 118.075 ;
        RECT 101.220 118.030 101.510 118.075 ;
        RECT 99.360 117.890 101.510 118.030 ;
        RECT 99.360 117.845 99.650 117.890 ;
        RECT 101.220 117.845 101.510 117.890 ;
        RECT 104.840 118.030 105.130 118.075 ;
        RECT 105.810 118.030 106.130 118.090 ;
        RECT 108.100 118.030 108.390 118.075 ;
        RECT 104.840 117.890 108.390 118.030 ;
        RECT 104.840 117.845 105.130 117.890 ;
        RECT 89.265 117.690 89.555 117.735 ;
        RECT 90.645 117.690 90.935 117.735 ;
        RECT 89.265 117.550 90.935 117.690 ;
        RECT 89.265 117.505 89.555 117.550 ;
        RECT 90.645 117.505 90.935 117.550 ;
        RECT 97.040 117.690 97.330 117.735 ;
        RECT 99.360 117.690 99.575 117.845 ;
        RECT 105.810 117.830 106.130 117.890 ;
        RECT 108.100 117.845 108.390 117.890 ;
        RECT 109.020 118.030 109.310 118.075 ;
        RECT 110.880 118.030 111.170 118.075 ;
        RECT 118.230 118.030 118.550 118.090 ;
        RECT 109.020 117.890 111.170 118.030 ;
        RECT 109.020 117.845 109.310 117.890 ;
        RECT 110.880 117.845 111.170 117.890 ;
        RECT 114.180 117.890 118.550 118.030 ;
        RECT 97.040 117.550 99.575 117.690 ;
        RECT 106.700 117.690 106.990 117.735 ;
        RECT 109.020 117.690 109.235 117.845 ;
        RECT 106.700 117.550 109.235 117.690 ;
        RECT 97.040 117.505 97.330 117.550 ;
        RECT 106.700 117.505 106.990 117.550 ;
        RECT 109.950 117.490 110.270 117.750 ;
        RECT 111.790 117.490 112.110 117.750 ;
        RECT 114.180 117.735 114.320 117.890 ;
        RECT 118.230 117.830 118.550 117.890 ;
        RECT 114.105 117.505 114.395 117.735 ;
        RECT 115.470 117.490 115.790 117.750 ;
        RECT 93.850 117.350 94.170 117.410 ;
        RECT 87.040 117.210 94.170 117.350 ;
        RECT 22.060 117.010 22.350 117.055 ;
        RECT 24.840 117.010 25.130 117.055 ;
        RECT 26.700 117.010 26.990 117.055 ;
        RECT 22.060 116.870 26.990 117.010 ;
        RECT 22.060 116.825 22.350 116.870 ;
        RECT 24.840 116.825 25.130 116.870 ;
        RECT 26.700 116.825 26.990 116.870 ;
        RECT 28.090 117.010 28.380 117.055 ;
        RECT 29.950 117.010 30.240 117.055 ;
        RECT 32.730 117.010 33.020 117.055 ;
        RECT 28.090 116.870 33.020 117.010 ;
        RECT 28.090 116.825 28.380 116.870 ;
        RECT 29.950 116.825 30.240 116.870 ;
        RECT 32.730 116.825 33.020 116.870 ;
        RECT 41.840 117.010 42.130 117.055 ;
        RECT 44.620 117.010 44.910 117.055 ;
        RECT 46.480 117.010 46.770 117.055 ;
        RECT 41.840 116.870 46.770 117.010 ;
        RECT 41.840 116.825 42.130 116.870 ;
        RECT 44.620 116.825 44.910 116.870 ;
        RECT 46.480 116.825 46.770 116.870 ;
        RECT 51.500 117.010 51.790 117.055 ;
        RECT 54.280 117.010 54.570 117.055 ;
        RECT 56.140 117.010 56.430 117.055 ;
        RECT 51.500 116.870 56.430 117.010 ;
        RECT 51.500 116.825 51.790 116.870 ;
        RECT 54.280 116.825 54.570 116.870 ;
        RECT 56.140 116.825 56.430 116.870 ;
        RECT 67.600 117.010 67.890 117.055 ;
        RECT 70.380 117.010 70.670 117.055 ;
        RECT 72.240 117.010 72.530 117.055 ;
        RECT 67.600 116.870 72.530 117.010 ;
        RECT 67.600 116.825 67.890 116.870 ;
        RECT 70.380 116.825 70.670 116.870 ;
        RECT 72.240 116.825 72.530 116.870 ;
        RECT 77.260 117.010 77.550 117.055 ;
        RECT 80.040 117.010 80.330 117.055 ;
        RECT 81.900 117.010 82.190 117.055 ;
        RECT 77.260 116.870 82.190 117.010 ;
        RECT 77.260 116.825 77.550 116.870 ;
        RECT 80.040 116.825 80.330 116.870 ;
        RECT 81.900 116.825 82.190 116.870 ;
        RECT 83.730 117.010 84.050 117.070 ;
        RECT 86.120 117.010 86.260 117.165 ;
        RECT 93.850 117.150 94.170 117.210 ;
        RECT 100.290 117.150 100.610 117.410 ;
        RECT 102.145 117.350 102.435 117.395 ;
        RECT 111.880 117.350 112.020 117.490 ;
        RECT 102.145 117.210 112.020 117.350 ;
        RECT 102.145 117.165 102.435 117.210 ;
        RECT 83.730 116.870 86.260 117.010 ;
        RECT 97.040 117.010 97.330 117.055 ;
        RECT 99.820 117.010 100.110 117.055 ;
        RECT 101.680 117.010 101.970 117.055 ;
        RECT 97.040 116.870 101.970 117.010 ;
        RECT 83.730 116.810 84.050 116.870 ;
        RECT 97.040 116.825 97.330 116.870 ;
        RECT 99.820 116.825 100.110 116.870 ;
        RECT 101.680 116.825 101.970 116.870 ;
        RECT 106.700 117.010 106.990 117.055 ;
        RECT 109.480 117.010 109.770 117.055 ;
        RECT 111.340 117.010 111.630 117.055 ;
        RECT 106.700 116.870 111.630 117.010 ;
        RECT 106.700 116.825 106.990 116.870 ;
        RECT 109.480 116.825 109.770 116.870 ;
        RECT 111.340 116.825 111.630 116.870 ;
        RECT 17.045 116.670 17.335 116.715 ;
        RECT 28.530 116.670 28.850 116.730 ;
        RECT 17.045 116.530 28.850 116.670 ;
        RECT 17.045 116.485 17.335 116.530 ;
        RECT 28.530 116.470 28.850 116.530 ;
        RECT 46.010 116.670 46.330 116.730 ;
        RECT 47.635 116.670 47.925 116.715 ;
        RECT 46.010 116.530 47.925 116.670 ;
        RECT 46.010 116.470 46.330 116.530 ;
        RECT 47.635 116.485 47.925 116.530 ;
        RECT 88.330 116.470 88.650 116.730 ;
        RECT 91.090 116.470 91.410 116.730 ;
        RECT 14.660 115.850 127.820 116.330 ;
        RECT 23.025 115.650 23.315 115.695 ;
        RECT 23.470 115.650 23.790 115.710 ;
        RECT 23.025 115.510 23.790 115.650 ;
        RECT 23.025 115.465 23.315 115.510 ;
        RECT 23.470 115.450 23.790 115.510 ;
        RECT 30.830 115.650 31.150 115.710 ;
        RECT 33.835 115.650 34.125 115.695 ;
        RECT 30.830 115.510 34.125 115.650 ;
        RECT 30.830 115.450 31.150 115.510 ;
        RECT 33.835 115.465 34.125 115.510 ;
        RECT 35.430 115.450 35.750 115.710 ;
        RECT 37.730 115.450 38.050 115.710 ;
        RECT 39.110 115.450 39.430 115.710 ;
        RECT 43.250 115.650 43.570 115.710 ;
        RECT 44.645 115.650 44.935 115.695 ;
        RECT 43.250 115.510 44.935 115.650 ;
        RECT 43.250 115.450 43.570 115.510 ;
        RECT 44.645 115.465 44.935 115.510 ;
        RECT 45.550 115.450 45.870 115.710 ;
        RECT 53.385 115.650 53.675 115.695 ;
        RECT 54.750 115.650 55.070 115.710 ;
        RECT 53.385 115.510 55.070 115.650 ;
        RECT 53.385 115.465 53.675 115.510 ;
        RECT 54.750 115.450 55.070 115.510 ;
        RECT 66.710 115.450 67.030 115.710 ;
        RECT 69.025 115.650 69.315 115.695 ;
        RECT 70.850 115.650 71.170 115.710 ;
        RECT 69.025 115.510 71.170 115.650 ;
        RECT 69.025 115.465 69.315 115.510 ;
        RECT 70.850 115.450 71.170 115.510 ;
        RECT 71.310 115.650 71.630 115.710 ;
        RECT 73.610 115.650 73.930 115.710 ;
        RECT 71.310 115.510 73.930 115.650 ;
        RECT 71.310 115.450 71.630 115.510 ;
        RECT 73.610 115.450 73.930 115.510 ;
        RECT 77.535 115.650 77.825 115.695 ;
        RECT 79.590 115.650 79.910 115.710 ;
        RECT 77.535 115.510 79.910 115.650 ;
        RECT 77.535 115.465 77.825 115.510 ;
        RECT 79.590 115.450 79.910 115.510 ;
        RECT 93.850 115.650 94.170 115.710 ;
        RECT 96.395 115.650 96.685 115.695 ;
        RECT 93.850 115.510 96.685 115.650 ;
        RECT 93.850 115.450 94.170 115.510 ;
        RECT 96.395 115.465 96.685 115.510 ;
        RECT 100.290 115.450 100.610 115.710 ;
        RECT 109.045 115.650 109.335 115.695 ;
        RECT 109.950 115.650 110.270 115.710 ;
        RECT 109.045 115.510 110.270 115.650 ;
        RECT 109.045 115.465 109.335 115.510 ;
        RECT 109.950 115.450 110.270 115.510 ;
        RECT 115.025 115.650 115.315 115.695 ;
        RECT 115.470 115.650 115.790 115.710 ;
        RECT 115.025 115.510 115.790 115.650 ;
        RECT 115.025 115.465 115.315 115.510 ;
        RECT 115.470 115.450 115.790 115.510 ;
        RECT 22.105 115.125 22.395 115.355 ;
        RECT 25.330 115.310 25.620 115.355 ;
        RECT 27.190 115.310 27.480 115.355 ;
        RECT 29.970 115.310 30.260 115.355 ;
        RECT 25.330 115.170 30.260 115.310 ;
        RECT 25.330 115.125 25.620 115.170 ;
        RECT 27.190 115.125 27.480 115.170 ;
        RECT 29.970 115.125 30.260 115.170 ;
        RECT 43.710 115.310 44.030 115.370 ;
        RECT 81.400 115.310 81.690 115.355 ;
        RECT 84.180 115.310 84.470 115.355 ;
        RECT 86.040 115.310 86.330 115.355 ;
        RECT 43.710 115.170 48.540 115.310 ;
        RECT 19.790 114.970 20.110 115.030 ;
        RECT 22.180 114.970 22.320 115.125 ;
        RECT 43.710 115.110 44.030 115.170 ;
        RECT 24.865 114.970 25.155 115.015 ;
        RECT 25.770 114.970 26.090 115.030 ;
        RECT 46.010 114.970 46.330 115.030 ;
        RECT 48.400 115.015 48.540 115.170 ;
        RECT 81.400 115.170 86.330 115.310 ;
        RECT 81.400 115.125 81.690 115.170 ;
        RECT 84.180 115.125 84.470 115.170 ;
        RECT 86.040 115.125 86.330 115.170 ;
        RECT 87.890 115.310 88.180 115.355 ;
        RECT 89.750 115.310 90.040 115.355 ;
        RECT 92.530 115.310 92.820 115.355 ;
        RECT 113.170 115.310 113.490 115.370 ;
        RECT 87.890 115.170 92.820 115.310 ;
        RECT 87.890 115.125 88.180 115.170 ;
        RECT 89.750 115.125 90.040 115.170 ;
        RECT 92.530 115.125 92.820 115.170 ;
        RECT 112.340 115.170 113.490 115.310 ;
        RECT 47.865 114.970 48.155 115.015 ;
        RECT 19.790 114.830 21.860 114.970 ;
        RECT 22.180 114.830 24.620 114.970 ;
        RECT 19.790 114.770 20.110 114.830 ;
        RECT 21.170 114.430 21.490 114.690 ;
        RECT 21.720 114.630 21.860 114.830 ;
        RECT 23.485 114.630 23.775 114.675 ;
        RECT 24.480 114.630 24.620 114.830 ;
        RECT 24.865 114.830 26.090 114.970 ;
        RECT 24.865 114.785 25.155 114.830 ;
        RECT 25.770 114.770 26.090 114.830 ;
        RECT 35.980 114.830 45.320 114.970 ;
        RECT 35.980 114.690 36.120 114.830 ;
        RECT 26.705 114.630 26.995 114.675 ;
        RECT 29.970 114.630 30.260 114.675 ;
        RECT 21.720 114.490 24.160 114.630 ;
        RECT 24.480 114.490 26.995 114.630 ;
        RECT 23.485 114.445 23.775 114.490 ;
        RECT 24.020 113.950 24.160 114.490 ;
        RECT 26.705 114.445 26.995 114.490 ;
        RECT 27.725 114.490 30.260 114.630 ;
        RECT 27.725 114.335 27.940 114.490 ;
        RECT 29.970 114.445 30.260 114.490 ;
        RECT 35.890 114.430 36.210 114.690 ;
        RECT 36.810 114.430 37.130 114.690 ;
        RECT 40.030 114.430 40.350 114.690 ;
        RECT 45.180 114.675 45.320 114.830 ;
        RECT 46.010 114.830 48.155 114.970 ;
        RECT 46.010 114.770 46.330 114.830 ;
        RECT 47.865 114.785 48.155 114.830 ;
        RECT 48.325 114.785 48.615 115.015 ;
        RECT 50.150 114.970 50.470 115.030 ;
        RECT 69.470 114.970 69.790 115.030 ;
        RECT 49.320 114.830 50.470 114.970 ;
        RECT 45.105 114.630 45.395 114.675 ;
        RECT 49.320 114.630 49.460 114.830 ;
        RECT 50.150 114.770 50.470 114.830 ;
        RECT 66.340 114.830 69.790 114.970 ;
        RECT 45.105 114.490 49.460 114.630 ;
        RECT 49.690 114.630 50.010 114.690 ;
        RECT 66.340 114.675 66.480 114.830 ;
        RECT 69.470 114.770 69.790 114.830 ;
        RECT 84.650 114.770 84.970 115.030 ;
        RECT 85.570 114.970 85.890 115.030 ;
        RECT 86.490 114.970 86.810 115.030 ;
        RECT 87.425 114.970 87.715 115.015 ;
        RECT 85.570 114.830 87.715 114.970 ;
        RECT 85.570 114.770 85.890 114.830 ;
        RECT 86.490 114.770 86.810 114.830 ;
        RECT 87.425 114.785 87.715 114.830 ;
        RECT 88.330 114.970 88.650 115.030 ;
        RECT 112.340 115.015 112.480 115.170 ;
        RECT 113.170 115.110 113.490 115.170 ;
        RECT 89.265 114.970 89.555 115.015 ;
        RECT 88.330 114.830 89.555 114.970 ;
        RECT 88.330 114.770 88.650 114.830 ;
        RECT 89.265 114.785 89.555 114.830 ;
        RECT 112.265 114.785 112.555 115.015 ;
        RECT 112.710 114.770 113.030 115.030 ;
        RECT 52.465 114.630 52.755 114.675 ;
        RECT 49.690 114.490 52.755 114.630 ;
        RECT 45.105 114.445 45.395 114.490 ;
        RECT 49.690 114.430 50.010 114.490 ;
        RECT 52.465 114.445 52.755 114.490 ;
        RECT 66.265 114.445 66.555 114.675 ;
        RECT 68.090 114.430 68.410 114.690 ;
        RECT 81.400 114.630 81.690 114.675 ;
        RECT 92.530 114.630 92.820 114.675 ;
        RECT 81.400 114.490 83.935 114.630 ;
        RECT 81.400 114.445 81.690 114.490 ;
        RECT 25.790 114.290 26.080 114.335 ;
        RECT 27.650 114.290 27.940 114.335 ;
        RECT 25.790 114.150 27.940 114.290 ;
        RECT 25.790 114.105 26.080 114.150 ;
        RECT 27.650 114.105 27.940 114.150 ;
        RECT 28.530 114.335 28.850 114.350 ;
        RECT 28.530 114.290 28.860 114.335 ;
        RECT 31.830 114.290 32.120 114.335 ;
        RECT 28.530 114.150 32.120 114.290 ;
        RECT 28.530 114.105 28.860 114.150 ;
        RECT 31.830 114.105 32.120 114.150 ;
        RECT 42.330 114.290 42.650 114.350 ;
        RECT 82.810 114.335 83.130 114.350 ;
        RECT 47.405 114.290 47.695 114.335 ;
        RECT 42.330 114.150 47.695 114.290 ;
        RECT 28.530 114.090 28.850 114.105 ;
        RECT 42.330 114.090 42.650 114.150 ;
        RECT 47.405 114.105 47.695 114.150 ;
        RECT 79.540 114.290 79.830 114.335 ;
        RECT 82.800 114.290 83.130 114.335 ;
        RECT 79.540 114.150 83.130 114.290 ;
        RECT 79.540 114.105 79.830 114.150 ;
        RECT 82.800 114.105 83.130 114.150 ;
        RECT 83.720 114.335 83.935 114.490 ;
        RECT 90.285 114.490 92.820 114.630 ;
        RECT 90.285 114.335 90.500 114.490 ;
        RECT 92.530 114.445 92.820 114.490 ;
        RECT 101.210 114.430 101.530 114.690 ;
        RECT 108.125 114.630 108.415 114.675 ;
        RECT 109.030 114.630 109.350 114.690 ;
        RECT 108.125 114.490 109.350 114.630 ;
        RECT 108.125 114.445 108.415 114.490 ;
        RECT 109.030 114.430 109.350 114.490 ;
        RECT 109.490 114.630 109.810 114.690 ;
        RECT 113.185 114.630 113.475 114.675 ;
        RECT 109.490 114.490 113.475 114.630 ;
        RECT 109.490 114.430 109.810 114.490 ;
        RECT 113.185 114.445 113.475 114.490 ;
        RECT 83.720 114.290 84.010 114.335 ;
        RECT 85.580 114.290 85.870 114.335 ;
        RECT 83.720 114.150 85.870 114.290 ;
        RECT 83.720 114.105 84.010 114.150 ;
        RECT 85.580 114.105 85.870 114.150 ;
        RECT 88.350 114.290 88.640 114.335 ;
        RECT 90.210 114.290 90.500 114.335 ;
        RECT 88.350 114.150 90.500 114.290 ;
        RECT 88.350 114.105 88.640 114.150 ;
        RECT 90.210 114.105 90.500 114.150 ;
        RECT 91.090 114.335 91.410 114.350 ;
        RECT 91.090 114.290 91.420 114.335 ;
        RECT 94.390 114.290 94.680 114.335 ;
        RECT 91.090 114.150 94.680 114.290 ;
        RECT 91.090 114.105 91.420 114.150 ;
        RECT 94.390 114.105 94.680 114.150 ;
        RECT 82.810 114.090 83.130 114.105 ;
        RECT 91.090 114.090 91.410 114.105 ;
        RECT 35.890 113.950 36.210 114.010 ;
        RECT 24.020 113.810 36.210 113.950 ;
        RECT 35.890 113.750 36.210 113.810 ;
        RECT 101.670 113.950 101.990 114.010 ;
        RECT 121.910 113.950 122.230 114.010 ;
        RECT 101.670 113.810 122.230 113.950 ;
        RECT 101.670 113.750 101.990 113.810 ;
        RECT 121.910 113.750 122.230 113.810 ;
        RECT 14.660 113.130 127.820 113.610 ;
        RECT 34.525 112.930 34.815 112.975 ;
        RECT 34.970 112.930 35.290 112.990 ;
        RECT 34.525 112.790 35.290 112.930 ;
        RECT 34.525 112.745 34.815 112.790 ;
        RECT 34.970 112.730 35.290 112.790 ;
        RECT 103.065 112.930 103.355 112.975 ;
        RECT 111.790 112.930 112.110 112.990 ;
        RECT 103.065 112.790 112.110 112.930 ;
        RECT 103.065 112.745 103.355 112.790 ;
        RECT 18.985 112.590 19.275 112.635 ;
        RECT 21.170 112.590 21.490 112.650 ;
        RECT 22.225 112.590 22.875 112.635 ;
        RECT 18.985 112.450 22.875 112.590 ;
        RECT 18.985 112.405 19.575 112.450 ;
        RECT 19.285 112.090 19.575 112.405 ;
        RECT 21.170 112.390 21.490 112.450 ;
        RECT 22.225 112.405 22.875 112.450 ;
        RECT 46.945 112.590 47.235 112.635 ;
        RECT 49.230 112.590 49.550 112.650 ;
        RECT 46.945 112.450 49.550 112.590 ;
        RECT 46.945 112.405 47.235 112.450 ;
        RECT 49.230 112.390 49.550 112.450 ;
        RECT 92.930 112.390 93.250 112.650 ;
        RECT 101.685 112.590 101.975 112.635 ;
        RECT 103.140 112.590 103.280 112.745 ;
        RECT 111.790 112.730 112.110 112.790 ;
        RECT 117.310 112.930 117.630 112.990 ;
        RECT 121.005 112.930 121.295 112.975 ;
        RECT 117.310 112.790 121.295 112.930 ;
        RECT 117.310 112.730 117.630 112.790 ;
        RECT 121.005 112.745 121.295 112.790 ;
        RECT 122.385 112.745 122.675 112.975 ;
        RECT 101.685 112.450 103.280 112.590 ;
        RECT 119.150 112.590 119.470 112.650 ;
        RECT 122.460 112.590 122.600 112.745 ;
        RECT 119.150 112.450 122.600 112.590 ;
        RECT 101.685 112.405 101.975 112.450 ;
        RECT 119.150 112.390 119.470 112.450 ;
        RECT 20.365 112.250 20.655 112.295 ;
        RECT 23.945 112.250 24.235 112.295 ;
        RECT 25.780 112.250 26.070 112.295 ;
        RECT 20.365 112.110 26.070 112.250 ;
        RECT 20.365 112.065 20.655 112.110 ;
        RECT 23.945 112.065 24.235 112.110 ;
        RECT 25.780 112.065 26.070 112.110 ;
        RECT 26.230 112.050 26.550 112.310 ;
        RECT 34.985 112.250 35.275 112.295 ;
        RECT 35.890 112.250 36.210 112.310 ;
        RECT 34.985 112.110 36.210 112.250 ;
        RECT 34.985 112.065 35.275 112.110 ;
        RECT 35.890 112.050 36.210 112.110 ;
        RECT 78.210 112.250 78.530 112.310 ;
        RECT 81.430 112.250 81.750 112.310 ;
        RECT 78.210 112.110 81.750 112.250 ;
        RECT 78.210 112.050 78.530 112.110 ;
        RECT 81.430 112.050 81.750 112.110 ;
        RECT 119.610 112.050 119.930 112.310 ;
        RECT 121.910 112.050 122.230 112.310 ;
        RECT 123.305 112.065 123.595 112.295 ;
        RECT 14.270 111.910 14.590 111.970 ;
        RECT 16.125 111.910 16.415 111.955 ;
        RECT 14.270 111.770 16.415 111.910 ;
        RECT 14.270 111.710 14.590 111.770 ;
        RECT 16.125 111.725 16.415 111.770 ;
        RECT 20.365 111.570 20.655 111.615 ;
        RECT 23.485 111.570 23.775 111.615 ;
        RECT 25.375 111.570 25.665 111.615 ;
        RECT 20.365 111.430 25.665 111.570 ;
        RECT 26.320 111.570 26.460 112.050 ;
        RECT 50.610 111.910 50.930 111.970 ;
        RECT 43.340 111.770 50.930 111.910 ;
        RECT 36.810 111.570 37.130 111.630 ;
        RECT 40.505 111.570 40.795 111.615 ;
        RECT 43.340 111.570 43.480 111.770 ;
        RECT 50.610 111.710 50.930 111.770 ;
        RECT 80.985 111.910 81.275 111.955 ;
        RECT 81.890 111.910 82.210 111.970 ;
        RECT 80.985 111.770 82.210 111.910 ;
        RECT 80.985 111.725 81.275 111.770 ;
        RECT 81.890 111.710 82.210 111.770 ;
        RECT 104.430 111.910 104.750 111.970 ;
        RECT 104.430 111.770 119.840 111.910 ;
        RECT 104.430 111.710 104.750 111.770 ;
        RECT 26.320 111.430 43.480 111.570 ;
        RECT 119.700 111.570 119.840 111.770 ;
        RECT 120.070 111.710 120.390 111.970 ;
        RECT 123.380 111.910 123.520 112.065 ;
        RECT 120.620 111.770 123.520 111.910 ;
        RECT 120.620 111.570 120.760 111.770 ;
        RECT 119.700 111.430 120.760 111.570 ;
        RECT 20.365 111.385 20.655 111.430 ;
        RECT 23.485 111.385 23.775 111.430 ;
        RECT 25.375 111.385 25.665 111.430 ;
        RECT 36.810 111.370 37.130 111.430 ;
        RECT 40.505 111.385 40.795 111.430 ;
        RECT 24.960 111.230 25.250 111.275 ;
        RECT 27.610 111.230 27.930 111.290 ;
        RECT 24.960 111.090 27.930 111.230 ;
        RECT 24.960 111.045 25.250 111.090 ;
        RECT 27.610 111.030 27.930 111.090 ;
        RECT 14.660 110.410 127.820 110.890 ;
        RECT 21.170 110.010 21.490 110.270 ;
        RECT 27.610 110.010 27.930 110.270 ;
        RECT 74.070 110.210 74.390 110.270 ;
        RECT 78.225 110.210 78.515 110.255 ;
        RECT 74.070 110.070 78.515 110.210 ;
        RECT 74.070 110.010 74.390 110.070 ;
        RECT 78.225 110.025 78.515 110.070 ;
        RECT 107.205 109.870 107.495 109.915 ;
        RECT 110.870 109.870 111.190 109.930 ;
        RECT 107.205 109.730 111.190 109.870 ;
        RECT 107.205 109.685 107.495 109.730 ;
        RECT 110.870 109.670 111.190 109.730 ;
        RECT 111.790 109.670 112.110 109.930 ;
        RECT 116.815 109.870 117.105 109.915 ;
        RECT 118.705 109.870 118.995 109.915 ;
        RECT 121.825 109.870 122.115 109.915 ;
        RECT 116.815 109.730 122.115 109.870 ;
        RECT 116.815 109.685 117.105 109.730 ;
        RECT 118.705 109.685 118.995 109.730 ;
        RECT 121.825 109.685 122.115 109.730 ;
        RECT 31.290 109.530 31.610 109.590 ;
        RECT 81.430 109.530 81.750 109.590 ;
        RECT 111.880 109.530 112.020 109.670 ;
        RECT 115.945 109.530 116.235 109.575 ;
        RECT 31.290 109.390 33.360 109.530 ;
        RECT 31.290 109.330 31.610 109.390 ;
        RECT 21.645 109.190 21.935 109.235 ;
        RECT 23.945 109.190 24.235 109.235 ;
        RECT 21.645 109.050 24.235 109.190 ;
        RECT 21.645 109.005 21.935 109.050 ;
        RECT 23.945 109.005 24.235 109.050 ;
        RECT 28.545 109.190 28.835 109.235 ;
        RECT 29.450 109.190 29.770 109.250 ;
        RECT 33.220 109.235 33.360 109.390 ;
        RECT 59.900 109.390 79.820 109.530 ;
        RECT 59.900 109.250 60.040 109.390 ;
        RECT 28.545 109.050 29.770 109.190 ;
        RECT 28.545 109.005 28.835 109.050 ;
        RECT 24.020 108.850 24.160 109.005 ;
        RECT 29.450 108.990 29.770 109.050 ;
        RECT 31.765 109.005 32.055 109.235 ;
        RECT 33.145 109.005 33.435 109.235 ;
        RECT 34.510 109.190 34.830 109.250 ;
        RECT 35.445 109.190 35.735 109.235 ;
        RECT 34.510 109.050 35.735 109.190 ;
        RECT 27.610 108.850 27.930 108.910 ;
        RECT 31.840 108.850 31.980 109.005 ;
        RECT 34.510 108.990 34.830 109.050 ;
        RECT 35.445 109.005 35.735 109.050 ;
        RECT 51.085 109.190 51.375 109.235 ;
        RECT 51.990 109.190 52.310 109.250 ;
        RECT 51.085 109.050 52.310 109.190 ;
        RECT 51.085 109.005 51.375 109.050 ;
        RECT 51.990 108.990 52.310 109.050 ;
        RECT 57.050 108.990 57.370 109.250 ;
        RECT 59.810 108.990 60.130 109.250 ;
        RECT 60.270 109.190 60.590 109.250 ;
        RECT 61.205 109.190 61.495 109.235 ;
        RECT 64.885 109.190 65.175 109.235 ;
        RECT 60.270 109.050 65.175 109.190 ;
        RECT 60.270 108.990 60.590 109.050 ;
        RECT 61.205 109.005 61.495 109.050 ;
        RECT 64.885 109.005 65.175 109.050 ;
        RECT 68.565 109.190 68.855 109.235 ;
        RECT 69.010 109.190 69.330 109.250 ;
        RECT 68.565 109.050 69.330 109.190 ;
        RECT 68.565 109.005 68.855 109.050 ;
        RECT 69.010 108.990 69.330 109.050 ;
        RECT 77.305 109.190 77.595 109.235 ;
        RECT 78.210 109.190 78.530 109.250 ;
        RECT 77.305 109.050 78.530 109.190 ;
        RECT 77.305 109.005 77.595 109.050 ;
        RECT 78.210 108.990 78.530 109.050 ;
        RECT 78.685 109.190 78.975 109.235 ;
        RECT 79.130 109.190 79.450 109.250 ;
        RECT 78.685 109.050 79.450 109.190 ;
        RECT 79.680 109.190 79.820 109.390 ;
        RECT 81.430 109.390 87.640 109.530 ;
        RECT 111.880 109.390 116.235 109.530 ;
        RECT 81.430 109.330 81.750 109.390 ;
        RECT 87.500 109.235 87.640 109.390 ;
        RECT 115.945 109.345 116.235 109.390 ;
        RECT 117.325 109.530 117.615 109.575 ;
        RECT 119.150 109.530 119.470 109.590 ;
        RECT 117.325 109.390 119.470 109.530 ;
        RECT 117.325 109.345 117.615 109.390 ;
        RECT 119.150 109.330 119.470 109.390 ;
        RECT 80.065 109.190 80.355 109.235 ;
        RECT 79.680 109.050 80.355 109.190 ;
        RECT 78.685 109.005 78.975 109.050 ;
        RECT 79.130 108.990 79.450 109.050 ;
        RECT 80.065 109.005 80.355 109.050 ;
        RECT 82.825 109.005 83.115 109.235 ;
        RECT 87.425 109.190 87.715 109.235 ;
        RECT 92.485 109.190 92.775 109.235 ;
        RECT 87.425 109.050 92.775 109.190 ;
        RECT 87.425 109.005 87.715 109.050 ;
        RECT 92.485 109.005 92.775 109.050 ;
        RECT 93.865 109.190 94.155 109.235 ;
        RECT 94.770 109.190 95.090 109.250 ;
        RECT 93.865 109.050 95.090 109.190 ;
        RECT 93.865 109.005 94.155 109.050 ;
        RECT 40.950 108.850 41.270 108.910 ;
        RECT 24.020 108.710 41.270 108.850 ;
        RECT 27.610 108.650 27.930 108.710 ;
        RECT 40.950 108.650 41.270 108.710 ;
        RECT 75.910 108.850 76.230 108.910 ;
        RECT 82.900 108.850 83.040 109.005 ;
        RECT 75.910 108.710 83.040 108.850 ;
        RECT 92.560 108.850 92.700 109.005 ;
        RECT 94.770 108.990 95.090 109.050 ;
        RECT 99.830 109.190 100.150 109.250 ;
        RECT 101.225 109.190 101.515 109.235 ;
        RECT 99.830 109.050 101.515 109.190 ;
        RECT 99.830 108.990 100.150 109.050 ;
        RECT 101.225 109.005 101.515 109.050 ;
        RECT 103.510 109.190 103.830 109.250 ;
        RECT 106.285 109.190 106.575 109.235 ;
        RECT 103.510 109.050 106.575 109.190 ;
        RECT 103.510 108.990 103.830 109.050 ;
        RECT 106.285 109.005 106.575 109.050 ;
        RECT 109.965 109.005 110.255 109.235 ;
        RECT 102.590 108.850 102.910 108.910 ;
        RECT 110.040 108.850 110.180 109.005 ;
        RECT 110.410 108.990 110.730 109.250 ;
        RECT 111.330 109.190 111.650 109.250 ;
        RECT 111.805 109.190 112.095 109.235 ;
        RECT 111.330 109.050 112.095 109.190 ;
        RECT 111.330 108.990 111.650 109.050 ;
        RECT 111.805 109.005 112.095 109.050 ;
        RECT 114.565 109.005 114.855 109.235 ;
        RECT 116.410 109.190 116.700 109.235 ;
        RECT 118.245 109.190 118.535 109.235 ;
        RECT 121.825 109.190 122.115 109.235 ;
        RECT 116.410 109.050 122.115 109.190 ;
        RECT 116.410 109.005 116.700 109.050 ;
        RECT 118.245 109.005 118.535 109.050 ;
        RECT 121.825 109.005 122.115 109.050 ;
        RECT 114.640 108.850 114.780 109.005 ;
        RECT 120.070 108.895 120.390 108.910 ;
        RECT 119.605 108.850 120.390 108.895 ;
        RECT 122.905 108.895 123.195 109.210 ;
        RECT 122.905 108.850 123.495 108.895 ;
        RECT 92.560 108.710 119.380 108.850 ;
        RECT 75.910 108.650 76.230 108.710 ;
        RECT 102.590 108.650 102.910 108.710 ;
        RECT 119.240 108.570 119.380 108.710 ;
        RECT 119.605 108.710 123.495 108.850 ;
        RECT 119.605 108.665 120.390 108.710 ;
        RECT 123.205 108.665 123.495 108.710 ;
        RECT 126.065 108.850 126.355 108.895 ;
        RECT 127.890 108.850 128.210 108.910 ;
        RECT 126.065 108.710 128.210 108.850 ;
        RECT 126.065 108.665 126.355 108.710 ;
        RECT 120.070 108.650 120.390 108.665 ;
        RECT 127.890 108.650 128.210 108.710 ;
        RECT 23.470 108.310 23.790 108.570 ;
        RECT 31.305 108.510 31.595 108.555 ;
        RECT 31.750 108.510 32.070 108.570 ;
        RECT 31.305 108.370 32.070 108.510 ;
        RECT 31.305 108.325 31.595 108.370 ;
        RECT 31.750 108.310 32.070 108.370 ;
        RECT 32.210 108.310 32.530 108.570 ;
        RECT 34.050 108.510 34.370 108.570 ;
        RECT 34.525 108.510 34.815 108.555 ;
        RECT 34.050 108.370 34.815 108.510 ;
        RECT 34.050 108.310 34.370 108.370 ;
        RECT 34.525 108.325 34.815 108.370 ;
        RECT 52.005 108.510 52.295 108.555 ;
        RECT 55.670 108.510 55.990 108.570 ;
        RECT 52.005 108.370 55.990 108.510 ;
        RECT 52.005 108.325 52.295 108.370 ;
        RECT 55.670 108.310 55.990 108.370 ;
        RECT 57.970 108.310 58.290 108.570 ;
        RECT 65.330 108.310 65.650 108.570 ;
        RECT 69.485 108.510 69.775 108.555 ;
        RECT 72.230 108.510 72.550 108.570 ;
        RECT 69.485 108.370 72.550 108.510 ;
        RECT 69.485 108.325 69.775 108.370 ;
        RECT 72.230 108.310 72.550 108.370 ;
        RECT 76.845 108.510 77.135 108.555 ;
        RECT 79.590 108.510 79.910 108.570 ;
        RECT 76.845 108.370 79.910 108.510 ;
        RECT 76.845 108.325 77.135 108.370 ;
        RECT 79.590 108.310 79.910 108.370 ;
        RECT 83.730 108.310 84.050 108.570 ;
        RECT 87.870 108.310 88.190 108.570 ;
        RECT 92.930 108.310 93.250 108.570 ;
        RECT 94.785 108.510 95.075 108.555 ;
        RECT 97.990 108.510 98.310 108.570 ;
        RECT 94.785 108.370 98.310 108.510 ;
        RECT 94.785 108.325 95.075 108.370 ;
        RECT 97.990 108.310 98.310 108.370 ;
        RECT 99.830 108.510 100.150 108.570 ;
        RECT 100.305 108.510 100.595 108.555 ;
        RECT 99.830 108.370 100.595 108.510 ;
        RECT 99.830 108.310 100.150 108.370 ;
        RECT 100.305 108.325 100.595 108.370 ;
        RECT 109.490 108.310 109.810 108.570 ;
        RECT 111.330 108.310 111.650 108.570 ;
        RECT 112.725 108.510 113.015 108.555 ;
        RECT 114.090 108.510 114.410 108.570 ;
        RECT 112.725 108.370 114.410 108.510 ;
        RECT 112.725 108.325 113.015 108.370 ;
        RECT 114.090 108.310 114.410 108.370 ;
        RECT 115.025 108.510 115.315 108.555 ;
        RECT 116.390 108.510 116.710 108.570 ;
        RECT 115.025 108.370 116.710 108.510 ;
        RECT 115.025 108.325 115.315 108.370 ;
        RECT 116.390 108.310 116.710 108.370 ;
        RECT 119.150 108.310 119.470 108.570 ;
        RECT 14.660 107.690 127.820 108.170 ;
        RECT 32.210 107.490 32.530 107.550 ;
        RECT 24.940 107.350 32.530 107.490 ;
        RECT 18.985 107.150 19.275 107.195 ;
        RECT 22.225 107.150 22.875 107.195 ;
        RECT 23.470 107.150 23.790 107.210 ;
        RECT 24.940 107.195 25.080 107.350 ;
        RECT 32.210 107.290 32.530 107.350 ;
        RECT 37.745 107.305 38.035 107.535 ;
        RECT 93.850 107.490 94.170 107.550 ;
        RECT 109.030 107.490 109.350 107.550 ;
        RECT 89.340 107.350 94.170 107.490 ;
        RECT 18.985 107.010 23.790 107.150 ;
        RECT 18.985 106.965 19.575 107.010 ;
        RECT 22.225 106.965 22.875 107.010 ;
        RECT 19.285 106.650 19.575 106.965 ;
        RECT 23.470 106.950 23.790 107.010 ;
        RECT 24.865 106.965 25.155 107.195 ;
        RECT 29.565 107.150 29.855 107.195 ;
        RECT 31.750 107.150 32.070 107.210 ;
        RECT 32.805 107.150 33.455 107.195 ;
        RECT 29.565 107.010 33.455 107.150 ;
        RECT 29.565 106.965 30.155 107.010 ;
        RECT 20.365 106.810 20.655 106.855 ;
        RECT 23.945 106.810 24.235 106.855 ;
        RECT 25.780 106.810 26.070 106.855 ;
        RECT 20.365 106.670 26.070 106.810 ;
        RECT 20.365 106.625 20.655 106.670 ;
        RECT 23.945 106.625 24.235 106.670 ;
        RECT 25.780 106.625 26.070 106.670 ;
        RECT 26.705 106.810 26.995 106.855 ;
        RECT 26.705 106.670 29.680 106.810 ;
        RECT 26.705 106.625 26.995 106.670 ;
        RECT 16.125 106.470 16.415 106.515 ;
        RECT 18.870 106.470 19.190 106.530 ;
        RECT 16.125 106.330 19.190 106.470 ;
        RECT 16.125 106.285 16.415 106.330 ;
        RECT 18.870 106.270 19.190 106.330 ;
        RECT 26.245 106.470 26.535 106.515 ;
        RECT 28.990 106.470 29.310 106.530 ;
        RECT 26.245 106.330 29.310 106.470 ;
        RECT 29.540 106.470 29.680 106.670 ;
        RECT 29.865 106.650 30.155 106.965 ;
        RECT 31.750 106.950 32.070 107.010 ;
        RECT 32.805 106.965 33.455 107.010 ;
        RECT 35.445 107.150 35.735 107.195 ;
        RECT 37.820 107.150 37.960 107.305 ;
        RECT 35.445 107.010 37.960 107.150 ;
        RECT 40.950 107.150 41.270 107.210 ;
        RECT 49.805 107.150 50.095 107.195 ;
        RECT 53.045 107.150 53.695 107.195 ;
        RECT 40.950 107.010 45.320 107.150 ;
        RECT 35.445 106.965 35.735 107.010 ;
        RECT 40.950 106.950 41.270 107.010 ;
        RECT 30.945 106.810 31.235 106.855 ;
        RECT 34.525 106.810 34.815 106.855 ;
        RECT 36.360 106.810 36.650 106.855 ;
        RECT 30.945 106.670 36.650 106.810 ;
        RECT 30.945 106.625 31.235 106.670 ;
        RECT 34.525 106.625 34.815 106.670 ;
        RECT 36.360 106.625 36.650 106.670 ;
        RECT 36.810 106.610 37.130 106.870 ;
        RECT 38.650 106.610 38.970 106.870 ;
        RECT 40.505 106.810 40.795 106.855 ;
        RECT 41.040 106.810 41.180 106.950 ;
        RECT 40.505 106.670 41.180 106.810 ;
        RECT 41.410 106.810 41.730 106.870 ;
        RECT 45.180 106.855 45.320 107.010 ;
        RECT 49.805 107.010 53.695 107.150 ;
        RECT 49.805 106.965 50.395 107.010 ;
        RECT 53.045 106.965 53.695 107.010 ;
        RECT 50.105 106.870 50.395 106.965 ;
        RECT 55.670 106.950 55.990 107.210 ;
        RECT 65.330 107.150 65.650 107.210 ;
        RECT 66.365 107.150 66.655 107.195 ;
        RECT 69.605 107.150 70.255 107.195 ;
        RECT 65.330 107.010 70.255 107.150 ;
        RECT 65.330 106.950 65.650 107.010 ;
        RECT 66.365 106.965 66.955 107.010 ;
        RECT 69.605 106.965 70.255 107.010 ;
        RECT 43.265 106.810 43.555 106.855 ;
        RECT 41.410 106.670 43.555 106.810 ;
        RECT 40.505 106.625 40.795 106.670 ;
        RECT 41.410 106.610 41.730 106.670 ;
        RECT 43.265 106.625 43.555 106.670 ;
        RECT 45.105 106.625 45.395 106.855 ;
        RECT 45.565 106.810 45.855 106.855 ;
        RECT 46.010 106.810 46.330 106.870 ;
        RECT 45.565 106.670 46.330 106.810 ;
        RECT 45.565 106.625 45.855 106.670 ;
        RECT 30.370 106.470 30.690 106.530 ;
        RECT 29.540 106.330 30.690 106.470 ;
        RECT 26.245 106.285 26.535 106.330 ;
        RECT 28.990 106.270 29.310 106.330 ;
        RECT 30.370 106.270 30.690 106.330 ;
        RECT 35.430 106.470 35.750 106.530 ;
        RECT 35.430 106.330 42.560 106.470 ;
        RECT 35.430 106.270 35.750 106.330 ;
        RECT 42.420 106.175 42.560 106.330 ;
        RECT 20.365 106.130 20.655 106.175 ;
        RECT 23.485 106.130 23.775 106.175 ;
        RECT 25.375 106.130 25.665 106.175 ;
        RECT 20.365 105.990 25.665 106.130 ;
        RECT 20.365 105.945 20.655 105.990 ;
        RECT 23.485 105.945 23.775 105.990 ;
        RECT 25.375 105.945 25.665 105.990 ;
        RECT 30.945 106.130 31.235 106.175 ;
        RECT 34.065 106.130 34.355 106.175 ;
        RECT 35.955 106.130 36.245 106.175 ;
        RECT 30.945 105.990 36.245 106.130 ;
        RECT 30.945 105.945 31.235 105.990 ;
        RECT 34.065 105.945 34.355 105.990 ;
        RECT 35.955 105.945 36.245 105.990 ;
        RECT 42.345 105.945 42.635 106.175 ;
        RECT 45.180 106.130 45.320 106.625 ;
        RECT 46.010 106.610 46.330 106.670 ;
        RECT 50.105 106.650 50.470 106.870 ;
        RECT 50.150 106.610 50.470 106.650 ;
        RECT 51.185 106.810 51.475 106.855 ;
        RECT 54.765 106.810 55.055 106.855 ;
        RECT 56.600 106.810 56.890 106.855 ;
        RECT 51.185 106.670 56.890 106.810 ;
        RECT 51.185 106.625 51.475 106.670 ;
        RECT 54.765 106.625 55.055 106.670 ;
        RECT 56.600 106.625 56.890 106.670 ;
        RECT 58.445 106.810 58.735 106.855 ;
        RECT 60.270 106.810 60.590 106.870 ;
        RECT 58.445 106.670 60.590 106.810 ;
        RECT 58.445 106.625 58.735 106.670 ;
        RECT 46.945 106.470 47.235 106.515 ;
        RECT 49.690 106.470 50.010 106.530 ;
        RECT 52.450 106.470 52.770 106.530 ;
        RECT 46.945 106.330 50.010 106.470 ;
        RECT 46.945 106.285 47.235 106.330 ;
        RECT 49.690 106.270 50.010 106.330 ;
        RECT 50.470 106.330 56.820 106.470 ;
        RECT 50.470 106.130 50.610 106.330 ;
        RECT 52.450 106.270 52.770 106.330 ;
        RECT 45.180 105.990 50.610 106.130 ;
        RECT 51.185 106.130 51.475 106.175 ;
        RECT 54.305 106.130 54.595 106.175 ;
        RECT 56.195 106.130 56.485 106.175 ;
        RECT 51.185 105.990 56.485 106.130 ;
        RECT 56.680 106.130 56.820 106.330 ;
        RECT 57.050 106.270 57.370 106.530 ;
        RECT 58.520 106.130 58.660 106.625 ;
        RECT 60.270 106.610 60.590 106.670 ;
        RECT 60.730 106.810 61.050 106.870 ;
        RECT 61.665 106.810 61.955 106.855 ;
        RECT 60.730 106.670 61.955 106.810 ;
        RECT 60.730 106.610 61.050 106.670 ;
        RECT 61.665 106.625 61.955 106.670 ;
        RECT 66.665 106.650 66.955 106.965 ;
        RECT 72.230 106.950 72.550 107.210 ;
        RECT 79.245 107.150 79.535 107.195 ;
        RECT 81.890 107.150 82.210 107.210 ;
        RECT 82.485 107.150 83.135 107.195 ;
        RECT 79.245 107.010 83.135 107.150 ;
        RECT 79.245 106.965 79.835 107.010 ;
        RECT 67.745 106.810 68.035 106.855 ;
        RECT 71.325 106.810 71.615 106.855 ;
        RECT 73.160 106.810 73.450 106.855 ;
        RECT 67.745 106.670 73.450 106.810 ;
        RECT 67.745 106.625 68.035 106.670 ;
        RECT 71.325 106.625 71.615 106.670 ;
        RECT 73.160 106.625 73.450 106.670 ;
        RECT 74.990 106.610 75.310 106.870 ;
        RECT 79.545 106.650 79.835 106.965 ;
        RECT 81.890 106.950 82.210 107.010 ;
        RECT 82.485 106.965 83.135 107.010 ;
        RECT 83.730 107.150 84.050 107.210 ;
        RECT 89.340 107.195 89.480 107.350 ;
        RECT 93.850 107.290 94.170 107.350 ;
        RECT 104.060 107.350 109.350 107.490 ;
        RECT 85.125 107.150 85.415 107.195 ;
        RECT 83.730 107.010 85.415 107.150 ;
        RECT 83.730 106.950 84.050 107.010 ;
        RECT 85.125 106.965 85.415 107.010 ;
        RECT 89.265 106.965 89.555 107.195 ;
        RECT 92.125 107.150 92.415 107.195 ;
        RECT 92.930 107.150 93.250 107.210 ;
        RECT 95.365 107.150 96.015 107.195 ;
        RECT 92.125 107.010 96.015 107.150 ;
        RECT 92.125 106.965 92.715 107.010 ;
        RECT 80.625 106.810 80.915 106.855 ;
        RECT 84.205 106.810 84.495 106.855 ;
        RECT 86.040 106.810 86.330 106.855 ;
        RECT 80.625 106.670 86.330 106.810 ;
        RECT 80.625 106.625 80.915 106.670 ;
        RECT 84.205 106.625 84.495 106.670 ;
        RECT 86.040 106.625 86.330 106.670 ;
        RECT 86.950 106.810 87.270 106.870 ;
        RECT 87.425 106.810 87.715 106.855 ;
        RECT 86.950 106.670 87.715 106.810 ;
        RECT 86.950 106.610 87.270 106.670 ;
        RECT 87.425 106.625 87.715 106.670 ;
        RECT 92.425 106.650 92.715 106.965 ;
        RECT 92.930 106.950 93.250 107.010 ;
        RECT 95.365 106.965 96.015 107.010 ;
        RECT 97.990 106.950 98.310 107.210 ;
        RECT 104.060 107.195 104.200 107.350 ;
        RECT 109.030 107.290 109.350 107.350 ;
        RECT 103.985 106.965 104.275 107.195 ;
        RECT 106.845 107.150 107.135 107.195 ;
        RECT 109.490 107.150 109.810 107.210 ;
        RECT 110.085 107.150 110.735 107.195 ;
        RECT 106.845 107.010 110.735 107.150 ;
        RECT 106.845 106.965 107.435 107.010 ;
        RECT 93.505 106.810 93.795 106.855 ;
        RECT 97.085 106.810 97.375 106.855 ;
        RECT 98.920 106.810 99.210 106.855 ;
        RECT 93.505 106.670 99.210 106.810 ;
        RECT 93.505 106.625 93.795 106.670 ;
        RECT 97.085 106.625 97.375 106.670 ;
        RECT 98.920 106.625 99.210 106.670 ;
        RECT 100.765 106.810 101.055 106.855 ;
        RECT 102.590 106.810 102.910 106.870 ;
        RECT 100.765 106.670 102.910 106.810 ;
        RECT 100.765 106.625 101.055 106.670 ;
        RECT 102.590 106.610 102.910 106.670 ;
        RECT 107.145 106.650 107.435 106.965 ;
        RECT 109.490 106.950 109.810 107.010 ;
        RECT 110.085 106.965 110.735 107.010 ;
        RECT 111.330 107.150 111.650 107.210 ;
        RECT 112.725 107.150 113.015 107.195 ;
        RECT 111.330 107.010 113.015 107.150 ;
        RECT 111.330 106.950 111.650 107.010 ;
        RECT 112.725 106.965 113.015 107.010 ;
        RECT 117.310 106.950 117.630 107.210 ;
        RECT 120.070 107.195 120.390 107.210 ;
        RECT 119.605 107.150 120.390 107.195 ;
        RECT 123.205 107.150 123.495 107.195 ;
        RECT 119.605 107.010 123.495 107.150 ;
        RECT 119.605 106.965 120.390 107.010 ;
        RECT 120.070 106.950 120.390 106.965 ;
        RECT 122.905 106.965 123.495 107.010 ;
        RECT 108.225 106.810 108.515 106.855 ;
        RECT 111.805 106.810 112.095 106.855 ;
        RECT 113.640 106.810 113.930 106.855 ;
        RECT 108.225 106.670 113.930 106.810 ;
        RECT 108.225 106.625 108.515 106.670 ;
        RECT 111.805 106.625 112.095 106.670 ;
        RECT 113.640 106.625 113.930 106.670 ;
        RECT 116.410 106.810 116.700 106.855 ;
        RECT 118.245 106.810 118.535 106.855 ;
        RECT 121.825 106.810 122.115 106.855 ;
        RECT 116.410 106.670 122.115 106.810 ;
        RECT 116.410 106.625 116.700 106.670 ;
        RECT 118.245 106.625 118.535 106.670 ;
        RECT 121.825 106.625 122.115 106.670 ;
        RECT 122.905 106.650 123.195 106.965 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 63.505 106.470 63.795 106.515 ;
        RECT 68.550 106.470 68.870 106.530 ;
        RECT 63.505 106.330 68.870 106.470 ;
        RECT 63.505 106.285 63.795 106.330 ;
        RECT 68.550 106.270 68.870 106.330 ;
        RECT 73.610 106.270 73.930 106.530 ;
        RECT 76.385 106.470 76.675 106.515 ;
        RECT 80.050 106.470 80.370 106.530 ;
        RECT 76.385 106.330 80.370 106.470 ;
        RECT 76.385 106.285 76.675 106.330 ;
        RECT 80.050 106.270 80.370 106.330 ;
        RECT 86.490 106.470 86.810 106.530 ;
        RECT 99.370 106.470 99.690 106.530 ;
        RECT 112.250 106.470 112.570 106.530 ;
        RECT 114.105 106.470 114.395 106.515 ;
        RECT 115.945 106.470 116.235 106.515 ;
        RECT 86.490 106.330 116.235 106.470 ;
        RECT 86.490 106.270 86.810 106.330 ;
        RECT 99.370 106.270 99.690 106.330 ;
        RECT 112.250 106.270 112.570 106.330 ;
        RECT 114.105 106.285 114.395 106.330 ;
        RECT 115.945 106.285 116.235 106.330 ;
        RECT 120.990 106.470 121.310 106.530 ;
        RECT 126.065 106.470 126.355 106.515 ;
        RECT 120.990 106.330 126.355 106.470 ;
        RECT 120.990 106.270 121.310 106.330 ;
        RECT 126.065 106.285 126.355 106.330 ;
        RECT 56.680 105.990 58.660 106.130 ;
        RECT 60.745 106.130 61.035 106.175 ;
        RECT 64.410 106.130 64.730 106.190 ;
        RECT 60.745 105.990 64.730 106.130 ;
        RECT 51.185 105.945 51.475 105.990 ;
        RECT 54.305 105.945 54.595 105.990 ;
        RECT 56.195 105.945 56.485 105.990 ;
        RECT 60.745 105.945 61.035 105.990 ;
        RECT 64.410 105.930 64.730 105.990 ;
        RECT 67.745 106.130 68.035 106.175 ;
        RECT 70.865 106.130 71.155 106.175 ;
        RECT 72.755 106.130 73.045 106.175 ;
        RECT 67.745 105.990 73.045 106.130 ;
        RECT 67.745 105.945 68.035 105.990 ;
        RECT 70.865 105.945 71.155 105.990 ;
        RECT 72.755 105.945 73.045 105.990 ;
        RECT 80.625 106.130 80.915 106.175 ;
        RECT 83.745 106.130 84.035 106.175 ;
        RECT 85.635 106.130 85.925 106.175 ;
        RECT 80.625 105.990 85.925 106.130 ;
        RECT 80.625 105.945 80.915 105.990 ;
        RECT 83.745 105.945 84.035 105.990 ;
        RECT 85.635 105.945 85.925 105.990 ;
        RECT 93.505 106.130 93.795 106.175 ;
        RECT 96.625 106.130 96.915 106.175 ;
        RECT 98.515 106.130 98.805 106.175 ;
        RECT 93.505 105.990 98.805 106.130 ;
        RECT 93.505 105.945 93.795 105.990 ;
        RECT 96.625 105.945 96.915 105.990 ;
        RECT 98.515 105.945 98.805 105.990 ;
        RECT 108.225 106.130 108.515 106.175 ;
        RECT 111.345 106.130 111.635 106.175 ;
        RECT 113.235 106.130 113.525 106.175 ;
        RECT 108.225 105.990 113.525 106.130 ;
        RECT 108.225 105.945 108.515 105.990 ;
        RECT 111.345 105.945 111.635 105.990 ;
        RECT 113.235 105.945 113.525 105.990 ;
        RECT 116.815 106.130 117.105 106.175 ;
        RECT 118.705 106.130 118.995 106.175 ;
        RECT 121.825 106.130 122.115 106.175 ;
        RECT 116.815 105.990 122.115 106.130 ;
        RECT 116.815 105.945 117.105 105.990 ;
        RECT 118.705 105.945 118.995 105.990 ;
        RECT 121.825 105.945 122.115 105.990 ;
        RECT 36.350 105.790 36.670 105.850 ;
        RECT 40.045 105.790 40.335 105.835 ;
        RECT 36.350 105.650 40.335 105.790 ;
        RECT 36.350 105.590 36.670 105.650 ;
        RECT 40.045 105.605 40.335 105.650 ;
        RECT 43.250 105.790 43.570 105.850 ;
        RECT 44.645 105.790 44.935 105.835 ;
        RECT 43.250 105.650 44.935 105.790 ;
        RECT 43.250 105.590 43.570 105.650 ;
        RECT 44.645 105.605 44.935 105.650 ;
        RECT 46.485 105.790 46.775 105.835 ;
        RECT 48.310 105.790 48.630 105.850 ;
        RECT 46.485 105.650 48.630 105.790 ;
        RECT 46.485 105.605 46.775 105.650 ;
        RECT 48.310 105.590 48.630 105.650 ;
        RECT 57.050 105.790 57.370 105.850 ;
        RECT 57.985 105.790 58.275 105.835 ;
        RECT 57.050 105.650 58.275 105.790 ;
        RECT 57.050 105.590 57.370 105.650 ;
        RECT 57.985 105.605 58.275 105.650 ;
        RECT 62.585 105.790 62.875 105.835 ;
        RECT 63.950 105.790 64.270 105.850 ;
        RECT 62.585 105.650 64.270 105.790 ;
        RECT 62.585 105.605 62.875 105.650 ;
        RECT 63.950 105.590 64.270 105.650 ;
        RECT 75.910 105.590 76.230 105.850 ;
        RECT 88.330 105.590 88.650 105.850 ;
        RECT 97.530 105.790 97.850 105.850 ;
        RECT 100.305 105.790 100.595 105.835 ;
        RECT 97.530 105.650 100.595 105.790 ;
        RECT 97.530 105.590 97.850 105.650 ;
        RECT 100.305 105.605 100.595 105.650 ;
        RECT 103.065 105.790 103.355 105.835 ;
        RECT 104.430 105.790 104.750 105.850 ;
        RECT 103.065 105.650 104.750 105.790 ;
        RECT 103.065 105.605 103.355 105.650 ;
        RECT 104.430 105.590 104.750 105.650 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 14.660 104.970 127.820 105.450 ;
        RECT 28.990 104.770 29.310 104.830 ;
        RECT 36.810 104.770 37.130 104.830 ;
        RECT 28.990 104.630 37.130 104.770 ;
        RECT 28.990 104.570 29.310 104.630 ;
        RECT 36.810 104.570 37.130 104.630 ;
        RECT 50.150 104.770 50.470 104.830 ;
        RECT 52.005 104.770 52.295 104.815 ;
        RECT 50.150 104.630 52.295 104.770 ;
        RECT 50.150 104.570 50.470 104.630 ;
        RECT 52.005 104.585 52.295 104.630 ;
        RECT 56.590 104.770 56.910 104.830 ;
        RECT 73.610 104.770 73.930 104.830 ;
        RECT 56.590 104.630 73.930 104.770 ;
        RECT 56.590 104.570 56.910 104.630 ;
        RECT 29.080 104.135 29.220 104.570 ;
        RECT 29.875 104.430 30.165 104.475 ;
        RECT 31.765 104.430 32.055 104.475 ;
        RECT 34.885 104.430 35.175 104.475 ;
        RECT 29.875 104.290 35.175 104.430 ;
        RECT 29.875 104.245 30.165 104.290 ;
        RECT 31.765 104.245 32.055 104.290 ;
        RECT 34.885 104.245 35.175 104.290 ;
        RECT 43.825 104.430 44.115 104.475 ;
        RECT 46.945 104.430 47.235 104.475 ;
        RECT 48.835 104.430 49.125 104.475 ;
        RECT 50.610 104.430 50.930 104.490 ;
        RECT 56.680 104.430 56.820 104.570 ;
        RECT 43.825 104.290 49.125 104.430 ;
        RECT 43.825 104.245 44.115 104.290 ;
        RECT 46.945 104.245 47.235 104.290 ;
        RECT 48.835 104.245 49.125 104.290 ;
        RECT 50.470 104.290 56.820 104.430 ;
        RECT 57.165 104.430 57.455 104.475 ;
        RECT 60.285 104.430 60.575 104.475 ;
        RECT 62.175 104.430 62.465 104.475 ;
        RECT 57.165 104.290 62.465 104.430 ;
        RECT 50.470 104.230 50.930 104.290 ;
        RECT 57.165 104.245 57.455 104.290 ;
        RECT 60.285 104.245 60.575 104.290 ;
        RECT 62.175 104.245 62.465 104.290 ;
        RECT 29.005 103.905 29.295 104.135 ;
        RECT 30.385 104.090 30.675 104.135 ;
        RECT 35.430 104.090 35.750 104.150 ;
        RECT 36.350 104.090 36.670 104.150 ;
        RECT 30.385 103.950 35.750 104.090 ;
        RECT 30.385 103.905 30.675 103.950 ;
        RECT 35.430 103.890 35.750 103.950 ;
        RECT 35.980 103.950 36.670 104.090 ;
        RECT 27.610 103.550 27.930 103.810 ;
        RECT 29.470 103.750 29.760 103.795 ;
        RECT 31.305 103.750 31.595 103.795 ;
        RECT 34.885 103.750 35.175 103.795 ;
        RECT 35.980 103.770 36.120 103.950 ;
        RECT 36.350 103.890 36.670 103.950 ;
        RECT 48.310 103.890 48.630 104.150 ;
        RECT 49.705 104.090 49.995 104.135 ;
        RECT 50.470 104.090 50.610 104.230 ;
        RECT 49.705 103.950 50.610 104.090 ;
        RECT 57.970 104.090 58.290 104.150 ;
        RECT 63.120 104.135 63.260 104.630 ;
        RECT 73.610 104.570 73.930 104.630 ;
        RECT 79.130 104.770 79.450 104.830 ;
        RECT 125.145 104.770 125.435 104.815 ;
        RECT 79.130 104.630 125.435 104.770 ;
        RECT 79.130 104.570 79.450 104.630 ;
        RECT 125.145 104.585 125.435 104.630 ;
        RECT 67.745 104.430 68.035 104.475 ;
        RECT 70.865 104.430 71.155 104.475 ;
        RECT 72.755 104.430 73.045 104.475 ;
        RECT 67.745 104.290 73.045 104.430 ;
        RECT 67.745 104.245 68.035 104.290 ;
        RECT 70.865 104.245 71.155 104.290 ;
        RECT 72.755 104.245 73.045 104.290 ;
        RECT 80.625 104.430 80.915 104.475 ;
        RECT 83.745 104.430 84.035 104.475 ;
        RECT 85.635 104.430 85.925 104.475 ;
        RECT 80.625 104.290 85.925 104.430 ;
        RECT 80.625 104.245 80.915 104.290 ;
        RECT 83.745 104.245 84.035 104.290 ;
        RECT 85.635 104.245 85.925 104.290 ;
        RECT 91.205 104.430 91.495 104.475 ;
        RECT 94.325 104.430 94.615 104.475 ;
        RECT 96.215 104.430 96.505 104.475 ;
        RECT 91.205 104.290 96.505 104.430 ;
        RECT 91.205 104.245 91.495 104.290 ;
        RECT 94.325 104.245 94.615 104.290 ;
        RECT 96.215 104.245 96.505 104.290 ;
        RECT 106.385 104.430 106.675 104.475 ;
        RECT 109.505 104.430 109.795 104.475 ;
        RECT 111.395 104.430 111.685 104.475 ;
        RECT 106.385 104.290 111.685 104.430 ;
        RECT 106.385 104.245 106.675 104.290 ;
        RECT 109.505 104.245 109.795 104.290 ;
        RECT 111.395 104.245 111.685 104.290 ;
        RECT 113.595 104.430 113.885 104.475 ;
        RECT 115.485 104.430 115.775 104.475 ;
        RECT 118.605 104.430 118.895 104.475 ;
        RECT 113.595 104.290 118.895 104.430 ;
        RECT 113.595 104.245 113.885 104.290 ;
        RECT 115.485 104.245 115.775 104.290 ;
        RECT 118.605 104.245 118.895 104.290 ;
        RECT 61.665 104.090 61.955 104.135 ;
        RECT 57.970 103.950 61.955 104.090 ;
        RECT 49.705 103.905 49.995 103.950 ;
        RECT 57.970 103.890 58.290 103.950 ;
        RECT 61.665 103.905 61.955 103.950 ;
        RECT 63.045 103.905 63.335 104.135 ;
        RECT 63.950 104.090 64.270 104.150 ;
        RECT 72.245 104.090 72.535 104.135 ;
        RECT 63.950 103.950 72.535 104.090 ;
        RECT 63.950 103.890 64.270 103.950 ;
        RECT 72.245 103.905 72.535 103.950 ;
        RECT 73.610 103.890 73.930 104.150 ;
        RECT 75.910 104.090 76.230 104.150 ;
        RECT 85.125 104.090 85.415 104.135 ;
        RECT 75.910 103.950 85.415 104.090 ;
        RECT 75.910 103.890 76.230 103.950 ;
        RECT 85.125 103.905 85.415 103.950 ;
        RECT 86.490 103.890 86.810 104.150 ;
        RECT 88.330 104.090 88.650 104.150 ;
        RECT 95.705 104.090 95.995 104.135 ;
        RECT 88.330 103.950 95.995 104.090 ;
        RECT 88.330 103.890 88.650 103.950 ;
        RECT 95.705 103.905 95.995 103.950 ;
        RECT 97.085 104.090 97.375 104.135 ;
        RECT 99.370 104.090 99.690 104.150 ;
        RECT 97.085 103.950 99.690 104.090 ;
        RECT 97.085 103.905 97.375 103.950 ;
        RECT 99.370 103.890 99.690 103.950 ;
        RECT 110.870 103.890 111.190 104.150 ;
        RECT 112.250 104.090 112.570 104.150 ;
        RECT 112.725 104.090 113.015 104.135 ;
        RECT 112.250 103.950 113.015 104.090 ;
        RECT 112.250 103.890 112.570 103.950 ;
        RECT 112.725 103.905 113.015 103.950 ;
        RECT 114.090 103.890 114.410 104.150 ;
        RECT 115.930 104.090 116.250 104.150 ;
        RECT 122.845 104.090 123.135 104.135 ;
        RECT 115.930 103.950 123.135 104.090 ;
        RECT 115.930 103.890 116.250 103.950 ;
        RECT 122.845 103.905 123.135 103.950 ;
        RECT 29.470 103.610 35.175 103.750 ;
        RECT 29.470 103.565 29.760 103.610 ;
        RECT 31.305 103.565 31.595 103.610 ;
        RECT 34.885 103.565 35.175 103.610 ;
        RECT 35.965 103.455 36.255 103.770 ;
        RECT 32.665 103.410 33.315 103.455 ;
        RECT 35.965 103.410 36.555 103.455 ;
        RECT 32.665 103.270 36.555 103.410 ;
        RECT 32.665 103.225 33.315 103.270 ;
        RECT 36.265 103.225 36.555 103.270 ;
        RECT 39.110 103.210 39.430 103.470 ;
        RECT 42.745 103.455 43.035 103.770 ;
        RECT 43.825 103.750 44.115 103.795 ;
        RECT 47.405 103.750 47.695 103.795 ;
        RECT 49.240 103.750 49.530 103.795 ;
        RECT 43.825 103.610 49.530 103.750 ;
        RECT 43.825 103.565 44.115 103.610 ;
        RECT 47.405 103.565 47.695 103.610 ;
        RECT 49.240 103.565 49.530 103.610 ;
        RECT 52.450 103.550 52.770 103.810 ;
        RECT 39.585 103.225 39.875 103.455 ;
        RECT 42.445 103.410 43.035 103.455 ;
        RECT 43.250 103.410 43.570 103.470 ;
        RECT 45.685 103.410 46.335 103.455 ;
        RECT 42.445 103.270 46.335 103.410 ;
        RECT 42.445 103.225 42.735 103.270 ;
        RECT 28.070 102.870 28.390 103.130 ;
        RECT 39.660 103.070 39.800 103.225 ;
        RECT 43.250 103.210 43.570 103.270 ;
        RECT 45.685 103.225 46.335 103.270 ;
        RECT 52.925 103.410 53.215 103.455 ;
        RECT 54.750 103.410 55.070 103.470 ;
        RECT 56.085 103.455 56.375 103.770 ;
        RECT 57.165 103.750 57.455 103.795 ;
        RECT 60.745 103.750 61.035 103.795 ;
        RECT 62.580 103.750 62.870 103.795 ;
        RECT 57.165 103.610 62.870 103.750 ;
        RECT 57.165 103.565 57.455 103.610 ;
        RECT 60.745 103.565 61.035 103.610 ;
        RECT 62.580 103.565 62.870 103.610 ;
        RECT 52.925 103.270 55.070 103.410 ;
        RECT 52.925 103.225 53.215 103.270 ;
        RECT 54.750 103.210 55.070 103.270 ;
        RECT 55.785 103.410 56.375 103.455 ;
        RECT 56.590 103.410 56.910 103.470 ;
        RECT 59.025 103.410 59.675 103.455 ;
        RECT 55.785 103.270 59.675 103.410 ;
        RECT 55.785 103.225 56.075 103.270 ;
        RECT 56.590 103.210 56.910 103.270 ;
        RECT 59.025 103.225 59.675 103.270 ;
        RECT 61.190 103.410 61.510 103.470 ;
        RECT 63.505 103.410 63.795 103.455 ;
        RECT 61.190 103.270 63.795 103.410 ;
        RECT 61.190 103.210 61.510 103.270 ;
        RECT 63.505 103.225 63.795 103.270 ;
        RECT 64.410 103.410 64.730 103.470 ;
        RECT 66.665 103.455 66.955 103.770 ;
        RECT 67.745 103.750 68.035 103.795 ;
        RECT 71.325 103.750 71.615 103.795 ;
        RECT 73.160 103.750 73.450 103.795 ;
        RECT 79.590 103.770 79.910 103.810 ;
        RECT 67.745 103.610 73.450 103.750 ;
        RECT 67.745 103.565 68.035 103.610 ;
        RECT 71.325 103.565 71.615 103.610 ;
        RECT 73.160 103.565 73.450 103.610 ;
        RECT 79.545 103.550 79.910 103.770 ;
        RECT 80.625 103.750 80.915 103.795 ;
        RECT 84.205 103.750 84.495 103.795 ;
        RECT 86.040 103.750 86.330 103.795 ;
        RECT 80.625 103.610 86.330 103.750 ;
        RECT 80.625 103.565 80.915 103.610 ;
        RECT 84.205 103.565 84.495 103.610 ;
        RECT 86.040 103.565 86.330 103.610 ;
        RECT 66.365 103.410 66.955 103.455 ;
        RECT 69.605 103.410 70.255 103.455 ;
        RECT 64.410 103.270 70.255 103.410 ;
        RECT 64.410 103.210 64.730 103.270 ;
        RECT 66.365 103.225 66.655 103.270 ;
        RECT 69.605 103.225 70.255 103.270 ;
        RECT 74.070 103.410 74.390 103.470 ;
        RECT 79.545 103.455 79.835 103.550 ;
        RECT 76.385 103.410 76.675 103.455 ;
        RECT 74.070 103.270 76.675 103.410 ;
        RECT 74.070 103.210 74.390 103.270 ;
        RECT 76.385 103.225 76.675 103.270 ;
        RECT 79.245 103.410 79.835 103.455 ;
        RECT 82.485 103.410 83.135 103.455 ;
        RECT 79.245 103.270 83.135 103.410 ;
        RECT 79.245 103.225 79.535 103.270 ;
        RECT 82.485 103.225 83.135 103.270 ;
        RECT 86.950 103.210 87.270 103.470 ;
        RECT 87.870 103.410 88.190 103.470 ;
        RECT 90.125 103.455 90.415 103.770 ;
        RECT 91.205 103.750 91.495 103.795 ;
        RECT 94.785 103.750 95.075 103.795 ;
        RECT 96.620 103.750 96.910 103.795 ;
        RECT 91.205 103.610 96.910 103.750 ;
        RECT 91.205 103.565 91.495 103.610 ;
        RECT 94.785 103.565 95.075 103.610 ;
        RECT 96.620 103.565 96.910 103.610 ;
        RECT 89.825 103.410 90.415 103.455 ;
        RECT 93.065 103.410 93.715 103.455 ;
        RECT 87.870 103.270 93.715 103.410 ;
        RECT 87.870 103.210 88.190 103.270 ;
        RECT 89.825 103.225 90.115 103.270 ;
        RECT 93.065 103.225 93.715 103.270 ;
        RECT 102.145 103.410 102.435 103.455 ;
        RECT 103.970 103.410 104.290 103.470 ;
        RECT 102.145 103.270 104.290 103.410 ;
        RECT 102.145 103.225 102.435 103.270 ;
        RECT 103.970 103.210 104.290 103.270 ;
        RECT 104.430 103.410 104.750 103.470 ;
        RECT 105.305 103.455 105.595 103.770 ;
        RECT 106.385 103.750 106.675 103.795 ;
        RECT 109.965 103.750 110.255 103.795 ;
        RECT 111.800 103.750 112.090 103.795 ;
        RECT 106.385 103.610 112.090 103.750 ;
        RECT 106.385 103.565 106.675 103.610 ;
        RECT 109.965 103.565 110.255 103.610 ;
        RECT 111.800 103.565 112.090 103.610 ;
        RECT 113.190 103.750 113.480 103.795 ;
        RECT 115.025 103.750 115.315 103.795 ;
        RECT 118.605 103.750 118.895 103.795 ;
        RECT 113.190 103.610 118.895 103.750 ;
        RECT 113.190 103.565 113.480 103.610 ;
        RECT 115.025 103.565 115.315 103.610 ;
        RECT 118.605 103.565 118.895 103.610 ;
        RECT 116.390 103.455 116.710 103.470 ;
        RECT 119.685 103.455 119.975 103.770 ;
        RECT 126.050 103.550 126.370 103.810 ;
        RECT 105.005 103.410 105.595 103.455 ;
        RECT 108.245 103.410 108.895 103.455 ;
        RECT 104.430 103.270 108.895 103.410 ;
        RECT 104.430 103.210 104.750 103.270 ;
        RECT 105.005 103.225 105.295 103.270 ;
        RECT 108.245 103.225 108.895 103.270 ;
        RECT 116.385 103.410 117.035 103.455 ;
        RECT 119.685 103.410 120.275 103.455 ;
        RECT 116.385 103.270 120.275 103.410 ;
        RECT 116.385 103.225 117.035 103.270 ;
        RECT 119.985 103.225 120.275 103.270 ;
        RECT 116.390 103.210 116.710 103.225 ;
        RECT 44.170 103.070 44.490 103.130 ;
        RECT 39.660 102.930 44.490 103.070 ;
        RECT 44.170 102.870 44.490 102.930 ;
        RECT 14.660 102.250 127.820 102.730 ;
        RECT 120.070 101.850 120.390 102.110 ;
        RECT 27.725 101.710 28.015 101.755 ;
        RECT 30.965 101.710 31.615 101.755 ;
        RECT 27.725 101.570 31.615 101.710 ;
        RECT 27.725 101.525 28.315 101.570 ;
        RECT 30.965 101.525 31.615 101.570 ;
        RECT 33.605 101.710 33.895 101.755 ;
        RECT 34.050 101.710 34.370 101.770 ;
        RECT 97.530 101.755 97.850 101.770 ;
        RECT 33.605 101.570 34.370 101.710 ;
        RECT 33.605 101.525 33.895 101.570 ;
        RECT 28.025 101.430 28.315 101.525 ;
        RECT 34.050 101.510 34.370 101.570 ;
        RECT 93.965 101.710 94.255 101.755 ;
        RECT 97.205 101.710 97.855 101.755 ;
        RECT 93.965 101.570 97.855 101.710 ;
        RECT 93.965 101.525 94.555 101.570 ;
        RECT 97.205 101.525 97.855 101.570 ;
        RECT 28.025 101.210 28.390 101.430 ;
        RECT 28.070 101.170 28.390 101.210 ;
        RECT 29.105 101.370 29.395 101.415 ;
        RECT 32.685 101.370 32.975 101.415 ;
        RECT 34.520 101.370 34.810 101.415 ;
        RECT 29.105 101.230 34.810 101.370 ;
        RECT 29.105 101.185 29.395 101.230 ;
        RECT 32.685 101.185 32.975 101.230 ;
        RECT 34.520 101.185 34.810 101.230 ;
        RECT 34.985 101.370 35.275 101.415 ;
        RECT 36.810 101.370 37.130 101.430 ;
        RECT 34.985 101.230 37.130 101.370 ;
        RECT 34.985 101.185 35.275 101.230 ;
        RECT 36.810 101.170 37.130 101.230 ;
        RECT 94.265 101.210 94.555 101.525 ;
        RECT 97.530 101.510 97.850 101.525 ;
        RECT 99.830 101.510 100.150 101.770 ;
        RECT 95.345 101.370 95.635 101.415 ;
        RECT 98.925 101.370 99.215 101.415 ;
        RECT 100.760 101.370 101.050 101.415 ;
        RECT 95.345 101.230 101.050 101.370 ;
        RECT 95.345 101.185 95.635 101.230 ;
        RECT 98.925 101.185 99.215 101.230 ;
        RECT 100.760 101.185 101.050 101.230 ;
        RECT 119.610 101.170 119.930 101.430 ;
        RECT 24.865 101.030 25.155 101.075 ;
        RECT 26.230 101.030 26.550 101.090 ;
        RECT 24.865 100.890 26.550 101.030 ;
        RECT 24.865 100.845 25.155 100.890 ;
        RECT 26.230 100.830 26.550 100.890 ;
        RECT 91.105 101.030 91.395 101.075 ;
        RECT 97.990 101.030 98.310 101.090 ;
        RECT 91.105 100.890 98.310 101.030 ;
        RECT 91.105 100.845 91.395 100.890 ;
        RECT 97.990 100.830 98.310 100.890 ;
        RECT 99.370 101.030 99.690 101.090 ;
        RECT 101.225 101.030 101.515 101.075 ;
        RECT 99.370 100.890 101.515 101.030 ;
        RECT 99.370 100.830 99.690 100.890 ;
        RECT 101.225 100.845 101.515 100.890 ;
        RECT 29.105 100.690 29.395 100.735 ;
        RECT 32.225 100.690 32.515 100.735 ;
        RECT 34.115 100.690 34.405 100.735 ;
        RECT 29.105 100.550 34.405 100.690 ;
        RECT 29.105 100.505 29.395 100.550 ;
        RECT 32.225 100.505 32.515 100.550 ;
        RECT 34.115 100.505 34.405 100.550 ;
        RECT 95.345 100.690 95.635 100.735 ;
        RECT 98.465 100.690 98.755 100.735 ;
        RECT 100.355 100.690 100.645 100.735 ;
        RECT 95.345 100.550 100.645 100.690 ;
        RECT 95.345 100.505 95.635 100.550 ;
        RECT 98.465 100.505 98.755 100.550 ;
        RECT 100.355 100.505 100.645 100.550 ;
        RECT 14.660 99.530 127.820 100.010 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 16.880 211.105 18.760 211.475 ;
        RECT 46.880 211.105 48.760 211.475 ;
        RECT 76.880 211.105 78.760 211.475 ;
        RECT 106.880 211.105 108.760 211.475 ;
        RECT 31.880 208.385 33.760 208.755 ;
        RECT 61.880 208.385 63.760 208.755 ;
        RECT 91.880 208.385 93.760 208.755 ;
        RECT 121.880 208.385 123.760 208.755 ;
        RECT 73.640 207.560 73.900 207.880 ;
        RECT 66.280 206.880 66.540 207.200 ;
        RECT 73.180 206.880 73.440 207.200 ;
        RECT 16.880 205.665 18.760 206.035 ;
        RECT 46.880 205.665 48.760 206.035 ;
        RECT 66.340 204.820 66.480 206.880 ;
        RECT 66.280 204.500 66.540 204.820 ;
        RECT 63.980 204.160 64.240 204.480 ;
        RECT 31.880 202.945 33.760 203.315 ;
        RECT 61.880 202.945 63.760 203.315 ;
        RECT 64.040 202.780 64.180 204.160 ;
        RECT 64.900 203.480 65.160 203.800 ;
        RECT 63.980 202.460 64.240 202.780 ;
        RECT 61.220 201.780 61.480 202.100 ;
        RECT 16.880 200.225 18.760 200.595 ;
        RECT 46.880 200.225 48.760 200.595 ;
        RECT 61.280 200.060 61.420 201.780 ;
        RECT 61.220 199.740 61.480 200.060 ;
        RECT 31.880 197.505 33.760 197.875 ;
        RECT 61.880 197.505 63.760 197.875 ;
        RECT 50.640 196.340 50.900 196.660 ;
        RECT 49.260 196.000 49.520 196.320 ;
        RECT 16.880 194.785 18.760 195.155 ;
        RECT 46.880 194.785 48.760 195.155 ;
        RECT 49.320 194.280 49.460 196.000 ;
        RECT 50.700 194.620 50.840 196.340 ;
        RECT 53.400 195.320 53.660 195.640 ;
        RECT 58.000 195.320 58.260 195.640 ;
        RECT 50.640 194.530 50.900 194.620 ;
        RECT 49.780 194.390 50.900 194.530 ;
        RECT 49.260 193.960 49.520 194.280 ;
        RECT 46.040 193.620 46.300 193.940 ;
        RECT 31.880 192.065 33.760 192.435 ;
        RECT 41.440 190.900 41.700 191.220 ;
        RECT 39.140 190.220 39.400 190.540 ;
        RECT 16.880 189.345 18.760 189.715 ;
        RECT 28.560 187.840 28.820 188.160 ;
        RECT 36.380 187.840 36.640 188.160 ;
        RECT 23.040 185.460 23.300 185.780 ;
        RECT 16.880 183.905 18.760 184.275 ;
        RECT 23.100 183.740 23.240 185.460 ;
        RECT 28.620 185.100 28.760 187.840 ;
        RECT 31.880 186.625 33.760 186.995 ;
        RECT 36.440 185.440 36.580 187.840 ;
        RECT 37.760 187.160 38.020 187.480 ;
        RECT 36.380 185.120 36.640 185.440 ;
        RECT 28.560 184.780 28.820 185.100 ;
        RECT 29.940 184.440 30.200 184.760 ;
        RECT 30.400 184.440 30.660 184.760 ;
        RECT 23.040 183.420 23.300 183.740 ;
        RECT 30.000 183.060 30.140 184.440 ;
        RECT 30.460 183.740 30.600 184.440 ;
        RECT 30.400 183.420 30.660 183.740 ;
        RECT 34.080 183.080 34.340 183.400 ;
        RECT 29.940 182.740 30.200 183.060 ;
        RECT 31.880 181.185 33.760 181.555 ;
        RECT 34.140 179.660 34.280 183.080 ;
        RECT 35.920 182.740 36.180 183.060 ;
        RECT 26.260 179.340 26.520 179.660 ;
        RECT 27.640 179.340 27.900 179.660 ;
        RECT 34.080 179.340 34.340 179.660 ;
        RECT 35.000 179.340 35.260 179.660 ;
        RECT 16.880 178.465 18.760 178.835 ;
        RECT 26.320 175.580 26.460 179.340 ;
        RECT 27.700 178.300 27.840 179.340 ;
        RECT 27.640 177.980 27.900 178.300 ;
        RECT 30.400 176.960 30.660 177.280 ;
        RECT 28.100 176.280 28.360 176.600 ;
        RECT 26.260 175.260 26.520 175.580 ;
        RECT 28.160 174.220 28.300 176.280 ;
        RECT 28.100 173.900 28.360 174.220 ;
        RECT 16.880 173.025 18.760 173.395 ;
        RECT 30.460 169.120 30.600 176.960 ;
        RECT 31.880 175.745 33.760 176.115 ;
        RECT 34.140 174.220 34.280 179.340 ;
        RECT 34.540 176.280 34.800 176.600 ;
        RECT 34.600 174.560 34.740 176.280 ;
        RECT 34.540 174.240 34.800 174.560 ;
        RECT 34.080 173.900 34.340 174.220 ;
        RECT 31.880 170.305 33.760 170.675 ;
        RECT 30.400 168.800 30.660 169.120 ;
        RECT 29.940 168.120 30.200 168.440 ;
        RECT 34.080 168.120 34.340 168.440 ;
        RECT 16.880 167.585 18.760 167.955 ;
        RECT 30.000 167.080 30.140 168.120 ;
        RECT 24.880 166.760 25.140 167.080 ;
        RECT 29.940 166.760 30.200 167.080 ;
        RECT 24.940 164.700 25.080 166.760 ;
        RECT 27.180 166.080 27.440 166.400 ;
        RECT 24.880 164.380 25.140 164.700 ;
        RECT 27.240 163.680 27.380 166.080 ;
        RECT 29.940 165.740 30.200 166.060 ;
        RECT 28.560 165.400 28.820 165.720 ;
        RECT 28.620 164.020 28.760 165.400 ;
        RECT 28.560 163.700 28.820 164.020 ;
        RECT 29.020 163.700 29.280 164.020 ;
        RECT 26.720 163.360 26.980 163.680 ;
        RECT 27.180 163.360 27.440 163.680 ;
        RECT 16.880 162.145 18.760 162.515 ;
        RECT 26.780 161.980 26.920 163.360 ;
        RECT 29.080 163.340 29.220 163.700 ;
        RECT 29.020 163.020 29.280 163.340 ;
        RECT 26.720 161.660 26.980 161.980 ;
        RECT 18.900 161.320 19.160 161.640 ;
        RECT 18.960 159.260 19.100 161.320 ;
        RECT 29.080 161.300 29.220 163.020 ;
        RECT 30.000 161.980 30.140 165.740 ;
        RECT 31.880 164.865 33.760 165.235 ;
        RECT 34.140 163.680 34.280 168.120 ;
        RECT 34.540 166.420 34.800 166.740 ;
        RECT 34.080 163.360 34.340 163.680 ;
        RECT 34.600 161.980 34.740 166.420 ;
        RECT 29.940 161.660 30.200 161.980 ;
        RECT 34.540 161.660 34.800 161.980 ;
        RECT 31.320 161.320 31.580 161.640 ;
        RECT 35.060 161.380 35.200 179.340 ;
        RECT 35.460 176.960 35.720 177.280 ;
        RECT 35.520 172.860 35.660 176.960 ;
        RECT 35.460 172.540 35.720 172.860 ;
        RECT 35.980 171.840 36.120 182.740 ;
        RECT 35.920 171.520 36.180 171.840 ;
        RECT 35.460 170.840 35.720 171.160 ;
        RECT 36.440 170.900 36.580 185.120 ;
        RECT 37.820 185.100 37.960 187.160 ;
        RECT 39.200 186.460 39.340 190.220 ;
        RECT 39.140 186.140 39.400 186.460 ;
        RECT 41.500 185.780 41.640 190.900 ;
        RECT 45.120 190.560 45.380 190.880 ;
        RECT 44.660 187.840 44.920 188.160 ;
        RECT 44.720 186.120 44.860 187.840 ;
        RECT 44.660 185.800 44.920 186.120 ;
        RECT 38.220 185.460 38.480 185.780 ;
        RECT 41.440 185.460 41.700 185.780 ;
        RECT 37.760 184.780 38.020 185.100 ;
        RECT 37.820 183.060 37.960 184.780 ;
        RECT 37.760 182.740 38.020 183.060 ;
        RECT 37.300 179.680 37.560 180.000 ;
        RECT 36.840 179.000 37.100 179.320 ;
        RECT 36.900 177.280 37.040 179.000 ;
        RECT 36.840 176.960 37.100 177.280 ;
        RECT 27.180 160.980 27.440 161.300 ;
        RECT 29.020 160.980 29.280 161.300 ;
        RECT 25.800 160.640 26.060 160.960 ;
        RECT 21.660 159.960 21.920 160.280 ;
        RECT 18.900 158.940 19.160 159.260 ;
        RECT 21.720 158.580 21.860 159.960 ;
        RECT 25.860 159.260 26.000 160.640 ;
        RECT 25.800 158.940 26.060 159.260 ;
        RECT 21.200 158.260 21.460 158.580 ;
        RECT 21.660 158.260 21.920 158.580 ;
        RECT 19.360 157.240 19.620 157.560 ;
        RECT 16.880 156.705 18.760 157.075 ;
        RECT 19.420 156.200 19.560 157.240 ;
        RECT 19.360 155.880 19.620 156.200 ;
        RECT 21.260 153.140 21.400 158.260 ;
        RECT 22.120 157.240 22.380 157.560 ;
        RECT 22.180 156.540 22.320 157.240 ;
        RECT 22.120 156.220 22.380 156.540 ;
        RECT 22.180 153.140 22.320 156.220 ;
        RECT 27.240 155.860 27.380 160.980 ;
        RECT 30.860 160.640 31.120 160.960 ;
        RECT 30.920 158.920 31.060 160.640 ;
        RECT 31.380 159.260 31.520 161.320 ;
        RECT 34.080 160.980 34.340 161.300 ;
        RECT 34.600 161.240 35.200 161.380 ;
        RECT 34.140 160.280 34.280 160.980 ;
        RECT 34.080 159.960 34.340 160.280 ;
        RECT 31.880 159.425 33.760 159.795 ;
        RECT 31.320 158.940 31.580 159.260 ;
        RECT 30.860 158.600 31.120 158.920 ;
        RECT 29.940 158.260 30.200 158.580 ;
        RECT 27.180 155.540 27.440 155.860 ;
        RECT 27.640 155.540 27.900 155.860 ;
        RECT 27.700 153.820 27.840 155.540 ;
        RECT 27.640 153.500 27.900 153.820 ;
        RECT 21.200 152.820 21.460 153.140 ;
        RECT 22.120 152.820 22.380 153.140 ;
        RECT 16.880 151.265 18.760 151.635 ;
        RECT 20.280 150.440 20.540 150.760 ;
        RECT 16.880 145.825 18.760 146.195 ;
        RECT 20.340 145.660 20.480 150.440 ;
        RECT 21.260 147.700 21.400 152.820 ;
        RECT 22.580 151.800 22.840 152.120 ;
        RECT 22.640 150.080 22.780 151.800 ;
        RECT 30.000 150.420 30.140 158.260 ;
        RECT 30.920 155.520 31.060 158.600 ;
        RECT 32.240 157.920 32.500 158.240 ;
        RECT 31.320 155.540 31.580 155.860 ;
        RECT 30.860 155.200 31.120 155.520 ;
        RECT 31.380 152.120 31.520 155.540 ;
        RECT 32.300 155.180 32.440 157.920 ;
        RECT 33.620 156.220 33.880 156.540 ;
        RECT 33.680 155.860 33.820 156.220 ;
        RECT 33.620 155.540 33.880 155.860 ;
        RECT 34.080 155.200 34.340 155.520 ;
        RECT 32.240 154.860 32.500 155.180 ;
        RECT 31.880 153.985 33.760 154.355 ;
        RECT 33.620 152.140 33.880 152.460 ;
        RECT 31.320 151.800 31.580 152.120 ;
        RECT 31.380 150.760 31.520 151.800 ;
        RECT 33.680 151.100 33.820 152.140 ;
        RECT 33.620 150.780 33.880 151.100 ;
        RECT 31.320 150.440 31.580 150.760 ;
        RECT 29.940 150.100 30.200 150.420 ;
        RECT 22.580 149.760 22.840 150.080 ;
        RECT 24.880 149.760 25.140 150.080 ;
        RECT 21.200 147.380 21.460 147.700 ;
        RECT 22.640 146.680 22.780 149.760 ;
        RECT 24.940 148.380 25.080 149.760 ;
        RECT 24.880 148.060 25.140 148.380 ;
        RECT 28.560 147.720 28.820 148.040 ;
        RECT 23.040 146.700 23.300 147.020 ;
        RECT 22.580 146.360 22.840 146.680 ;
        RECT 23.100 145.660 23.240 146.700 ;
        RECT 28.620 146.680 28.760 147.720 ;
        RECT 28.560 146.360 28.820 146.680 ;
        RECT 29.020 146.360 29.280 146.680 ;
        RECT 20.280 145.340 20.540 145.660 ;
        RECT 23.040 145.340 23.300 145.660 ;
        RECT 29.080 144.640 29.220 146.360 ;
        RECT 30.000 145.060 30.140 150.100 ;
        RECT 31.380 147.360 31.520 150.440 ;
        RECT 31.880 148.545 33.760 148.915 ;
        RECT 34.140 147.700 34.280 155.200 ;
        RECT 34.080 147.380 34.340 147.700 ;
        RECT 31.320 147.040 31.580 147.360 ;
        RECT 30.000 144.980 30.600 145.060 ;
        RECT 30.000 144.920 30.660 144.980 ;
        RECT 29.020 144.320 29.280 144.640 ;
        RECT 30.000 143.960 30.140 144.920 ;
        RECT 30.400 144.660 30.660 144.920 ;
        RECT 29.940 143.640 30.200 143.960 ;
        RECT 31.880 143.105 33.760 143.475 ;
        RECT 34.600 142.260 34.740 161.240 ;
        RECT 35.000 159.960 35.260 160.280 ;
        RECT 35.060 157.560 35.200 159.960 ;
        RECT 35.000 157.240 35.260 157.560 ;
        RECT 35.060 156.540 35.200 157.240 ;
        RECT 35.000 156.220 35.260 156.540 ;
        RECT 35.000 151.800 35.260 152.120 ;
        RECT 34.540 141.940 34.800 142.260 ;
        RECT 35.060 141.920 35.200 151.800 ;
        RECT 35.000 141.600 35.260 141.920 ;
        RECT 29.480 140.920 29.740 141.240 ;
        RECT 16.880 140.385 18.760 140.755 ;
        RECT 19.360 139.560 19.620 139.880 ;
        RECT 18.900 135.480 19.160 135.800 ;
        RECT 16.880 134.945 18.760 135.315 ;
        RECT 18.960 134.100 19.100 135.480 ;
        RECT 19.420 134.780 19.560 139.560 ;
        RECT 23.500 138.880 23.760 139.200 ;
        RECT 22.580 138.200 22.840 138.520 ;
        RECT 21.660 136.500 21.920 136.820 ;
        RECT 19.360 134.460 19.620 134.780 ;
        RECT 21.720 134.180 21.860 136.500 ;
        RECT 22.640 136.480 22.780 138.200 ;
        RECT 22.580 136.160 22.840 136.480 ;
        RECT 22.120 135.480 22.380 135.800 ;
        RECT 22.180 134.780 22.320 135.480 ;
        RECT 22.120 134.460 22.380 134.780 ;
        RECT 18.900 133.780 19.160 134.100 ;
        RECT 21.720 134.040 22.320 134.180 ;
        RECT 22.180 133.760 22.320 134.040 ;
        RECT 19.820 133.440 20.080 133.760 ;
        RECT 22.120 133.440 22.380 133.760 ;
        RECT 16.880 129.505 18.760 129.875 ;
        RECT 19.880 125.940 20.020 133.440 ;
        RECT 22.180 131.380 22.320 133.440 ;
        RECT 22.120 131.060 22.380 131.380 ;
        RECT 21.200 128.680 21.460 129.000 ;
        RECT 19.820 125.620 20.080 125.940 ;
        RECT 16.880 124.065 18.760 124.435 ;
        RECT 16.880 118.625 18.760 118.995 ;
        RECT 19.880 117.860 20.020 125.620 ;
        RECT 21.260 125.600 21.400 128.680 ;
        RECT 21.200 125.280 21.460 125.600 ;
        RECT 22.180 122.880 22.320 131.060 ;
        RECT 22.640 130.360 22.780 136.160 ;
        RECT 23.560 133.420 23.700 138.880 ;
        RECT 28.560 135.480 28.820 135.800 ;
        RECT 23.500 133.100 23.760 133.420 ;
        RECT 28.620 131.040 28.760 135.480 ;
        RECT 29.020 133.440 29.280 133.760 ;
        RECT 29.080 132.060 29.220 133.440 ;
        RECT 29.020 131.740 29.280 132.060 ;
        RECT 28.560 130.720 28.820 131.040 ;
        RECT 23.500 130.380 23.760 130.700 ;
        RECT 22.580 130.040 22.840 130.360 ;
        RECT 23.040 130.040 23.300 130.360 ;
        RECT 22.640 127.640 22.780 130.040 ;
        RECT 22.580 127.320 22.840 127.640 ;
        RECT 23.100 125.600 23.240 130.040 ;
        RECT 23.560 129.340 23.700 130.380 ;
        RECT 23.500 129.020 23.760 129.340 ;
        RECT 23.040 125.280 23.300 125.600 ;
        RECT 23.560 123.900 23.700 129.020 ;
        RECT 23.960 128.000 24.220 128.320 ;
        RECT 24.020 126.620 24.160 128.000 ;
        RECT 23.960 126.300 24.220 126.620 ;
        RECT 22.580 123.580 22.840 123.900 ;
        RECT 23.500 123.580 23.760 123.900 ;
        RECT 22.120 122.560 22.380 122.880 ;
        RECT 22.180 120.840 22.320 122.560 ;
        RECT 22.120 120.520 22.380 120.840 ;
        RECT 22.640 120.500 22.780 123.580 ;
        RECT 26.720 121.880 26.980 122.200 ;
        RECT 22.580 120.180 22.840 120.500 ;
        RECT 21.200 119.160 21.460 119.480 ;
        RECT 19.420 117.780 20.020 117.860 ;
        RECT 19.360 117.720 20.020 117.780 ;
        RECT 19.360 117.460 19.620 117.720 ;
        RECT 19.880 115.060 20.020 117.720 ;
        RECT 19.820 114.740 20.080 115.060 ;
        RECT 21.260 114.720 21.400 119.160 ;
        RECT 22.640 118.460 22.780 120.180 ;
        RECT 26.780 120.160 26.920 121.880 ;
        RECT 26.720 119.840 26.980 120.160 ;
        RECT 25.340 119.160 25.600 119.480 ;
        RECT 22.580 118.140 22.840 118.460 ;
        RECT 23.500 117.800 23.760 118.120 ;
        RECT 23.560 115.740 23.700 117.800 ;
        RECT 25.400 117.780 25.540 119.160 ;
        RECT 25.340 117.460 25.600 117.780 ;
        RECT 25.800 117.120 26.060 117.440 ;
        RECT 23.500 115.420 23.760 115.740 ;
        RECT 25.860 115.140 26.000 117.120 ;
        RECT 28.560 116.440 28.820 116.760 ;
        RECT 25.860 115.060 26.460 115.140 ;
        RECT 25.800 115.000 26.460 115.060 ;
        RECT 25.800 114.740 26.060 115.000 ;
        RECT 21.200 114.400 21.460 114.720 ;
        RECT 16.880 113.185 18.760 113.555 ;
        RECT 21.200 112.360 21.460 112.680 ;
        RECT 14.300 111.680 14.560 112.000 ;
        RECT 14.360 89.420 14.500 111.680 ;
        RECT 21.260 110.300 21.400 112.360 ;
        RECT 26.320 112.340 26.460 115.000 ;
        RECT 28.620 114.380 28.760 116.440 ;
        RECT 28.560 114.060 28.820 114.380 ;
        RECT 26.260 112.020 26.520 112.340 ;
        RECT 27.640 111.000 27.900 111.320 ;
        RECT 27.700 110.300 27.840 111.000 ;
        RECT 21.200 109.980 21.460 110.300 ;
        RECT 27.640 109.980 27.900 110.300 ;
        RECT 29.540 109.280 29.680 140.920 ;
        RECT 35.000 139.220 35.260 139.540 ;
        RECT 29.940 138.880 30.200 139.200 ;
        RECT 30.400 138.880 30.660 139.200 ;
        RECT 30.000 134.100 30.140 138.880 ;
        RECT 30.460 136.140 30.600 138.880 ;
        RECT 34.540 138.200 34.800 138.520 ;
        RECT 31.880 137.665 33.760 138.035 ;
        RECT 34.600 137.500 34.740 138.200 ;
        RECT 34.540 137.180 34.800 137.500 ;
        RECT 34.080 136.840 34.340 137.160 ;
        RECT 31.320 136.500 31.580 136.820 ;
        RECT 30.400 135.820 30.660 136.140 ;
        RECT 30.860 135.480 31.120 135.800 ;
        RECT 29.940 133.780 30.200 134.100 ;
        RECT 30.000 128.660 30.140 133.780 ;
        RECT 30.920 132.060 31.060 135.480 ;
        RECT 31.380 134.100 31.520 136.500 ;
        RECT 33.620 136.160 33.880 136.480 ;
        RECT 32.700 135.480 32.960 135.800 ;
        RECT 32.760 134.100 32.900 135.480 ;
        RECT 31.320 133.780 31.580 134.100 ;
        RECT 32.240 133.780 32.500 134.100 ;
        RECT 32.700 133.780 32.960 134.100 ;
        RECT 32.300 133.500 32.440 133.780 ;
        RECT 33.680 133.500 33.820 136.160 ;
        RECT 34.140 134.780 34.280 136.840 ;
        RECT 35.060 136.480 35.200 139.220 ;
        RECT 35.520 136.820 35.660 170.840 ;
        RECT 35.980 170.760 36.580 170.900 ;
        RECT 35.980 169.120 36.120 170.760 ;
        RECT 35.920 168.800 36.180 169.120 ;
        RECT 35.980 167.080 36.120 168.800 ;
        RECT 36.900 168.440 37.040 176.960 ;
        RECT 37.360 172.520 37.500 179.680 ;
        RECT 37.820 174.900 37.960 182.740 ;
        RECT 38.280 182.720 38.420 185.460 ;
        RECT 38.220 182.400 38.480 182.720 ;
        RECT 38.280 177.280 38.420 182.400 ;
        RECT 39.600 181.720 39.860 182.040 ;
        RECT 39.660 178.300 39.800 181.720 ;
        RECT 40.980 179.910 41.240 180.000 ;
        RECT 41.500 179.910 41.640 185.460 ;
        RECT 43.740 184.440 44.000 184.760 ;
        RECT 44.200 184.440 44.460 184.760 ;
        RECT 43.800 182.720 43.940 184.440 ;
        RECT 44.260 183.060 44.400 184.440 ;
        RECT 45.180 183.740 45.320 190.560 ;
        RECT 46.100 186.460 46.240 193.620 ;
        RECT 49.260 193.280 49.520 193.600 ;
        RECT 46.500 190.900 46.760 191.220 ;
        RECT 46.560 187.900 46.700 190.900 ;
        RECT 49.320 190.540 49.460 193.280 ;
        RECT 49.260 190.220 49.520 190.540 ;
        RECT 46.880 189.345 48.760 189.715 ;
        RECT 46.960 187.900 47.220 188.160 ;
        RECT 46.560 187.840 47.220 187.900 ;
        RECT 46.560 187.760 47.160 187.840 ;
        RECT 49.320 187.820 49.460 190.220 ;
        RECT 46.040 186.140 46.300 186.460 ;
        RECT 46.560 186.120 46.700 187.760 ;
        RECT 49.260 187.500 49.520 187.820 ;
        RECT 46.500 185.800 46.760 186.120 ;
        RECT 45.580 185.120 45.840 185.440 ;
        RECT 45.120 183.420 45.380 183.740 ;
        RECT 44.200 182.740 44.460 183.060 ;
        RECT 43.740 182.400 44.000 182.720 ;
        RECT 45.640 181.020 45.780 185.120 ;
        RECT 46.040 184.440 46.300 184.760 ;
        RECT 46.500 184.440 46.760 184.760 ;
        RECT 46.100 182.040 46.240 184.440 ;
        RECT 46.560 183.060 46.700 184.440 ;
        RECT 46.880 183.905 48.760 184.275 ;
        RECT 46.500 182.740 46.760 183.060 ;
        RECT 46.040 181.720 46.300 182.040 ;
        RECT 45.580 180.700 45.840 181.020 ;
        RECT 46.560 180.340 46.700 182.740 ;
        RECT 47.420 181.720 47.680 182.040 ;
        RECT 46.960 180.700 47.220 181.020 ;
        RECT 47.020 180.340 47.160 180.700 ;
        RECT 47.480 180.340 47.620 181.720 ;
        RECT 46.500 180.020 46.760 180.340 ;
        RECT 46.960 180.020 47.220 180.340 ;
        RECT 47.420 180.020 47.680 180.340 ;
        RECT 40.510 179.485 40.790 179.855 ;
        RECT 40.980 179.770 41.640 179.910 ;
        RECT 40.980 179.680 41.240 179.770 ;
        RECT 41.890 179.485 42.170 179.855 ;
        RECT 44.200 179.680 44.460 180.000 ;
        RECT 45.580 179.680 45.840 180.000 ;
        RECT 40.580 179.320 40.720 179.485 ;
        RECT 40.060 179.000 40.320 179.320 ;
        RECT 40.520 179.000 40.780 179.320 ;
        RECT 40.980 179.000 41.240 179.320 ;
        RECT 39.600 177.980 39.860 178.300 ;
        RECT 38.220 176.960 38.480 177.280 ;
        RECT 38.280 175.580 38.420 176.960 ;
        RECT 38.220 175.260 38.480 175.580 ;
        RECT 40.120 175.095 40.260 179.000 ;
        RECT 41.040 175.580 41.180 179.000 ;
        RECT 40.980 175.260 41.240 175.580 ;
        RECT 37.760 174.580 38.020 174.900 ;
        RECT 40.050 174.725 40.330 175.095 ;
        RECT 40.520 174.920 40.780 175.240 ;
        RECT 40.120 174.560 40.260 174.725 ;
        RECT 38.220 174.240 38.480 174.560 ;
        RECT 40.060 174.240 40.320 174.560 ;
        RECT 37.300 172.200 37.560 172.520 ;
        RECT 38.280 172.180 38.420 174.240 ;
        RECT 39.140 173.900 39.400 174.220 ;
        RECT 39.600 173.900 39.860 174.220 ;
        RECT 38.220 171.860 38.480 172.180 ;
        RECT 36.840 168.120 37.100 168.440 ;
        RECT 35.920 166.760 36.180 167.080 ;
        RECT 36.900 166.740 37.040 168.120 ;
        RECT 36.840 166.420 37.100 166.740 ;
        RECT 36.900 164.020 37.040 166.420 ;
        RECT 38.220 165.400 38.480 165.720 ;
        RECT 36.840 163.700 37.100 164.020 ;
        RECT 38.280 163.680 38.420 165.400 ;
        RECT 38.220 163.360 38.480 163.680 ;
        RECT 35.920 162.680 36.180 163.000 ;
        RECT 36.380 162.680 36.640 163.000 ;
        RECT 35.980 158.240 36.120 162.680 ;
        RECT 36.440 161.640 36.580 162.680 ;
        RECT 36.380 161.320 36.640 161.640 ;
        RECT 35.920 157.920 36.180 158.240 ;
        RECT 36.440 157.900 36.580 161.320 ;
        RECT 37.760 160.300 38.020 160.620 ;
        RECT 36.380 157.580 36.640 157.900 ;
        RECT 35.920 154.520 36.180 154.840 ;
        RECT 35.980 150.420 36.120 154.520 ;
        RECT 37.820 153.140 37.960 160.300 ;
        RECT 37.300 152.820 37.560 153.140 ;
        RECT 37.760 152.820 38.020 153.140 ;
        RECT 36.840 152.710 37.100 152.800 ;
        RECT 36.440 152.570 37.100 152.710 ;
        RECT 35.920 150.100 36.180 150.420 ;
        RECT 36.440 150.080 36.580 152.570 ;
        RECT 36.840 152.480 37.100 152.570 ;
        RECT 37.360 151.100 37.500 152.820 ;
        RECT 37.300 150.780 37.560 151.100 ;
        RECT 36.380 149.760 36.640 150.080 ;
        RECT 35.920 148.060 36.180 148.380 ;
        RECT 35.980 147.360 36.120 148.060 ;
        RECT 35.920 147.040 36.180 147.360 ;
        RECT 36.440 144.640 36.580 149.760 ;
        RECT 36.840 146.360 37.100 146.680 ;
        RECT 38.680 146.360 38.940 146.680 ;
        RECT 36.380 144.320 36.640 144.640 ;
        RECT 35.920 142.620 36.180 142.940 ;
        RECT 35.980 140.220 36.120 142.620 ;
        RECT 35.920 139.900 36.180 140.220 ;
        RECT 35.920 139.220 36.180 139.540 ;
        RECT 35.460 136.500 35.720 136.820 ;
        RECT 35.000 136.160 35.260 136.480 ;
        RECT 34.540 135.480 34.800 135.800 ;
        RECT 34.080 134.460 34.340 134.780 ;
        RECT 32.300 133.360 34.280 133.500 ;
        RECT 31.320 132.760 31.580 133.080 ;
        RECT 30.860 131.740 31.120 132.060 ;
        RECT 29.940 128.340 30.200 128.660 ;
        RECT 30.400 128.340 30.660 128.660 ;
        RECT 30.460 125.940 30.600 128.340 ;
        RECT 30.400 125.620 30.660 125.940 ;
        RECT 30.860 119.500 31.120 119.820 ;
        RECT 30.920 115.740 31.060 119.500 ;
        RECT 30.860 115.420 31.120 115.740 ;
        RECT 31.380 109.620 31.520 132.760 ;
        RECT 31.880 132.225 33.760 132.595 ;
        RECT 34.140 132.060 34.280 133.360 ;
        RECT 34.080 131.740 34.340 132.060 ;
        RECT 34.080 130.380 34.340 130.700 ;
        RECT 34.140 129.340 34.280 130.380 ;
        RECT 34.080 129.020 34.340 129.340 ;
        RECT 31.880 126.785 33.760 127.155 ;
        RECT 31.880 121.345 33.760 121.715 ;
        RECT 31.880 115.905 33.760 116.275 ;
        RECT 31.880 110.465 33.760 110.835 ;
        RECT 31.320 109.300 31.580 109.620 ;
        RECT 34.600 109.280 34.740 135.480 ;
        RECT 35.000 133.100 35.260 133.420 ;
        RECT 35.060 123.220 35.200 133.100 ;
        RECT 35.980 133.080 36.120 139.220 ;
        RECT 36.440 134.440 36.580 144.320 ;
        RECT 36.900 136.480 37.040 146.360 ;
        RECT 38.220 137.180 38.480 137.500 ;
        RECT 36.840 136.160 37.100 136.480 ;
        RECT 36.380 134.120 36.640 134.440 ;
        RECT 35.920 132.760 36.180 133.080 ;
        RECT 36.440 131.380 36.580 134.120 ;
        RECT 36.380 131.060 36.640 131.380 ;
        RECT 37.760 131.060 38.020 131.380 ;
        RECT 37.820 129.340 37.960 131.060 ;
        RECT 37.760 129.020 38.020 129.340 ;
        RECT 35.920 125.620 36.180 125.940 ;
        RECT 35.000 122.900 35.260 123.220 ;
        RECT 35.060 121.180 35.200 122.900 ;
        RECT 35.000 120.860 35.260 121.180 ;
        RECT 35.980 120.500 36.120 125.620 ;
        RECT 38.280 125.600 38.420 137.180 ;
        RECT 38.740 136.480 38.880 146.360 ;
        RECT 39.200 136.820 39.340 173.900 ;
        RECT 39.660 172.180 39.800 173.900 ;
        RECT 39.600 171.860 39.860 172.180 ;
        RECT 40.060 154.520 40.320 154.840 ;
        RECT 39.600 141.260 39.860 141.580 ;
        RECT 39.660 140.220 39.800 141.260 ;
        RECT 39.600 139.900 39.860 140.220 ;
        RECT 40.120 139.200 40.260 154.520 ;
        RECT 40.060 138.880 40.320 139.200 ;
        RECT 39.140 136.500 39.400 136.820 ;
        RECT 38.680 136.160 38.940 136.480 ;
        RECT 38.680 135.480 38.940 135.800 ;
        RECT 36.840 125.280 37.100 125.600 ;
        RECT 38.220 125.280 38.480 125.600 ;
        RECT 36.900 122.880 37.040 125.280 ;
        RECT 36.840 122.790 37.100 122.880 ;
        RECT 36.440 122.650 37.100 122.790 ;
        RECT 35.920 120.180 36.180 120.500 ;
        RECT 35.000 119.500 35.260 119.820 ;
        RECT 35.060 113.020 35.200 119.500 ;
        RECT 36.440 118.460 36.580 122.650 ;
        RECT 36.840 122.560 37.100 122.650 ;
        RECT 36.840 121.880 37.100 122.200 ;
        RECT 36.380 118.140 36.640 118.460 ;
        RECT 35.460 117.800 35.720 118.120 ;
        RECT 35.520 115.740 35.660 117.800 ;
        RECT 35.460 115.420 35.720 115.740 ;
        RECT 36.900 114.720 37.040 121.880 ;
        RECT 37.760 119.840 38.020 120.160 ;
        RECT 37.820 115.740 37.960 119.840 ;
        RECT 37.760 115.420 38.020 115.740 ;
        RECT 35.920 114.400 36.180 114.720 ;
        RECT 36.840 114.400 37.100 114.720 ;
        RECT 35.980 114.040 36.120 114.400 ;
        RECT 35.920 113.720 36.180 114.040 ;
        RECT 35.000 112.700 35.260 113.020 ;
        RECT 35.980 112.340 36.120 113.720 ;
        RECT 35.920 112.020 36.180 112.340 ;
        RECT 36.840 111.340 37.100 111.660 ;
        RECT 29.480 108.960 29.740 109.280 ;
        RECT 34.540 108.960 34.800 109.280 ;
        RECT 27.640 108.620 27.900 108.940 ;
        RECT 23.500 108.280 23.760 108.600 ;
        RECT 16.880 107.745 18.760 108.115 ;
        RECT 23.560 107.240 23.700 108.280 ;
        RECT 23.500 106.920 23.760 107.240 ;
        RECT 18.900 106.240 19.160 106.560 ;
        RECT 16.880 102.305 18.760 102.675 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 18.960 88.620 19.100 106.240 ;
        RECT 27.700 103.840 27.840 108.620 ;
        RECT 31.780 108.280 32.040 108.600 ;
        RECT 32.240 108.280 32.500 108.600 ;
        RECT 34.080 108.280 34.340 108.600 ;
        RECT 31.840 107.240 31.980 108.280 ;
        RECT 32.300 107.580 32.440 108.280 ;
        RECT 32.240 107.260 32.500 107.580 ;
        RECT 31.780 106.920 32.040 107.240 ;
        RECT 29.020 106.240 29.280 106.560 ;
        RECT 30.400 106.240 30.660 106.560 ;
        RECT 29.080 104.860 29.220 106.240 ;
        RECT 29.020 104.540 29.280 104.860 ;
        RECT 27.640 103.520 27.900 103.840 ;
        RECT 28.100 102.840 28.360 103.160 ;
        RECT 28.160 101.460 28.300 102.840 ;
        RECT 28.100 101.140 28.360 101.460 ;
        RECT 26.260 100.800 26.520 101.120 ;
        RECT 19.910 88.620 21.130 89.850 ;
        RECT 26.320 89.170 26.460 100.800 ;
        RECT 26.250 88.990 26.530 89.170 ;
        RECT 18.960 88.480 21.130 88.620 ;
        RECT 19.910 85.980 21.130 88.480 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 30.460 88.620 30.600 106.240 ;
        RECT 31.880 105.025 33.760 105.395 ;
        RECT 34.140 101.800 34.280 108.280 ;
        RECT 36.900 106.900 37.040 111.340 ;
        RECT 38.740 106.900 38.880 135.480 ;
        RECT 40.580 134.100 40.720 174.920 ;
        RECT 41.040 172.180 41.180 175.260 ;
        RECT 41.960 174.220 42.100 179.485 ;
        RECT 42.360 179.000 42.620 179.320 ;
        RECT 41.900 173.900 42.160 174.220 ;
        RECT 40.980 171.860 41.240 172.180 ;
        RECT 41.040 169.800 41.180 171.860 ;
        RECT 41.440 170.840 41.700 171.160 ;
        RECT 40.980 169.480 41.240 169.800 ;
        RECT 41.040 156.200 41.180 169.480 ;
        RECT 40.980 155.880 41.240 156.200 ;
        RECT 40.980 149.080 41.240 149.400 ;
        RECT 41.040 134.100 41.180 149.080 ;
        RECT 41.500 139.880 41.640 170.840 ;
        RECT 42.420 160.140 42.560 179.000 ;
        RECT 43.740 177.300 44.000 177.620 ;
        RECT 42.820 176.280 43.080 176.600 ;
        RECT 42.880 172.180 43.020 176.280 ;
        RECT 43.800 174.560 43.940 177.300 ;
        RECT 44.260 174.560 44.400 179.680 ;
        RECT 44.660 179.000 44.920 179.320 ;
        RECT 44.720 174.560 44.860 179.000 ;
        RECT 45.640 177.620 45.780 179.680 ;
        RECT 47.020 179.570 47.160 180.020 ;
        RECT 46.560 179.430 47.160 179.570 ;
        RECT 46.040 179.000 46.300 179.320 ;
        RECT 46.100 178.300 46.240 179.000 ;
        RECT 46.040 177.980 46.300 178.300 ;
        RECT 45.580 177.300 45.840 177.620 ;
        RECT 45.640 174.900 45.780 177.300 ;
        RECT 46.560 175.580 46.700 179.430 ;
        RECT 46.880 178.465 48.760 178.835 ;
        RECT 47.880 177.300 48.140 177.620 ;
        RECT 49.260 177.300 49.520 177.620 ;
        RECT 46.500 175.260 46.760 175.580 ;
        RECT 45.580 174.580 45.840 174.900 ;
        RECT 43.740 174.240 44.000 174.560 ;
        RECT 44.200 174.240 44.460 174.560 ;
        RECT 44.660 174.240 44.920 174.560 ;
        RECT 44.720 172.860 44.860 174.240 ;
        RECT 47.940 174.220 48.080 177.300 ;
        RECT 45.580 173.900 45.840 174.220 ;
        RECT 47.880 173.900 48.140 174.220 ;
        RECT 44.660 172.540 44.920 172.860 ;
        RECT 42.820 171.860 43.080 172.180 ;
        RECT 44.190 169.285 44.470 169.655 ;
        RECT 44.260 169.120 44.400 169.285 ;
        RECT 44.200 168.800 44.460 169.120 ;
        RECT 43.280 166.080 43.540 166.400 ;
        RECT 42.820 165.400 43.080 165.720 ;
        RECT 42.880 161.980 43.020 165.400 ;
        RECT 42.820 161.660 43.080 161.980 ;
        RECT 42.420 160.000 43.020 160.140 ;
        RECT 41.900 157.920 42.160 158.240 ;
        RECT 41.960 156.540 42.100 157.920 ;
        RECT 42.360 157.240 42.620 157.560 ;
        RECT 41.900 156.220 42.160 156.540 ;
        RECT 41.890 155.685 42.170 156.055 ;
        RECT 41.900 155.540 42.160 155.685 ;
        RECT 41.900 151.800 42.160 152.120 ;
        RECT 41.960 150.420 42.100 151.800 ;
        RECT 41.900 150.100 42.160 150.420 ;
        RECT 41.960 146.680 42.100 150.100 ;
        RECT 41.900 146.360 42.160 146.680 ;
        RECT 41.440 139.560 41.700 139.880 ;
        RECT 42.420 136.480 42.560 157.240 ;
        RECT 42.360 136.160 42.620 136.480 ;
        RECT 42.880 134.100 43.020 160.000 ;
        RECT 43.340 158.240 43.480 166.080 ;
        RECT 43.280 157.920 43.540 158.240 ;
        RECT 45.120 157.920 45.380 158.240 ;
        RECT 43.280 157.240 43.540 157.560 ;
        RECT 43.340 156.055 43.480 157.240 ;
        RECT 45.180 156.540 45.320 157.920 ;
        RECT 45.120 156.220 45.380 156.540 ;
        RECT 43.270 155.685 43.550 156.055 ;
        RECT 43.340 155.430 43.480 155.685 ;
        RECT 43.740 155.430 44.000 155.520 ;
        RECT 43.340 155.290 44.000 155.430 ;
        RECT 43.740 155.200 44.000 155.290 ;
        RECT 43.740 154.520 44.000 154.840 ;
        RECT 45.120 154.520 45.380 154.840 ;
        RECT 43.280 152.140 43.540 152.460 ;
        RECT 43.340 150.420 43.480 152.140 ;
        RECT 43.280 150.100 43.540 150.420 ;
        RECT 43.340 147.020 43.480 150.100 ;
        RECT 43.280 146.700 43.540 147.020 ;
        RECT 43.800 134.100 43.940 154.520 ;
        RECT 44.660 152.655 44.920 152.800 ;
        RECT 44.650 152.285 44.930 152.655 ;
        RECT 44.200 149.080 44.460 149.400 ;
        RECT 40.520 133.780 40.780 134.100 ;
        RECT 40.980 133.780 41.240 134.100 ;
        RECT 42.820 133.780 43.080 134.100 ;
        RECT 43.740 133.780 44.000 134.100 ;
        RECT 44.260 133.500 44.400 149.080 ;
        RECT 44.720 147.360 44.860 152.285 ;
        RECT 45.180 150.420 45.320 154.520 ;
        RECT 45.120 150.100 45.380 150.420 ;
        RECT 44.660 147.040 44.920 147.360 ;
        RECT 45.120 142.280 45.380 142.600 ;
        RECT 44.660 137.180 44.920 137.500 ;
        RECT 43.800 133.360 44.400 133.500 ;
        RECT 39.600 132.760 39.860 133.080 ;
        RECT 40.520 132.760 40.780 133.080 ;
        RECT 41.440 132.760 41.700 133.080 ;
        RECT 43.280 132.760 43.540 133.080 ;
        RECT 39.660 128.660 39.800 132.760 ;
        RECT 40.060 131.400 40.320 131.720 ;
        RECT 39.600 128.340 39.860 128.660 ;
        RECT 40.120 125.260 40.260 131.400 ;
        RECT 40.580 125.600 40.720 132.760 ;
        RECT 40.520 125.280 40.780 125.600 ;
        RECT 40.060 124.940 40.320 125.260 ;
        RECT 40.060 119.160 40.320 119.480 ;
        RECT 39.140 117.120 39.400 117.440 ;
        RECT 39.200 115.740 39.340 117.120 ;
        RECT 39.140 115.420 39.400 115.740 ;
        RECT 40.120 114.720 40.260 119.160 ;
        RECT 40.060 114.400 40.320 114.720 ;
        RECT 40.980 108.620 41.240 108.940 ;
        RECT 41.040 107.240 41.180 108.620 ;
        RECT 40.980 106.920 41.240 107.240 ;
        RECT 41.500 106.900 41.640 132.760 ;
        RECT 42.820 130.040 43.080 130.360 ;
        RECT 42.880 129.000 43.020 130.040 ;
        RECT 42.820 128.680 43.080 129.000 ;
        RECT 42.820 128.000 43.080 128.320 ;
        RECT 42.360 125.280 42.620 125.600 ;
        RECT 41.900 122.560 42.160 122.880 ;
        RECT 41.960 120.160 42.100 122.560 ;
        RECT 41.900 119.840 42.160 120.160 ;
        RECT 42.420 119.480 42.560 125.280 ;
        RECT 42.880 123.900 43.020 128.000 ;
        RECT 43.340 125.260 43.480 132.760 ;
        RECT 43.800 129.340 43.940 133.360 ;
        RECT 44.200 132.760 44.460 133.080 ;
        RECT 43.740 129.020 44.000 129.340 ;
        RECT 43.280 124.940 43.540 125.260 ;
        RECT 42.820 123.580 43.080 123.900 ;
        RECT 43.740 122.220 44.000 122.540 ;
        RECT 43.800 120.500 43.940 122.220 ;
        RECT 43.740 120.180 44.000 120.500 ;
        RECT 42.360 119.160 42.620 119.480 ;
        RECT 42.420 118.460 42.560 119.160 ;
        RECT 42.360 118.140 42.620 118.460 ;
        RECT 42.420 114.380 42.560 118.140 ;
        RECT 43.280 117.800 43.540 118.120 ;
        RECT 43.340 115.740 43.480 117.800 ;
        RECT 43.280 115.420 43.540 115.740 ;
        RECT 43.800 115.400 43.940 120.180 ;
        RECT 43.740 115.080 44.000 115.400 ;
        RECT 42.360 114.060 42.620 114.380 ;
        RECT 44.260 111.840 44.400 132.760 ;
        RECT 44.720 125.600 44.860 137.180 ;
        RECT 45.180 129.340 45.320 142.280 ;
        RECT 45.640 136.820 45.780 173.900 ;
        RECT 46.880 173.025 48.760 173.395 ;
        RECT 49.320 172.860 49.460 177.300 ;
        RECT 49.780 172.860 49.920 194.390 ;
        RECT 50.640 194.300 50.900 194.390 ;
        RECT 53.460 194.280 53.600 195.320 ;
        RECT 53.400 193.960 53.660 194.280 ;
        RECT 50.640 193.280 50.900 193.600 ;
        RECT 50.700 191.900 50.840 193.280 ;
        RECT 54.320 192.600 54.580 192.920 ;
        RECT 50.640 191.580 50.900 191.900 ;
        RECT 52.480 190.900 52.740 191.220 ;
        RECT 50.180 187.160 50.440 187.480 ;
        RECT 50.240 183.740 50.380 187.160 ;
        RECT 50.180 183.420 50.440 183.740 ;
        RECT 50.180 182.400 50.440 182.720 ;
        RECT 50.240 181.020 50.380 182.400 ;
        RECT 50.180 180.700 50.440 181.020 ;
        RECT 52.540 180.340 52.680 190.900 ;
        RECT 54.380 190.880 54.520 192.600 ;
        RECT 54.320 190.560 54.580 190.880 ;
        RECT 58.060 190.200 58.200 195.320 ;
        RECT 61.880 192.065 63.760 192.435 ;
        RECT 64.040 191.560 64.180 202.460 ;
        RECT 64.960 201.420 65.100 203.480 ;
        RECT 64.900 201.100 65.160 201.420 ;
        RECT 64.900 198.040 65.160 198.360 ;
        RECT 63.980 191.240 64.240 191.560 ;
        RECT 59.380 190.900 59.640 191.220 ;
        RECT 58.000 189.880 58.260 190.200 ;
        RECT 58.060 189.180 58.200 189.880 ;
        RECT 58.000 188.860 58.260 189.180 ;
        RECT 55.700 188.180 55.960 188.500 ;
        RECT 56.620 188.180 56.880 188.500 ;
        RECT 55.760 188.015 55.900 188.180 ;
        RECT 55.690 187.645 55.970 188.015 ;
        RECT 56.160 181.720 56.420 182.040 ;
        RECT 52.480 180.020 52.740 180.340 ;
        RECT 54.320 180.020 54.580 180.340 ;
        RECT 50.640 179.000 50.900 179.320 ;
        RECT 50.700 177.620 50.840 179.000 ;
        RECT 52.540 177.960 52.680 180.020 ;
        RECT 53.860 179.340 54.120 179.660 ;
        RECT 53.920 178.300 54.060 179.340 ;
        RECT 53.860 177.980 54.120 178.300 ;
        RECT 52.480 177.640 52.740 177.960 ;
        RECT 50.640 177.300 50.900 177.620 ;
        RECT 51.100 176.620 51.360 176.940 ;
        RECT 50.180 176.280 50.440 176.600 ;
        RECT 49.260 172.540 49.520 172.860 ;
        RECT 49.720 172.540 49.980 172.860 ;
        RECT 49.320 172.180 49.460 172.540 ;
        RECT 47.420 171.860 47.680 172.180 ;
        RECT 49.260 171.860 49.520 172.180 ;
        RECT 49.720 171.860 49.980 172.180 ;
        RECT 46.040 170.840 46.300 171.160 ;
        RECT 46.100 160.140 46.240 170.840 ;
        RECT 47.480 170.140 47.620 171.860 ;
        RECT 49.780 171.500 49.920 171.860 ;
        RECT 49.720 171.180 49.980 171.500 ;
        RECT 47.420 169.820 47.680 170.140 ;
        RECT 46.880 167.585 48.760 167.955 ;
        RECT 49.720 165.400 49.980 165.720 ;
        RECT 49.260 163.360 49.520 163.680 ;
        RECT 46.500 163.020 46.760 163.340 ;
        RECT 46.560 161.980 46.700 163.020 ;
        RECT 46.880 162.145 48.760 162.515 ;
        RECT 49.320 161.980 49.460 163.360 ;
        RECT 49.780 161.980 49.920 165.400 ;
        RECT 46.500 161.660 46.760 161.980 ;
        RECT 49.260 161.660 49.520 161.980 ;
        RECT 49.720 161.660 49.980 161.980 ;
        RECT 49.720 160.980 49.980 161.300 ;
        RECT 49.260 160.640 49.520 160.960 ;
        RECT 46.100 160.000 46.700 160.140 ;
        RECT 46.040 157.240 46.300 157.560 ;
        RECT 46.100 141.920 46.240 157.240 ;
        RECT 46.560 142.260 46.700 160.000 ;
        RECT 46.880 156.705 48.760 157.075 ;
        RECT 49.320 156.540 49.460 160.640 ;
        RECT 49.780 159.260 49.920 160.980 ;
        RECT 49.720 158.940 49.980 159.260 ;
        RECT 50.240 157.980 50.380 176.280 ;
        RECT 51.160 172.860 51.300 176.620 ;
        RECT 54.380 175.580 54.520 180.020 ;
        RECT 56.220 177.960 56.360 181.720 ;
        RECT 56.680 180.680 56.820 188.180 ;
        RECT 59.440 187.820 59.580 190.900 ;
        RECT 60.300 190.220 60.560 190.540 ;
        RECT 60.360 189.180 60.500 190.220 ;
        RECT 62.140 189.880 62.400 190.200 ;
        RECT 60.300 188.860 60.560 189.180 ;
        RECT 62.200 188.160 62.340 189.880 ;
        RECT 62.140 187.840 62.400 188.160 ;
        RECT 59.380 187.500 59.640 187.820 ;
        RECT 59.440 185.780 59.580 187.500 ;
        RECT 64.960 187.220 65.100 198.040 ;
        RECT 66.340 193.940 66.480 204.500 ;
        RECT 73.240 203.800 73.380 206.880 ;
        RECT 73.180 203.480 73.440 203.800 ;
        RECT 66.740 202.460 67.000 202.780 ;
        RECT 66.280 193.620 66.540 193.940 ;
        RECT 65.820 192.600 66.080 192.920 ;
        RECT 65.880 190.540 66.020 192.600 ;
        RECT 65.820 190.220 66.080 190.540 ;
        RECT 66.340 190.200 66.480 193.620 ;
        RECT 66.280 189.880 66.540 190.200 ;
        RECT 65.820 187.840 66.080 188.160 ;
        RECT 64.500 187.080 65.100 187.220 ;
        RECT 61.880 186.625 63.760 186.995 ;
        RECT 60.760 185.800 61.020 186.120 ;
        RECT 59.380 185.460 59.640 185.780 ;
        RECT 58.000 184.780 58.260 185.100 ;
        RECT 58.060 183.740 58.200 184.780 ;
        RECT 58.000 183.420 58.260 183.740 ;
        RECT 59.440 183.060 59.580 185.460 ;
        RECT 60.820 183.060 60.960 185.800 ;
        RECT 59.380 182.740 59.640 183.060 ;
        RECT 60.760 182.740 61.020 183.060 ;
        RECT 56.620 180.360 56.880 180.680 ;
        RECT 56.160 177.640 56.420 177.960 ;
        RECT 54.320 175.260 54.580 175.580 ;
        RECT 54.380 174.900 54.520 175.260 ;
        RECT 53.860 174.580 54.120 174.900 ;
        RECT 54.320 174.580 54.580 174.900 ;
        RECT 53.400 173.900 53.660 174.220 ;
        RECT 51.100 172.540 51.360 172.860 ;
        RECT 51.160 172.180 51.300 172.540 ;
        RECT 53.460 172.180 53.600 173.900 ;
        RECT 53.920 172.180 54.060 174.580 ;
        RECT 56.680 174.560 56.820 180.360 ;
        RECT 58.000 179.000 58.260 179.320 ;
        RECT 58.060 174.900 58.200 179.000 ;
        RECT 59.440 177.280 59.580 182.740 ;
        RECT 59.380 176.960 59.640 177.280 ;
        RECT 58.000 174.580 58.260 174.900 ;
        RECT 54.770 174.045 55.050 174.415 ;
        RECT 56.620 174.240 56.880 174.560 ;
        RECT 54.840 172.860 54.980 174.045 ;
        RECT 57.080 173.560 57.340 173.880 ;
        RECT 54.780 172.540 55.040 172.860 ;
        RECT 54.840 172.180 54.980 172.540 ;
        RECT 57.140 172.520 57.280 173.560 ;
        RECT 57.080 172.200 57.340 172.520 ;
        RECT 60.820 172.180 60.960 182.740 ;
        RECT 61.880 181.185 63.760 181.555 ;
        RECT 61.280 178.300 62.340 178.380 ;
        RECT 61.280 178.240 62.400 178.300 ;
        RECT 61.280 177.960 61.420 178.240 ;
        RECT 62.140 177.980 62.400 178.240 ;
        RECT 61.220 177.640 61.480 177.960 ;
        RECT 63.980 176.960 64.240 177.280 ;
        RECT 61.880 175.745 63.760 176.115 ;
        RECT 64.040 175.580 64.180 176.960 ;
        RECT 63.980 175.260 64.240 175.580 ;
        RECT 61.220 173.900 61.480 174.220 ;
        RECT 63.050 174.045 63.330 174.415 ;
        RECT 61.280 172.860 61.420 173.900 ;
        RECT 63.120 173.880 63.260 174.045 ;
        RECT 63.060 173.560 63.320 173.880 ;
        RECT 61.220 172.540 61.480 172.860 ;
        RECT 51.100 171.860 51.360 172.180 ;
        RECT 53.400 171.860 53.660 172.180 ;
        RECT 53.860 171.860 54.120 172.180 ;
        RECT 54.780 171.860 55.040 172.180 ;
        RECT 60.760 171.860 61.020 172.180 ;
        RECT 52.480 170.840 52.740 171.160 ;
        RECT 51.100 166.760 51.360 167.080 ;
        RECT 51.160 164.700 51.300 166.760 ;
        RECT 51.100 164.380 51.360 164.700 ;
        RECT 50.640 158.940 50.900 159.260 ;
        RECT 50.700 158.580 50.840 158.940 ;
        RECT 50.640 158.260 50.900 158.580 ;
        RECT 49.780 157.840 50.380 157.980 ;
        RECT 49.260 156.220 49.520 156.540 ;
        RECT 46.960 155.540 47.220 155.860 ;
        RECT 47.020 155.180 47.160 155.540 ;
        RECT 46.960 154.860 47.220 155.180 ;
        RECT 49.260 154.520 49.520 154.840 ;
        RECT 46.880 151.265 48.760 151.635 ;
        RECT 49.320 150.500 49.460 154.520 ;
        RECT 48.860 150.360 49.460 150.500 ;
        RECT 49.780 150.420 49.920 157.840 ;
        RECT 50.180 157.240 50.440 157.560 ;
        RECT 50.240 150.420 50.380 157.240 ;
        RECT 50.640 156.220 50.900 156.540 ;
        RECT 50.700 152.120 50.840 156.220 ;
        RECT 51.100 152.480 51.360 152.800 ;
        RECT 50.640 151.800 50.900 152.120 ;
        RECT 48.860 147.360 49.000 150.360 ;
        RECT 49.720 150.100 49.980 150.420 ;
        RECT 50.180 150.100 50.440 150.420 ;
        RECT 50.640 149.760 50.900 150.080 ;
        RECT 50.700 148.380 50.840 149.760 ;
        RECT 49.260 148.060 49.520 148.380 ;
        RECT 50.640 148.060 50.900 148.380 ;
        RECT 48.800 147.040 49.060 147.360 ;
        RECT 46.880 145.825 48.760 146.195 ;
        RECT 49.320 144.380 49.460 148.060 ;
        RECT 49.720 146.360 49.980 146.680 ;
        RECT 49.780 144.980 49.920 146.360 ;
        RECT 51.160 145.660 51.300 152.480 ;
        RECT 51.560 149.080 51.820 149.400 ;
        RECT 51.620 147.020 51.760 149.080 ;
        RECT 52.540 147.700 52.680 170.840 ;
        RECT 53.400 166.760 53.660 167.080 ;
        RECT 53.460 163.680 53.600 166.760 ;
        RECT 54.320 166.080 54.580 166.400 ;
        RECT 54.780 166.080 55.040 166.400 ;
        RECT 57.540 166.080 57.800 166.400 ;
        RECT 53.400 163.360 53.660 163.680 ;
        RECT 52.940 162.680 53.200 163.000 ;
        RECT 53.000 159.260 53.140 162.680 ;
        RECT 54.380 161.980 54.520 166.080 ;
        RECT 54.840 164.700 54.980 166.080 ;
        RECT 54.780 164.380 55.040 164.700 ;
        RECT 57.600 164.360 57.740 166.080 ;
        RECT 58.920 165.400 59.180 165.720 ;
        RECT 57.540 164.040 57.800 164.360 ;
        RECT 58.980 163.340 59.120 165.400 ;
        RECT 60.820 164.020 60.960 171.860 ;
        RECT 61.880 170.305 63.760 170.675 ;
        RECT 61.680 166.420 61.940 166.740 ;
        RECT 61.740 166.140 61.880 166.420 ;
        RECT 61.280 166.000 61.880 166.140 ;
        RECT 63.980 166.080 64.240 166.400 ;
        RECT 61.280 164.100 61.420 166.000 ;
        RECT 61.880 164.865 63.760 165.235 ;
        RECT 61.680 164.380 61.940 164.700 ;
        RECT 61.740 164.100 61.880 164.380 ;
        RECT 60.760 163.700 61.020 164.020 ;
        RECT 61.280 163.960 61.880 164.100 ;
        RECT 58.920 163.020 59.180 163.340 ;
        RECT 54.320 161.660 54.580 161.980 ;
        RECT 53.400 160.300 53.660 160.620 ;
        RECT 52.940 158.940 53.200 159.260 ;
        RECT 53.000 158.240 53.140 158.940 ;
        RECT 52.940 157.920 53.200 158.240 ;
        RECT 53.460 157.560 53.600 160.300 ;
        RECT 53.860 157.920 54.120 158.240 ;
        RECT 57.080 157.920 57.340 158.240 ;
        RECT 61.280 158.150 61.420 163.960 ;
        RECT 64.040 163.680 64.180 166.080 ;
        RECT 63.980 163.360 64.240 163.680 ;
        RECT 62.600 163.020 62.860 163.340 ;
        RECT 62.660 161.980 62.800 163.020 ;
        RECT 62.600 161.660 62.860 161.980 ;
        RECT 61.880 159.425 63.760 159.795 ;
        RECT 63.060 158.150 63.320 158.240 ;
        RECT 61.280 158.010 63.320 158.150 ;
        RECT 63.060 157.920 63.320 158.010 ;
        RECT 53.400 157.240 53.660 157.560 ;
        RECT 53.460 156.200 53.600 157.240 ;
        RECT 53.400 155.880 53.660 156.200 ;
        RECT 53.920 155.860 54.060 157.920 ;
        RECT 53.860 155.540 54.120 155.860 ;
        RECT 53.860 154.520 54.120 154.840 ;
        RECT 54.320 154.520 54.580 154.840 ;
        RECT 53.920 150.420 54.060 154.520 ;
        RECT 54.380 153.480 54.520 154.520 ;
        RECT 54.320 153.160 54.580 153.480 ;
        RECT 57.140 152.800 57.280 157.920 ;
        RECT 58.920 157.240 59.180 157.560 ;
        RECT 58.980 156.200 59.120 157.240 ;
        RECT 58.920 155.880 59.180 156.200 ;
        RECT 64.040 155.860 64.180 163.360 ;
        RECT 63.980 155.540 64.240 155.860 ;
        RECT 61.220 155.200 61.480 155.520 ;
        RECT 57.080 152.480 57.340 152.800 ;
        RECT 58.920 151.800 59.180 152.120 ;
        RECT 58.980 150.420 59.120 151.800 ;
        RECT 61.280 151.100 61.420 155.200 ;
        RECT 61.880 153.985 63.760 154.355 ;
        RECT 64.500 153.140 64.640 187.080 ;
        RECT 65.880 180.000 66.020 187.840 ;
        RECT 65.820 179.680 66.080 180.000 ;
        RECT 66.280 179.000 66.540 179.320 ;
        RECT 66.340 177.815 66.480 179.000 ;
        RECT 66.270 177.445 66.550 177.815 ;
        RECT 65.360 176.620 65.620 176.940 ;
        RECT 64.900 176.280 65.160 176.600 ;
        RECT 64.960 174.900 65.100 176.280 ;
        RECT 65.420 175.095 65.560 176.620 ;
        RECT 66.280 175.260 66.540 175.580 ;
        RECT 64.900 174.580 65.160 174.900 ;
        RECT 65.350 174.725 65.630 175.095 ;
        RECT 66.340 174.900 66.480 175.260 ;
        RECT 66.280 174.580 66.540 174.900 ;
        RECT 64.900 173.900 65.160 174.220 ;
        RECT 64.960 172.860 65.100 173.900 ;
        RECT 64.900 172.540 65.160 172.860 ;
        RECT 66.800 166.400 66.940 202.460 ;
        RECT 73.240 202.100 73.380 203.480 ;
        RECT 73.180 201.780 73.440 202.100 ;
        RECT 71.800 200.760 72.060 201.080 ;
        RECT 72.720 200.760 72.980 201.080 ;
        RECT 71.860 199.380 72.000 200.760 ;
        RECT 68.580 199.060 68.840 199.380 ;
        RECT 71.800 199.060 72.060 199.380 ;
        RECT 68.640 197.340 68.780 199.060 ;
        RECT 72.780 198.360 72.920 200.760 ;
        RECT 73.700 198.700 73.840 207.560 ;
        RECT 79.620 207.220 79.880 207.540 ;
        RECT 74.100 206.200 74.360 206.520 ;
        RECT 75.940 206.200 76.200 206.520 ;
        RECT 74.160 205.500 74.300 206.200 ;
        RECT 74.100 205.180 74.360 205.500 ;
        RECT 76.000 205.160 76.140 206.200 ;
        RECT 76.880 205.665 78.760 206.035 ;
        RECT 75.940 204.840 76.200 205.160 ;
        RECT 74.100 203.480 74.360 203.800 ;
        RECT 74.160 201.760 74.300 203.480 ;
        RECT 76.400 202.120 76.660 202.440 ;
        RECT 74.560 201.780 74.820 202.100 ;
        RECT 74.100 201.440 74.360 201.760 ;
        RECT 74.160 200.060 74.300 201.440 ;
        RECT 74.100 199.740 74.360 200.060 ;
        RECT 74.620 199.720 74.760 201.780 ;
        RECT 75.020 201.100 75.280 201.420 ;
        RECT 75.480 201.100 75.740 201.420 ;
        RECT 75.080 200.060 75.220 201.100 ;
        RECT 75.020 199.740 75.280 200.060 ;
        RECT 74.560 199.400 74.820 199.720 ;
        RECT 73.180 198.380 73.440 198.700 ;
        RECT 73.640 198.380 73.900 198.700 ;
        RECT 72.720 198.040 72.980 198.360 ;
        RECT 68.580 197.020 68.840 197.340 ;
        RECT 69.960 197.020 70.220 197.340 ;
        RECT 69.040 196.000 69.300 196.320 ;
        RECT 69.100 193.940 69.240 196.000 ;
        RECT 69.040 193.620 69.300 193.940 ;
        RECT 70.020 190.620 70.160 197.020 ;
        RECT 72.780 196.660 72.920 198.040 ;
        RECT 73.240 196.660 73.380 198.380 ;
        RECT 73.700 197.340 73.840 198.380 ;
        RECT 73.640 197.020 73.900 197.340 ;
        RECT 70.420 196.340 70.680 196.660 ;
        RECT 72.720 196.340 72.980 196.660 ;
        RECT 73.180 196.340 73.440 196.660 ;
        RECT 70.480 192.920 70.620 196.340 ;
        RECT 71.800 195.660 72.060 195.980 ;
        RECT 71.860 194.620 72.000 195.660 ;
        RECT 71.800 194.300 72.060 194.620 ;
        RECT 72.780 194.280 72.920 196.340 ;
        RECT 72.720 193.960 72.980 194.280 ;
        RECT 73.240 193.940 73.380 196.340 ;
        RECT 73.180 193.620 73.440 193.940 ;
        RECT 70.420 192.600 70.680 192.920 ;
        RECT 72.720 192.830 72.980 192.920 ;
        RECT 72.320 192.690 72.980 192.830 ;
        RECT 71.340 190.900 71.600 191.220 ;
        RECT 71.400 190.620 71.540 190.900 ;
        RECT 70.020 190.480 71.540 190.620 ;
        RECT 69.960 189.880 70.220 190.200 ;
        RECT 68.120 185.460 68.380 185.780 ;
        RECT 68.180 183.060 68.320 185.460 ;
        RECT 68.120 182.740 68.380 183.060 ;
        RECT 69.500 181.720 69.760 182.040 ;
        RECT 67.660 180.360 67.920 180.680 ;
        RECT 67.720 179.855 67.860 180.360 ;
        RECT 67.650 179.485 67.930 179.855 ;
        RECT 68.580 179.740 68.840 180.000 ;
        RECT 68.580 179.680 69.240 179.740 ;
        RECT 68.640 179.600 69.240 179.680 ;
        RECT 69.100 177.620 69.240 179.600 ;
        RECT 69.560 177.620 69.700 181.720 ;
        RECT 69.040 177.300 69.300 177.620 ;
        RECT 69.500 177.300 69.760 177.620 ;
        RECT 69.100 176.600 69.240 177.300 ;
        RECT 68.120 176.280 68.380 176.600 ;
        RECT 69.040 176.280 69.300 176.600 ;
        RECT 68.180 175.580 68.320 176.280 ;
        RECT 68.120 175.260 68.380 175.580 ;
        RECT 70.020 174.900 70.160 189.880 ;
        RECT 72.320 188.160 72.460 192.690 ;
        RECT 72.720 192.600 72.980 192.690 ;
        RECT 73.240 191.300 73.380 193.620 ;
        RECT 72.780 191.160 73.380 191.300 ;
        RECT 72.260 187.840 72.520 188.160 ;
        RECT 71.340 185.800 71.600 186.120 ;
        RECT 71.400 183.740 71.540 185.800 ;
        RECT 71.340 183.420 71.600 183.740 ;
        RECT 71.800 183.420 72.060 183.740 ;
        RECT 71.860 183.060 72.000 183.420 ;
        RECT 71.800 182.740 72.060 183.060 ;
        RECT 72.320 182.970 72.460 187.840 ;
        RECT 72.780 185.100 72.920 191.160 ;
        RECT 73.180 190.560 73.440 190.880 ;
        RECT 73.240 189.180 73.380 190.560 ;
        RECT 73.700 190.540 73.840 197.020 ;
        RECT 74.620 196.320 74.760 199.400 ;
        RECT 74.560 196.000 74.820 196.320 ;
        RECT 74.620 190.880 74.760 196.000 ;
        RECT 75.540 195.980 75.680 201.100 ;
        RECT 75.940 200.760 76.200 201.080 ;
        RECT 76.000 199.040 76.140 200.760 ;
        RECT 76.460 200.060 76.600 202.120 ;
        RECT 79.160 201.780 79.420 202.100 ;
        RECT 76.880 200.225 78.760 200.595 ;
        RECT 76.400 199.740 76.660 200.060 ;
        RECT 79.220 199.380 79.360 201.780 ;
        RECT 79.680 201.420 79.820 207.220 ;
        RECT 106.880 205.665 108.760 206.035 ;
        RECT 83.760 204.840 84.020 205.160 ;
        RECT 79.620 201.100 79.880 201.420 ;
        RECT 79.680 200.060 79.820 201.100 ;
        RECT 83.820 200.060 83.960 204.840 ;
        RECT 88.360 204.160 88.620 204.480 ;
        RECT 84.680 201.780 84.940 202.100 ;
        RECT 84.740 200.060 84.880 201.780 ;
        RECT 88.420 201.760 88.560 204.160 ;
        RECT 91.880 202.945 93.760 203.315 ;
        RECT 121.880 202.945 123.760 203.315 ;
        RECT 88.360 201.440 88.620 201.760 ;
        RECT 96.640 201.440 96.900 201.760 ;
        RECT 85.600 201.100 85.860 201.420 ;
        RECT 85.660 200.060 85.800 201.100 ;
        RECT 79.620 199.740 79.880 200.060 ;
        RECT 83.760 199.740 84.020 200.060 ;
        RECT 84.680 199.740 84.940 200.060 ;
        RECT 85.600 199.740 85.860 200.060 ;
        RECT 81.000 199.400 81.260 199.720 ;
        RECT 79.160 199.060 79.420 199.380 ;
        RECT 80.080 199.060 80.340 199.380 ;
        RECT 75.940 198.720 76.200 199.040 ;
        RECT 80.140 197.000 80.280 199.060 ;
        RECT 81.060 198.360 81.200 199.400 ;
        RECT 86.980 199.060 87.240 199.380 ;
        RECT 81.000 198.040 81.260 198.360 ;
        RECT 80.080 196.680 80.340 197.000 ;
        RECT 75.480 195.660 75.740 195.980 ;
        RECT 76.880 194.785 78.760 195.155 ;
        RECT 76.400 193.620 76.660 193.940 ;
        RECT 74.560 190.560 74.820 190.880 ;
        RECT 73.640 190.220 73.900 190.540 ;
        RECT 73.180 188.860 73.440 189.180 ;
        RECT 73.700 185.780 73.840 190.220 ;
        RECT 73.640 185.460 73.900 185.780 ;
        RECT 72.720 184.780 72.980 185.100 ;
        RECT 72.780 183.740 72.920 184.780 ;
        RECT 72.720 183.420 72.980 183.740 ;
        RECT 73.700 183.400 73.840 185.460 ;
        RECT 74.620 185.440 74.760 190.560 ;
        RECT 76.460 190.200 76.600 193.620 ;
        RECT 80.140 191.220 80.280 196.680 ;
        RECT 85.600 195.320 85.860 195.640 ;
        RECT 85.660 194.620 85.800 195.320 ;
        RECT 85.600 194.300 85.860 194.620 ;
        RECT 85.140 193.280 85.400 193.600 ;
        RECT 80.080 190.900 80.340 191.220 ;
        RECT 76.400 189.880 76.660 190.200 ;
        RECT 76.460 186.120 76.600 189.880 ;
        RECT 76.880 189.345 78.760 189.715 ;
        RECT 76.400 185.800 76.660 186.120 ;
        RECT 74.560 185.120 74.820 185.440 ;
        RECT 75.940 184.780 76.200 185.100 ;
        RECT 74.560 184.440 74.820 184.760 ;
        RECT 74.100 183.420 74.360 183.740 ;
        RECT 73.640 183.310 73.900 183.400 ;
        RECT 73.240 183.170 73.900 183.310 ;
        RECT 72.720 182.970 72.980 183.060 ;
        RECT 72.320 182.830 72.980 182.970 ;
        RECT 72.720 182.740 72.980 182.830 ;
        RECT 72.720 182.060 72.980 182.380 ;
        RECT 72.780 180.340 72.920 182.060 ;
        RECT 73.240 180.340 73.380 183.170 ;
        RECT 73.640 183.080 73.900 183.170 ;
        RECT 73.640 182.400 73.900 182.720 ;
        RECT 72.720 180.020 72.980 180.340 ;
        RECT 73.180 180.020 73.440 180.340 ;
        RECT 71.340 179.680 71.600 180.000 ;
        RECT 70.410 177.445 70.690 177.815 ;
        RECT 69.960 174.580 70.220 174.900 ;
        RECT 69.040 174.240 69.300 174.560 ;
        RECT 69.100 172.180 69.240 174.240 ;
        RECT 69.040 171.860 69.300 172.180 ;
        RECT 67.660 169.820 67.920 170.140 ;
        RECT 66.740 166.080 67.000 166.400 ;
        RECT 66.800 161.300 66.940 166.080 ;
        RECT 67.200 162.680 67.460 163.000 ;
        RECT 66.740 160.980 67.000 161.300 ;
        RECT 67.260 160.960 67.400 162.680 ;
        RECT 67.200 160.640 67.460 160.960 ;
        RECT 67.200 159.960 67.460 160.280 ;
        RECT 67.260 156.540 67.400 159.960 ;
        RECT 67.200 156.220 67.460 156.540 ;
        RECT 65.820 155.375 66.080 155.520 ;
        RECT 65.810 155.005 66.090 155.375 ;
        RECT 64.440 152.820 64.700 153.140 ;
        RECT 65.820 152.480 66.080 152.800 ;
        RECT 65.880 151.100 66.020 152.480 ;
        RECT 61.220 150.780 61.480 151.100 ;
        RECT 65.820 150.780 66.080 151.100 ;
        RECT 53.400 150.100 53.660 150.420 ;
        RECT 53.860 150.100 54.120 150.420 ;
        RECT 56.620 150.100 56.880 150.420 ;
        RECT 58.920 150.100 59.180 150.420 ;
        RECT 63.980 150.100 64.240 150.420 ;
        RECT 53.460 147.700 53.600 150.100 ;
        RECT 52.480 147.380 52.740 147.700 ;
        RECT 53.400 147.380 53.660 147.700 ;
        RECT 52.020 147.040 52.280 147.360 ;
        RECT 51.560 146.700 51.820 147.020 ;
        RECT 52.080 145.660 52.220 147.040 ;
        RECT 51.100 145.340 51.360 145.660 ;
        RECT 52.020 145.340 52.280 145.660 ;
        RECT 49.720 144.660 49.980 144.980 ;
        RECT 49.320 144.240 49.920 144.380 ;
        RECT 50.640 144.320 50.900 144.640 ;
        RECT 46.500 141.940 46.760 142.260 ;
        RECT 46.040 141.600 46.300 141.920 ;
        RECT 46.880 140.385 48.760 140.755 ;
        RECT 47.880 138.200 48.140 138.520 ;
        RECT 45.580 136.500 45.840 136.820 ;
        RECT 47.940 136.480 48.080 138.200 ;
        RECT 48.340 137.180 48.600 137.500 ;
        RECT 48.400 136.480 48.540 137.180 ;
        RECT 47.880 136.390 48.140 136.480 ;
        RECT 46.560 136.250 48.140 136.390 ;
        RECT 46.560 134.100 46.700 136.250 ;
        RECT 47.880 136.160 48.140 136.250 ;
        RECT 48.340 136.160 48.600 136.480 ;
        RECT 49.260 135.820 49.520 136.140 ;
        RECT 46.880 134.945 48.760 135.315 ;
        RECT 46.500 133.780 46.760 134.100 ;
        RECT 49.320 133.760 49.460 135.820 ;
        RECT 49.260 133.440 49.520 133.760 ;
        RECT 49.250 131.885 49.530 132.255 ;
        RECT 49.320 130.700 49.460 131.885 ;
        RECT 49.260 130.380 49.520 130.700 ;
        RECT 46.880 129.505 48.760 129.875 ;
        RECT 45.120 129.020 45.380 129.340 ;
        RECT 46.040 128.340 46.300 128.660 ;
        RECT 46.100 125.600 46.240 128.340 ;
        RECT 44.660 125.280 44.920 125.600 ;
        RECT 46.040 125.280 46.300 125.600 ;
        RECT 46.500 125.280 46.760 125.600 ;
        RECT 46.040 124.600 46.300 124.920 ;
        RECT 46.100 122.540 46.240 124.600 ;
        RECT 46.040 122.220 46.300 122.540 ;
        RECT 46.560 120.500 46.700 125.280 ;
        RECT 46.880 124.065 48.760 124.435 ;
        RECT 46.960 122.220 47.220 122.540 ;
        RECT 47.020 120.500 47.160 122.220 ;
        RECT 46.500 120.410 46.760 120.500 ;
        RECT 46.100 120.270 46.760 120.410 ;
        RECT 45.580 119.840 45.840 120.160 ;
        RECT 45.120 119.160 45.380 119.480 ;
        RECT 45.180 117.780 45.320 119.160 ;
        RECT 45.120 117.460 45.380 117.780 ;
        RECT 45.640 115.740 45.780 119.840 ;
        RECT 46.100 116.760 46.240 120.270 ;
        RECT 46.500 120.180 46.760 120.270 ;
        RECT 46.960 120.180 47.220 120.500 ;
        RECT 46.500 119.500 46.760 119.820 ;
        RECT 46.560 117.780 46.700 119.500 ;
        RECT 46.880 118.625 48.760 118.995 ;
        RECT 46.500 117.460 46.760 117.780 ;
        RECT 46.040 116.440 46.300 116.760 ;
        RECT 45.580 115.420 45.840 115.740 ;
        RECT 46.100 115.060 46.240 116.440 ;
        RECT 46.040 114.740 46.300 115.060 ;
        RECT 46.880 113.185 48.760 113.555 ;
        RECT 49.320 112.680 49.460 130.380 ;
        RECT 49.780 129.340 49.920 144.240 ;
        RECT 50.180 138.200 50.440 138.520 ;
        RECT 50.240 134.100 50.380 138.200 ;
        RECT 50.700 136.820 50.840 144.320 ;
        RECT 53.460 142.260 53.600 147.380 ;
        RECT 53.920 145.660 54.060 150.100 ;
        RECT 54.320 149.820 54.580 150.080 ;
        RECT 54.320 149.760 54.980 149.820 ;
        RECT 54.380 149.680 54.980 149.760 ;
        RECT 54.840 148.380 54.980 149.680 ;
        RECT 54.780 148.060 55.040 148.380 ;
        RECT 54.840 147.360 54.980 148.060 ;
        RECT 56.680 147.360 56.820 150.100 ;
        RECT 57.080 147.720 57.340 148.040 ;
        RECT 54.780 147.270 55.040 147.360 ;
        RECT 56.620 147.270 56.880 147.360 ;
        RECT 54.380 147.130 55.040 147.270 ;
        RECT 53.860 145.340 54.120 145.660 ;
        RECT 54.380 142.340 54.520 147.130 ;
        RECT 54.780 147.040 55.040 147.130 ;
        RECT 56.220 147.130 56.880 147.270 ;
        RECT 55.240 145.000 55.500 145.320 ;
        RECT 54.780 144.320 55.040 144.640 ;
        RECT 53.400 141.940 53.660 142.260 ;
        RECT 53.920 142.200 54.520 142.340 ;
        RECT 53.460 137.500 53.600 141.940 ;
        RECT 53.920 141.920 54.060 142.200 ;
        RECT 53.860 141.600 54.120 141.920 ;
        RECT 53.920 138.520 54.060 141.600 ;
        RECT 53.860 138.200 54.120 138.520 ;
        RECT 51.100 137.180 51.360 137.500 ;
        RECT 53.400 137.180 53.660 137.500 ;
        RECT 50.640 136.500 50.900 136.820 ;
        RECT 50.640 135.820 50.900 136.140 ;
        RECT 50.700 134.780 50.840 135.820 ;
        RECT 50.640 134.460 50.900 134.780 ;
        RECT 51.160 134.180 51.300 137.180 ;
        RECT 54.840 136.820 54.980 144.320 ;
        RECT 55.300 139.200 55.440 145.000 ;
        RECT 56.220 141.920 56.360 147.130 ;
        RECT 56.620 147.040 56.880 147.130 ;
        RECT 56.160 141.600 56.420 141.920 ;
        RECT 56.220 140.300 56.360 141.600 ;
        RECT 55.760 140.160 56.360 140.300 ;
        RECT 55.240 138.880 55.500 139.200 ;
        RECT 54.780 136.500 55.040 136.820 ;
        RECT 52.480 135.820 52.740 136.140 ;
        RECT 52.020 135.480 52.280 135.800 ;
        RECT 50.700 134.100 51.300 134.180 ;
        RECT 50.180 133.780 50.440 134.100 ;
        RECT 50.640 134.040 51.300 134.100 ;
        RECT 50.640 133.780 50.900 134.040 ;
        RECT 50.700 133.080 50.840 133.780 ;
        RECT 50.640 132.760 50.900 133.080 ;
        RECT 49.720 129.020 49.980 129.340 ;
        RECT 50.180 119.840 50.440 120.160 ;
        RECT 49.720 119.160 49.980 119.480 ;
        RECT 49.780 114.720 49.920 119.160 ;
        RECT 50.240 115.060 50.380 119.840 ;
        RECT 51.100 119.160 51.360 119.480 ;
        RECT 51.160 118.120 51.300 119.160 ;
        RECT 51.100 117.800 51.360 118.120 ;
        RECT 50.180 114.740 50.440 115.060 ;
        RECT 49.720 114.400 49.980 114.720 ;
        RECT 49.260 112.360 49.520 112.680 ;
        RECT 44.260 111.700 46.240 111.840 ;
        RECT 46.100 106.900 46.240 111.700 ;
        RECT 50.640 111.680 50.900 112.000 ;
        RECT 46.880 107.745 48.760 108.115 ;
        RECT 36.840 106.580 37.100 106.900 ;
        RECT 38.680 106.580 38.940 106.900 ;
        RECT 41.440 106.580 41.700 106.900 ;
        RECT 46.040 106.580 46.300 106.900 ;
        RECT 50.180 106.580 50.440 106.900 ;
        RECT 35.460 106.240 35.720 106.560 ;
        RECT 35.520 104.180 35.660 106.240 ;
        RECT 36.380 105.560 36.640 105.880 ;
        RECT 36.440 104.180 36.580 105.560 ;
        RECT 36.900 104.860 37.040 106.580 ;
        RECT 49.720 106.240 49.980 106.560 ;
        RECT 43.280 105.560 43.540 105.880 ;
        RECT 48.340 105.560 48.600 105.880 ;
        RECT 36.840 104.540 37.100 104.860 ;
        RECT 35.460 103.860 35.720 104.180 ;
        RECT 36.380 103.860 36.640 104.180 ;
        RECT 34.080 101.480 34.340 101.800 ;
        RECT 36.900 101.460 37.040 104.540 ;
        RECT 43.340 103.500 43.480 105.560 ;
        RECT 48.400 104.180 48.540 105.560 ;
        RECT 49.780 104.260 49.920 106.240 ;
        RECT 50.240 104.860 50.380 106.580 ;
        RECT 50.180 104.540 50.440 104.860 ;
        RECT 50.700 104.520 50.840 111.680 ;
        RECT 52.080 109.280 52.220 135.480 ;
        RECT 52.540 134.100 52.680 135.820 ;
        RECT 52.480 133.780 52.740 134.100 ;
        RECT 54.840 128.320 54.980 136.500 ;
        RECT 55.760 136.140 55.900 140.160 ;
        RECT 56.160 139.220 56.420 139.540 ;
        RECT 55.700 135.820 55.960 136.140 ;
        RECT 56.220 134.440 56.360 139.220 ;
        RECT 56.620 135.480 56.880 135.800 ;
        RECT 56.680 134.780 56.820 135.480 ;
        RECT 56.620 134.460 56.880 134.780 ;
        RECT 56.160 134.120 56.420 134.440 ;
        RECT 55.700 133.100 55.960 133.420 ;
        RECT 55.760 129.340 55.900 133.100 ;
        RECT 56.680 129.340 56.820 134.460 ;
        RECT 55.700 129.020 55.960 129.340 ;
        RECT 56.620 129.020 56.880 129.340 ;
        RECT 54.780 128.000 55.040 128.320 ;
        RECT 54.840 125.940 54.980 128.000 ;
        RECT 55.760 126.280 55.900 129.020 ;
        RECT 55.700 125.960 55.960 126.280 ;
        RECT 54.780 125.620 55.040 125.940 ;
        RECT 55.760 123.900 55.900 125.960 ;
        RECT 55.700 123.580 55.960 123.900 ;
        RECT 54.780 117.460 55.040 117.780 ;
        RECT 54.840 115.740 54.980 117.460 ;
        RECT 56.620 117.120 56.880 117.440 ;
        RECT 54.780 115.420 55.040 115.740 ;
        RECT 52.020 108.960 52.280 109.280 ;
        RECT 55.700 108.280 55.960 108.600 ;
        RECT 55.760 107.240 55.900 108.280 ;
        RECT 55.700 106.920 55.960 107.240 ;
        RECT 52.480 106.240 52.740 106.560 ;
        RECT 56.680 106.470 56.820 117.120 ;
        RECT 57.140 109.280 57.280 147.720 ;
        RECT 58.980 147.020 59.120 150.100 ;
        RECT 60.300 149.420 60.560 149.740 ;
        RECT 58.920 146.700 59.180 147.020 ;
        RECT 59.380 146.360 59.640 146.680 ;
        RECT 59.440 145.320 59.580 146.360 ;
        RECT 59.380 145.000 59.640 145.320 ;
        RECT 58.920 143.640 59.180 143.960 ;
        RECT 58.980 141.580 59.120 143.640 ;
        RECT 59.440 142.940 59.580 145.000 ;
        RECT 59.380 142.620 59.640 142.940 ;
        RECT 58.920 141.260 59.180 141.580 ;
        RECT 59.840 135.480 60.100 135.800 ;
        RECT 59.900 134.100 60.040 135.480 ;
        RECT 59.840 133.780 60.100 134.100 ;
        RECT 60.360 133.500 60.500 149.420 ;
        RECT 61.880 148.545 63.760 148.915 ;
        RECT 64.040 146.680 64.180 150.100 ;
        RECT 65.820 149.760 66.080 150.080 ;
        RECT 64.900 149.420 65.160 149.740 ;
        RECT 64.960 147.700 65.100 149.420 ;
        RECT 65.360 149.080 65.620 149.400 ;
        RECT 64.900 147.380 65.160 147.700 ;
        RECT 63.980 146.360 64.240 146.680 ;
        RECT 64.960 144.640 65.100 147.380 ;
        RECT 64.900 144.320 65.160 144.640 ;
        RECT 63.980 143.980 64.240 144.300 ;
        RECT 61.880 143.105 63.760 143.475 ;
        RECT 64.040 141.240 64.180 143.980 ;
        RECT 63.980 140.920 64.240 141.240 ;
        RECT 61.220 139.900 61.480 140.220 ;
        RECT 60.760 139.220 61.020 139.540 ;
        RECT 60.820 137.500 60.960 139.220 ;
        RECT 60.760 137.180 61.020 137.500 ;
        RECT 60.760 135.820 61.020 136.140 ;
        RECT 59.900 133.360 60.500 133.500 ;
        RECT 58.000 127.320 58.260 127.640 ;
        RECT 58.060 125.600 58.200 127.320 ;
        RECT 58.000 125.280 58.260 125.600 ;
        RECT 57.540 123.240 57.800 123.560 ;
        RECT 57.600 121.180 57.740 123.240 ;
        RECT 59.900 122.620 60.040 133.360 ;
        RECT 60.820 125.600 60.960 135.820 ;
        RECT 61.280 135.800 61.420 139.900 ;
        RECT 61.880 137.665 63.760 138.035 ;
        RECT 61.220 135.480 61.480 135.800 ;
        RECT 64.040 134.100 64.180 140.920 ;
        RECT 65.420 139.540 65.560 149.080 ;
        RECT 65.880 147.360 66.020 149.760 ;
        RECT 65.820 147.040 66.080 147.360 ;
        RECT 65.820 144.660 66.080 144.980 ;
        RECT 65.880 140.220 66.020 144.660 ;
        RECT 65.820 139.900 66.080 140.220 ;
        RECT 65.360 139.220 65.620 139.540 ;
        RECT 64.440 138.540 64.700 138.860 ;
        RECT 64.500 136.480 64.640 138.540 ;
        RECT 65.420 137.500 65.560 139.220 ;
        RECT 65.360 137.180 65.620 137.500 ;
        RECT 65.420 136.900 65.560 137.180 ;
        RECT 64.960 136.760 65.560 136.900 ;
        RECT 65.880 136.820 66.020 139.900 ;
        RECT 66.280 139.220 66.540 139.540 ;
        RECT 64.440 136.160 64.700 136.480 ;
        RECT 64.500 134.440 64.640 136.160 ;
        RECT 64.440 134.120 64.700 134.440 ;
        RECT 64.960 134.100 65.100 136.760 ;
        RECT 65.820 136.500 66.080 136.820 ;
        RECT 65.360 135.820 65.620 136.140 ;
        RECT 65.420 134.100 65.560 135.820 ;
        RECT 63.980 133.780 64.240 134.100 ;
        RECT 64.900 133.780 65.160 134.100 ;
        RECT 65.360 133.780 65.620 134.100 ;
        RECT 65.820 133.780 66.080 134.100 ;
        RECT 61.880 132.225 63.760 132.595 ;
        RECT 64.040 129.000 64.180 133.780 ;
        RECT 64.900 131.060 65.160 131.380 ;
        RECT 64.440 130.380 64.700 130.700 ;
        RECT 63.980 128.680 64.240 129.000 ;
        RECT 64.040 128.320 64.180 128.680 ;
        RECT 63.980 128.000 64.240 128.320 ;
        RECT 61.880 126.785 63.760 127.155 ;
        RECT 60.760 125.280 61.020 125.600 ;
        RECT 60.300 124.600 60.560 124.920 ;
        RECT 60.360 123.220 60.500 124.600 ;
        RECT 60.820 123.900 60.960 125.280 ;
        RECT 60.760 123.580 61.020 123.900 ;
        RECT 60.300 122.900 60.560 123.220 ;
        RECT 59.900 122.480 60.500 122.620 ;
        RECT 57.540 120.860 57.800 121.180 ;
        RECT 58.000 119.840 58.260 120.160 ;
        RECT 58.060 117.780 58.200 119.840 ;
        RECT 58.000 117.460 58.260 117.780 ;
        RECT 59.840 117.460 60.100 117.780 ;
        RECT 59.900 109.280 60.040 117.460 ;
        RECT 60.360 111.840 60.500 122.480 ;
        RECT 60.820 121.180 60.960 123.580 ;
        RECT 64.040 123.220 64.180 128.000 ;
        RECT 64.500 123.220 64.640 130.380 ;
        RECT 63.980 122.900 64.240 123.220 ;
        RECT 64.440 122.900 64.700 123.220 ;
        RECT 61.880 121.345 63.760 121.715 ;
        RECT 60.760 120.860 61.020 121.180 ;
        RECT 62.140 119.500 62.400 119.820 ;
        RECT 62.200 118.460 62.340 119.500 ;
        RECT 64.500 118.460 64.640 122.900 ;
        RECT 64.960 122.880 65.100 131.060 ;
        RECT 65.880 130.700 66.020 133.780 ;
        RECT 65.820 130.380 66.080 130.700 ;
        RECT 66.340 130.360 66.480 139.220 ;
        RECT 67.720 138.860 67.860 169.820 ;
        RECT 68.580 166.420 68.840 166.740 ;
        RECT 68.640 163.680 68.780 166.420 ;
        RECT 69.100 165.720 69.240 171.860 ;
        RECT 70.480 169.120 70.620 177.445 ;
        RECT 70.880 173.560 71.140 173.880 ;
        RECT 70.940 170.140 71.080 173.560 ;
        RECT 70.880 169.820 71.140 170.140 ;
        RECT 70.420 168.800 70.680 169.120 ;
        RECT 70.480 167.420 70.620 168.800 ;
        RECT 70.420 167.100 70.680 167.420 ;
        RECT 69.040 165.400 69.300 165.720 ;
        RECT 68.580 163.360 68.840 163.680 ;
        RECT 68.110 158.405 68.390 158.775 ;
        RECT 68.180 152.655 68.320 158.405 ;
        RECT 68.110 152.285 68.390 152.655 ;
        RECT 68.580 152.480 68.840 152.800 ;
        RECT 68.180 139.540 68.320 152.285 ;
        RECT 68.640 142.260 68.780 152.480 ;
        RECT 69.100 144.300 69.240 165.400 ;
        RECT 69.960 159.960 70.220 160.280 ;
        RECT 69.500 157.920 69.760 158.240 ;
        RECT 69.560 153.140 69.700 157.920 ;
        RECT 70.020 154.840 70.160 159.960 ;
        RECT 70.480 158.240 70.620 167.100 ;
        RECT 71.400 166.820 71.540 179.680 ;
        RECT 73.180 179.340 73.440 179.660 ;
        RECT 73.240 178.300 73.380 179.340 ;
        RECT 71.800 177.980 72.060 178.300 ;
        RECT 73.180 177.980 73.440 178.300 ;
        RECT 71.860 177.135 72.000 177.980 ;
        RECT 72.710 177.445 72.990 177.815 ;
        RECT 72.720 177.300 72.980 177.445 ;
        RECT 71.790 176.765 72.070 177.135 ;
        RECT 72.780 174.560 72.920 177.300 ;
        RECT 72.720 174.240 72.980 174.560 ;
        RECT 73.700 171.580 73.840 182.400 ;
        RECT 74.160 180.000 74.300 183.420 ;
        RECT 74.100 179.680 74.360 180.000 ;
        RECT 74.100 177.300 74.360 177.620 ;
        RECT 70.940 166.740 71.540 166.820 ;
        RECT 70.880 166.680 71.540 166.740 ;
        RECT 70.880 166.420 71.140 166.680 ;
        RECT 71.400 161.300 71.540 166.680 ;
        RECT 72.780 171.440 73.840 171.580 ;
        RECT 71.340 160.980 71.600 161.300 ;
        RECT 70.880 160.300 71.140 160.620 ;
        RECT 70.940 158.920 71.080 160.300 ;
        RECT 71.800 158.940 72.060 159.260 ;
        RECT 70.880 158.600 71.140 158.920 ;
        RECT 71.860 158.775 72.000 158.940 ;
        RECT 71.790 158.405 72.070 158.775 ;
        RECT 70.420 157.920 70.680 158.240 ;
        RECT 69.960 154.520 70.220 154.840 ;
        RECT 70.020 153.480 70.160 154.520 ;
        RECT 70.420 153.500 70.680 153.820 ;
        RECT 69.960 153.160 70.220 153.480 ;
        RECT 69.500 152.820 69.760 153.140 ;
        RECT 69.560 150.420 69.700 152.820 ;
        RECT 70.480 152.120 70.620 153.500 ;
        RECT 70.880 152.540 71.140 152.800 ;
        RECT 71.800 152.540 72.060 152.800 ;
        RECT 70.880 152.480 72.060 152.540 ;
        RECT 70.940 152.400 72.000 152.480 ;
        RECT 70.420 151.800 70.680 152.120 ;
        RECT 69.500 150.100 69.760 150.420 ;
        RECT 69.500 144.320 69.760 144.640 ;
        RECT 69.040 143.980 69.300 144.300 ;
        RECT 69.040 142.280 69.300 142.600 ;
        RECT 68.580 141.940 68.840 142.260 ;
        RECT 68.640 141.240 68.780 141.940 ;
        RECT 68.580 140.920 68.840 141.240 ;
        RECT 68.120 139.220 68.380 139.540 ;
        RECT 67.660 138.540 67.920 138.860 ;
        RECT 66.740 138.200 67.000 138.520 ;
        RECT 66.800 136.140 66.940 138.200 ;
        RECT 66.740 135.820 67.000 136.140 ;
        RECT 68.120 130.380 68.380 130.700 ;
        RECT 66.280 130.040 66.540 130.360 ;
        RECT 66.340 129.340 66.480 130.040 ;
        RECT 66.280 129.020 66.540 129.340 ;
        RECT 68.180 128.660 68.320 130.380 ;
        RECT 68.580 128.680 68.840 129.000 ;
        RECT 68.120 128.340 68.380 128.660 ;
        RECT 68.640 125.600 68.780 128.680 ;
        RECT 68.580 125.280 68.840 125.600 ;
        RECT 64.900 122.560 65.160 122.880 ;
        RECT 68.120 121.880 68.380 122.200 ;
        RECT 62.140 118.140 62.400 118.460 ;
        RECT 64.440 118.140 64.700 118.460 ;
        RECT 66.740 117.800 67.000 118.120 ;
        RECT 61.880 115.905 63.760 116.275 ;
        RECT 66.800 115.740 66.940 117.800 ;
        RECT 66.740 115.420 67.000 115.740 ;
        RECT 68.180 114.720 68.320 121.880 ;
        RECT 68.120 114.400 68.380 114.720 ;
        RECT 60.360 111.700 60.960 111.840 ;
        RECT 57.080 108.960 57.340 109.280 ;
        RECT 59.840 108.960 60.100 109.280 ;
        RECT 60.300 108.960 60.560 109.280 ;
        RECT 58.000 108.280 58.260 108.600 ;
        RECT 57.080 106.470 57.340 106.560 ;
        RECT 56.680 106.330 57.340 106.470 ;
        RECT 48.340 103.860 48.600 104.180 ;
        RECT 49.780 104.120 50.380 104.260 ;
        RECT 50.640 104.200 50.900 104.520 ;
        RECT 39.140 103.180 39.400 103.500 ;
        RECT 43.280 103.180 43.540 103.500 ;
        RECT 36.840 101.140 37.100 101.460 ;
        RECT 31.880 99.585 33.760 99.955 ;
        RECT 31.780 88.620 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 30.460 88.480 33.000 88.620 ;
        RECT 31.780 85.510 33.000 88.480 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 39.200 88.620 39.340 103.180 ;
        RECT 44.200 102.840 44.460 103.160 ;
        RECT 44.260 89.530 44.400 102.840 ;
        RECT 46.880 102.305 48.760 102.675 ;
        RECT 37.680 88.480 39.340 88.620 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 50.240 89.170 50.380 104.120 ;
        RECT 52.540 103.840 52.680 106.240 ;
        RECT 56.680 104.860 56.820 106.330 ;
        RECT 57.080 106.240 57.340 106.330 ;
        RECT 57.080 105.560 57.340 105.880 ;
        RECT 56.620 104.540 56.880 104.860 ;
        RECT 57.140 104.260 57.280 105.560 ;
        RECT 56.680 104.120 57.280 104.260 ;
        RECT 58.060 104.180 58.200 108.280 ;
        RECT 60.360 106.900 60.500 108.960 ;
        RECT 60.820 106.900 60.960 111.700 ;
        RECT 61.880 110.465 63.760 110.835 ;
        RECT 69.100 109.280 69.240 142.280 ;
        RECT 69.560 136.480 69.700 144.320 ;
        RECT 69.960 143.640 70.220 143.960 ;
        RECT 70.020 141.920 70.160 143.640 ;
        RECT 69.960 141.600 70.220 141.920 ;
        RECT 70.480 139.200 70.620 151.800 ;
        RECT 70.940 150.420 71.080 152.400 ;
        RECT 72.260 152.140 72.520 152.460 ;
        RECT 70.880 150.100 71.140 150.420 ;
        RECT 70.940 147.700 71.080 150.100 ;
        RECT 70.880 147.380 71.140 147.700 ;
        RECT 72.320 147.360 72.460 152.140 ;
        RECT 72.260 147.040 72.520 147.360 ;
        RECT 70.880 143.980 71.140 144.300 ;
        RECT 70.940 141.920 71.080 143.980 ;
        RECT 70.880 141.600 71.140 141.920 ;
        RECT 70.420 138.880 70.680 139.200 ;
        RECT 69.500 136.160 69.760 136.480 ;
        RECT 69.560 131.380 69.700 136.160 ;
        RECT 69.500 131.060 69.760 131.380 ;
        RECT 70.940 130.780 71.080 141.600 ;
        RECT 72.260 140.920 72.520 141.240 ;
        RECT 72.320 139.880 72.460 140.920 ;
        RECT 72.260 139.560 72.520 139.880 ;
        RECT 72.780 131.040 72.920 171.440 ;
        RECT 74.160 166.400 74.300 177.300 ;
        RECT 74.100 166.080 74.360 166.400 ;
        RECT 73.180 165.400 73.440 165.720 ;
        RECT 73.240 163.680 73.380 165.400 ;
        RECT 73.180 163.360 73.440 163.680 ;
        RECT 73.240 158.240 73.380 163.360 ;
        RECT 74.620 161.210 74.760 184.440 ;
        RECT 76.000 183.060 76.140 184.780 ;
        RECT 75.940 182.740 76.200 183.060 ;
        RECT 76.000 182.380 76.140 182.740 ;
        RECT 75.940 182.060 76.200 182.380 ;
        RECT 75.020 181.720 75.280 182.040 ;
        RECT 76.460 181.780 76.600 185.800 ;
        RECT 85.200 185.780 85.340 193.280 ;
        RECT 85.660 191.900 85.800 194.300 ;
        RECT 87.040 194.280 87.180 199.060 ;
        RECT 91.880 197.505 93.760 197.875 ;
        RECT 93.880 196.340 94.140 196.660 ;
        RECT 90.200 195.660 90.460 195.980 ;
        RECT 90.260 194.620 90.400 195.660 ;
        RECT 90.200 194.300 90.460 194.620 ;
        RECT 86.980 193.960 87.240 194.280 ;
        RECT 86.060 193.620 86.320 193.940 ;
        RECT 90.200 193.620 90.460 193.940 ;
        RECT 85.600 191.580 85.860 191.900 ;
        RECT 85.140 185.460 85.400 185.780 ;
        RECT 76.880 183.905 78.760 184.275 ;
        RECT 76.860 182.740 77.120 183.060 ;
        RECT 76.920 181.780 77.060 182.740 ;
        RECT 85.200 182.040 85.340 185.460 ;
        RECT 75.080 177.620 75.220 181.720 ;
        RECT 76.000 181.640 77.060 181.780 ;
        RECT 79.620 181.720 79.880 182.040 ;
        RECT 85.140 181.720 85.400 182.040 ;
        RECT 76.000 180.340 76.140 181.640 ;
        RECT 79.160 180.360 79.420 180.680 ;
        RECT 75.940 180.020 76.200 180.340 ;
        RECT 76.400 179.680 76.660 180.000 ;
        RECT 76.460 177.620 76.600 179.680 ;
        RECT 78.690 179.485 78.970 179.855 ;
        RECT 78.760 179.320 78.900 179.485 ;
        RECT 78.700 179.000 78.960 179.320 ;
        RECT 76.880 178.465 78.760 178.835 ;
        RECT 75.020 177.300 75.280 177.620 ;
        RECT 76.400 177.300 76.660 177.620 ;
        RECT 77.780 177.300 78.040 177.620 ;
        RECT 78.240 177.300 78.500 177.620 ;
        RECT 75.080 176.600 75.220 177.300 ;
        RECT 75.020 176.280 75.280 176.600 ;
        RECT 76.460 175.240 76.600 177.300 ;
        RECT 77.840 175.580 77.980 177.300 ;
        RECT 78.300 177.135 78.440 177.300 ;
        RECT 79.220 177.280 79.360 180.360 ;
        RECT 79.680 180.340 79.820 181.720 ;
        RECT 82.380 180.700 82.640 181.020 ;
        RECT 79.620 180.020 79.880 180.340 ;
        RECT 81.460 179.680 81.720 180.000 ;
        RECT 81.920 179.680 82.180 180.000 ;
        RECT 79.620 177.640 79.880 177.960 ;
        RECT 78.230 176.765 78.510 177.135 ;
        RECT 79.160 176.960 79.420 177.280 ;
        RECT 77.780 175.260 78.040 175.580 ;
        RECT 76.400 174.920 76.660 175.240 ;
        RECT 78.300 174.560 78.440 176.765 ;
        RECT 78.240 174.240 78.500 174.560 ;
        RECT 76.880 173.025 78.760 173.395 ;
        RECT 76.400 168.120 76.660 168.440 ;
        RECT 79.160 168.120 79.420 168.440 ;
        RECT 75.020 166.080 75.280 166.400 ;
        RECT 73.700 161.070 74.760 161.210 ;
        RECT 73.180 157.920 73.440 158.240 ;
        RECT 73.170 156.365 73.450 156.735 ;
        RECT 70.020 130.640 71.080 130.780 ;
        RECT 72.720 130.720 72.980 131.040 ;
        RECT 70.020 125.600 70.160 130.640 ;
        RECT 70.420 130.040 70.680 130.360 ;
        RECT 71.800 130.040 72.060 130.360 ;
        RECT 70.480 125.600 70.620 130.040 ;
        RECT 71.860 125.600 72.000 130.040 ;
        RECT 72.260 128.340 72.520 128.660 ;
        RECT 72.320 126.620 72.460 128.340 ;
        RECT 72.260 126.300 72.520 126.620 ;
        RECT 69.960 125.510 70.220 125.600 ;
        RECT 69.560 125.370 70.220 125.510 ;
        RECT 69.560 117.440 69.700 125.370 ;
        RECT 69.960 125.280 70.220 125.370 ;
        RECT 70.420 125.280 70.680 125.600 ;
        RECT 71.800 125.280 72.060 125.600 ;
        RECT 69.960 124.600 70.220 124.920 ;
        RECT 70.020 120.160 70.160 124.600 ;
        RECT 73.240 123.220 73.380 156.365 ;
        RECT 73.700 153.820 73.840 161.070 ;
        RECT 74.100 159.960 74.360 160.280 ;
        RECT 74.160 158.240 74.300 159.960 ;
        RECT 74.100 157.920 74.360 158.240 ;
        RECT 74.160 157.560 74.300 157.920 ;
        RECT 74.100 157.240 74.360 157.560 ;
        RECT 74.160 156.200 74.300 157.240 ;
        RECT 74.100 155.880 74.360 156.200 ;
        RECT 74.560 155.540 74.820 155.860 ;
        RECT 74.620 155.375 74.760 155.540 ;
        RECT 74.550 155.005 74.830 155.375 ;
        RECT 73.640 153.500 73.900 153.820 ;
        RECT 73.700 152.460 73.840 153.500 ;
        RECT 74.100 153.050 74.360 153.140 ;
        RECT 75.080 153.050 75.220 166.080 ;
        RECT 75.480 163.020 75.740 163.340 ;
        RECT 75.540 156.735 75.680 163.020 ;
        RECT 76.460 158.580 76.600 168.120 ;
        RECT 76.880 167.585 78.760 167.955 ;
        RECT 78.700 165.740 78.960 166.060 ;
        RECT 78.760 164.020 78.900 165.740 ;
        RECT 78.700 163.700 78.960 164.020 ;
        RECT 79.220 163.340 79.360 168.120 ;
        RECT 79.160 163.020 79.420 163.340 ;
        RECT 76.880 162.145 78.760 162.515 ;
        RECT 76.400 158.260 76.660 158.580 ;
        RECT 79.160 157.920 79.420 158.240 ;
        RECT 76.400 157.580 76.660 157.900 ;
        RECT 75.940 157.240 76.200 157.560 ;
        RECT 75.470 156.365 75.750 156.735 ;
        RECT 74.100 152.910 75.220 153.050 ;
        RECT 74.100 152.820 74.360 152.910 ;
        RECT 73.640 152.140 73.900 152.460 ;
        RECT 73.640 148.060 73.900 148.380 ;
        RECT 73.700 146.680 73.840 148.060 ;
        RECT 73.640 146.360 73.900 146.680 ;
        RECT 74.160 136.820 74.300 152.820 ;
        RECT 75.020 151.800 75.280 152.120 ;
        RECT 75.080 150.760 75.220 151.800 ;
        RECT 75.020 150.440 75.280 150.760 ;
        RECT 76.000 150.420 76.140 157.240 ;
        RECT 76.460 155.520 76.600 157.580 ;
        RECT 76.880 156.705 78.760 157.075 ;
        RECT 79.220 156.450 79.360 157.920 ;
        RECT 78.300 156.310 79.360 156.450 ;
        RECT 78.300 155.860 78.440 156.310 ;
        RECT 78.240 155.540 78.500 155.860 ;
        RECT 78.700 155.540 78.960 155.860 ;
        RECT 76.400 155.200 76.660 155.520 ;
        RECT 78.760 155.180 78.900 155.540 ;
        RECT 78.700 154.860 78.960 155.180 ;
        RECT 76.400 154.520 76.660 154.840 ;
        RECT 75.940 150.100 76.200 150.420 ;
        RECT 75.940 149.080 76.200 149.400 ;
        RECT 75.480 143.980 75.740 144.300 ;
        RECT 75.020 138.880 75.280 139.200 ;
        RECT 75.080 137.500 75.220 138.880 ;
        RECT 75.020 137.180 75.280 137.500 ;
        RECT 74.560 136.840 74.820 137.160 ;
        RECT 74.100 136.500 74.360 136.820 ;
        RECT 74.160 131.380 74.300 136.500 ;
        RECT 74.620 134.780 74.760 136.840 ;
        RECT 74.560 134.460 74.820 134.780 ;
        RECT 74.100 131.060 74.360 131.380 ;
        RECT 73.180 122.900 73.440 123.220 ;
        RECT 73.240 120.160 73.380 122.900 ;
        RECT 69.960 119.840 70.220 120.160 ;
        RECT 73.180 119.840 73.440 120.160 ;
        RECT 70.880 119.500 71.140 119.820 ;
        RECT 70.940 118.540 71.080 119.500 ;
        RECT 70.940 118.400 71.540 118.540 ;
        RECT 71.400 117.440 71.540 118.400 ;
        RECT 69.500 117.120 69.760 117.440 ;
        RECT 70.880 117.120 71.140 117.440 ;
        RECT 71.340 117.120 71.600 117.440 ;
        RECT 69.560 115.060 69.700 117.120 ;
        RECT 70.940 115.740 71.080 117.120 ;
        RECT 71.400 115.740 71.540 117.120 ;
        RECT 70.880 115.420 71.140 115.740 ;
        RECT 71.340 115.420 71.600 115.740 ;
        RECT 73.640 115.420 73.900 115.740 ;
        RECT 69.500 114.740 69.760 115.060 ;
        RECT 69.040 108.960 69.300 109.280 ;
        RECT 65.360 108.280 65.620 108.600 ;
        RECT 72.260 108.280 72.520 108.600 ;
        RECT 65.420 107.240 65.560 108.280 ;
        RECT 72.320 107.240 72.460 108.280 ;
        RECT 65.360 106.920 65.620 107.240 ;
        RECT 72.260 106.920 72.520 107.240 ;
        RECT 60.300 106.580 60.560 106.900 ;
        RECT 60.760 106.580 61.020 106.900 ;
        RECT 73.700 106.560 73.840 115.420 ;
        RECT 74.160 110.300 74.300 131.060 ;
        RECT 75.020 130.040 75.280 130.360 ;
        RECT 75.080 128.660 75.220 130.040 ;
        RECT 75.020 128.340 75.280 128.660 ;
        RECT 75.540 128.060 75.680 143.980 ;
        RECT 75.080 127.920 75.680 128.060 ;
        RECT 74.100 109.980 74.360 110.300 ;
        RECT 75.080 106.900 75.220 127.920 ;
        RECT 75.480 119.160 75.740 119.480 ;
        RECT 75.540 118.120 75.680 119.160 ;
        RECT 75.480 117.800 75.740 118.120 ;
        RECT 76.000 108.940 76.140 149.080 ;
        RECT 76.460 136.480 76.600 154.520 ;
        RECT 76.880 151.265 78.760 151.635 ;
        RECT 79.680 150.080 79.820 177.640 ;
        RECT 81.520 177.530 81.660 179.680 ;
        RECT 81.980 178.300 82.120 179.680 ;
        RECT 82.440 178.300 82.580 180.700 ;
        RECT 85.200 180.340 85.340 181.720 ;
        RECT 85.660 180.680 85.800 191.580 ;
        RECT 86.120 190.200 86.260 193.620 ;
        RECT 87.900 190.220 88.160 190.540 ;
        RECT 86.060 189.880 86.320 190.200 ;
        RECT 86.120 184.760 86.260 189.880 ;
        RECT 87.960 189.180 88.100 190.220 ;
        RECT 87.900 188.860 88.160 189.180 ;
        RECT 89.280 188.180 89.540 188.500 ;
        RECT 89.340 186.460 89.480 188.180 ;
        RECT 90.260 188.160 90.400 193.620 ;
        RECT 91.120 192.600 91.380 192.920 ;
        RECT 91.180 190.880 91.320 192.600 ;
        RECT 91.880 192.065 93.760 192.435 ;
        RECT 93.940 191.900 94.080 196.340 ;
        RECT 96.700 196.320 96.840 201.440 ;
        RECT 106.880 200.225 108.760 200.595 ;
        RECT 98.020 199.400 98.280 199.720 ;
        RECT 96.640 196.000 96.900 196.320 ;
        RECT 96.700 194.280 96.840 196.000 ;
        RECT 98.080 194.620 98.220 199.400 ;
        RECT 104.460 198.720 104.720 199.040 ;
        RECT 105.840 198.720 106.100 199.040 ;
        RECT 98.480 198.040 98.740 198.360 ;
        RECT 98.540 196.320 98.680 198.040 ;
        RECT 98.480 196.000 98.740 196.320 ;
        RECT 98.020 194.300 98.280 194.620 ;
        RECT 96.640 193.960 96.900 194.280 ;
        RECT 94.800 193.620 95.060 193.940 ;
        RECT 93.880 191.580 94.140 191.900 ;
        RECT 93.880 190.900 94.140 191.220 ;
        RECT 90.660 190.560 90.920 190.880 ;
        RECT 91.120 190.560 91.380 190.880 ;
        RECT 90.720 189.180 90.860 190.560 ;
        RECT 90.660 188.860 90.920 189.180 ;
        RECT 90.200 187.840 90.460 188.160 ;
        RECT 91.120 187.840 91.380 188.160 ;
        RECT 89.280 186.140 89.540 186.460 ;
        RECT 91.180 186.120 91.320 187.840 ;
        RECT 91.880 186.625 93.760 186.995 ;
        RECT 91.120 185.800 91.380 186.120 ;
        RECT 86.060 184.440 86.320 184.760 ;
        RECT 86.520 184.440 86.780 184.760 ;
        RECT 85.600 180.360 85.860 180.680 ;
        RECT 85.140 180.020 85.400 180.340 ;
        RECT 85.200 179.855 85.340 180.020 ;
        RECT 85.130 179.485 85.410 179.855 ;
        RECT 82.840 179.000 83.100 179.320 ;
        RECT 83.760 179.000 84.020 179.320 ;
        RECT 81.920 177.980 82.180 178.300 ;
        RECT 82.380 177.980 82.640 178.300 ;
        RECT 82.900 177.620 83.040 179.000 ;
        RECT 81.920 177.530 82.180 177.620 ;
        RECT 81.520 177.390 82.180 177.530 ;
        RECT 81.920 177.300 82.180 177.390 ;
        RECT 82.840 177.300 83.100 177.620 ;
        RECT 80.540 176.960 80.800 177.280 ;
        RECT 80.080 169.140 80.340 169.460 ;
        RECT 80.140 165.720 80.280 169.140 ;
        RECT 80.080 165.400 80.340 165.720 ;
        RECT 80.140 160.960 80.280 165.400 ;
        RECT 80.080 160.640 80.340 160.960 ;
        RECT 80.070 159.085 80.350 159.455 ;
        RECT 80.080 158.940 80.340 159.085 ;
        RECT 80.600 155.260 80.740 176.960 ;
        RECT 81.980 175.580 82.120 177.300 ;
        RECT 81.920 175.260 82.180 175.580 ;
        RECT 81.920 173.900 82.180 174.220 ;
        RECT 81.000 162.680 81.260 163.000 ;
        RECT 81.980 162.740 82.120 173.900 ;
        RECT 83.300 168.120 83.560 168.440 ;
        RECT 82.840 166.080 83.100 166.400 ;
        RECT 82.900 164.700 83.040 166.080 ;
        RECT 82.840 164.380 83.100 164.700 ;
        RECT 83.360 163.680 83.500 168.120 ;
        RECT 83.820 166.140 83.960 179.000 ;
        RECT 86.120 177.960 86.260 184.440 ;
        RECT 86.580 179.660 86.720 184.440 ;
        RECT 91.180 183.060 91.320 185.800 ;
        RECT 91.120 182.740 91.380 183.060 ;
        RECT 89.740 182.060 90.000 182.380 ;
        RECT 89.800 181.020 89.940 182.060 ;
        RECT 89.740 180.700 90.000 181.020 ;
        RECT 91.180 180.000 91.320 182.740 ;
        RECT 93.940 182.720 94.080 190.900 ;
        RECT 94.860 188.015 95.000 193.620 ;
        RECT 96.700 190.880 96.840 193.960 ;
        RECT 98.020 190.900 98.280 191.220 ;
        RECT 96.640 190.560 96.900 190.880 ;
        RECT 94.790 187.645 95.070 188.015 ;
        RECT 97.560 184.440 97.820 184.760 ;
        RECT 97.620 183.740 97.760 184.440 ;
        RECT 97.560 183.420 97.820 183.740 ;
        RECT 96.180 182.740 96.440 183.060 ;
        RECT 93.880 182.400 94.140 182.720 ;
        RECT 91.880 181.185 93.760 181.555 ;
        RECT 90.660 179.680 90.920 180.000 ;
        RECT 91.120 179.680 91.380 180.000 ;
        RECT 86.520 179.340 86.780 179.660 ;
        RECT 87.440 179.000 87.700 179.320 ;
        RECT 89.280 179.000 89.540 179.320 ;
        RECT 86.060 177.640 86.320 177.960 ;
        RECT 84.220 177.300 84.480 177.620 ;
        RECT 84.280 174.560 84.420 177.300 ;
        RECT 87.500 174.900 87.640 179.000 ;
        RECT 89.340 177.620 89.480 179.000 ;
        RECT 90.720 178.300 90.860 179.680 ;
        RECT 90.660 177.980 90.920 178.300 ;
        RECT 89.280 177.300 89.540 177.620 ;
        RECT 87.440 174.580 87.700 174.900 ;
        RECT 84.220 174.240 84.480 174.560 ;
        RECT 91.180 172.860 91.320 179.680 ;
        RECT 96.240 179.320 96.380 182.740 ;
        RECT 98.080 182.720 98.220 190.900 ;
        RECT 98.020 182.400 98.280 182.720 ;
        RECT 98.540 182.380 98.680 196.000 ;
        RECT 101.240 195.320 101.500 195.640 ;
        RECT 101.300 191.220 101.440 195.320 ;
        RECT 104.520 191.900 104.660 198.720 ;
        RECT 105.900 194.280 106.040 198.720 ;
        RECT 121.880 197.505 123.760 197.875 ;
        RECT 115.500 195.660 115.760 195.980 ;
        RECT 117.800 195.660 118.060 195.980 ;
        RECT 118.260 195.660 118.520 195.980 ;
        RECT 109.060 195.320 109.320 195.640 ;
        RECT 106.880 194.785 108.760 195.155 ;
        RECT 105.840 193.960 106.100 194.280 ;
        RECT 108.140 193.280 108.400 193.600 ;
        RECT 104.460 191.580 104.720 191.900 ;
        RECT 108.200 191.560 108.340 193.280 ;
        RECT 108.140 191.240 108.400 191.560 ;
        RECT 101.240 190.900 101.500 191.220 ;
        RECT 106.300 190.900 106.560 191.220 ;
        RECT 106.360 189.180 106.500 190.900 ;
        RECT 106.880 189.345 108.760 189.715 ;
        RECT 106.300 188.860 106.560 189.180 ;
        RECT 100.320 188.520 100.580 188.840 ;
        RECT 99.400 187.160 99.660 187.480 ;
        RECT 99.860 187.160 100.120 187.480 ;
        RECT 99.460 185.780 99.600 187.160 ;
        RECT 99.920 186.460 100.060 187.160 ;
        RECT 100.380 186.460 100.520 188.520 ;
        RECT 99.860 186.140 100.120 186.460 ;
        RECT 100.320 186.140 100.580 186.460 ;
        RECT 109.120 185.780 109.260 195.320 ;
        RECT 115.560 194.620 115.700 195.660 ;
        RECT 112.740 194.300 113.000 194.620 ;
        RECT 115.500 194.300 115.760 194.620 ;
        RECT 110.900 193.280 111.160 193.600 ;
        RECT 109.520 192.600 109.780 192.920 ;
        RECT 109.580 190.540 109.720 192.600 ;
        RECT 109.980 190.900 110.240 191.220 ;
        RECT 109.520 190.220 109.780 190.540 ;
        RECT 110.040 188.500 110.180 190.900 ;
        RECT 109.980 188.180 110.240 188.500 ;
        RECT 99.400 185.460 99.660 185.780 ;
        RECT 105.380 185.460 105.640 185.780 ;
        RECT 109.060 185.460 109.320 185.780 ;
        RECT 99.460 183.060 99.600 185.460 ;
        RECT 99.400 182.740 99.660 183.060 ;
        RECT 98.480 182.060 98.740 182.380 ;
        RECT 96.180 179.000 96.440 179.320 ;
        RECT 99.460 177.620 99.600 182.740 ;
        RECT 104.460 182.460 104.720 182.720 ;
        RECT 103.600 182.400 104.720 182.460 ;
        RECT 103.600 182.320 104.660 182.400 ;
        RECT 99.860 179.340 100.120 179.660 ;
        RECT 102.160 179.340 102.420 179.660 ;
        RECT 99.920 178.300 100.060 179.340 ;
        RECT 99.860 177.980 100.120 178.300 ;
        RECT 102.220 177.620 102.360 179.340 ;
        RECT 98.480 177.300 98.740 177.620 ;
        RECT 99.400 177.300 99.660 177.620 ;
        RECT 102.160 177.300 102.420 177.620 ;
        RECT 91.880 175.745 93.760 176.115 ;
        RECT 98.540 174.560 98.680 177.300 ;
        RECT 100.780 176.280 101.040 176.600 ;
        RECT 102.160 176.280 102.420 176.600 ;
        RECT 98.480 174.240 98.740 174.560 ;
        RECT 98.540 173.880 98.680 174.240 ;
        RECT 98.480 173.560 98.740 173.880 ;
        RECT 91.120 172.540 91.380 172.860 ;
        RECT 98.480 171.520 98.740 171.840 ;
        RECT 89.740 170.840 90.000 171.160 ;
        RECT 89.800 169.800 89.940 170.840 ;
        RECT 91.880 170.305 93.760 170.675 ;
        RECT 98.540 170.140 98.680 171.520 ;
        RECT 98.480 169.820 98.740 170.140 ;
        RECT 89.740 169.480 90.000 169.800 ;
        RECT 92.040 169.140 92.300 169.460 ;
        RECT 87.900 168.800 88.160 169.120 ;
        RECT 91.120 168.800 91.380 169.120 ;
        RECT 84.220 168.460 84.480 168.780 ;
        RECT 84.280 167.080 84.420 168.460 ;
        RECT 84.220 166.760 84.480 167.080 ;
        RECT 83.820 166.000 84.420 166.140 ;
        RECT 83.300 163.360 83.560 163.680 ;
        RECT 81.060 160.620 81.200 162.680 ;
        RECT 81.980 162.600 83.960 162.740 ;
        RECT 82.840 161.660 83.100 161.980 ;
        RECT 81.000 160.300 81.260 160.620 ;
        RECT 81.060 159.260 81.200 160.300 ;
        RECT 81.000 158.940 81.260 159.260 ;
        RECT 81.450 159.085 81.730 159.455 ;
        RECT 81.060 156.200 81.200 158.940 ;
        RECT 81.000 155.880 81.260 156.200 ;
        RECT 80.600 155.120 81.200 155.260 ;
        RECT 80.540 154.520 80.800 154.840 ;
        RECT 80.080 150.100 80.340 150.420 ;
        RECT 79.620 149.760 79.880 150.080 ;
        RECT 78.240 149.420 78.500 149.740 ;
        RECT 78.300 148.040 78.440 149.420 ;
        RECT 80.140 148.380 80.280 150.100 ;
        RECT 80.080 148.060 80.340 148.380 ;
        RECT 78.240 147.720 78.500 148.040 ;
        RECT 78.240 147.040 78.500 147.360 ;
        RECT 80.080 147.040 80.340 147.360 ;
        RECT 78.300 146.680 78.440 147.040 ;
        RECT 78.240 146.360 78.500 146.680 ;
        RECT 79.620 146.360 79.880 146.680 ;
        RECT 76.880 145.825 78.760 146.195 ;
        RECT 79.680 145.320 79.820 146.360 ;
        RECT 79.620 145.000 79.880 145.320 ;
        RECT 76.880 140.385 78.760 140.755 ;
        RECT 80.140 139.880 80.280 147.040 ;
        RECT 80.080 139.560 80.340 139.880 ;
        RECT 79.620 138.200 79.880 138.520 ;
        RECT 79.680 136.480 79.820 138.200 ;
        RECT 80.080 137.180 80.340 137.500 ;
        RECT 76.400 136.160 76.660 136.480 ;
        RECT 79.620 136.160 79.880 136.480 ;
        RECT 79.160 135.480 79.420 135.800 ;
        RECT 76.880 134.945 78.760 135.315 ;
        RECT 79.220 134.440 79.360 135.480 ;
        RECT 79.160 134.120 79.420 134.440 ;
        RECT 80.140 132.060 80.280 137.180 ;
        RECT 80.600 134.100 80.740 154.520 ;
        RECT 81.060 145.660 81.200 155.120 ;
        RECT 81.000 145.340 81.260 145.660 ;
        RECT 81.520 144.980 81.660 159.085 ;
        RECT 81.920 157.920 82.180 158.240 ;
        RECT 81.980 155.860 82.120 157.920 ;
        RECT 82.380 157.580 82.640 157.900 ;
        RECT 82.440 155.860 82.580 157.580 ;
        RECT 82.900 155.860 83.040 161.660 ;
        RECT 83.300 159.960 83.560 160.280 ;
        RECT 83.360 157.900 83.500 159.960 ;
        RECT 83.300 157.580 83.560 157.900 ;
        RECT 81.920 155.540 82.180 155.860 ;
        RECT 82.380 155.540 82.640 155.860 ;
        RECT 82.840 155.540 83.100 155.860 ;
        RECT 82.440 155.180 82.580 155.540 ;
        RECT 82.380 154.860 82.640 155.180 ;
        RECT 81.920 149.080 82.180 149.400 ;
        RECT 81.460 144.660 81.720 144.980 ;
        RECT 81.000 143.640 81.260 143.960 ;
        RECT 80.540 133.780 80.800 134.100 ;
        RECT 81.060 133.500 81.200 143.640 ;
        RECT 81.460 139.900 81.720 140.220 ;
        RECT 81.520 136.480 81.660 139.900 ;
        RECT 81.460 136.160 81.720 136.480 ;
        RECT 80.600 133.360 81.200 133.500 ;
        RECT 80.080 131.740 80.340 132.060 ;
        RECT 80.080 130.720 80.340 131.040 ;
        RECT 76.880 129.505 78.760 129.875 ;
        RECT 78.700 128.000 78.960 128.320 ;
        RECT 78.760 126.620 78.900 128.000 ;
        RECT 79.160 127.660 79.420 127.980 ;
        RECT 79.220 126.620 79.360 127.660 ;
        RECT 78.700 126.300 78.960 126.620 ;
        RECT 79.160 126.300 79.420 126.620 ;
        RECT 76.880 124.065 78.760 124.435 ;
        RECT 79.220 119.480 79.360 126.300 ;
        RECT 79.620 125.620 79.880 125.940 ;
        RECT 79.680 120.500 79.820 125.620 ;
        RECT 79.620 120.180 79.880 120.500 ;
        RECT 79.620 119.730 79.880 119.820 ;
        RECT 80.140 119.730 80.280 130.720 ;
        RECT 80.600 129.000 80.740 133.360 ;
        RECT 80.540 128.680 80.800 129.000 ;
        RECT 80.540 128.000 80.800 128.320 ;
        RECT 80.600 126.620 80.740 128.000 ;
        RECT 81.980 127.640 82.120 149.080 ;
        RECT 83.300 147.720 83.560 148.040 ;
        RECT 83.360 147.360 83.500 147.720 ;
        RECT 82.380 147.040 82.640 147.360 ;
        RECT 83.300 147.040 83.560 147.360 ;
        RECT 82.440 146.680 82.580 147.040 ;
        RECT 82.840 146.700 83.100 147.020 ;
        RECT 82.380 146.360 82.640 146.680 ;
        RECT 82.380 139.110 82.640 139.200 ;
        RECT 82.900 139.110 83.040 146.700 ;
        RECT 83.360 139.200 83.500 147.040 ;
        RECT 82.380 138.970 83.040 139.110 ;
        RECT 82.380 138.880 82.640 138.970 ;
        RECT 83.300 138.880 83.560 139.200 ;
        RECT 82.440 137.160 82.580 138.880 ;
        RECT 82.380 136.840 82.640 137.160 ;
        RECT 83.360 136.480 83.500 138.880 ;
        RECT 83.300 136.160 83.560 136.480 ;
        RECT 83.820 133.760 83.960 162.600 ;
        RECT 84.280 136.140 84.420 166.000 ;
        RECT 87.960 164.700 88.100 168.800 ;
        RECT 88.820 166.420 89.080 166.740 ;
        RECT 87.900 164.380 88.160 164.700 ;
        RECT 88.880 160.620 89.020 166.420 ;
        RECT 91.180 166.400 91.320 168.800 ;
        RECT 92.100 166.400 92.240 169.140 ;
        RECT 100.320 166.760 100.580 167.080 ;
        RECT 91.120 166.080 91.380 166.400 ;
        RECT 92.040 166.080 92.300 166.400 ;
        RECT 93.880 166.080 94.140 166.400 ;
        RECT 94.800 166.080 95.060 166.400 ;
        RECT 98.480 166.080 98.740 166.400 ;
        RECT 91.180 163.000 91.320 166.080 ;
        RECT 92.100 165.720 92.240 166.080 ;
        RECT 92.040 165.400 92.300 165.720 ;
        RECT 91.880 164.865 93.760 165.235 ;
        RECT 93.940 164.020 94.080 166.080 ;
        RECT 93.880 163.700 94.140 164.020 ;
        RECT 91.120 162.680 91.380 163.000 ;
        RECT 88.820 160.300 89.080 160.620 ;
        RECT 88.360 159.960 88.620 160.280 ;
        RECT 84.670 158.405 84.950 158.775 ;
        RECT 88.420 158.580 88.560 159.960 ;
        RECT 88.880 158.580 89.020 160.300 ;
        RECT 84.740 155.860 84.880 158.405 ;
        RECT 88.360 158.260 88.620 158.580 ;
        RECT 88.820 158.260 89.080 158.580 ;
        RECT 91.180 158.240 91.320 162.680 ;
        RECT 94.860 161.980 95.000 166.080 ;
        RECT 96.640 165.400 96.900 165.720 ;
        RECT 94.800 161.660 95.060 161.980 ;
        RECT 94.340 161.320 94.600 161.640 ;
        RECT 91.880 159.425 93.760 159.795 ;
        RECT 94.400 159.260 94.540 161.320 ;
        RECT 94.340 158.940 94.600 159.260 ;
        RECT 96.700 158.240 96.840 165.400 ;
        RECT 98.540 163.340 98.680 166.080 ;
        RECT 98.480 163.020 98.740 163.340 ;
        RECT 97.560 162.680 97.820 163.000 ;
        RECT 97.620 161.300 97.760 162.680 ;
        RECT 97.560 160.980 97.820 161.300 ;
        RECT 97.100 160.640 97.360 160.960 ;
        RECT 97.160 159.260 97.300 160.640 ;
        RECT 97.100 158.940 97.360 159.260 ;
        RECT 91.120 157.920 91.380 158.240 ;
        RECT 96.640 157.920 96.900 158.240 ;
        RECT 84.680 155.540 84.940 155.860 ;
        RECT 91.180 153.730 91.320 157.920 ;
        RECT 95.260 157.580 95.520 157.900 ;
        RECT 91.880 153.985 93.760 154.355 ;
        RECT 91.180 153.590 92.240 153.730 ;
        RECT 92.100 153.140 92.240 153.590 ;
        RECT 92.040 152.820 92.300 153.140 ;
        RECT 93.880 153.050 94.140 153.140 ;
        RECT 93.480 152.910 94.140 153.050 ;
        RECT 87.900 152.140 88.160 152.460 ;
        RECT 86.520 151.800 86.780 152.120 ;
        RECT 86.580 151.100 86.720 151.800 ;
        RECT 86.520 150.780 86.780 151.100 ;
        RECT 86.060 150.100 86.320 150.420 ;
        RECT 85.140 149.760 85.400 150.080 ;
        RECT 85.200 148.380 85.340 149.760 ;
        RECT 85.140 148.060 85.400 148.380 ;
        RECT 84.680 144.660 84.940 144.980 ;
        RECT 84.740 140.220 84.880 144.660 ;
        RECT 85.200 144.640 85.340 148.060 ;
        RECT 86.120 146.680 86.260 150.100 ;
        RECT 86.580 147.700 86.720 150.780 ;
        RECT 87.960 150.615 88.100 152.140 ;
        RECT 93.480 151.100 93.620 152.910 ;
        RECT 93.880 152.820 94.140 152.910 ;
        RECT 93.880 151.800 94.140 152.120 ;
        RECT 93.940 151.100 94.080 151.800 ;
        RECT 93.420 150.780 93.680 151.100 ;
        RECT 93.880 150.780 94.140 151.100 ;
        RECT 87.890 150.245 88.170 150.615 ;
        RECT 93.880 149.420 94.140 149.740 ;
        RECT 94.340 149.420 94.600 149.740 ;
        RECT 90.660 149.080 90.920 149.400 ;
        RECT 86.520 147.380 86.780 147.700 ;
        RECT 90.720 147.020 90.860 149.080 ;
        RECT 91.880 148.545 93.760 148.915 ;
        RECT 91.120 147.380 91.380 147.700 ;
        RECT 90.660 146.700 90.920 147.020 ;
        RECT 86.060 146.360 86.320 146.680 ;
        RECT 86.120 145.660 86.260 146.360 ;
        RECT 91.180 145.660 91.320 147.380 ;
        RECT 93.940 147.020 94.080 149.420 ;
        RECT 94.400 147.360 94.540 149.420 ;
        RECT 95.320 147.360 95.460 157.580 ;
        RECT 98.540 155.860 98.680 163.020 ;
        RECT 100.380 159.260 100.520 166.760 ;
        RECT 100.320 158.940 100.580 159.260 ;
        RECT 98.480 155.540 98.740 155.860 ;
        RECT 98.940 155.540 99.200 155.860 ;
        RECT 99.000 153.820 99.140 155.540 ;
        RECT 99.860 154.520 100.120 154.840 ;
        RECT 98.940 153.500 99.200 153.820 ;
        RECT 95.720 150.440 95.980 150.760 ;
        RECT 95.780 148.380 95.920 150.440 ;
        RECT 99.390 150.245 99.670 150.615 ;
        RECT 96.640 149.080 96.900 149.400 ;
        RECT 96.700 148.380 96.840 149.080 ;
        RECT 95.720 148.060 95.980 148.380 ;
        RECT 96.640 148.060 96.900 148.380 ;
        RECT 94.340 147.040 94.600 147.360 ;
        RECT 95.260 147.040 95.520 147.360 ;
        RECT 93.880 146.700 94.140 147.020 ;
        RECT 86.060 145.340 86.320 145.660 ;
        RECT 91.120 145.340 91.380 145.660 ;
        RECT 85.140 144.320 85.400 144.640 ;
        RECT 84.680 139.900 84.940 140.220 ;
        RECT 84.740 137.500 84.880 139.900 ;
        RECT 85.200 139.200 85.340 144.320 ;
        RECT 91.880 143.105 93.760 143.475 ;
        RECT 86.520 139.220 86.780 139.540 ;
        RECT 85.140 138.880 85.400 139.200 ;
        RECT 85.200 137.500 85.340 138.880 ;
        RECT 84.680 137.180 84.940 137.500 ;
        RECT 85.140 137.180 85.400 137.500 ;
        RECT 86.580 136.820 86.720 139.220 ;
        RECT 94.400 138.860 94.540 147.040 ;
        RECT 96.700 144.980 96.840 148.060 ;
        RECT 97.100 146.360 97.360 146.680 ;
        RECT 97.160 145.660 97.300 146.360 ;
        RECT 97.100 145.340 97.360 145.660 ;
        RECT 96.640 144.660 96.900 144.980 ;
        RECT 98.940 138.880 99.200 139.200 ;
        RECT 94.340 138.540 94.600 138.860 ;
        RECT 91.120 138.200 91.380 138.520 ;
        RECT 86.980 136.840 87.240 137.160 ;
        RECT 86.520 136.500 86.780 136.820 ;
        RECT 84.220 135.820 84.480 136.140 ;
        RECT 85.140 135.480 85.400 135.800 ;
        RECT 85.200 134.440 85.340 135.480 ;
        RECT 85.140 134.120 85.400 134.440 ;
        RECT 86.580 133.760 86.720 136.500 ;
        RECT 83.760 133.440 84.020 133.760 ;
        RECT 86.520 133.440 86.780 133.760 ;
        RECT 83.300 132.760 83.560 133.080 ;
        RECT 83.360 129.340 83.500 132.760 ;
        RECT 83.300 129.020 83.560 129.340 ;
        RECT 81.920 127.320 82.180 127.640 ;
        RECT 83.760 127.320 84.020 127.640 ;
        RECT 84.680 127.320 84.940 127.640 ;
        RECT 80.540 126.300 80.800 126.620 ;
        RECT 82.840 124.940 83.100 125.260 ;
        RECT 82.900 123.900 83.040 124.940 ;
        RECT 82.840 123.580 83.100 123.900 ;
        RECT 83.820 123.220 83.960 127.320 ;
        RECT 84.740 125.940 84.880 127.320 ;
        RECT 84.680 125.620 84.940 125.940 ;
        RECT 85.600 125.280 85.860 125.600 ;
        RECT 85.660 123.900 85.800 125.280 ;
        RECT 85.600 123.580 85.860 123.900 ;
        RECT 83.300 122.900 83.560 123.220 ;
        RECT 83.760 122.900 84.020 123.220 ;
        RECT 83.360 120.160 83.500 122.900 ;
        RECT 83.760 120.180 84.020 120.500 ;
        RECT 83.300 119.840 83.560 120.160 ;
        RECT 79.620 119.590 80.280 119.730 ;
        RECT 79.620 119.500 79.880 119.590 ;
        RECT 79.160 119.160 79.420 119.480 ;
        RECT 76.880 118.625 78.760 118.995 ;
        RECT 79.220 118.460 79.360 119.160 ;
        RECT 79.160 118.140 79.420 118.460 ;
        RECT 79.680 117.440 79.820 119.500 ;
        RECT 81.000 119.160 81.260 119.480 ;
        RECT 82.840 119.160 83.100 119.480 ;
        RECT 81.060 117.780 81.200 119.160 ;
        RECT 81.000 117.460 81.260 117.780 ;
        RECT 79.620 117.120 79.880 117.440 ;
        RECT 79.680 115.740 79.820 117.120 ;
        RECT 79.620 115.420 79.880 115.740 ;
        RECT 82.900 114.380 83.040 119.160 ;
        RECT 83.360 118.120 83.500 119.840 ;
        RECT 83.300 117.800 83.560 118.120 ;
        RECT 83.820 117.100 83.960 120.180 ;
        RECT 84.220 119.840 84.480 120.160 ;
        RECT 84.280 118.460 84.420 119.840 ;
        RECT 84.680 119.160 84.940 119.480 ;
        RECT 84.220 118.140 84.480 118.460 ;
        RECT 83.760 116.780 84.020 117.100 ;
        RECT 84.740 115.060 84.880 119.160 ;
        RECT 85.600 117.120 85.860 117.440 ;
        RECT 85.660 115.060 85.800 117.120 ;
        RECT 84.680 114.740 84.940 115.060 ;
        RECT 85.600 114.740 85.860 115.060 ;
        RECT 86.520 114.740 86.780 115.060 ;
        RECT 82.840 114.060 83.100 114.380 ;
        RECT 76.880 113.185 78.760 113.555 ;
        RECT 78.240 112.020 78.500 112.340 ;
        RECT 81.460 112.020 81.720 112.340 ;
        RECT 78.300 109.280 78.440 112.020 ;
        RECT 81.520 109.620 81.660 112.020 ;
        RECT 81.920 111.680 82.180 112.000 ;
        RECT 81.460 109.300 81.720 109.620 ;
        RECT 78.240 108.960 78.500 109.280 ;
        RECT 79.160 108.960 79.420 109.280 ;
        RECT 75.940 108.620 76.200 108.940 ;
        RECT 76.880 107.745 78.760 108.115 ;
        RECT 75.020 106.580 75.280 106.900 ;
        RECT 68.580 106.470 68.840 106.560 ;
        RECT 68.180 106.330 68.840 106.470 ;
        RECT 64.440 105.900 64.700 106.220 ;
        RECT 63.980 105.560 64.240 105.880 ;
        RECT 61.880 105.025 63.760 105.395 ;
        RECT 64.040 104.180 64.180 105.560 ;
        RECT 52.480 103.520 52.740 103.840 ;
        RECT 56.680 103.500 56.820 104.120 ;
        RECT 58.000 103.860 58.260 104.180 ;
        RECT 63.980 103.860 64.240 104.180 ;
        RECT 64.500 103.500 64.640 105.900 ;
        RECT 54.780 103.180 55.040 103.500 ;
        RECT 56.620 103.180 56.880 103.500 ;
        RECT 61.220 103.180 61.480 103.500 ;
        RECT 64.440 103.180 64.700 103.500 ;
        RECT 50.170 89.040 50.450 89.170 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.480 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 54.840 88.620 54.980 103.180 ;
        RECT 61.280 98.820 61.420 103.180 ;
        RECT 61.880 99.585 63.760 99.955 ;
        RECT 61.280 98.680 62.340 98.820 ;
        RECT 55.530 88.620 56.750 89.190 ;
        RECT 62.200 89.170 62.340 98.680 ;
        RECT 68.180 89.840 68.320 106.330 ;
        RECT 68.580 106.240 68.840 106.330 ;
        RECT 73.640 106.240 73.900 106.560 ;
        RECT 73.700 104.860 73.840 106.240 ;
        RECT 75.940 105.560 76.200 105.880 ;
        RECT 73.640 104.540 73.900 104.860 ;
        RECT 73.700 104.180 73.840 104.540 ;
        RECT 76.000 104.180 76.140 105.560 ;
        RECT 79.220 104.860 79.360 108.960 ;
        RECT 79.620 108.280 79.880 108.600 ;
        RECT 79.160 104.540 79.420 104.860 ;
        RECT 73.640 103.860 73.900 104.180 ;
        RECT 75.940 103.860 76.200 104.180 ;
        RECT 79.680 103.840 79.820 108.280 ;
        RECT 81.980 107.240 82.120 111.680 ;
        RECT 83.760 108.280 84.020 108.600 ;
        RECT 83.820 107.240 83.960 108.280 ;
        RECT 81.920 106.920 82.180 107.240 ;
        RECT 83.760 106.920 84.020 107.240 ;
        RECT 86.580 106.560 86.720 114.740 ;
        RECT 87.040 106.900 87.180 136.840 ;
        RECT 91.180 136.820 91.320 138.200 ;
        RECT 91.880 137.665 93.760 138.035 ;
        RECT 91.120 136.500 91.380 136.820 ;
        RECT 91.580 136.500 91.840 136.820 ;
        RECT 88.360 135.820 88.620 136.140 ;
        RECT 88.420 134.780 88.560 135.820 ;
        RECT 88.360 134.460 88.620 134.780 ;
        RECT 90.660 134.120 90.920 134.440 ;
        RECT 88.360 133.780 88.620 134.100 ;
        RECT 88.420 131.040 88.560 133.780 ;
        RECT 90.720 132.060 90.860 134.120 ;
        RECT 91.640 133.760 91.780 136.500 ;
        RECT 93.420 136.390 93.680 136.480 ;
        RECT 93.020 136.250 93.680 136.390 ;
        RECT 93.020 135.800 93.160 136.250 ;
        RECT 93.420 136.160 93.680 136.250 ;
        RECT 94.400 136.140 94.540 138.540 ;
        RECT 98.480 138.200 98.740 138.520 ;
        RECT 98.020 136.160 98.280 136.480 ;
        RECT 94.340 135.820 94.600 136.140 ;
        RECT 92.960 135.480 93.220 135.800 ;
        RECT 93.880 135.480 94.140 135.800 ;
        RECT 91.580 133.440 91.840 133.760 ;
        RECT 91.880 132.225 93.760 132.595 ;
        RECT 90.660 131.740 90.920 132.060 ;
        RECT 88.360 130.720 88.620 131.040 ;
        RECT 91.120 130.720 91.380 131.040 ;
        RECT 88.360 129.020 88.620 129.340 ;
        RECT 88.420 125.940 88.560 129.020 ;
        RECT 88.360 125.620 88.620 125.940 ;
        RECT 91.180 123.220 91.320 130.720 ;
        RECT 93.940 128.660 94.080 135.480 ;
        RECT 98.080 134.100 98.220 136.160 ;
        RECT 98.540 136.140 98.680 138.200 ;
        RECT 99.000 136.480 99.140 138.880 ;
        RECT 99.460 136.480 99.600 150.245 ;
        RECT 98.940 136.160 99.200 136.480 ;
        RECT 99.400 136.160 99.660 136.480 ;
        RECT 98.480 135.820 98.740 136.140 ;
        RECT 98.540 134.100 98.680 135.820 ;
        RECT 99.460 134.295 99.600 136.160 ;
        RECT 98.020 133.780 98.280 134.100 ;
        RECT 98.480 133.780 98.740 134.100 ;
        RECT 99.390 133.925 99.670 134.295 ;
        RECT 99.920 134.100 100.060 154.520 ;
        RECT 100.320 136.160 100.580 136.480 ;
        RECT 100.380 134.780 100.520 136.160 ;
        RECT 100.320 134.460 100.580 134.780 ;
        RECT 99.860 133.780 100.120 134.100 ;
        RECT 95.260 133.440 95.520 133.760 ;
        RECT 94.800 132.760 95.060 133.080 ;
        RECT 93.880 128.340 94.140 128.660 ;
        RECT 91.640 127.980 94.080 128.060 ;
        RECT 91.580 127.920 94.080 127.980 ;
        RECT 91.580 127.660 91.840 127.920 ;
        RECT 91.880 126.785 93.760 127.155 ;
        RECT 93.420 124.940 93.680 125.260 ;
        RECT 93.480 123.900 93.620 124.940 ;
        RECT 93.420 123.580 93.680 123.900 ;
        RECT 91.120 122.900 91.380 123.220 ;
        RECT 91.880 121.345 93.760 121.715 ;
        RECT 93.420 119.840 93.680 120.160 ;
        RECT 87.440 119.160 87.700 119.480 ;
        RECT 87.500 117.780 87.640 119.160 ;
        RECT 93.480 118.460 93.620 119.840 ;
        RECT 93.940 119.480 94.080 127.920 ;
        RECT 93.880 119.160 94.140 119.480 ;
        RECT 93.420 118.140 93.680 118.460 ;
        RECT 87.440 117.460 87.700 117.780 ;
        RECT 93.940 117.440 94.080 119.160 ;
        RECT 93.880 117.120 94.140 117.440 ;
        RECT 88.360 116.440 88.620 116.760 ;
        RECT 91.120 116.440 91.380 116.760 ;
        RECT 88.420 115.060 88.560 116.440 ;
        RECT 88.360 114.740 88.620 115.060 ;
        RECT 91.180 114.380 91.320 116.440 ;
        RECT 91.880 115.905 93.760 116.275 ;
        RECT 93.940 115.740 94.080 117.120 ;
        RECT 93.880 115.420 94.140 115.740 ;
        RECT 91.120 114.060 91.380 114.380 ;
        RECT 92.950 112.845 93.230 113.215 ;
        RECT 93.020 112.680 93.160 112.845 ;
        RECT 92.960 112.360 93.220 112.680 ;
        RECT 91.880 110.465 93.760 110.835 ;
        RECT 94.860 109.280 95.000 132.760 ;
        RECT 95.320 129.340 95.460 133.440 ;
        RECT 98.540 131.040 98.680 133.780 ;
        RECT 100.840 133.760 100.980 176.280 ;
        RECT 101.230 163.845 101.510 164.215 ;
        RECT 101.300 163.680 101.440 163.845 ;
        RECT 101.240 163.360 101.500 163.680 ;
        RECT 101.700 151.800 101.960 152.120 ;
        RECT 101.240 135.480 101.500 135.800 ;
        RECT 101.300 134.440 101.440 135.480 ;
        RECT 101.240 134.120 101.500 134.440 ;
        RECT 100.780 133.440 101.040 133.760 ;
        RECT 99.860 132.760 100.120 133.080 ;
        RECT 101.240 132.760 101.500 133.080 ;
        RECT 98.480 130.720 98.740 131.040 ;
        RECT 95.260 129.020 95.520 129.340 ;
        RECT 95.710 129.165 95.990 129.535 ;
        RECT 98.540 129.340 98.680 130.720 ;
        RECT 95.780 129.000 95.920 129.165 ;
        RECT 98.480 129.020 98.740 129.340 ;
        RECT 95.720 128.680 95.980 129.000 ;
        RECT 98.540 125.940 98.680 129.020 ;
        RECT 98.940 128.000 99.200 128.320 ;
        RECT 99.000 126.620 99.140 128.000 ;
        RECT 98.940 126.300 99.200 126.620 ;
        RECT 98.480 125.620 98.740 125.940 ;
        RECT 99.400 125.280 99.660 125.600 ;
        RECT 99.460 120.160 99.600 125.280 ;
        RECT 99.400 119.840 99.660 120.160 ;
        RECT 99.920 109.280 100.060 132.760 ;
        RECT 100.320 131.400 100.580 131.720 ;
        RECT 100.380 128.660 100.520 131.400 ;
        RECT 100.320 128.340 100.580 128.660 ;
        RECT 100.380 125.600 100.520 128.340 ;
        RECT 101.300 125.600 101.440 132.760 ;
        RECT 100.320 125.280 100.580 125.600 ;
        RECT 101.240 125.280 101.500 125.600 ;
        RECT 100.320 122.900 100.580 123.220 ;
        RECT 100.380 120.160 100.520 122.900 ;
        RECT 100.320 119.840 100.580 120.160 ;
        RECT 101.240 119.160 101.500 119.480 ;
        RECT 100.320 117.120 100.580 117.440 ;
        RECT 100.380 115.740 100.520 117.120 ;
        RECT 100.320 115.420 100.580 115.740 ;
        RECT 101.300 114.720 101.440 119.160 ;
        RECT 101.240 114.400 101.500 114.720 ;
        RECT 101.760 114.040 101.900 151.800 ;
        RECT 102.220 133.760 102.360 176.280 ;
        RECT 102.620 168.120 102.880 168.440 ;
        RECT 102.680 161.300 102.820 168.120 ;
        RECT 102.620 160.980 102.880 161.300 ;
        RECT 102.680 160.140 102.820 160.980 ;
        RECT 102.680 160.000 103.280 160.140 ;
        RECT 102.620 156.220 102.880 156.540 ;
        RECT 102.680 155.180 102.820 156.220 ;
        RECT 103.140 156.200 103.280 160.000 ;
        RECT 103.080 155.880 103.340 156.200 ;
        RECT 102.620 154.860 102.880 155.180 ;
        RECT 103.080 153.730 103.340 153.820 ;
        RECT 102.680 153.590 103.340 153.730 ;
        RECT 102.680 147.100 102.820 153.590 ;
        RECT 103.080 153.500 103.340 153.590 ;
        RECT 103.600 151.180 103.740 182.320 ;
        RECT 104.920 181.720 105.180 182.040 ;
        RECT 104.980 180.340 105.120 181.720 ;
        RECT 104.920 180.020 105.180 180.340 ;
        RECT 104.920 174.470 105.180 174.560 ;
        RECT 105.440 174.470 105.580 185.460 ;
        RECT 105.840 185.120 106.100 185.440 ;
        RECT 105.900 183.740 106.040 185.120 ;
        RECT 106.880 183.905 108.760 184.275 ;
        RECT 105.840 183.420 106.100 183.740 ;
        RECT 105.840 182.740 106.100 183.060 ;
        RECT 106.300 182.740 106.560 183.060 ;
        RECT 108.140 182.740 108.400 183.060 ;
        RECT 109.520 182.740 109.780 183.060 ;
        RECT 105.900 181.020 106.040 182.740 ;
        RECT 105.840 180.700 106.100 181.020 ;
        RECT 105.840 180.020 106.100 180.340 ;
        RECT 105.900 177.280 106.040 180.020 ;
        RECT 106.360 177.530 106.500 182.740 ;
        RECT 108.200 180.340 108.340 182.740 ;
        RECT 108.140 180.020 108.400 180.340 ;
        RECT 109.060 179.680 109.320 180.000 ;
        RECT 106.880 178.465 108.760 178.835 ;
        RECT 109.120 177.960 109.260 179.680 ;
        RECT 109.060 177.640 109.320 177.960 ;
        RECT 109.580 177.620 109.720 182.740 ;
        RECT 106.760 177.530 107.020 177.620 ;
        RECT 106.360 177.390 107.020 177.530 ;
        RECT 106.760 177.300 107.020 177.390 ;
        RECT 108.140 177.300 108.400 177.620 ;
        RECT 109.520 177.300 109.780 177.620 ;
        RECT 105.840 176.960 106.100 177.280 ;
        RECT 105.900 174.560 106.040 176.960 ;
        RECT 106.300 175.260 106.560 175.580 ;
        RECT 104.920 174.330 105.580 174.470 ;
        RECT 104.920 174.240 105.180 174.330 ;
        RECT 105.840 174.240 106.100 174.560 ;
        RECT 104.460 173.900 104.720 174.220 ;
        RECT 104.000 154.520 104.260 154.840 ;
        RECT 103.140 151.040 103.740 151.180 ;
        RECT 103.140 147.700 103.280 151.040 ;
        RECT 103.540 150.440 103.800 150.760 ;
        RECT 103.600 148.380 103.740 150.440 ;
        RECT 103.540 148.060 103.800 148.380 ;
        RECT 103.080 147.380 103.340 147.700 ;
        RECT 102.680 146.960 103.280 147.100 ;
        RECT 102.620 139.560 102.880 139.880 ;
        RECT 102.680 134.780 102.820 139.560 ;
        RECT 102.620 134.460 102.880 134.780 ;
        RECT 102.620 133.780 102.880 134.100 ;
        RECT 102.160 133.440 102.420 133.760 ;
        RECT 102.680 131.720 102.820 133.780 ;
        RECT 102.620 131.400 102.880 131.720 ;
        RECT 103.140 127.980 103.280 146.960 ;
        RECT 104.060 134.100 104.200 154.520 ;
        RECT 104.520 153.140 104.660 173.900 ;
        RECT 106.360 172.520 106.500 175.260 ;
        RECT 106.820 174.900 106.960 177.300 ;
        RECT 108.200 175.580 108.340 177.300 ;
        RECT 108.140 175.260 108.400 175.580 ;
        RECT 109.060 174.920 109.320 175.240 ;
        RECT 106.760 174.580 107.020 174.900 ;
        RECT 106.880 173.025 108.760 173.395 ;
        RECT 106.300 172.200 106.560 172.520 ;
        RECT 105.840 171.520 106.100 171.840 ;
        RECT 105.900 166.400 106.040 171.520 ;
        RECT 107.220 170.840 107.480 171.160 ;
        RECT 107.280 168.780 107.420 170.840 ;
        RECT 107.220 168.460 107.480 168.780 ;
        RECT 106.880 167.585 108.760 167.955 ;
        RECT 104.920 166.080 105.180 166.400 ;
        RECT 105.840 166.080 106.100 166.400 ;
        RECT 104.980 159.260 105.120 166.080 ;
        RECT 105.380 162.680 105.640 163.000 ;
        RECT 104.920 158.940 105.180 159.260 ;
        RECT 105.440 158.240 105.580 162.680 ;
        RECT 105.900 160.960 106.040 166.080 ;
        RECT 109.120 166.060 109.260 174.920 ;
        RECT 110.040 174.560 110.180 188.180 ;
        RECT 110.440 185.120 110.700 185.440 ;
        RECT 110.500 182.380 110.640 185.120 ;
        RECT 110.960 182.720 111.100 193.280 ;
        RECT 112.280 192.940 112.540 193.260 ;
        RECT 112.340 185.100 112.480 192.940 ;
        RECT 112.800 191.900 112.940 194.300 ;
        RECT 115.960 193.620 116.220 193.940 ;
        RECT 112.740 191.580 113.000 191.900 ;
        RECT 113.200 189.880 113.460 190.200 ;
        RECT 113.260 188.500 113.400 189.880 ;
        RECT 113.200 188.180 113.460 188.500 ;
        RECT 112.280 184.780 112.540 185.100 ;
        RECT 111.820 184.440 112.080 184.760 ;
        RECT 111.880 183.060 112.020 184.440 ;
        RECT 111.820 182.740 112.080 183.060 ;
        RECT 110.900 182.400 111.160 182.720 ;
        RECT 110.440 182.060 110.700 182.380 ;
        RECT 109.520 174.240 109.780 174.560 ;
        RECT 109.980 174.240 110.240 174.560 ;
        RECT 109.580 172.180 109.720 174.240 ;
        RECT 109.980 173.560 110.240 173.880 ;
        RECT 110.040 172.180 110.180 173.560 ;
        RECT 110.500 172.520 110.640 182.060 ;
        RECT 110.960 177.280 111.100 182.400 ;
        RECT 111.880 178.300 112.020 182.740 ;
        RECT 112.340 178.300 112.480 184.780 ;
        RECT 116.020 180.340 116.160 193.620 ;
        RECT 117.860 191.900 118.000 195.660 ;
        RECT 118.320 194.280 118.460 195.660 ;
        RECT 118.260 193.960 118.520 194.280 ;
        RECT 117.800 191.580 118.060 191.900 ;
        RECT 118.320 190.880 118.460 193.960 ;
        RECT 119.180 192.600 119.440 192.920 ;
        RECT 119.240 190.880 119.380 192.600 ;
        RECT 121.880 192.065 123.760 192.435 ;
        RECT 118.260 190.560 118.520 190.880 ;
        RECT 119.180 190.560 119.440 190.880 ;
        RECT 116.420 190.220 116.680 190.540 ;
        RECT 116.480 189.180 116.620 190.220 ;
        RECT 116.420 188.860 116.680 189.180 ;
        RECT 118.320 188.160 118.460 190.560 ;
        RECT 118.260 187.840 118.520 188.160 ;
        RECT 117.800 182.740 118.060 183.060 ;
        RECT 116.880 181.720 117.140 182.040 ;
        RECT 115.960 180.020 116.220 180.340 ;
        RECT 111.820 177.980 112.080 178.300 ;
        RECT 112.280 177.980 112.540 178.300 ;
        RECT 116.940 177.620 117.080 181.720 ;
        RECT 117.860 181.020 118.000 182.740 ;
        RECT 118.320 182.720 118.460 187.840 ;
        RECT 121.880 186.625 123.760 186.995 ;
        RECT 124.700 183.080 124.960 183.400 ;
        RECT 118.260 182.400 118.520 182.720 ;
        RECT 117.800 180.700 118.060 181.020 ;
        RECT 118.320 179.320 118.460 182.400 ;
        RECT 121.880 181.185 123.760 181.555 ;
        RECT 124.760 181.020 124.900 183.080 ;
        RECT 124.700 180.700 124.960 181.020 ;
        RECT 121.940 179.680 122.200 180.000 ;
        RECT 118.720 179.340 118.980 179.660 ;
        RECT 118.260 179.000 118.520 179.320 ;
        RECT 118.780 178.300 118.920 179.340 ;
        RECT 118.720 177.980 118.980 178.300 ;
        RECT 122.000 177.960 122.140 179.680 ;
        RECT 121.940 177.640 122.200 177.960 ;
        RECT 116.880 177.300 117.140 177.620 ;
        RECT 110.900 176.960 111.160 177.280 ;
        RECT 121.880 175.745 123.760 176.115 ;
        RECT 119.180 174.240 119.440 174.560 ;
        RECT 118.260 173.560 118.520 173.880 ;
        RECT 118.320 172.520 118.460 173.560 ;
        RECT 119.240 172.860 119.380 174.240 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 119.180 172.540 119.440 172.860 ;
        RECT 110.440 172.200 110.700 172.520 ;
        RECT 118.260 172.200 118.520 172.520 ;
        RECT 109.520 171.860 109.780 172.180 ;
        RECT 109.980 171.860 110.240 172.180 ;
        RECT 114.580 171.180 114.840 171.500 ;
        RECT 111.360 170.840 111.620 171.160 ;
        RECT 113.660 170.840 113.920 171.160 ;
        RECT 109.980 169.140 110.240 169.460 ;
        RECT 109.060 165.740 109.320 166.060 ;
        RECT 110.040 164.780 110.180 169.140 ;
        RECT 110.440 168.460 110.700 168.780 ;
        RECT 110.500 167.420 110.640 168.460 ;
        RECT 110.900 168.120 111.160 168.440 ;
        RECT 110.440 167.100 110.700 167.420 ;
        RECT 110.960 166.740 111.100 168.120 ;
        RECT 110.900 166.420 111.160 166.740 ;
        RECT 110.900 165.740 111.160 166.060 ;
        RECT 109.580 164.640 110.180 164.780 ;
        RECT 109.060 164.040 109.320 164.360 ;
        RECT 106.300 163.020 106.560 163.340 ;
        RECT 106.360 161.980 106.500 163.020 ;
        RECT 106.880 162.145 108.760 162.515 ;
        RECT 106.300 161.660 106.560 161.980 ;
        RECT 105.840 160.640 106.100 160.960 ;
        RECT 109.120 158.240 109.260 164.040 ;
        RECT 109.580 158.920 109.720 164.640 ;
        RECT 110.440 163.700 110.700 164.020 ;
        RECT 109.980 162.680 110.240 163.000 ;
        RECT 110.040 161.980 110.180 162.680 ;
        RECT 109.980 161.660 110.240 161.980 ;
        RECT 110.500 161.300 110.640 163.700 ;
        RECT 110.440 160.980 110.700 161.300 ;
        RECT 110.960 160.700 111.100 165.740 ;
        RECT 110.500 160.560 111.100 160.700 ;
        RECT 109.520 158.600 109.780 158.920 ;
        RECT 105.380 157.920 105.640 158.240 ;
        RECT 109.060 157.920 109.320 158.240 ;
        RECT 109.520 157.920 109.780 158.240 ;
        RECT 109.980 157.920 110.240 158.240 ;
        RECT 109.060 157.240 109.320 157.560 ;
        RECT 106.880 156.705 108.760 157.075 ;
        RECT 108.600 156.220 108.860 156.540 ;
        RECT 105.380 155.540 105.640 155.860 ;
        RECT 105.440 153.480 105.580 155.540 ;
        RECT 106.760 154.520 107.020 154.840 ;
        RECT 105.380 153.160 105.640 153.480 ;
        RECT 104.460 152.820 104.720 153.140 ;
        RECT 106.820 152.800 106.960 154.520 ;
        RECT 108.140 153.160 108.400 153.480 ;
        RECT 106.760 152.480 107.020 152.800 ;
        RECT 107.680 152.710 107.940 152.800 ;
        RECT 108.200 152.710 108.340 153.160 ;
        RECT 108.660 152.800 108.800 156.220 ;
        RECT 107.680 152.570 108.340 152.710 ;
        RECT 107.680 152.480 107.940 152.570 ;
        RECT 108.600 152.480 108.860 152.800 ;
        RECT 104.920 152.140 105.180 152.460 ;
        RECT 104.980 151.100 105.120 152.140 ;
        RECT 108.660 152.120 108.800 152.480 ;
        RECT 105.380 151.800 105.640 152.120 ;
        RECT 108.600 151.800 108.860 152.120 ;
        RECT 104.920 150.780 105.180 151.100 ;
        RECT 104.460 148.060 104.720 148.380 ;
        RECT 104.000 133.780 104.260 134.100 ;
        RECT 103.540 132.760 103.800 133.080 ;
        RECT 103.080 127.660 103.340 127.980 ;
        RECT 102.620 119.500 102.880 119.820 ;
        RECT 102.680 118.460 102.820 119.500 ;
        RECT 102.620 118.140 102.880 118.460 ;
        RECT 101.700 113.720 101.960 114.040 ;
        RECT 103.600 109.280 103.740 132.760 ;
        RECT 104.520 112.000 104.660 148.060 ;
        RECT 105.440 147.360 105.580 151.800 ;
        RECT 106.880 151.265 108.760 151.635 ;
        RECT 107.670 150.245 107.950 150.615 ;
        RECT 107.740 150.080 107.880 150.245 ;
        RECT 108.140 150.100 108.400 150.420 ;
        RECT 107.680 149.760 107.940 150.080 ;
        RECT 106.300 148.060 106.560 148.380 ;
        RECT 105.380 147.040 105.640 147.360 ;
        RECT 105.380 138.880 105.640 139.200 ;
        RECT 105.440 137.500 105.580 138.880 ;
        RECT 105.380 137.180 105.640 137.500 ;
        RECT 104.920 132.760 105.180 133.080 ;
        RECT 104.980 129.340 105.120 132.760 ;
        RECT 106.360 129.340 106.500 148.060 ;
        RECT 107.740 147.700 107.880 149.760 ;
        RECT 107.680 147.380 107.940 147.700 ;
        RECT 108.200 147.360 108.340 150.100 ;
        RECT 108.140 147.040 108.400 147.360 ;
        RECT 108.200 146.680 108.340 147.040 ;
        RECT 108.140 146.360 108.400 146.680 ;
        RECT 106.880 145.825 108.760 146.195 ;
        RECT 109.120 144.980 109.260 157.240 ;
        RECT 109.580 155.860 109.720 157.920 ;
        RECT 109.520 155.540 109.780 155.860 ;
        RECT 109.580 152.800 109.720 155.540 ;
        RECT 110.040 153.820 110.180 157.920 ;
        RECT 109.980 153.500 110.240 153.820 ;
        RECT 110.040 153.140 110.180 153.500 ;
        RECT 109.980 152.820 110.240 153.140 ;
        RECT 109.520 152.480 109.780 152.800 ;
        RECT 109.980 150.100 110.240 150.420 ;
        RECT 110.040 147.360 110.180 150.100 ;
        RECT 109.980 147.040 110.240 147.360 ;
        RECT 109.520 146.360 109.780 146.680 ;
        RECT 109.580 144.980 109.720 146.360 ;
        RECT 109.060 144.660 109.320 144.980 ;
        RECT 109.520 144.660 109.780 144.980 ;
        RECT 110.040 144.380 110.180 147.040 ;
        RECT 110.500 144.640 110.640 160.560 ;
        RECT 110.900 159.960 111.160 160.280 ;
        RECT 110.960 156.200 111.100 159.960 ;
        RECT 110.900 155.880 111.160 156.200 ;
        RECT 110.900 154.520 111.160 154.840 ;
        RECT 109.060 143.980 109.320 144.300 ;
        RECT 109.580 144.240 110.180 144.380 ;
        RECT 110.440 144.320 110.700 144.640 ;
        RECT 109.120 142.940 109.260 143.980 ;
        RECT 109.060 142.620 109.320 142.940 ;
        RECT 106.880 140.385 108.760 140.755 ;
        RECT 109.580 139.540 109.720 144.240 ;
        RECT 109.980 143.640 110.240 143.960 ;
        RECT 110.440 143.640 110.700 143.960 ;
        RECT 109.520 139.220 109.780 139.540 ;
        RECT 109.060 135.820 109.320 136.140 ;
        RECT 106.880 134.945 108.760 135.315 ;
        RECT 108.130 133.925 108.410 134.295 ;
        RECT 109.120 134.100 109.260 135.820 ;
        RECT 109.580 134.100 109.720 139.220 ;
        RECT 108.140 133.780 108.400 133.925 ;
        RECT 109.060 133.780 109.320 134.100 ;
        RECT 109.520 133.780 109.780 134.100 ;
        RECT 110.040 132.060 110.180 143.640 ;
        RECT 110.500 139.880 110.640 143.640 ;
        RECT 110.440 139.560 110.700 139.880 ;
        RECT 110.500 134.440 110.640 139.560 ;
        RECT 110.440 134.120 110.700 134.440 ;
        RECT 110.960 134.100 111.100 154.520 ;
        RECT 111.420 134.100 111.560 170.840 ;
        RECT 112.740 169.140 113.000 169.460 ;
        RECT 111.820 168.800 112.080 169.120 ;
        RECT 111.880 166.400 112.020 168.800 ;
        RECT 112.280 166.420 112.540 166.740 ;
        RECT 111.820 166.080 112.080 166.400 ;
        RECT 112.340 166.060 112.480 166.420 ;
        RECT 112.280 165.740 112.540 166.060 ;
        RECT 111.820 163.020 112.080 163.340 ;
        RECT 111.880 158.660 112.020 163.020 ;
        RECT 112.340 159.260 112.480 165.740 ;
        RECT 112.800 163.680 112.940 169.140 ;
        RECT 113.200 168.120 113.460 168.440 ;
        RECT 113.260 164.700 113.400 168.120 ;
        RECT 113.200 164.380 113.460 164.700 ;
        RECT 113.260 163.680 113.400 164.380 ;
        RECT 112.740 163.360 113.000 163.680 ;
        RECT 113.200 163.360 113.460 163.680 ;
        RECT 112.800 160.960 112.940 163.360 ;
        RECT 112.740 160.640 113.000 160.960 ;
        RECT 112.280 158.940 112.540 159.260 ;
        RECT 111.880 158.520 112.480 158.660 ;
        RECT 111.820 157.920 112.080 158.240 ;
        RECT 111.880 156.540 112.020 157.920 ;
        RECT 112.340 157.900 112.480 158.520 ;
        RECT 112.280 157.580 112.540 157.900 ;
        RECT 111.820 156.220 112.080 156.540 ;
        RECT 112.340 152.120 112.480 157.580 ;
        RECT 113.260 155.860 113.400 163.360 ;
        RECT 113.720 163.340 113.860 170.840 ;
        RECT 114.640 169.120 114.780 171.180 ;
        RECT 117.340 170.840 117.600 171.160 ;
        RECT 117.400 169.460 117.540 170.840 ;
        RECT 117.340 169.140 117.600 169.460 ;
        RECT 114.580 168.800 114.840 169.120 ;
        RECT 114.120 165.400 114.380 165.720 ;
        RECT 113.660 163.020 113.920 163.340 ;
        RECT 114.180 161.300 114.320 165.400 ;
        RECT 114.120 160.980 114.380 161.300 ;
        RECT 113.200 155.540 113.460 155.860 ;
        RECT 114.640 153.480 114.780 168.800 ;
        RECT 117.400 161.980 117.540 169.140 ;
        RECT 116.420 161.660 116.680 161.980 ;
        RECT 117.340 161.660 117.600 161.980 ;
        RECT 114.580 153.160 114.840 153.480 ;
        RECT 116.480 153.140 116.620 161.660 ;
        RECT 119.240 161.300 119.380 172.540 ;
        RECT 121.480 171.520 121.740 171.840 ;
        RECT 124.700 171.520 124.960 171.840 ;
        RECT 121.540 170.140 121.680 171.520 ;
        RECT 121.880 170.305 123.760 170.675 ;
        RECT 121.480 169.820 121.740 170.140 ;
        RECT 119.640 166.760 119.900 167.080 ;
        RECT 119.700 161.980 119.840 166.760 ;
        RECT 124.760 166.740 124.900 171.520 ;
        RECT 127.910 171.325 128.190 171.695 ;
        RECT 127.980 169.120 128.120 171.325 ;
        RECT 129.290 170.560 133.760 172.150 ;
        RECT 127.920 168.800 128.180 169.120 ;
        RECT 124.700 166.420 124.960 166.740 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 121.480 165.400 121.740 165.720 ;
        RECT 121.540 161.980 121.680 165.400 ;
        RECT 121.880 164.865 123.760 165.235 ;
        RECT 124.760 164.020 124.900 166.420 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 124.700 163.700 124.960 164.020 ;
        RECT 123.780 163.360 124.040 163.680 ;
        RECT 119.640 161.660 119.900 161.980 ;
        RECT 121.480 161.660 121.740 161.980 ;
        RECT 123.840 161.640 123.980 163.360 ;
        RECT 123.780 161.320 124.040 161.640 ;
        RECT 119.180 160.980 119.440 161.300 ;
        RECT 121.020 160.980 121.280 161.300 ;
        RECT 116.880 159.960 117.140 160.280 ;
        RECT 116.940 158.580 117.080 159.960 ;
        RECT 121.080 159.260 121.220 160.980 ;
        RECT 121.880 159.425 123.760 159.795 ;
        RECT 121.020 158.940 121.280 159.260 ;
        RECT 116.880 158.260 117.140 158.580 ;
        RECT 117.800 155.200 118.060 155.520 ;
        RECT 116.420 152.820 116.680 153.140 ;
        RECT 115.960 152.140 116.220 152.460 ;
        RECT 112.280 151.800 112.540 152.120 ;
        RECT 111.820 149.420 112.080 149.740 ;
        RECT 111.880 144.980 112.020 149.420 ;
        RECT 114.120 149.080 114.380 149.400 ;
        RECT 113.200 147.380 113.460 147.700 ;
        RECT 112.280 147.040 112.540 147.360 ;
        RECT 111.820 144.660 112.080 144.980 ;
        RECT 112.340 144.890 112.480 147.040 ;
        RECT 112.740 144.890 113.000 144.980 ;
        RECT 112.340 144.750 113.000 144.890 ;
        RECT 112.740 144.660 113.000 144.750 ;
        RECT 111.880 143.700 112.020 144.660 ;
        RECT 113.260 144.550 113.400 147.380 ;
        RECT 114.180 146.680 114.320 149.080 ;
        RECT 116.020 148.380 116.160 152.140 ;
        RECT 116.880 150.670 117.140 150.760 ;
        RECT 117.860 150.670 118.000 155.200 ;
        RECT 121.880 153.985 123.760 154.355 ;
        RECT 119.640 152.480 119.900 152.800 ;
        RECT 118.260 151.800 118.520 152.120 ;
        RECT 118.320 150.760 118.460 151.800 ;
        RECT 116.880 150.530 118.000 150.670 ;
        RECT 116.880 150.440 117.140 150.530 ;
        RECT 115.960 148.060 116.220 148.380 ;
        RECT 117.860 147.610 118.000 150.530 ;
        RECT 118.260 150.440 118.520 150.760 ;
        RECT 117.860 147.470 118.460 147.610 ;
        RECT 117.800 146.700 118.060 147.020 ;
        RECT 114.120 146.360 114.380 146.680 ;
        RECT 117.340 146.360 117.600 146.680 ;
        RECT 117.400 145.660 117.540 146.360 ;
        RECT 117.340 145.340 117.600 145.660 ;
        RECT 117.860 144.640 118.000 146.700 ;
        RECT 113.660 144.550 113.920 144.640 ;
        RECT 113.260 144.410 113.920 144.550 ;
        RECT 111.880 143.560 112.940 143.700 ;
        RECT 111.820 142.620 112.080 142.940 ;
        RECT 110.900 133.780 111.160 134.100 ;
        RECT 111.360 133.780 111.620 134.100 ;
        RECT 110.440 132.760 110.700 133.080 ;
        RECT 111.360 132.760 111.620 133.080 ;
        RECT 109.980 131.740 110.240 132.060 ;
        RECT 106.880 129.505 108.760 129.875 ;
        RECT 104.920 129.020 105.180 129.340 ;
        RECT 106.300 129.020 106.560 129.340 ;
        RECT 106.300 128.340 106.560 128.660 ;
        RECT 105.380 128.000 105.640 128.320 ;
        RECT 105.440 125.600 105.580 128.000 ;
        RECT 105.380 125.280 105.640 125.600 ;
        RECT 105.380 122.560 105.640 122.880 ;
        RECT 105.440 120.500 105.580 122.560 ;
        RECT 105.380 120.180 105.640 120.500 ;
        RECT 106.360 119.820 106.500 128.340 ;
        RECT 109.520 128.000 109.780 128.320 ;
        RECT 106.880 124.065 108.760 124.435 ;
        RECT 109.580 120.500 109.720 128.000 ;
        RECT 109.520 120.180 109.780 120.500 ;
        RECT 106.300 119.500 106.560 119.820 ;
        RECT 105.840 119.160 106.100 119.480 ;
        RECT 109.060 119.160 109.320 119.480 ;
        RECT 105.900 118.120 106.040 119.160 ;
        RECT 106.880 118.625 108.760 118.995 ;
        RECT 105.840 117.800 106.100 118.120 ;
        RECT 109.120 114.720 109.260 119.160 ;
        RECT 109.580 114.720 109.720 120.180 ;
        RECT 109.980 117.460 110.240 117.780 ;
        RECT 110.040 115.740 110.180 117.460 ;
        RECT 109.980 115.420 110.240 115.740 ;
        RECT 109.060 114.400 109.320 114.720 ;
        RECT 109.520 114.400 109.780 114.720 ;
        RECT 106.880 113.185 108.760 113.555 ;
        RECT 104.460 111.680 104.720 112.000 ;
        RECT 110.500 109.280 110.640 132.760 ;
        RECT 110.900 130.720 111.160 131.040 ;
        RECT 110.960 128.660 111.100 130.720 ;
        RECT 111.420 129.340 111.560 132.760 ;
        RECT 111.360 129.020 111.620 129.340 ;
        RECT 111.880 128.740 112.020 142.620 ;
        RECT 112.280 139.560 112.540 139.880 ;
        RECT 112.340 134.440 112.480 139.560 ;
        RECT 112.800 139.540 112.940 143.560 ;
        RECT 113.260 142.260 113.400 144.410 ;
        RECT 113.660 144.320 113.920 144.410 ;
        RECT 117.800 144.320 118.060 144.640 ;
        RECT 113.200 141.940 113.460 142.260 ;
        RECT 112.740 139.220 113.000 139.540 ;
        RECT 112.740 138.540 113.000 138.860 ;
        RECT 112.800 136.480 112.940 138.540 ;
        RECT 113.260 137.160 113.400 141.940 ;
        RECT 117.860 141.920 118.000 144.320 ;
        RECT 117.800 141.600 118.060 141.920 ;
        RECT 117.340 140.920 117.600 141.240 ;
        RECT 117.400 139.880 117.540 140.920 ;
        RECT 117.340 139.560 117.600 139.880 ;
        RECT 115.960 139.220 116.220 139.540 ;
        RECT 113.200 136.840 113.460 137.160 ;
        RECT 112.740 136.160 113.000 136.480 ;
        RECT 116.020 136.140 116.160 139.220 ;
        RECT 115.960 135.820 116.220 136.140 ;
        RECT 113.200 135.480 113.460 135.800 ;
        RECT 112.280 134.120 112.540 134.440 ;
        RECT 113.260 134.100 113.400 135.480 ;
        RECT 113.200 133.780 113.460 134.100 ;
        RECT 118.320 131.720 118.460 147.470 ;
        RECT 119.700 144.980 119.840 152.480 ;
        RECT 123.320 151.800 123.580 152.120 ;
        RECT 123.380 150.760 123.520 151.800 ;
        RECT 123.320 150.440 123.580 150.760 ;
        RECT 126.080 149.760 126.340 150.080 ;
        RECT 121.880 148.545 123.760 148.915 ;
        RECT 126.140 147.360 126.280 149.760 ;
        RECT 123.780 147.040 124.040 147.360 ;
        RECT 126.080 147.040 126.340 147.360 ;
        RECT 120.100 146.700 120.360 147.020 ;
        RECT 120.160 145.660 120.300 146.700 ;
        RECT 123.840 145.660 123.980 147.040 ;
        RECT 120.100 145.340 120.360 145.660 ;
        RECT 123.780 145.340 124.040 145.660 ;
        RECT 119.640 144.660 119.900 144.980 ;
        RECT 119.700 141.920 119.840 144.660 ;
        RECT 121.880 143.105 123.760 143.475 ;
        RECT 119.640 141.660 119.900 141.920 ;
        RECT 119.640 141.600 120.300 141.660 ;
        RECT 119.700 141.520 120.300 141.600 ;
        RECT 119.640 140.920 119.900 141.240 ;
        RECT 119.700 137.500 119.840 140.920 ;
        RECT 120.160 138.860 120.300 141.520 ;
        RECT 120.560 140.920 120.820 141.240 ;
        RECT 120.620 139.880 120.760 140.920 ;
        RECT 120.560 139.560 120.820 139.880 ;
        RECT 124.240 139.220 124.500 139.540 ;
        RECT 120.100 138.540 120.360 138.860 ;
        RECT 121.480 138.200 121.740 138.520 ;
        RECT 119.640 137.180 119.900 137.500 ;
        RECT 121.540 136.820 121.680 138.200 ;
        RECT 121.880 137.665 123.760 138.035 ;
        RECT 124.300 137.500 124.440 139.220 ;
        RECT 126.140 139.200 126.280 147.040 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 126.080 138.880 126.340 139.200 ;
        RECT 124.700 138.200 124.960 138.520 ;
        RECT 124.240 137.180 124.500 137.500 ;
        RECT 121.480 136.500 121.740 136.820 ;
        RECT 121.020 136.160 121.280 136.480 ;
        RECT 121.080 134.780 121.220 136.160 ;
        RECT 121.020 134.460 121.280 134.780 ;
        RECT 121.880 132.225 123.760 132.595 ;
        RECT 118.260 131.400 118.520 131.720 ;
        RECT 112.280 130.720 112.540 131.040 ;
        RECT 110.900 128.340 111.160 128.660 ;
        RECT 111.420 128.600 112.020 128.740 ;
        RECT 110.900 109.640 111.160 109.960 ;
        RECT 94.800 108.960 95.060 109.280 ;
        RECT 99.860 108.960 100.120 109.280 ;
        RECT 103.540 108.960 103.800 109.280 ;
        RECT 110.440 108.960 110.700 109.280 ;
        RECT 102.620 108.620 102.880 108.940 ;
        RECT 87.900 108.280 88.160 108.600 ;
        RECT 92.960 108.280 93.220 108.600 ;
        RECT 98.020 108.280 98.280 108.600 ;
        RECT 99.860 108.280 100.120 108.600 ;
        RECT 86.980 106.580 87.240 106.900 ;
        RECT 80.080 106.240 80.340 106.560 ;
        RECT 86.520 106.240 86.780 106.560 ;
        RECT 79.620 103.520 79.880 103.840 ;
        RECT 74.100 103.180 74.360 103.500 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 62.130 88.870 62.410 89.170 ;
        RECT 54.840 88.480 56.750 88.620 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 88.480 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 74.160 89.170 74.300 103.180 ;
        RECT 76.880 102.305 78.760 102.675 ;
        RECT 80.140 89.170 80.280 106.240 ;
        RECT 86.580 104.180 86.720 106.240 ;
        RECT 86.520 103.860 86.780 104.180 ;
        RECT 87.960 103.500 88.100 108.280 ;
        RECT 93.020 107.240 93.160 108.280 ;
        RECT 93.880 107.260 94.140 107.580 ;
        RECT 92.960 106.920 93.220 107.240 ;
        RECT 88.360 105.560 88.620 105.880 ;
        RECT 88.420 104.180 88.560 105.560 ;
        RECT 91.880 105.025 93.760 105.395 ;
        RECT 88.360 103.860 88.620 104.180 ;
        RECT 86.980 103.180 87.240 103.500 ;
        RECT 87.900 103.180 88.160 103.500 ;
        RECT 74.090 88.160 74.370 89.170 ;
        RECT 80.070 88.180 80.350 89.170 ;
        RECT 86.050 88.620 86.330 89.170 ;
        RECT 87.040 88.620 87.180 103.180 ;
        RECT 91.880 99.585 93.760 99.955 ;
        RECT 86.050 88.480 87.180 88.620 ;
        RECT 92.030 88.620 92.310 89.170 ;
        RECT 93.940 88.620 94.080 107.260 ;
        RECT 98.080 107.240 98.220 108.280 ;
        RECT 98.020 106.920 98.280 107.240 ;
        RECT 99.400 106.240 99.660 106.560 ;
        RECT 97.560 105.560 97.820 105.880 ;
        RECT 97.620 101.800 97.760 105.560 ;
        RECT 99.460 104.180 99.600 106.240 ;
        RECT 99.400 103.860 99.660 104.180 ;
        RECT 97.560 101.480 97.820 101.800 ;
        RECT 99.460 101.120 99.600 103.860 ;
        RECT 99.920 101.800 100.060 108.280 ;
        RECT 102.680 106.900 102.820 108.620 ;
        RECT 109.520 108.280 109.780 108.600 ;
        RECT 106.880 107.745 108.760 108.115 ;
        RECT 109.060 107.260 109.320 107.580 ;
        RECT 102.620 106.580 102.880 106.900 ;
        RECT 104.460 105.560 104.720 105.880 ;
        RECT 104.520 103.500 104.660 105.560 ;
        RECT 104.000 103.180 104.260 103.500 ;
        RECT 104.460 103.180 104.720 103.500 ;
        RECT 99.860 101.480 100.120 101.800 ;
        RECT 98.020 100.800 98.280 101.120 ;
        RECT 99.400 100.800 99.660 101.120 ;
        RECT 98.080 89.170 98.220 100.800 ;
        RECT 104.060 89.170 104.200 103.180 ;
        RECT 106.880 102.305 108.760 102.675 ;
        RECT 109.120 98.140 109.260 107.260 ;
        RECT 109.580 107.240 109.720 108.280 ;
        RECT 109.520 106.920 109.780 107.240 ;
        RECT 110.960 104.180 111.100 109.640 ;
        RECT 111.420 109.280 111.560 128.600 ;
        RECT 112.340 125.510 112.480 130.720 ;
        RECT 118.320 128.660 118.460 131.400 ;
        RECT 113.200 128.340 113.460 128.660 ;
        RECT 118.260 128.340 118.520 128.660 ;
        RECT 112.340 125.370 112.940 125.510 ;
        RECT 112.800 123.220 112.940 125.370 ;
        RECT 113.260 124.920 113.400 128.340 ;
        RECT 115.040 128.000 115.300 128.320 ;
        RECT 115.100 126.620 115.240 128.000 ;
        RECT 115.040 126.300 115.300 126.620 ;
        RECT 113.660 125.620 113.920 125.940 ;
        RECT 113.200 124.600 113.460 124.920 ;
        RECT 113.260 123.560 113.400 124.600 ;
        RECT 113.200 123.240 113.460 123.560 ;
        RECT 112.740 122.900 113.000 123.220 ;
        RECT 111.820 119.160 112.080 119.480 ;
        RECT 111.880 117.780 112.020 119.160 ;
        RECT 111.820 117.460 112.080 117.780 ;
        RECT 111.880 113.020 112.020 117.460 ;
        RECT 112.800 115.060 112.940 122.900 ;
        RECT 113.720 122.880 113.860 125.620 ;
        RECT 113.660 122.790 113.920 122.880 ;
        RECT 113.260 122.650 113.920 122.790 ;
        RECT 113.260 115.400 113.400 122.650 ;
        RECT 113.660 122.560 113.920 122.650 ;
        RECT 116.420 119.840 116.680 120.160 ;
        RECT 118.320 120.070 118.460 128.340 ;
        RECT 118.720 127.320 118.980 127.640 ;
        RECT 120.560 127.320 120.820 127.640 ;
        RECT 118.780 125.260 118.920 127.320 ;
        RECT 120.620 125.940 120.760 127.320 ;
        RECT 121.880 126.785 123.760 127.155 ;
        RECT 120.560 125.620 120.820 125.940 ;
        RECT 124.760 125.600 124.900 138.200 ;
        RECT 129.140 138.175 134.100 139.455 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 124.700 125.280 124.960 125.600 ;
        RECT 118.720 124.940 118.980 125.260 ;
        RECT 119.180 123.240 119.440 123.560 ;
        RECT 119.240 121.180 119.380 123.240 ;
        RECT 124.760 123.220 124.900 125.280 ;
        RECT 124.700 122.900 124.960 123.220 ;
        RECT 121.480 122.560 121.740 122.880 ;
        RECT 120.560 121.880 120.820 122.200 ;
        RECT 119.180 120.860 119.440 121.180 ;
        RECT 120.620 120.160 120.760 121.880 ;
        RECT 121.540 121.180 121.680 122.560 ;
        RECT 121.880 121.345 123.760 121.715 ;
        RECT 121.480 120.860 121.740 121.180 ;
        RECT 118.720 120.070 118.980 120.160 ;
        RECT 118.320 119.930 118.980 120.070 ;
        RECT 113.660 119.500 113.920 119.820 ;
        RECT 113.720 118.460 113.860 119.500 ;
        RECT 116.480 118.460 116.620 119.840 ;
        RECT 113.660 118.140 113.920 118.460 ;
        RECT 116.420 118.140 116.680 118.460 ;
        RECT 118.320 118.120 118.460 119.930 ;
        RECT 118.720 119.840 118.980 119.930 ;
        RECT 120.560 119.840 120.820 120.160 ;
        RECT 118.260 117.800 118.520 118.120 ;
        RECT 115.500 117.460 115.760 117.780 ;
        RECT 115.560 115.740 115.700 117.460 ;
        RECT 121.880 115.905 123.760 116.275 ;
        RECT 115.500 115.420 115.760 115.740 ;
        RECT 113.200 115.080 113.460 115.400 ;
        RECT 112.740 114.740 113.000 115.060 ;
        RECT 121.940 113.720 122.200 114.040 ;
        RECT 111.820 112.700 112.080 113.020 ;
        RECT 117.340 112.700 117.600 113.020 ;
        RECT 111.880 109.960 112.020 112.700 ;
        RECT 111.820 109.640 112.080 109.960 ;
        RECT 111.360 108.960 111.620 109.280 ;
        RECT 111.360 108.280 111.620 108.600 ;
        RECT 111.420 107.240 111.560 108.280 ;
        RECT 111.360 106.920 111.620 107.240 ;
        RECT 111.880 106.980 112.020 109.640 ;
        RECT 114.120 108.280 114.380 108.600 ;
        RECT 116.420 108.280 116.680 108.600 ;
        RECT 111.880 106.840 112.480 106.980 ;
        RECT 112.340 106.560 112.480 106.840 ;
        RECT 112.280 106.240 112.540 106.560 ;
        RECT 112.340 104.180 112.480 106.240 ;
        RECT 114.180 104.180 114.320 108.280 ;
        RECT 110.900 103.860 111.160 104.180 ;
        RECT 112.280 103.860 112.540 104.180 ;
        RECT 114.120 103.860 114.380 104.180 ;
        RECT 115.960 103.860 116.220 104.180 ;
        RECT 109.120 98.000 110.180 98.140 ;
        RECT 110.040 89.290 110.180 98.000 ;
        RECT 116.020 89.570 116.160 103.860 ;
        RECT 116.480 103.500 116.620 108.280 ;
        RECT 117.400 107.240 117.540 112.700 ;
        RECT 119.180 112.360 119.440 112.680 ;
        RECT 119.240 109.620 119.380 112.360 ;
        RECT 122.000 112.340 122.140 113.720 ;
        RECT 119.640 112.020 119.900 112.340 ;
        RECT 121.940 112.020 122.200 112.340 ;
        RECT 119.180 109.300 119.440 109.620 ;
        RECT 119.180 108.510 119.440 108.600 ;
        RECT 119.700 108.510 119.840 112.020 ;
        RECT 120.100 111.680 120.360 112.000 ;
        RECT 120.160 108.940 120.300 111.680 ;
        RECT 121.880 110.465 123.760 110.835 ;
        RECT 120.100 108.620 120.360 108.940 ;
        RECT 127.920 108.620 128.180 108.940 ;
        RECT 119.180 108.370 119.840 108.510 ;
        RECT 119.180 108.280 119.440 108.370 ;
        RECT 117.340 106.920 117.600 107.240 ;
        RECT 116.420 103.180 116.680 103.500 ;
        RECT 119.700 101.460 119.840 108.370 ;
        RECT 120.100 106.920 120.360 107.240 ;
        RECT 120.160 102.140 120.300 106.920 ;
        RECT 121.020 106.240 121.280 106.560 ;
        RECT 120.100 101.820 120.360 102.140 ;
        RECT 119.640 101.140 119.900 101.460 ;
        RECT 121.080 98.820 121.220 106.240 ;
        RECT 126.070 106.045 126.350 106.415 ;
        RECT 121.880 105.025 123.760 105.395 ;
        RECT 126.140 103.840 126.280 106.045 ;
        RECT 126.080 103.520 126.340 103.840 ;
        RECT 121.880 99.585 123.760 99.955 ;
        RECT 121.080 98.680 122.140 98.820 ;
        RECT 122.000 89.570 122.140 98.680 ;
        RECT 92.030 88.480 94.080 88.620 ;
        RECT 98.010 88.500 98.290 89.170 ;
        RECT 103.990 88.610 104.270 89.170 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 86.050 87.970 86.330 88.480 ;
        RECT 92.030 88.320 92.310 88.480 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.500 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 127.980 89.380 128.120 108.620 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 16.830 211.125 18.810 211.455 ;
        RECT 46.830 211.125 48.810 211.455 ;
        RECT 76.830 211.125 78.810 211.455 ;
        RECT 106.830 211.125 108.810 211.455 ;
        RECT 31.830 208.405 33.810 208.735 ;
        RECT 61.830 208.405 63.810 208.735 ;
        RECT 91.830 208.405 93.810 208.735 ;
        RECT 121.830 208.405 123.810 208.735 ;
        RECT 16.830 205.685 18.810 206.015 ;
        RECT 46.830 205.685 48.810 206.015 ;
        RECT 76.830 205.685 78.810 206.015 ;
        RECT 106.830 205.685 108.810 206.015 ;
        RECT 31.830 202.965 33.810 203.295 ;
        RECT 61.830 202.965 63.810 203.295 ;
        RECT 91.830 202.965 93.810 203.295 ;
        RECT 121.830 202.965 123.810 203.295 ;
        RECT 16.830 200.245 18.810 200.575 ;
        RECT 46.830 200.245 48.810 200.575 ;
        RECT 76.830 200.245 78.810 200.575 ;
        RECT 106.830 200.245 108.810 200.575 ;
        RECT 31.830 197.525 33.810 197.855 ;
        RECT 61.830 197.525 63.810 197.855 ;
        RECT 91.830 197.525 93.810 197.855 ;
        RECT 121.830 197.525 123.810 197.855 ;
        RECT 16.830 194.805 18.810 195.135 ;
        RECT 46.830 194.805 48.810 195.135 ;
        RECT 76.830 194.805 78.810 195.135 ;
        RECT 106.830 194.805 108.810 195.135 ;
        RECT 31.830 192.085 33.810 192.415 ;
        RECT 61.830 192.085 63.810 192.415 ;
        RECT 91.830 192.085 93.810 192.415 ;
        RECT 121.830 192.085 123.810 192.415 ;
        RECT 16.830 189.365 18.810 189.695 ;
        RECT 46.830 189.365 48.810 189.695 ;
        RECT 76.830 189.365 78.810 189.695 ;
        RECT 106.830 189.365 108.810 189.695 ;
        RECT 44.370 187.980 44.750 187.990 ;
        RECT 55.665 187.980 55.995 187.995 ;
        RECT 44.370 187.680 55.995 187.980 ;
        RECT 44.370 187.670 44.750 187.680 ;
        RECT 55.665 187.665 55.995 187.680 ;
        RECT 94.765 187.980 95.095 187.995 ;
        RECT 98.650 187.980 99.030 187.990 ;
        RECT 94.765 187.680 99.030 187.980 ;
        RECT 94.765 187.665 95.095 187.680 ;
        RECT 98.650 187.670 99.030 187.680 ;
        RECT 31.830 186.645 33.810 186.975 ;
        RECT 61.830 186.645 63.810 186.975 ;
        RECT 91.830 186.645 93.810 186.975 ;
        RECT 121.830 186.645 123.810 186.975 ;
        RECT 16.830 183.925 18.810 184.255 ;
        RECT 46.830 183.925 48.810 184.255 ;
        RECT 76.830 183.925 78.810 184.255 ;
        RECT 106.830 183.925 108.810 184.255 ;
        RECT 31.830 181.205 33.810 181.535 ;
        RECT 61.830 181.205 63.810 181.535 ;
        RECT 91.830 181.205 93.810 181.535 ;
        RECT 121.830 181.205 123.810 181.535 ;
        RECT 40.485 179.820 40.815 179.835 ;
        RECT 41.865 179.820 42.195 179.835 ;
        RECT 67.625 179.820 67.955 179.835 ;
        RECT 40.485 179.520 67.955 179.820 ;
        RECT 40.485 179.505 40.815 179.520 ;
        RECT 41.865 179.505 42.195 179.520 ;
        RECT 67.625 179.505 67.955 179.520 ;
        RECT 78.665 179.820 78.995 179.835 ;
        RECT 85.105 179.820 85.435 179.835 ;
        RECT 78.665 179.520 85.435 179.820 ;
        RECT 78.665 179.505 78.995 179.520 ;
        RECT 85.105 179.505 85.435 179.520 ;
        RECT 16.830 178.485 18.810 178.815 ;
        RECT 46.830 178.485 48.810 178.815 ;
        RECT 76.830 178.485 78.810 178.815 ;
        RECT 106.830 178.485 108.810 178.815 ;
        RECT 66.245 177.780 66.575 177.795 ;
        RECT 70.385 177.780 70.715 177.795 ;
        RECT 72.685 177.780 73.015 177.795 ;
        RECT 66.245 177.480 73.015 177.780 ;
        RECT 66.245 177.465 66.575 177.480 ;
        RECT 70.385 177.465 70.715 177.480 ;
        RECT 72.685 177.465 73.015 177.480 ;
        RECT 71.765 177.100 72.095 177.115 ;
        RECT 78.205 177.100 78.535 177.115 ;
        RECT 71.765 176.800 78.535 177.100 ;
        RECT 71.765 176.785 72.095 176.800 ;
        RECT 78.205 176.785 78.535 176.800 ;
        RECT 31.830 175.765 33.810 176.095 ;
        RECT 61.830 175.765 63.810 176.095 ;
        RECT 91.830 175.765 93.810 176.095 ;
        RECT 121.830 175.765 123.810 176.095 ;
        RECT 40.025 175.060 40.355 175.075 ;
        RECT 65.325 175.060 65.655 175.075 ;
        RECT 40.025 174.760 65.655 175.060 ;
        RECT 40.025 174.745 40.355 174.760 ;
        RECT 65.325 174.745 65.655 174.760 ;
        RECT 54.745 174.380 55.075 174.395 ;
        RECT 63.025 174.380 63.355 174.395 ;
        RECT 54.745 174.080 63.355 174.380 ;
        RECT 54.745 174.065 55.075 174.080 ;
        RECT 63.025 174.065 63.355 174.080 ;
        RECT 16.830 173.045 18.810 173.375 ;
        RECT 46.830 173.045 48.810 173.375 ;
        RECT 76.830 173.045 78.810 173.375 ;
        RECT 106.830 173.045 108.810 173.375 ;
        RECT 127.885 171.660 128.215 171.675 ;
        RECT 129.240 171.660 133.810 172.125 ;
        RECT 127.885 171.360 133.810 171.660 ;
        RECT 127.885 171.345 128.215 171.360 ;
        RECT 31.830 170.325 33.810 170.655 ;
        RECT 61.830 170.325 63.810 170.655 ;
        RECT 91.830 170.325 93.810 170.655 ;
        RECT 121.830 170.325 123.810 170.655 ;
        RECT 129.240 170.585 133.810 171.360 ;
        RECT 44.165 169.630 44.495 169.635 ;
        RECT 44.165 169.620 44.750 169.630 ;
        RECT 43.940 169.320 44.750 169.620 ;
        RECT 44.165 169.310 44.750 169.320 ;
        RECT 44.165 169.305 44.495 169.310 ;
        RECT 16.830 167.605 18.810 167.935 ;
        RECT 46.830 167.605 48.810 167.935 ;
        RECT 76.830 167.605 78.810 167.935 ;
        RECT 106.830 167.605 108.810 167.935 ;
        RECT 31.830 164.885 33.810 165.215 ;
        RECT 61.830 164.885 63.810 165.215 ;
        RECT 91.830 164.885 93.810 165.215 ;
        RECT 121.830 164.885 123.810 165.215 ;
        RECT 94.970 164.180 95.350 164.190 ;
        RECT 98.650 164.180 99.030 164.190 ;
        RECT 101.205 164.180 101.535 164.195 ;
        RECT 94.970 163.880 101.535 164.180 ;
        RECT 94.970 163.870 95.350 163.880 ;
        RECT 98.650 163.870 99.030 163.880 ;
        RECT 101.205 163.865 101.535 163.880 ;
        RECT 16.830 162.165 18.810 162.495 ;
        RECT 46.830 162.165 48.810 162.495 ;
        RECT 76.830 162.165 78.810 162.495 ;
        RECT 106.830 162.165 108.810 162.495 ;
        RECT 31.830 159.445 33.810 159.775 ;
        RECT 61.830 159.445 63.810 159.775 ;
        RECT 91.830 159.445 93.810 159.775 ;
        RECT 121.830 159.445 123.810 159.775 ;
        RECT 80.045 159.420 80.375 159.435 ;
        RECT 81.425 159.420 81.755 159.435 ;
        RECT 80.045 159.120 81.755 159.420 ;
        RECT 80.045 159.105 80.375 159.120 ;
        RECT 81.425 159.105 81.755 159.120 ;
        RECT 68.085 158.740 68.415 158.755 ;
        RECT 71.765 158.740 72.095 158.755 ;
        RECT 84.645 158.740 84.975 158.755 ;
        RECT 68.085 158.440 84.975 158.740 ;
        RECT 68.085 158.425 68.415 158.440 ;
        RECT 71.765 158.425 72.095 158.440 ;
        RECT 84.645 158.425 84.975 158.440 ;
        RECT 16.830 156.725 18.810 157.055 ;
        RECT 46.830 156.725 48.810 157.055 ;
        RECT 76.830 156.725 78.810 157.055 ;
        RECT 106.830 156.725 108.810 157.055 ;
        RECT 73.145 156.700 73.475 156.715 ;
        RECT 75.445 156.700 75.775 156.715 ;
        RECT 73.145 156.400 75.775 156.700 ;
        RECT 73.145 156.385 73.475 156.400 ;
        RECT 75.445 156.385 75.775 156.400 ;
        RECT 41.865 156.020 42.195 156.035 ;
        RECT 43.245 156.020 43.575 156.035 ;
        RECT 94.970 156.020 95.350 156.030 ;
        RECT 41.865 155.720 43.575 156.020 ;
        RECT 41.865 155.705 42.195 155.720 ;
        RECT 43.245 155.705 43.575 155.720 ;
        RECT 71.090 155.720 95.350 156.020 ;
        RECT 44.370 155.340 44.750 155.350 ;
        RECT 65.785 155.340 66.115 155.355 ;
        RECT 71.090 155.340 71.390 155.720 ;
        RECT 94.970 155.710 95.350 155.720 ;
        RECT 44.370 155.040 71.390 155.340 ;
        RECT 74.525 155.340 74.855 155.355 ;
        RECT 112.450 155.340 112.830 155.350 ;
        RECT 74.525 155.040 112.830 155.340 ;
        RECT 44.370 155.030 44.750 155.040 ;
        RECT 65.785 155.025 66.115 155.040 ;
        RECT 74.525 155.025 74.855 155.040 ;
        RECT 112.450 155.030 112.830 155.040 ;
        RECT 31.830 154.005 33.810 154.335 ;
        RECT 61.830 154.005 63.810 154.335 ;
        RECT 91.830 154.005 93.810 154.335 ;
        RECT 121.830 154.005 123.810 154.335 ;
        RECT 44.625 152.620 44.955 152.635 ;
        RECT 68.085 152.620 68.415 152.635 ;
        RECT 44.625 152.320 68.415 152.620 ;
        RECT 44.625 152.305 44.955 152.320 ;
        RECT 68.085 152.305 68.415 152.320 ;
        RECT 16.830 151.285 18.810 151.615 ;
        RECT 46.830 151.285 48.810 151.615 ;
        RECT 76.830 151.285 78.810 151.615 ;
        RECT 106.830 151.285 108.810 151.615 ;
        RECT 87.865 150.580 88.195 150.595 ;
        RECT 99.365 150.580 99.695 150.595 ;
        RECT 107.645 150.580 107.975 150.595 ;
        RECT 87.865 150.280 107.975 150.580 ;
        RECT 87.865 150.265 88.195 150.280 ;
        RECT 99.365 150.265 99.695 150.280 ;
        RECT 107.645 150.265 107.975 150.280 ;
        RECT 31.830 148.565 33.810 148.895 ;
        RECT 61.830 148.565 63.810 148.895 ;
        RECT 91.830 148.565 93.810 148.895 ;
        RECT 121.830 148.565 123.810 148.895 ;
        RECT 16.830 145.845 18.810 146.175 ;
        RECT 46.830 145.845 48.810 146.175 ;
        RECT 76.830 145.845 78.810 146.175 ;
        RECT 106.830 145.845 108.810 146.175 ;
        RECT 31.830 143.125 33.810 143.455 ;
        RECT 61.830 143.125 63.810 143.455 ;
        RECT 91.830 143.125 93.810 143.455 ;
        RECT 121.830 143.125 123.810 143.455 ;
        RECT 16.830 140.405 18.810 140.735 ;
        RECT 46.830 140.405 48.810 140.735 ;
        RECT 76.830 140.405 78.810 140.735 ;
        RECT 106.830 140.405 108.810 140.735 ;
        RECT 112.450 139.020 112.830 139.030 ;
        RECT 129.090 139.020 134.150 139.430 ;
        RECT 112.450 138.720 134.150 139.020 ;
        RECT 112.450 138.710 112.830 138.720 ;
        RECT 129.090 138.200 134.150 138.720 ;
        RECT 31.830 137.685 33.810 138.015 ;
        RECT 61.830 137.685 63.810 138.015 ;
        RECT 91.830 137.685 93.810 138.015 ;
        RECT 121.830 137.685 123.810 138.015 ;
        RECT 16.830 134.965 18.810 135.295 ;
        RECT 46.830 134.965 48.810 135.295 ;
        RECT 76.830 134.965 78.810 135.295 ;
        RECT 106.830 134.965 108.810 135.295 ;
        RECT 99.365 134.260 99.695 134.275 ;
        RECT 108.105 134.260 108.435 134.275 ;
        RECT 99.365 133.960 108.435 134.260 ;
        RECT 99.365 133.945 99.695 133.960 ;
        RECT 108.105 133.945 108.435 133.960 ;
        RECT 31.830 132.245 33.810 132.575 ;
        RECT 61.830 132.245 63.810 132.575 ;
        RECT 91.830 132.245 93.810 132.575 ;
        RECT 121.830 132.245 123.810 132.575 ;
        RECT 44.370 132.220 44.750 132.230 ;
        RECT 49.225 132.220 49.555 132.235 ;
        RECT 44.370 131.920 49.555 132.220 ;
        RECT 44.370 131.910 44.750 131.920 ;
        RECT 49.225 131.905 49.555 131.920 ;
        RECT 16.830 129.525 18.810 129.855 ;
        RECT 46.830 129.525 48.810 129.855 ;
        RECT 76.830 129.525 78.810 129.855 ;
        RECT 106.830 129.525 108.810 129.855 ;
        RECT 94.970 129.500 95.350 129.510 ;
        RECT 95.685 129.500 96.015 129.515 ;
        RECT 94.970 129.200 96.015 129.500 ;
        RECT 94.970 129.190 95.350 129.200 ;
        RECT 95.685 129.185 96.015 129.200 ;
        RECT 31.830 126.805 33.810 127.135 ;
        RECT 61.830 126.805 63.810 127.135 ;
        RECT 91.830 126.805 93.810 127.135 ;
        RECT 121.830 126.805 123.810 127.135 ;
        RECT 16.830 124.085 18.810 124.415 ;
        RECT 46.830 124.085 48.810 124.415 ;
        RECT 76.830 124.085 78.810 124.415 ;
        RECT 106.830 124.085 108.810 124.415 ;
        RECT 31.830 121.365 33.810 121.695 ;
        RECT 61.830 121.365 63.810 121.695 ;
        RECT 91.830 121.365 93.810 121.695 ;
        RECT 121.830 121.365 123.810 121.695 ;
        RECT 16.830 118.645 18.810 118.975 ;
        RECT 46.830 118.645 48.810 118.975 ;
        RECT 76.830 118.645 78.810 118.975 ;
        RECT 106.830 118.645 108.810 118.975 ;
        RECT 31.830 115.925 33.810 116.255 ;
        RECT 61.830 115.925 63.810 116.255 ;
        RECT 91.830 115.925 93.810 116.255 ;
        RECT 121.830 115.925 123.810 116.255 ;
        RECT 16.830 113.205 18.810 113.535 ;
        RECT 46.830 113.205 48.810 113.535 ;
        RECT 76.830 113.205 78.810 113.535 ;
        RECT 106.830 113.205 108.810 113.535 ;
        RECT 92.925 113.180 93.255 113.195 ;
        RECT 94.970 113.180 95.350 113.190 ;
        RECT 92.925 112.880 95.350 113.180 ;
        RECT 92.925 112.865 93.255 112.880 ;
        RECT 94.970 112.870 95.350 112.880 ;
        RECT 31.830 110.485 33.810 110.815 ;
        RECT 61.830 110.485 63.810 110.815 ;
        RECT 91.830 110.485 93.810 110.815 ;
        RECT 121.830 110.485 123.810 110.815 ;
        RECT 16.830 107.765 18.810 108.095 ;
        RECT 46.830 107.765 48.810 108.095 ;
        RECT 76.830 107.765 78.810 108.095 ;
        RECT 106.830 107.765 108.810 108.095 ;
        RECT 129.700 106.530 133.210 106.625 ;
        RECT 126.045 106.380 126.375 106.395 ;
        RECT 129.700 106.380 133.340 106.530 ;
        RECT 126.045 106.080 133.340 106.380 ;
        RECT 126.045 106.065 126.375 106.080 ;
        RECT 129.700 105.930 133.340 106.080 ;
        RECT 129.700 105.605 133.210 105.930 ;
        RECT 31.830 105.045 33.810 105.375 ;
        RECT 61.830 105.045 63.810 105.375 ;
        RECT 91.830 105.045 93.810 105.375 ;
        RECT 121.830 105.045 123.810 105.375 ;
        RECT 16.830 102.325 18.810 102.655 ;
        RECT 46.830 102.325 48.810 102.655 ;
        RECT 76.830 102.325 78.810 102.655 ;
        RECT 106.830 102.325 108.810 102.655 ;
        RECT 31.830 99.605 33.810 99.935 ;
        RECT 61.830 99.605 63.810 99.935 ;
        RECT 91.830 99.605 93.810 99.935 ;
        RECT 121.830 99.605 123.810 99.935 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 16.820 99.530 18.820 211.530 ;
        RECT 31.820 99.530 33.820 211.530 ;
        RECT 44.395 187.665 44.725 187.995 ;
        RECT 44.410 169.635 44.710 187.665 ;
        RECT 44.395 169.305 44.725 169.635 ;
        RECT 44.410 155.355 44.710 169.305 ;
        RECT 44.395 155.025 44.725 155.355 ;
        RECT 44.410 132.235 44.710 155.025 ;
        RECT 44.395 131.905 44.725 132.235 ;
        RECT 46.820 99.530 48.820 211.530 ;
        RECT 61.820 99.530 63.820 211.530 ;
        RECT 76.820 99.530 78.820 211.530 ;
        RECT 91.820 99.530 93.820 211.530 ;
        RECT 98.675 187.665 99.005 187.995 ;
        RECT 98.690 164.195 98.990 187.665 ;
        RECT 94.995 163.865 95.325 164.195 ;
        RECT 98.675 163.865 99.005 164.195 ;
        RECT 95.010 156.035 95.310 163.865 ;
        RECT 94.995 155.705 95.325 156.035 ;
        RECT 95.010 129.515 95.310 155.705 ;
        RECT 94.995 129.185 95.325 129.515 ;
        RECT 95.010 113.195 95.310 129.185 ;
        RECT 94.995 112.865 95.325 113.195 ;
        RECT 106.820 99.530 108.820 211.530 ;
        RECT 112.475 155.025 112.805 155.355 ;
        RECT 112.490 139.035 112.790 155.025 ;
        RECT 112.475 138.705 112.805 139.035 ;
        RECT 121.820 99.720 123.820 211.530 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

